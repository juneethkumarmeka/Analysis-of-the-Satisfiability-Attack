module basic_5000_50000_5000_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_476,In_706);
and U1 (N_1,In_635,In_964);
or U2 (N_2,In_1918,In_689);
nor U3 (N_3,In_3807,In_1105);
nor U4 (N_4,In_1397,In_4238);
and U5 (N_5,In_3370,In_2495);
xor U6 (N_6,In_3138,In_2188);
or U7 (N_7,In_857,In_3436);
nor U8 (N_8,In_2256,In_4511);
nand U9 (N_9,In_4298,In_3317);
nor U10 (N_10,In_1340,In_4290);
nor U11 (N_11,In_269,In_1400);
and U12 (N_12,In_4678,In_771);
and U13 (N_13,In_3506,In_4944);
and U14 (N_14,In_3028,In_4934);
or U15 (N_15,In_2328,In_553);
nor U16 (N_16,In_491,In_1941);
xor U17 (N_17,In_1141,In_32);
and U18 (N_18,In_1687,In_1963);
nand U19 (N_19,In_806,In_3795);
or U20 (N_20,In_4666,In_1878);
or U21 (N_21,In_1641,In_2402);
or U22 (N_22,In_4336,In_4959);
or U23 (N_23,In_236,In_3452);
or U24 (N_24,In_480,In_2194);
or U25 (N_25,In_4975,In_3832);
or U26 (N_26,In_4092,In_3803);
nor U27 (N_27,In_3380,In_4122);
and U28 (N_28,In_2906,In_3813);
nor U29 (N_29,In_2067,In_3220);
or U30 (N_30,In_4726,In_4854);
nor U31 (N_31,In_4228,In_636);
nor U32 (N_32,In_3110,In_1939);
nor U33 (N_33,In_3538,In_1143);
or U34 (N_34,In_2469,In_1860);
nand U35 (N_35,In_4328,In_240);
nand U36 (N_36,In_2204,In_3933);
xnor U37 (N_37,In_4019,In_2895);
nand U38 (N_38,In_3341,In_2455);
or U39 (N_39,In_2967,In_1311);
nor U40 (N_40,In_1779,In_2209);
nand U41 (N_41,In_2213,In_395);
nor U42 (N_42,In_1040,In_2387);
or U43 (N_43,In_472,In_902);
xnor U44 (N_44,In_1122,In_4299);
or U45 (N_45,In_270,In_4656);
xor U46 (N_46,In_452,In_2037);
nand U47 (N_47,In_330,In_3569);
and U48 (N_48,In_4296,In_844);
nand U49 (N_49,In_782,In_3804);
or U50 (N_50,In_1306,In_541);
or U51 (N_51,In_2656,In_4099);
nand U52 (N_52,In_1540,In_3109);
or U53 (N_53,In_1838,In_1415);
or U54 (N_54,In_1380,In_2480);
and U55 (N_55,In_4597,In_2279);
xor U56 (N_56,In_2274,In_2675);
and U57 (N_57,In_1693,In_4041);
and U58 (N_58,In_3505,In_4503);
nand U59 (N_59,In_3444,In_1383);
nand U60 (N_60,In_13,In_150);
or U61 (N_61,In_1926,In_2804);
xor U62 (N_62,In_781,In_246);
nor U63 (N_63,In_1973,In_2090);
or U64 (N_64,In_3197,In_744);
and U65 (N_65,In_2853,In_3327);
nand U66 (N_66,In_3481,In_2657);
nand U67 (N_67,In_302,In_3361);
nand U68 (N_68,In_2098,In_1901);
nand U69 (N_69,In_941,In_3586);
or U70 (N_70,In_83,In_1818);
xnor U71 (N_71,In_4512,In_3978);
xnor U72 (N_72,In_2169,In_226);
nor U73 (N_73,In_2710,In_4554);
xnor U74 (N_74,In_310,In_970);
or U75 (N_75,In_1822,In_4853);
nand U76 (N_76,In_2396,In_1549);
nor U77 (N_77,In_905,In_4948);
or U78 (N_78,In_2499,In_2549);
xnor U79 (N_79,In_2881,In_2702);
nor U80 (N_80,In_2034,In_3258);
nor U81 (N_81,In_1942,In_1735);
or U82 (N_82,In_3074,In_4356);
nor U83 (N_83,In_1757,In_2391);
nor U84 (N_84,In_1013,In_4060);
nand U85 (N_85,In_815,In_1534);
and U86 (N_86,In_4216,In_1845);
and U87 (N_87,In_3175,In_107);
and U88 (N_88,In_899,In_862);
nor U89 (N_89,In_3581,In_1153);
xor U90 (N_90,In_4237,In_2730);
nand U91 (N_91,In_2979,In_2844);
or U92 (N_92,In_758,In_897);
or U93 (N_93,In_2879,In_4081);
nand U94 (N_94,In_843,In_1676);
and U95 (N_95,In_8,In_3821);
and U96 (N_96,In_1607,In_3600);
nand U97 (N_97,In_776,In_4546);
nor U98 (N_98,In_2411,In_3130);
and U99 (N_99,In_45,In_1689);
and U100 (N_100,In_3720,In_872);
xnor U101 (N_101,In_4555,In_199);
or U102 (N_102,In_828,In_2557);
or U103 (N_103,In_4276,In_1185);
xor U104 (N_104,In_1323,In_4638);
nor U105 (N_105,In_2413,In_1982);
xnor U106 (N_106,In_2479,In_4493);
and U107 (N_107,In_365,In_3772);
nand U108 (N_108,In_1937,In_3364);
nor U109 (N_109,In_4773,In_4951);
or U110 (N_110,In_1189,In_3122);
or U111 (N_111,In_1423,In_2364);
nor U112 (N_112,In_455,In_4358);
nand U113 (N_113,In_529,In_1166);
xnor U114 (N_114,In_4892,In_2426);
or U115 (N_115,In_4365,In_2536);
nor U116 (N_116,In_1108,In_1571);
or U117 (N_117,In_3185,In_3292);
or U118 (N_118,In_2002,In_4942);
xnor U119 (N_119,In_2705,In_4603);
nand U120 (N_120,In_3542,In_1812);
or U121 (N_121,In_1979,In_438);
or U122 (N_122,In_1493,In_3412);
xor U123 (N_123,In_3771,In_3328);
nor U124 (N_124,In_4890,In_2636);
nand U125 (N_125,In_1039,In_1513);
nor U126 (N_126,In_4691,In_1191);
and U127 (N_127,In_1590,In_33);
nand U128 (N_128,In_304,In_1815);
or U129 (N_129,In_1900,In_2260);
and U130 (N_130,In_4132,In_3171);
xnor U131 (N_131,In_878,In_4794);
xor U132 (N_132,In_1770,In_4401);
or U133 (N_133,In_3209,In_2870);
nand U134 (N_134,In_3511,In_1242);
nor U135 (N_135,In_2239,In_850);
nor U136 (N_136,In_2872,In_4448);
nor U137 (N_137,In_4509,In_4725);
or U138 (N_138,In_313,In_4536);
nand U139 (N_139,In_170,In_3226);
and U140 (N_140,In_4883,In_2676);
and U141 (N_141,In_1318,In_2756);
and U142 (N_142,In_1624,In_4728);
nor U143 (N_143,In_1453,In_1849);
nand U144 (N_144,In_749,In_227);
and U145 (N_145,In_4158,In_1626);
nor U146 (N_146,In_2537,In_349);
nor U147 (N_147,In_3393,In_4592);
nor U148 (N_148,In_2379,In_4331);
nor U149 (N_149,In_3540,In_254);
nor U150 (N_150,In_2717,In_171);
or U151 (N_151,In_702,In_4736);
or U152 (N_152,In_954,In_1111);
xnor U153 (N_153,In_1581,In_2056);
xnor U154 (N_154,In_934,In_1281);
or U155 (N_155,In_2294,In_2024);
nor U156 (N_156,In_1562,In_698);
xnor U157 (N_157,In_2350,In_3354);
xnor U158 (N_158,In_3355,In_1649);
nor U159 (N_159,In_725,In_3023);
and U160 (N_160,In_4177,In_4961);
xor U161 (N_161,In_1042,In_3133);
nand U162 (N_162,In_3472,In_2227);
or U163 (N_163,In_1932,In_3667);
nand U164 (N_164,In_3950,In_62);
nor U165 (N_165,In_4413,In_3887);
xor U166 (N_166,In_4003,In_3627);
and U167 (N_167,In_1183,In_1091);
xor U168 (N_168,In_60,In_4861);
nand U169 (N_169,In_3104,In_223);
nor U170 (N_170,In_514,In_3866);
nor U171 (N_171,In_4306,In_3948);
xor U172 (N_172,In_2305,In_1407);
nand U173 (N_173,In_921,In_2613);
nor U174 (N_174,In_185,In_713);
nor U175 (N_175,In_3092,In_4841);
or U176 (N_176,In_1935,In_1519);
nor U177 (N_177,In_3943,In_2807);
xor U178 (N_178,In_4375,In_1269);
nor U179 (N_179,In_2370,In_235);
or U180 (N_180,In_3187,In_4540);
or U181 (N_181,In_4778,In_3683);
xor U182 (N_182,In_3124,In_4100);
xnor U183 (N_183,In_726,In_3874);
xnor U184 (N_184,In_2981,In_586);
and U185 (N_185,In_3811,In_3259);
nor U186 (N_186,In_3844,In_4250);
nor U187 (N_187,In_3886,In_943);
nand U188 (N_188,In_258,In_4325);
xnor U189 (N_189,In_3180,In_1221);
nand U190 (N_190,In_3075,In_1811);
and U191 (N_191,In_1328,In_1545);
nor U192 (N_192,In_539,In_4069);
nor U193 (N_193,In_1597,In_4095);
xnor U194 (N_194,In_3622,In_3806);
nand U195 (N_195,In_2538,In_3984);
or U196 (N_196,In_1637,In_1159);
or U197 (N_197,In_2437,In_3764);
or U198 (N_198,In_530,In_1120);
or U199 (N_199,In_383,In_1516);
nand U200 (N_200,In_63,In_3729);
and U201 (N_201,In_4741,In_3432);
or U202 (N_202,In_1241,In_2021);
nand U203 (N_203,In_1077,In_1988);
or U204 (N_204,In_204,In_4400);
or U205 (N_205,In_3402,In_4215);
nand U206 (N_206,In_1966,In_1686);
or U207 (N_207,In_1802,In_4247);
or U208 (N_208,In_648,In_1441);
and U209 (N_209,In_835,In_4478);
and U210 (N_210,In_1097,In_3789);
xnor U211 (N_211,In_4112,In_2162);
and U212 (N_212,In_1985,In_4192);
nand U213 (N_213,In_1448,In_2810);
nand U214 (N_214,In_238,In_1165);
nand U215 (N_215,In_111,In_3727);
nand U216 (N_216,In_1248,In_4538);
nand U217 (N_217,In_4836,In_149);
nand U218 (N_218,In_4779,In_4314);
and U219 (N_219,In_1186,In_2608);
or U220 (N_220,In_3006,In_1904);
and U221 (N_221,In_821,In_3993);
nand U222 (N_222,In_2755,In_1518);
nor U223 (N_223,In_2159,In_4798);
nor U224 (N_224,In_1222,In_1279);
nor U225 (N_225,In_1082,In_1007);
nand U226 (N_226,In_3952,In_4175);
or U227 (N_227,In_2514,In_2400);
nor U228 (N_228,In_1442,In_4915);
and U229 (N_229,In_1999,In_2569);
nand U230 (N_230,In_4024,In_2544);
nor U231 (N_231,In_3898,In_4991);
or U232 (N_232,In_4406,In_4548);
and U233 (N_233,In_230,In_4847);
nand U234 (N_234,In_1955,In_3639);
or U235 (N_235,In_4223,In_3188);
or U236 (N_236,In_3275,In_1520);
and U237 (N_237,In_4574,In_2018);
nand U238 (N_238,In_4218,In_3498);
nor U239 (N_239,In_3490,In_2088);
or U240 (N_240,In_677,In_3567);
nand U241 (N_241,In_181,In_1079);
and U242 (N_242,In_499,In_4838);
xor U243 (N_243,In_1215,In_2959);
and U244 (N_244,In_3514,In_1021);
xor U245 (N_245,In_3007,In_4360);
nor U246 (N_246,In_2956,In_1148);
nor U247 (N_247,In_4236,In_3775);
xnor U248 (N_248,In_3613,In_1219);
and U249 (N_249,In_4720,In_445);
xor U250 (N_250,In_3422,In_97);
or U251 (N_251,In_3616,In_601);
nor U252 (N_252,In_450,In_3946);
or U253 (N_253,In_3773,In_128);
or U254 (N_254,In_3920,In_913);
or U255 (N_255,In_4746,In_3815);
nand U256 (N_256,In_3870,In_3461);
nor U257 (N_257,In_217,In_94);
xor U258 (N_258,In_1156,In_3405);
nor U259 (N_259,In_1865,In_3283);
nand U260 (N_260,In_2697,In_1617);
and U261 (N_261,In_2834,In_4953);
or U262 (N_262,In_3636,In_3985);
nand U263 (N_263,In_858,In_2312);
xor U264 (N_264,In_2321,In_4050);
nor U265 (N_265,In_1911,In_2890);
nor U266 (N_266,In_3580,In_1214);
nor U267 (N_267,In_1876,In_2116);
or U268 (N_268,In_818,In_884);
nand U269 (N_269,In_1140,In_93);
or U270 (N_270,In_3375,In_2284);
nand U271 (N_271,In_66,In_2342);
and U272 (N_272,In_36,In_978);
nor U273 (N_273,In_3930,In_4186);
or U274 (N_274,In_82,In_443);
nand U275 (N_275,In_3377,In_4226);
and U276 (N_276,In_2992,In_1787);
and U277 (N_277,In_998,In_594);
nand U278 (N_278,In_2304,In_1868);
nor U279 (N_279,In_1987,In_72);
nor U280 (N_280,In_2818,In_192);
xnor U281 (N_281,In_1836,In_4895);
or U282 (N_282,In_3929,In_641);
nand U283 (N_283,In_2502,In_2242);
nand U284 (N_284,In_3239,In_3168);
or U285 (N_285,In_4026,In_3734);
nand U286 (N_286,In_947,In_1093);
or U287 (N_287,In_4542,In_2572);
and U288 (N_288,In_3923,In_2899);
nor U289 (N_289,In_4083,In_201);
and U290 (N_290,In_4197,In_1420);
nor U291 (N_291,In_4072,In_1043);
nor U292 (N_292,In_3536,In_699);
and U293 (N_293,In_4173,In_4008);
and U294 (N_294,In_183,In_1072);
or U295 (N_295,In_4471,In_1025);
nand U296 (N_296,In_1389,In_1605);
nand U297 (N_297,In_2798,In_1316);
or U298 (N_298,In_275,In_2443);
and U299 (N_299,In_1577,In_2078);
or U300 (N_300,In_2891,In_4430);
nor U301 (N_301,In_2662,In_2843);
xnor U302 (N_302,In_3382,In_1173);
xnor U303 (N_303,In_1983,In_1974);
xnor U304 (N_304,In_841,In_1862);
xnor U305 (N_305,In_95,In_3438);
nand U306 (N_306,In_2440,In_3421);
nor U307 (N_307,In_2434,In_1683);
nand U308 (N_308,In_622,In_3953);
nand U309 (N_309,In_1694,In_3647);
and U310 (N_310,In_1573,In_1743);
nor U311 (N_311,In_3853,In_3068);
and U312 (N_312,In_4234,In_2257);
and U313 (N_313,In_232,In_3704);
and U314 (N_314,In_4034,In_2679);
or U315 (N_315,In_4950,In_274);
nand U316 (N_316,In_2739,In_3424);
nor U317 (N_317,In_3052,In_4711);
or U318 (N_318,In_4229,In_3996);
and U319 (N_319,In_1890,In_2757);
and U320 (N_320,In_3686,In_2070);
and U321 (N_321,In_4823,In_2317);
nand U322 (N_322,In_487,In_3974);
xor U323 (N_323,In_1753,In_2471);
nor U324 (N_324,In_2000,In_697);
or U325 (N_325,In_3041,In_1413);
nor U326 (N_326,In_753,In_1629);
xor U327 (N_327,In_4149,In_669);
nor U328 (N_328,In_305,In_3169);
and U329 (N_329,In_396,In_1582);
nand U330 (N_330,In_4167,In_1633);
and U331 (N_331,In_103,In_271);
nor U332 (N_332,In_4363,In_4465);
nand U333 (N_333,In_1182,In_2991);
or U334 (N_334,In_3696,In_1895);
nand U335 (N_335,In_2190,In_653);
and U336 (N_336,In_2047,In_390);
nand U337 (N_337,In_4289,In_4202);
nand U338 (N_338,In_2850,In_566);
xnor U339 (N_339,In_1384,In_2822);
nand U340 (N_340,In_1579,In_3409);
nor U341 (N_341,In_4117,In_2029);
nand U342 (N_342,In_3918,In_1347);
or U343 (N_343,In_2545,In_168);
nand U344 (N_344,In_666,In_1919);
or U345 (N_345,In_1738,In_4687);
nand U346 (N_346,In_3280,In_3644);
nand U347 (N_347,In_521,In_2652);
and U348 (N_348,In_3423,In_3758);
nand U349 (N_349,In_2405,In_3570);
or U350 (N_350,In_2425,In_4402);
and U351 (N_351,In_21,In_1501);
nor U352 (N_352,In_2156,In_3598);
or U353 (N_353,In_2582,In_3206);
nor U354 (N_354,In_2735,In_4071);
nand U355 (N_355,In_4119,In_4379);
or U356 (N_356,In_2165,In_1555);
xnor U357 (N_357,In_531,In_2158);
or U358 (N_358,In_4923,In_2759);
or U359 (N_359,In_2362,In_4939);
nor U360 (N_360,In_3102,In_2193);
or U361 (N_361,In_827,In_986);
nand U362 (N_362,In_4452,In_4450);
xor U363 (N_363,In_422,In_879);
or U364 (N_364,In_4813,In_3013);
nand U365 (N_365,In_3332,In_4253);
xor U366 (N_366,In_1051,In_2408);
nand U367 (N_367,In_4749,In_705);
xnor U368 (N_368,In_757,In_4464);
nor U369 (N_369,In_626,In_163);
and U370 (N_370,In_4984,In_3396);
nand U371 (N_371,In_2310,In_3817);
or U372 (N_372,In_4333,In_4058);
nor U373 (N_373,In_1760,In_3491);
xor U374 (N_374,In_1533,In_939);
or U375 (N_375,In_4907,In_822);
xnor U376 (N_376,In_516,In_3040);
and U377 (N_377,In_4947,In_4433);
and U378 (N_378,In_3135,In_3851);
nor U379 (N_379,In_3414,In_3687);
xor U380 (N_380,In_1702,In_3043);
xor U381 (N_381,In_585,In_606);
or U382 (N_382,In_4272,In_2873);
nand U383 (N_383,In_3921,In_4482);
or U384 (N_384,In_1107,In_378);
nor U385 (N_385,In_1695,In_4013);
or U386 (N_386,In_4703,In_4805);
nand U387 (N_387,In_1038,In_4629);
nor U388 (N_388,In_392,In_4976);
nand U389 (N_389,In_4994,In_52);
nand U390 (N_390,In_4206,In_4302);
or U391 (N_391,In_3562,In_4874);
nand U392 (N_392,In_3493,In_3010);
nand U393 (N_393,In_4618,In_4563);
nand U394 (N_394,In_382,In_565);
xor U395 (N_395,In_715,In_89);
xor U396 (N_396,In_2752,In_1368);
nor U397 (N_397,In_3685,In_4270);
nor U398 (N_398,In_4801,In_3193);
or U399 (N_399,In_4369,In_4284);
nand U400 (N_400,In_1841,In_3208);
and U401 (N_401,In_2994,In_3891);
nor U402 (N_402,In_115,In_662);
and U403 (N_403,In_2688,In_9);
and U404 (N_404,In_2179,In_4098);
nor U405 (N_405,In_424,In_4374);
and U406 (N_406,In_583,In_267);
or U407 (N_407,In_4326,In_4475);
nor U408 (N_408,In_4431,In_1280);
and U409 (N_409,In_3750,In_2199);
nor U410 (N_410,In_2496,In_889);
nor U411 (N_411,In_1313,In_2394);
nand U412 (N_412,In_2973,In_239);
and U413 (N_413,In_4224,In_2417);
xnor U414 (N_414,In_4561,In_3822);
nand U415 (N_415,In_3583,In_3922);
or U416 (N_416,In_2222,In_3682);
nand U417 (N_417,In_2921,In_3033);
xnor U418 (N_418,In_4731,In_629);
nor U419 (N_419,In_2650,In_1833);
xnor U420 (N_420,In_3205,In_3352);
or U421 (N_421,In_888,In_1503);
nand U422 (N_422,In_214,In_2064);
xnor U423 (N_423,In_2949,In_1471);
and U424 (N_424,In_831,In_3417);
nand U425 (N_425,In_710,In_4172);
and U426 (N_426,In_2285,In_2847);
xnor U427 (N_427,In_647,In_2201);
and U428 (N_428,In_1485,In_2280);
xor U429 (N_429,In_724,In_1658);
nor U430 (N_430,In_3609,In_4665);
or U431 (N_431,In_1668,In_1056);
xnor U432 (N_432,In_2725,In_665);
or U433 (N_433,In_2237,In_1224);
nand U434 (N_434,In_1099,In_2039);
or U435 (N_435,In_3427,In_1132);
xnor U436 (N_436,In_965,In_4004);
nand U437 (N_437,In_4604,In_3190);
nand U438 (N_438,In_3016,In_1612);
and U439 (N_439,In_1490,In_4266);
nor U440 (N_440,In_3167,In_875);
nand U441 (N_441,In_2183,In_2344);
nand U442 (N_442,In_2205,In_4411);
or U443 (N_443,In_3961,In_4123);
xor U444 (N_444,In_4911,In_602);
xor U445 (N_445,In_2664,In_2111);
xor U446 (N_446,In_2628,In_4851);
nand U447 (N_447,In_754,In_4021);
or U448 (N_448,In_1664,In_4631);
nor U449 (N_449,In_1650,In_3534);
and U450 (N_450,In_167,In_4766);
and U451 (N_451,In_2011,In_1160);
and U452 (N_452,In_2773,In_524);
and U453 (N_453,In_3661,In_208);
xor U454 (N_454,In_4899,In_837);
and U455 (N_455,In_4040,In_3966);
nor U456 (N_456,In_3757,In_2858);
nand U457 (N_457,In_4639,In_3914);
xnor U458 (N_458,In_2678,In_2811);
nand U459 (N_459,In_3722,In_1619);
xnor U460 (N_460,In_381,In_1139);
nand U461 (N_461,In_2987,In_3501);
nor U462 (N_462,In_540,In_447);
and U463 (N_463,In_3294,In_1986);
xnor U464 (N_464,In_3854,In_4125);
nor U465 (N_465,In_2905,In_2734);
xnor U466 (N_466,In_4190,In_4097);
nor U467 (N_467,In_1741,In_4045);
or U468 (N_468,In_4865,In_4646);
nor U469 (N_469,In_1899,In_2916);
nor U470 (N_470,In_2917,In_1152);
nand U471 (N_471,In_4116,In_3499);
nor U472 (N_472,In_2290,In_2420);
xor U473 (N_473,In_1045,In_3211);
nand U474 (N_474,In_1925,In_2065);
nor U475 (N_475,In_960,In_3991);
or U476 (N_476,In_2030,In_130);
xor U477 (N_477,In_222,In_1526);
nand U478 (N_478,In_1290,In_2673);
nand U479 (N_479,In_1644,In_547);
and U480 (N_480,In_4259,In_621);
xnor U481 (N_481,In_3446,In_2711);
or U482 (N_482,In_3151,In_4064);
xnor U483 (N_483,In_3590,In_4101);
nand U484 (N_484,In_4622,In_3545);
nand U485 (N_485,In_794,In_478);
xor U486 (N_486,In_1334,In_2903);
nand U487 (N_487,In_2976,In_4789);
or U488 (N_488,In_785,In_709);
nand U489 (N_489,In_3248,In_4335);
nor U490 (N_490,In_2689,In_2839);
xnor U491 (N_491,In_3050,In_193);
nand U492 (N_492,In_338,In_3349);
nor U493 (N_493,In_4442,In_2123);
and U494 (N_494,In_681,In_1603);
xnor U495 (N_495,In_4420,In_2210);
nand U496 (N_496,In_4156,In_279);
nand U497 (N_497,In_1472,In_3728);
nor U498 (N_498,In_4900,In_2347);
xnor U499 (N_499,In_4579,In_312);
and U500 (N_500,In_3741,In_3262);
and U501 (N_501,In_628,In_400);
nor U502 (N_502,In_161,In_2597);
nor U503 (N_503,In_1237,In_2114);
or U504 (N_504,In_122,In_1906);
and U505 (N_505,In_2584,In_22);
or U506 (N_506,In_3855,In_4459);
nand U507 (N_507,In_1873,In_4565);
nand U508 (N_508,In_3219,In_1618);
nor U509 (N_509,In_323,In_3988);
xnor U510 (N_510,In_2505,In_3244);
or U511 (N_511,In_4393,In_421);
or U512 (N_512,In_4148,In_1814);
nand U513 (N_513,In_2244,In_4739);
xor U514 (N_514,In_3241,In_4373);
nand U515 (N_515,In_1151,In_931);
nand U516 (N_516,In_4107,In_3066);
xor U517 (N_517,In_2339,In_714);
xor U518 (N_518,In_1022,In_3340);
or U519 (N_519,In_2781,In_856);
xnor U520 (N_520,In_2232,In_54);
and U521 (N_521,In_2681,In_3312);
nor U522 (N_522,In_3108,In_4256);
and U523 (N_523,In_4648,In_588);
nor U524 (N_524,In_2319,In_1910);
or U525 (N_525,In_3433,In_1645);
nand U526 (N_526,In_169,In_3631);
and U527 (N_527,In_959,In_4388);
nor U528 (N_528,In_1940,In_436);
xor U529 (N_529,In_460,In_743);
xor U530 (N_530,In_3091,In_1721);
nor U531 (N_531,In_737,In_1733);
xor U532 (N_532,In_1285,In_2174);
or U533 (N_533,In_2786,In_1580);
or U534 (N_534,In_2511,In_1867);
nand U535 (N_535,In_2137,In_4962);
and U536 (N_536,In_2149,In_507);
or U537 (N_537,In_2696,In_4653);
nor U538 (N_538,In_4257,In_1848);
and U539 (N_539,In_2720,In_1391);
and U540 (N_540,In_4552,In_4614);
nand U541 (N_541,In_1850,In_973);
and U542 (N_542,In_4254,In_1700);
and U543 (N_543,In_2630,In_3698);
nand U544 (N_544,In_1419,In_4840);
nand U545 (N_545,In_4082,In_2320);
xnor U546 (N_546,In_545,In_2948);
and U547 (N_547,In_1444,In_2645);
nor U548 (N_548,In_2774,In_3415);
or U549 (N_549,In_4178,In_4709);
xnor U550 (N_550,In_1507,In_3677);
and U551 (N_551,In_1563,In_3873);
xor U552 (N_552,In_3621,In_1729);
or U553 (N_553,In_3526,In_1466);
nand U554 (N_554,In_3486,In_2955);
xnor U555 (N_555,In_4291,In_919);
xor U556 (N_556,In_55,In_3203);
or U557 (N_557,In_1259,In_2353);
nand U558 (N_558,In_658,In_4605);
nand U559 (N_559,In_930,In_4769);
nor U560 (N_560,In_1706,In_1325);
and U561 (N_561,In_4571,In_2574);
or U562 (N_562,In_91,In_3254);
xnor U563 (N_563,In_1611,In_4189);
or U564 (N_564,In_742,In_3909);
xnor U565 (N_565,In_2620,In_1364);
and U566 (N_566,In_4166,In_216);
xnor U567 (N_567,In_3346,In_2049);
nand U568 (N_568,In_4283,In_4395);
xor U569 (N_569,In_2969,In_1543);
nor U570 (N_570,In_1830,In_907);
xnor U571 (N_571,In_3945,In_1014);
xor U572 (N_572,In_587,In_4321);
or U573 (N_573,In_402,In_3127);
nand U574 (N_574,In_2936,In_2908);
nor U575 (N_575,In_3360,In_2750);
nor U576 (N_576,In_2918,In_175);
or U577 (N_577,In_4467,In_774);
xnor U578 (N_578,In_1871,In_457);
nand U579 (N_579,In_4111,In_2912);
nor U580 (N_580,In_1821,In_2336);
and U581 (N_581,In_4392,In_3554);
nor U582 (N_582,In_3132,In_2530);
or U583 (N_583,In_345,In_2016);
nand U584 (N_584,In_3084,In_3565);
nand U585 (N_585,In_1712,In_3746);
nor U586 (N_586,In_3478,In_205);
and U587 (N_587,In_679,In_2986);
and U588 (N_588,In_465,In_3604);
nand U589 (N_589,In_732,In_2586);
nand U590 (N_590,In_1630,In_1844);
nand U591 (N_591,In_494,In_2292);
and U592 (N_592,In_711,In_461);
or U593 (N_593,In_4184,In_2163);
xor U594 (N_594,In_427,In_3289);
xor U595 (N_595,In_3309,In_2238);
or U596 (N_596,In_631,In_261);
and U597 (N_597,In_2924,In_1263);
nor U598 (N_598,In_1517,In_2670);
or U599 (N_599,In_1158,In_1109);
and U600 (N_600,In_3136,In_1608);
nand U601 (N_601,In_2132,In_2288);
or U602 (N_602,In_4486,In_359);
nand U603 (N_603,In_3366,In_3708);
nand U604 (N_604,In_252,In_3488);
and U605 (N_605,In_3030,In_4722);
nand U606 (N_606,In_533,In_762);
and U607 (N_607,In_464,In_501);
and U608 (N_608,In_459,In_1326);
and U609 (N_609,In_3664,In_3522);
nor U610 (N_610,In_468,In_3015);
nand U611 (N_611,In_4383,In_3347);
nor U612 (N_612,In_272,In_4280);
xor U613 (N_613,In_3256,In_525);
nor U614 (N_614,In_2152,In_4398);
xor U615 (N_615,In_4384,In_1991);
nand U616 (N_616,In_1535,In_3926);
xnor U617 (N_617,In_1936,In_4935);
nor U618 (N_618,In_2564,In_2086);
nand U619 (N_619,In_2655,In_4515);
or U620 (N_620,In_290,In_2849);
nand U621 (N_621,In_3674,In_3739);
or U622 (N_622,In_0,In_4416);
nor U623 (N_623,In_2747,In_2087);
nand U624 (N_624,In_4550,In_3809);
xor U625 (N_625,In_1792,In_2352);
xnor U626 (N_626,In_1054,In_3736);
xor U627 (N_627,In_3120,In_3318);
and U628 (N_628,In_1314,In_4407);
or U629 (N_629,In_2197,In_2019);
nor U630 (N_630,In_81,In_484);
and U631 (N_631,In_4683,In_4444);
and U632 (N_632,In_1309,In_2296);
nor U633 (N_633,In_4906,In_4240);
or U634 (N_634,In_508,In_3814);
nand U635 (N_635,In_3507,In_1730);
and U636 (N_636,In_3673,In_135);
nand U637 (N_637,In_2801,In_1639);
or U638 (N_638,In_2966,In_3406);
nand U639 (N_639,In_3307,In_3048);
and U640 (N_640,In_3894,In_4998);
and U641 (N_641,In_2448,In_4278);
xor U642 (N_642,In_2787,In_2122);
or U643 (N_643,In_139,In_1750);
and U644 (N_644,In_4353,In_4533);
nand U645 (N_645,In_2771,In_4963);
xnor U646 (N_646,In_153,In_576);
xnor U647 (N_647,In_4322,In_3408);
nand U648 (N_648,In_914,In_4674);
nor U649 (N_649,In_2639,In_4608);
nor U650 (N_650,In_1255,In_4860);
nand U651 (N_651,In_2680,In_3039);
nor U652 (N_652,In_991,In_3761);
nor U653 (N_653,In_316,In_2497);
xnor U654 (N_654,In_4143,In_1546);
xor U655 (N_655,In_3229,In_3594);
nand U656 (N_656,In_2271,In_3004);
nand U657 (N_657,In_3496,In_1852);
nand U658 (N_658,In_2693,In_2331);
nand U659 (N_659,In_112,In_1226);
and U660 (N_660,In_4440,In_439);
nand U661 (N_661,In_4169,In_1909);
or U662 (N_662,In_4986,In_1230);
nand U663 (N_663,In_1623,In_4274);
and U664 (N_664,In_570,In_1216);
or U665 (N_665,In_1373,In_2603);
nor U666 (N_666,In_866,In_4759);
xnor U667 (N_667,In_4983,In_2519);
nor U668 (N_668,In_510,In_4317);
nand U669 (N_669,In_4334,In_2552);
nand U670 (N_670,In_4787,In_2376);
and U671 (N_671,In_509,In_3301);
or U672 (N_672,In_3612,In_1859);
nor U673 (N_673,In_4980,In_86);
and U674 (N_674,In_3217,In_1244);
and U675 (N_675,In_811,In_1720);
or U676 (N_676,In_4966,In_3392);
or U677 (N_677,In_3172,In_4399);
nor U678 (N_678,In_3204,In_3861);
xor U679 (N_679,In_4193,In_1995);
or U680 (N_680,In_4958,In_619);
or U681 (N_681,In_432,In_4757);
nor U682 (N_682,In_1288,In_876);
nand U683 (N_683,In_3207,In_2478);
or U684 (N_684,In_805,In_1195);
nor U685 (N_685,In_4514,In_4863);
nand U686 (N_686,In_3591,In_2713);
nor U687 (N_687,In_1390,In_4670);
xor U688 (N_688,In_1335,In_1589);
and U689 (N_689,In_1385,In_2343);
and U690 (N_690,In_3,In_2397);
nand U691 (N_691,In_2181,In_2813);
xor U692 (N_692,In_1424,In_1602);
nand U693 (N_693,In_4826,In_1967);
xor U694 (N_694,In_1476,In_125);
nand U695 (N_695,In_3668,In_649);
or U696 (N_696,In_2515,In_2961);
nand U697 (N_697,In_1406,In_3819);
nand U698 (N_698,In_4844,In_4564);
nand U699 (N_699,In_4517,In_3588);
or U700 (N_700,In_4086,In_3137);
and U701 (N_701,In_738,In_2857);
nand U702 (N_702,In_2825,In_687);
nor U703 (N_703,In_3298,In_4153);
or U704 (N_704,In_925,In_3529);
nor U705 (N_705,In_2449,In_3386);
nand U706 (N_706,In_2110,In_1924);
nand U707 (N_707,In_3463,In_2072);
and U708 (N_708,In_3725,In_577);
nor U709 (N_709,In_2803,In_1541);
nor U710 (N_710,In_1588,In_2351);
or U711 (N_711,In_58,In_3605);
and U712 (N_712,In_314,In_1308);
xnor U713 (N_713,In_337,In_3663);
and U714 (N_714,In_2432,In_3620);
and U715 (N_715,In_504,In_4577);
nor U716 (N_716,In_3281,In_1096);
xor U717 (N_717,In_3541,In_4418);
xor U718 (N_718,In_4842,In_668);
xor U719 (N_719,In_4210,In_984);
xnor U720 (N_720,In_2007,In_1277);
xnor U721 (N_721,In_2887,In_2802);
xnor U722 (N_722,In_4814,In_4837);
or U723 (N_723,In_1282,In_2154);
nor U724 (N_724,In_2531,In_3462);
and U725 (N_725,In_4775,In_134);
and U726 (N_726,In_4835,In_2965);
and U727 (N_727,In_4790,In_1382);
and U728 (N_728,In_1497,In_1047);
xor U729 (N_729,In_2840,In_4528);
nand U730 (N_730,In_3841,In_1992);
xor U731 (N_731,In_4707,In_1119);
nand U732 (N_732,In_3231,In_652);
nor U733 (N_733,In_3965,In_916);
nand U734 (N_734,In_361,In_1386);
and U735 (N_735,In_1494,In_3753);
nor U736 (N_736,In_2224,In_2382);
nand U737 (N_737,In_1068,In_1840);
and U738 (N_738,In_174,In_4342);
and U739 (N_739,In_368,In_1299);
or U740 (N_740,In_3756,In_1536);
or U741 (N_741,In_4636,In_3482);
nand U742 (N_742,In_3608,In_2790);
nand U743 (N_743,In_2789,In_3862);
and U744 (N_744,In_2031,In_1360);
and U745 (N_745,In_4628,In_24);
nor U746 (N_746,In_1677,In_3539);
xor U747 (N_747,In_3989,In_2649);
xor U748 (N_748,In_599,In_2837);
nor U749 (N_749,In_4199,In_1976);
nor U750 (N_750,In_1713,In_2272);
nand U751 (N_751,In_4251,In_772);
nor U752 (N_752,In_3212,In_3982);
nand U753 (N_753,In_4913,In_4088);
xor U754 (N_754,In_1268,In_426);
xor U755 (N_755,In_2185,In_927);
or U756 (N_756,In_283,In_1647);
or U757 (N_757,In_4920,In_4168);
or U758 (N_758,In_3876,In_159);
nand U759 (N_759,In_3157,In_1832);
nand U760 (N_760,In_4893,In_1291);
nor U761 (N_761,In_3263,In_1234);
nor U762 (N_762,In_4601,In_3240);
xnor U763 (N_763,In_3504,In_92);
nor U764 (N_764,In_2004,In_952);
nor U765 (N_765,In_4762,In_2334);
xor U766 (N_766,In_1616,In_2621);
nand U767 (N_767,In_116,In_2307);
nor U768 (N_768,In_1944,In_2498);
xor U769 (N_769,In_1351,In_4926);
or U770 (N_770,In_2267,In_2481);
nand U771 (N_771,In_2939,In_2097);
nor U772 (N_772,In_1240,In_1053);
xnor U773 (N_773,In_4598,In_891);
or U774 (N_774,In_881,In_1927);
nor U775 (N_775,In_1897,In_3551);
xor U776 (N_776,In_3260,In_898);
xnor U777 (N_777,In_4080,In_374);
nor U778 (N_778,In_2683,In_4831);
or U779 (N_779,In_538,In_4903);
xor U780 (N_780,In_764,In_4287);
or U781 (N_781,In_2882,In_2982);
nor U782 (N_782,In_3532,In_1437);
nand U783 (N_783,In_1508,In_2180);
nand U784 (N_784,In_19,In_2963);
nor U785 (N_785,In_479,In_4729);
and U786 (N_786,In_260,In_1635);
or U787 (N_787,In_1023,In_778);
and U788 (N_788,In_4364,In_1737);
xor U789 (N_789,In_4320,In_3650);
and U790 (N_790,In_2491,In_1716);
xnor U791 (N_791,In_4606,In_4567);
and U792 (N_792,In_2368,In_4527);
or U793 (N_793,In_598,In_4587);
or U794 (N_794,In_2403,In_3353);
xnor U795 (N_795,In_3177,In_2780);
nand U796 (N_796,In_4061,In_38);
xnor U797 (N_797,In_2145,In_2648);
nor U798 (N_798,In_2381,In_1569);
or U799 (N_799,In_528,In_3699);
nand U800 (N_800,In_2687,In_2512);
xnor U801 (N_801,In_219,In_833);
nand U802 (N_802,In_100,In_1474);
xor U803 (N_803,In_1060,In_4508);
nand U804 (N_804,In_1283,In_288);
nor U805 (N_805,In_4848,In_2775);
nor U806 (N_806,In_4553,In_1142);
xnor U807 (N_807,In_3801,In_4396);
xor U808 (N_808,In_4624,In_1764);
and U809 (N_809,In_644,In_160);
or U810 (N_810,In_2522,In_722);
or U811 (N_811,In_3365,In_1803);
nor U812 (N_812,In_3473,In_1921);
xor U813 (N_813,In_2767,In_1464);
and U814 (N_814,In_40,In_3899);
nor U815 (N_815,In_1050,In_2250);
xor U816 (N_816,In_3842,In_114);
or U817 (N_817,In_4425,In_2974);
or U818 (N_818,In_4144,In_4054);
nor U819 (N_819,In_448,In_559);
nand U820 (N_820,In_4164,In_4134);
xnor U821 (N_821,In_3986,In_1210);
or U822 (N_822,In_298,In_3037);
nand U823 (N_823,In_734,In_2091);
xnor U824 (N_824,In_1968,In_2900);
nor U825 (N_825,In_2622,In_1058);
and U826 (N_826,In_3838,In_2776);
or U827 (N_827,In_4642,In_1177);
xnor U828 (N_828,In_1359,In_4417);
xor U829 (N_829,In_241,In_4016);
nor U830 (N_830,In_2988,In_4690);
or U831 (N_831,In_4797,In_3411);
nand U832 (N_832,In_2454,In_4803);
nand U833 (N_833,In_4492,In_1454);
or U834 (N_834,In_2348,In_511);
nor U835 (N_835,In_3477,In_131);
xor U836 (N_836,In_4877,In_121);
xnor U837 (N_837,In_2329,In_730);
nor U838 (N_838,In_674,In_2054);
and U839 (N_839,In_3827,In_3014);
nor U840 (N_840,In_1118,In_2456);
nand U841 (N_841,In_2464,In_4109);
or U842 (N_842,In_485,In_3060);
or U843 (N_843,In_963,In_4908);
nand U844 (N_844,In_2732,In_912);
and U845 (N_845,In_3679,In_315);
nand U846 (N_846,In_282,In_3692);
and U847 (N_847,In_2602,In_4244);
or U848 (N_848,In_1303,In_3253);
or U849 (N_849,In_1614,In_1436);
nand U850 (N_850,In_2225,In_1435);
nand U851 (N_851,In_1062,In_2616);
and U852 (N_852,In_4505,In_4829);
or U853 (N_853,In_3793,In_2084);
nor U854 (N_854,In_3518,In_981);
and U855 (N_855,In_558,In_2428);
xnor U856 (N_856,In_393,In_3290);
and U857 (N_857,In_2719,In_3879);
nor U858 (N_858,In_2984,In_2475);
xor U859 (N_859,In_4750,In_874);
and U860 (N_860,In_2143,In_707);
xor U861 (N_861,In_1566,In_2896);
nand U862 (N_862,In_1302,In_3214);
or U863 (N_863,In_1661,In_416);
and U864 (N_864,In_1558,In_1575);
nor U865 (N_865,In_1636,In_1106);
and U866 (N_866,In_285,In_4161);
nand U867 (N_867,In_1484,In_2150);
nand U868 (N_868,In_187,In_4249);
xor U869 (N_869,In_1154,In_1798);
and U870 (N_870,In_4992,In_2746);
nand U871 (N_871,In_143,In_1892);
nand U872 (N_872,In_3237,In_1252);
xor U873 (N_873,In_2716,In_2533);
xnor U874 (N_874,In_1026,In_2332);
and U875 (N_875,In_1825,In_218);
nor U876 (N_876,In_2009,In_4001);
nand U877 (N_877,In_4704,In_2591);
xor U878 (N_878,In_760,In_1889);
xor U879 (N_879,In_2485,In_3654);
xnor U880 (N_880,In_4804,In_3859);
or U881 (N_881,In_4180,In_492);
nor U882 (N_882,In_1348,In_2527);
nor U883 (N_883,In_810,In_3645);
and U884 (N_884,In_2884,In_4706);
and U885 (N_885,In_3454,In_3025);
nor U886 (N_886,In_1804,In_347);
nand U887 (N_887,In_2392,In_2700);
and U888 (N_888,In_420,In_2541);
nor U889 (N_889,In_1367,In_2117);
and U890 (N_890,In_2824,In_3195);
and U891 (N_891,In_3778,In_3641);
and U892 (N_892,In_4743,In_676);
nor U893 (N_893,In_4094,In_1036);
nor U894 (N_894,In_3881,In_4352);
or U895 (N_895,In_3399,In_2492);
or U896 (N_896,In_1399,In_4917);
and U897 (N_897,In_2109,In_4596);
nor U898 (N_898,In_1642,In_245);
or U899 (N_899,In_2080,In_2465);
xnor U900 (N_900,In_3218,In_2919);
and U901 (N_901,In_4780,In_3893);
or U902 (N_902,In_2626,In_4269);
nand U903 (N_903,In_1856,In_2155);
xnor U904 (N_904,In_4047,In_2556);
nor U905 (N_905,In_2653,In_1917);
nor U906 (N_906,In_142,In_1257);
or U907 (N_907,In_3494,In_2427);
xnor U908 (N_908,In_1606,In_1460);
xor U909 (N_909,In_1902,In_4043);
and U910 (N_910,In_4513,In_985);
nor U911 (N_911,In_2892,In_929);
nand U912 (N_912,In_3625,In_2594);
nand U913 (N_913,In_247,In_2829);
nand U914 (N_914,In_158,In_4077);
and U915 (N_915,In_4241,In_2748);
nand U916 (N_916,In_3368,In_326);
nand U917 (N_917,In_146,In_894);
and U918 (N_918,In_4507,In_3903);
or U919 (N_919,In_343,In_2228);
xor U920 (N_920,In_2325,In_2036);
nand U921 (N_921,In_2298,In_3836);
nand U922 (N_922,In_958,In_3524);
nand U923 (N_923,In_3584,In_829);
or U924 (N_924,In_1176,In_3223);
nor U925 (N_925,In_2385,In_4162);
and U926 (N_926,In_3121,In_3549);
xor U927 (N_927,In_1144,In_1393);
and U928 (N_928,In_926,In_1576);
xnor U929 (N_929,In_2575,In_3805);
xnor U930 (N_930,In_1465,In_3090);
xnor U931 (N_931,In_3718,In_651);
nor U932 (N_932,In_1134,In_4621);
and U933 (N_933,In_2794,In_4815);
nor U934 (N_934,In_1353,In_3160);
or U935 (N_935,In_4458,In_3026);
nor U936 (N_936,In_4999,In_4035);
and U937 (N_937,In_1725,In_3550);
xnor U938 (N_938,In_3012,In_4936);
nand U939 (N_939,In_3111,In_505);
xnor U940 (N_940,In_4219,In_1012);
and U941 (N_941,In_1250,In_4827);
nor U942 (N_942,In_3796,In_3910);
and U943 (N_943,In_4338,In_1223);
nor U944 (N_944,In_2619,In_4382);
or U945 (N_945,In_3637,In_999);
or U946 (N_946,In_4689,In_3760);
xnor U947 (N_947,In_590,In_428);
nand U948 (N_948,In_1169,In_2866);
nand U949 (N_949,In_1515,In_4208);
or U950 (N_950,In_3021,In_4663);
nor U951 (N_951,In_4705,In_3780);
xnor U952 (N_952,In_4735,In_4927);
xnor U953 (N_953,In_3632,In_4537);
nand U954 (N_954,In_2944,In_4808);
nor U955 (N_955,In_3902,In_3045);
or U956 (N_956,In_1213,In_1886);
or U957 (N_957,In_3242,In_1427);
xor U958 (N_958,In_1067,In_3351);
xor U959 (N_959,In_3652,In_2015);
xnor U960 (N_960,In_2915,In_3963);
and U961 (N_961,In_4185,In_1765);
nand U962 (N_962,In_4498,In_4696);
nor U963 (N_963,In_3149,In_1920);
or U964 (N_964,In_4049,In_1376);
and U965 (N_965,In_3548,In_1723);
or U966 (N_966,In_4545,In_2131);
nor U967 (N_967,In_4160,In_967);
and U968 (N_968,In_105,In_1872);
xor U969 (N_969,In_2121,In_1229);
or U970 (N_970,In_493,In_3657);
xor U971 (N_971,In_4341,In_70);
nand U972 (N_972,In_3828,In_937);
xnor U973 (N_973,In_1394,In_502);
xor U974 (N_974,In_4385,In_2206);
and U975 (N_975,In_384,In_4869);
or U976 (N_976,In_1112,In_2395);
nor U977 (N_977,In_1137,In_2694);
or U978 (N_978,In_1488,In_2050);
or U979 (N_979,In_2612,In_1317);
nor U980 (N_980,In_4888,In_1324);
nor U981 (N_981,In_2871,In_437);
or U982 (N_982,In_2962,In_1912);
nand U983 (N_983,In_1136,In_2833);
and U984 (N_984,In_2184,In_4456);
or U985 (N_985,In_1675,In_1666);
and U986 (N_986,In_3818,In_503);
or U987 (N_987,In_453,In_1354);
or U988 (N_988,In_2214,In_4051);
nor U989 (N_989,In_3596,In_1080);
xor U990 (N_990,In_2607,In_3857);
nand U991 (N_991,In_2003,In_1657);
and U992 (N_992,In_4902,In_1301);
or U993 (N_993,In_4989,In_1015);
nor U994 (N_994,In_2904,In_3709);
or U995 (N_995,In_1714,In_2971);
nand U996 (N_996,In_1998,In_2535);
and U997 (N_997,In_1239,In_1128);
or U998 (N_998,In_4263,In_1669);
nor U999 (N_999,In_2315,In_2058);
nand U1000 (N_1000,In_895,In_955);
nor U1001 (N_1001,In_4085,In_1126);
or U1002 (N_1002,In_1330,In_2359);
nor U1003 (N_1003,In_1071,In_3555);
and U1004 (N_1004,In_1962,In_4015);
xor U1005 (N_1005,In_1113,In_3724);
or U1006 (N_1006,In_481,In_41);
and U1007 (N_1007,In_2187,In_2812);
and U1008 (N_1008,In_1344,In_1705);
nand U1009 (N_1009,In_3448,In_155);
xnor U1010 (N_1010,In_604,In_2708);
nor U1011 (N_1011,In_2598,In_2704);
xor U1012 (N_1012,In_3105,In_430);
xor U1013 (N_1013,In_1934,In_1477);
nor U1014 (N_1014,In_2186,In_2301);
nor U1015 (N_1015,In_4140,In_2468);
and U1016 (N_1016,In_4017,In_414);
xor U1017 (N_1017,In_663,In_488);
nand U1018 (N_1018,In_3981,In_4589);
and U1019 (N_1019,In_3779,In_1073);
xor U1020 (N_1020,In_3658,In_3983);
nand U1021 (N_1021,In_4232,In_3535);
and U1022 (N_1022,In_972,In_3672);
and U1023 (N_1023,In_4115,In_3480);
nand U1024 (N_1024,In_2120,In_2450);
nand U1025 (N_1025,In_4640,In_2472);
or U1026 (N_1026,In_1853,In_4580);
nor U1027 (N_1027,In_1742,In_2355);
nor U1028 (N_1028,In_4811,In_4439);
or U1029 (N_1029,In_4502,In_4052);
nand U1030 (N_1030,In_292,In_2561);
nand U1031 (N_1031,In_3046,In_10);
nor U1032 (N_1032,In_1646,In_1553);
nand U1033 (N_1033,In_1041,In_4501);
nand U1034 (N_1034,In_1527,In_4010);
and U1035 (N_1035,In_4377,In_4038);
nor U1036 (N_1036,In_3907,In_3002);
nand U1037 (N_1037,In_4595,In_2474);
nand U1038 (N_1038,In_1208,In_4127);
nand U1039 (N_1039,In_4183,In_4880);
xnor U1040 (N_1040,In_3101,In_328);
and U1041 (N_1041,In_1478,In_4886);
and U1042 (N_1042,In_1048,In_1387);
and U1043 (N_1043,In_1552,In_1509);
nand U1044 (N_1044,In_2092,In_104);
nand U1045 (N_1045,In_3829,In_2543);
or U1046 (N_1046,In_1514,In_4887);
nor U1047 (N_1047,In_4330,In_1483);
xnor U1048 (N_1048,In_4965,In_2318);
xnor U1049 (N_1049,In_4239,In_2327);
or U1050 (N_1050,In_2685,In_4896);
nand U1051 (N_1051,In_4568,In_1358);
or U1052 (N_1052,In_4524,In_3553);
xor U1053 (N_1053,In_2929,In_1321);
nand U1054 (N_1054,In_3878,In_4710);
nand U1055 (N_1055,In_4858,In_327);
nand U1056 (N_1056,In_2241,In_549);
nand U1057 (N_1057,In_700,In_4819);
nand U1058 (N_1058,In_1135,In_4784);
and U1059 (N_1059,In_300,In_3215);
and U1060 (N_1060,In_4593,In_4265);
nand U1061 (N_1061,In_4820,In_2635);
and U1062 (N_1062,In_4878,In_2920);
nor U1063 (N_1063,In_2129,In_4654);
or U1064 (N_1064,In_362,In_1548);
nand U1065 (N_1065,In_2253,In_2442);
nand U1066 (N_1066,In_989,In_4849);
nand U1067 (N_1067,In_1167,In_2265);
xnor U1068 (N_1068,In_4698,In_29);
or U1069 (N_1069,In_249,In_2095);
nand U1070 (N_1070,In_2215,In_2633);
and U1071 (N_1071,In_340,In_1707);
or U1072 (N_1072,In_731,In_4412);
xnor U1073 (N_1073,In_2311,In_4281);
nor U1074 (N_1074,In_1711,In_3194);
xor U1075 (N_1075,In_3247,In_910);
xnor U1076 (N_1076,In_3752,In_1004);
xnor U1077 (N_1077,In_4277,In_3546);
or U1078 (N_1078,In_729,In_3915);
nand U1079 (N_1079,In_593,In_4701);
and U1080 (N_1080,In_1001,In_1908);
xnor U1081 (N_1081,In_2978,In_369);
nand U1082 (N_1082,In_506,In_2972);
or U1083 (N_1083,In_3147,In_1377);
nor U1084 (N_1084,In_4872,In_2977);
xor U1085 (N_1085,In_477,In_4793);
and U1086 (N_1086,In_4227,In_1774);
and U1087 (N_1087,In_2526,In_191);
and U1088 (N_1088,In_3150,In_4964);
xor U1089 (N_1089,In_4409,In_1916);
nor U1090 (N_1090,In_2014,In_2053);
nor U1091 (N_1091,In_4260,In_2509);
nor U1092 (N_1092,In_3994,In_3418);
and U1093 (N_1093,In_3153,In_1928);
nor U1094 (N_1094,In_900,In_2451);
nand U1095 (N_1095,In_2660,In_2761);
nor U1096 (N_1096,In_2216,In_2669);
and U1097 (N_1097,In_735,In_4519);
nor U1098 (N_1098,In_3437,In_1749);
xor U1099 (N_1099,In_3450,In_4258);
or U1100 (N_1100,In_1457,In_627);
nor U1101 (N_1101,In_1379,In_303);
or U1102 (N_1102,In_147,In_1174);
nand U1103 (N_1103,In_704,In_2130);
nor U1104 (N_1104,In_610,In_1596);
or U1105 (N_1105,In_1834,In_1179);
nand U1106 (N_1106,In_3129,In_4391);
nor U1107 (N_1107,In_3916,In_1704);
or U1108 (N_1108,In_3707,In_1864);
or U1109 (N_1109,In_4386,In_1114);
nand U1110 (N_1110,In_1747,In_1278);
xor U1111 (N_1111,In_3363,In_3173);
nand U1112 (N_1112,In_3700,In_4447);
nand U1113 (N_1113,In_2414,In_4680);
and U1114 (N_1114,In_3348,In_3297);
xnor U1115 (N_1115,In_1506,In_953);
nor U1116 (N_1116,In_550,In_2553);
or U1117 (N_1117,In_198,In_3531);
and U1118 (N_1118,In_834,In_4677);
and U1119 (N_1119,In_2580,In_3928);
nor U1120 (N_1120,In_3018,In_791);
nor U1121 (N_1121,In_3561,In_4473);
nand U1122 (N_1122,In_2300,In_3924);
or U1123 (N_1123,In_2764,In_57);
nand U1124 (N_1124,In_1456,In_3139);
or U1125 (N_1125,In_2863,In_1613);
nor U1126 (N_1126,In_2282,In_1131);
or U1127 (N_1127,In_656,In_387);
or U1128 (N_1128,In_4267,In_2876);
xnor U1129 (N_1129,In_2234,In_4495);
and U1130 (N_1130,In_1475,In_2772);
nand U1131 (N_1131,In_4152,In_4301);
or U1132 (N_1132,In_3892,In_259);
xnor U1133 (N_1133,In_3675,In_2507);
or U1134 (N_1134,In_3067,In_2568);
and U1135 (N_1135,In_1307,In_3837);
nand U1136 (N_1136,In_12,In_4163);
xnor U1137 (N_1137,In_2742,In_148);
and U1138 (N_1138,In_2624,In_3343);
and U1139 (N_1139,In_2230,In_1212);
nor U1140 (N_1140,In_745,In_2125);
nand U1141 (N_1141,In_1198,In_2198);
and U1142 (N_1142,In_3362,In_2601);
xnor U1143 (N_1143,In_2452,In_969);
and U1144 (N_1144,In_4830,In_1500);
or U1145 (N_1145,In_3395,In_4754);
or U1146 (N_1146,In_1089,In_2782);
and U1147 (N_1147,In_4136,In_3502);
and U1148 (N_1148,In_4066,In_250);
nor U1149 (N_1149,In_690,In_1790);
or U1150 (N_1150,In_3964,In_3166);
and U1151 (N_1151,In_4438,In_4312);
and U1152 (N_1152,In_3181,In_1338);
or U1153 (N_1153,In_1100,In_1870);
or U1154 (N_1154,In_2749,In_655);
or U1155 (N_1155,In_2941,In_4556);
nand U1156 (N_1156,In_475,In_4468);
and U1157 (N_1157,In_2506,In_1593);
or U1158 (N_1158,In_4009,In_2302);
xnor U1159 (N_1159,In_335,In_2667);
or U1160 (N_1160,In_3269,In_2589);
and U1161 (N_1161,In_2671,In_890);
or U1162 (N_1162,In_3799,In_3054);
nor U1163 (N_1163,In_4772,In_4802);
and U1164 (N_1164,In_3134,In_2820);
and U1165 (N_1165,In_2457,In_2173);
nand U1166 (N_1166,In_2326,In_132);
nand U1167 (N_1167,In_1786,In_3512);
or U1168 (N_1168,In_4559,In_3249);
xnor U1169 (N_1169,In_4742,In_1164);
xor U1170 (N_1170,In_3336,In_3224);
or U1171 (N_1171,In_4873,In_4297);
xor U1172 (N_1172,In_901,In_2112);
xor U1173 (N_1173,In_3973,In_1083);
xor U1174 (N_1174,In_852,In_1970);
nor U1175 (N_1175,In_127,In_1404);
or U1176 (N_1176,In_1232,In_2642);
nand U1177 (N_1177,In_2151,In_2682);
and U1178 (N_1178,In_4018,In_1628);
nand U1179 (N_1179,In_1296,In_556);
and U1180 (N_1180,In_3749,In_617);
xnor U1181 (N_1181,In_1319,In_1620);
and U1182 (N_1182,In_4504,In_53);
or U1183 (N_1183,In_3900,In_4434);
nand U1184 (N_1184,In_466,In_807);
nor U1185 (N_1185,In_3510,In_4599);
nand U1186 (N_1186,In_1964,In_2778);
or U1187 (N_1187,In_3152,In_195);
nand U1188 (N_1188,In_4946,In_4520);
or U1189 (N_1189,In_126,In_2436);
or U1190 (N_1190,In_3833,In_860);
or U1191 (N_1191,In_4014,In_2830);
nand U1192 (N_1192,In_4738,In_2874);
and U1193 (N_1193,In_522,In_3234);
nand U1194 (N_1194,In_2672,In_2805);
nand U1195 (N_1195,In_1024,In_2659);
and U1196 (N_1196,In_331,In_354);
or U1197 (N_1197,In_2217,In_3762);
nand U1198 (N_1198,In_1550,In_4832);
nor U1199 (N_1199,In_2164,In_2869);
nand U1200 (N_1200,In_4059,In_4213);
and U1201 (N_1201,In_2268,In_680);
and U1202 (N_1202,In_4181,In_3458);
and U1203 (N_1203,In_2438,In_3931);
nor U1204 (N_1204,In_2249,In_1002);
xor U1205 (N_1205,In_2995,In_2147);
xnor U1206 (N_1206,In_1016,In_2062);
xnor U1207 (N_1207,In_1495,In_3723);
nor U1208 (N_1208,In_1175,In_2028);
and U1209 (N_1209,In_515,In_2954);
nor U1210 (N_1210,In_4931,In_2071);
nand U1211 (N_1211,In_1948,In_987);
or U1212 (N_1212,In_4969,In_3537);
xnor U1213 (N_1213,In_2940,In_1196);
nand U1214 (N_1214,In_194,In_4702);
and U1215 (N_1215,In_2898,In_2714);
and U1216 (N_1216,In_2646,In_294);
and U1217 (N_1217,In_4499,In_2167);
xnor U1218 (N_1218,In_31,In_1561);
nor U1219 (N_1219,In_2027,In_2985);
nor U1220 (N_1220,In_3064,In_1381);
nor U1221 (N_1221,In_3797,In_321);
nand U1222 (N_1222,In_3831,In_4057);
nor U1223 (N_1223,In_787,In_2383);
or U1224 (N_1224,In_1020,In_3282);
nand U1225 (N_1225,In_3047,In_4233);
nand U1226 (N_1226,In_1409,In_2721);
nand U1227 (N_1227,In_2248,In_408);
xor U1228 (N_1228,In_2341,In_4933);
or U1229 (N_1229,In_4211,In_784);
xnor U1230 (N_1230,In_364,In_3759);
nand U1231 (N_1231,In_412,In_2043);
and U1232 (N_1232,In_940,In_4525);
xnor U1233 (N_1233,In_79,In_4609);
xnor U1234 (N_1234,In_2684,In_557);
nor U1235 (N_1235,In_3638,In_2113);
nor U1236 (N_1236,In_4692,In_4782);
or U1237 (N_1237,In_3460,In_1149);
and U1238 (N_1238,In_2701,In_3848);
xor U1239 (N_1239,In_1253,In_2045);
or U1240 (N_1240,In_4981,In_1679);
nand U1241 (N_1241,In_1565,In_4042);
xor U1242 (N_1242,In_87,In_830);
nor U1243 (N_1243,In_2196,In_1101);
xor U1244 (N_1244,In_2208,In_3528);
or U1245 (N_1245,In_1363,In_3378);
nand U1246 (N_1246,In_280,In_864);
or U1247 (N_1247,In_720,In_1246);
and U1248 (N_1248,In_333,In_513);
and U1249 (N_1249,In_3019,In_2751);
nand U1250 (N_1250,In_3635,In_1059);
nor U1251 (N_1251,In_306,In_4510);
nand U1252 (N_1252,In_1146,In_759);
or U1253 (N_1253,In_3388,In_1194);
xor U1254 (N_1254,In_3888,In_1469);
and U1255 (N_1255,In_3689,In_2524);
and U1256 (N_1256,In_1331,In_4131);
nand U1257 (N_1257,In_1337,In_3520);
xnor U1258 (N_1258,In_3243,In_434);
and U1259 (N_1259,In_4938,In_1260);
nor U1260 (N_1260,In_3940,In_4056);
xor U1261 (N_1261,In_3733,In_2800);
xor U1262 (N_1262,In_2076,In_1820);
and U1263 (N_1263,In_120,In_3329);
xnor U1264 (N_1264,In_4812,In_4120);
xnor U1265 (N_1265,In_1502,In_1110);
nand U1266 (N_1266,In_1829,In_1933);
nor U1267 (N_1267,In_4643,In_353);
xor U1268 (N_1268,In_4000,In_2821);
and U1269 (N_1269,In_1461,In_2793);
nand U1270 (N_1270,In_3485,In_4868);
and U1271 (N_1271,In_956,In_3096);
nand U1272 (N_1272,In_2313,In_145);
or U1273 (N_1273,In_1600,In_596);
nor U1274 (N_1274,In_614,In_2583);
nand U1275 (N_1275,In_3314,In_2275);
nor U1276 (N_1276,In_892,In_670);
nor U1277 (N_1277,In_3261,In_297);
and U1278 (N_1278,In_3113,In_2220);
xor U1279 (N_1279,In_1063,In_2838);
xnor U1280 (N_1280,In_88,In_496);
nand U1281 (N_1281,In_4300,In_2127);
xor U1282 (N_1282,In_332,In_278);
or U1283 (N_1283,In_4796,In_4114);
nor U1284 (N_1284,In_3863,In_1547);
and U1285 (N_1285,In_3088,In_3617);
and U1286 (N_1286,In_630,In_4242);
and U1287 (N_1287,In_2783,In_933);
nand U1288 (N_1288,In_1997,In_4764);
nor U1289 (N_1289,In_3670,In_4315);
xor U1290 (N_1290,In_3872,In_4970);
or U1291 (N_1291,In_4139,In_4529);
xor U1292 (N_1292,In_1188,In_3158);
xnor U1293 (N_1293,In_3337,In_1622);
xnor U1294 (N_1294,In_1287,In_1969);
xor U1295 (N_1295,In_2587,In_3791);
nand U1296 (N_1296,In_3643,In_2226);
nand U1297 (N_1297,In_4637,In_308);
nand U1298 (N_1298,In_3404,In_2361);
or U1299 (N_1299,In_4572,In_2902);
nand U1300 (N_1300,In_966,In_3469);
xnor U1301 (N_1301,In_951,In_3476);
xnor U1302 (N_1302,In_3069,In_4252);
xor U1303 (N_1303,In_836,In_2458);
or U1304 (N_1304,In_1673,In_1320);
xnor U1305 (N_1305,In_4995,In_489);
and U1306 (N_1306,In_3324,In_2075);
nor U1307 (N_1307,In_1952,In_4048);
or U1308 (N_1308,In_4708,In_2139);
nand U1309 (N_1309,In_490,In_76);
nor U1310 (N_1310,In_3330,In_71);
nand U1311 (N_1311,In_3268,In_3655);
xor U1312 (N_1312,In_2528,In_2943);
and U1313 (N_1313,In_4641,In_18);
or U1314 (N_1314,In_1665,In_1766);
and U1315 (N_1315,In_982,In_3932);
and U1316 (N_1316,In_410,In_1591);
xor U1317 (N_1317,In_4682,In_4996);
and U1318 (N_1318,In_3955,In_1528);
or U1319 (N_1319,In_780,In_357);
nor U1320 (N_1320,In_4357,In_3868);
nand U1321 (N_1321,In_1791,In_355);
and U1322 (N_1322,In_75,In_1238);
nand U1323 (N_1323,In_2577,In_2421);
and U1324 (N_1324,In_4956,In_3210);
xor U1325 (N_1325,In_2202,In_632);
or U1326 (N_1326,In_3559,In_3467);
nand U1327 (N_1327,In_4346,In_1595);
nand U1328 (N_1328,In_2814,In_996);
nor U1329 (N_1329,In_3626,In_1557);
or U1330 (N_1330,In_4020,In_1709);
and U1331 (N_1331,In_2040,In_231);
or U1332 (N_1332,In_2093,In_336);
and U1333 (N_1333,In_4591,In_728);
nor U1334 (N_1334,In_1957,In_3885);
or U1335 (N_1335,In_2105,In_564);
and U1336 (N_1336,In_4968,In_595);
or U1337 (N_1337,In_2200,In_98);
or U1338 (N_1338,In_2136,In_4987);
or U1339 (N_1339,In_3186,In_1748);
nand U1340 (N_1340,In_2521,In_3783);
or U1341 (N_1341,In_741,In_380);
xnor U1342 (N_1342,In_4380,In_3869);
nor U1343 (N_1343,In_3162,In_2706);
nand U1344 (N_1344,In_2504,In_2901);
nor U1345 (N_1345,In_401,In_210);
and U1346 (N_1346,In_1449,In_1560);
nand U1347 (N_1347,In_106,In_1184);
or U1348 (N_1348,In_4108,In_2073);
and U1349 (N_1349,In_903,In_832);
nand U1350 (N_1350,In_2407,In_37);
and U1351 (N_1351,In_4752,In_3426);
nand U1352 (N_1352,In_2445,In_4940);
nand U1353 (N_1353,In_928,In_435);
nand U1354 (N_1354,In_3384,In_4972);
or U1355 (N_1355,In_1411,In_3935);
and U1356 (N_1356,In_4261,In_4340);
xor U1357 (N_1357,In_4667,In_3543);
or U1358 (N_1358,In_3937,In_2447);
xnor U1359 (N_1359,In_1339,In_1070);
or U1360 (N_1360,In_1010,In_4727);
nand U1361 (N_1361,In_3270,In_3578);
nand U1362 (N_1362,In_4774,In_909);
xor U1363 (N_1363,In_2513,In_4613);
xor U1364 (N_1364,In_2945,In_1439);
nand U1365 (N_1365,In_4957,In_2928);
or U1366 (N_1366,In_2958,In_3232);
nand U1367 (N_1367,In_2726,In_2729);
nand U1368 (N_1368,In_2308,In_1771);
or U1369 (N_1369,In_3697,In_3649);
xnor U1370 (N_1370,In_2638,In_2483);
nor U1371 (N_1371,In_1426,In_824);
nand U1372 (N_1372,In_2289,In_1117);
nor U1373 (N_1373,In_2835,In_4645);
xnor U1374 (N_1374,In_1537,In_992);
nand U1375 (N_1375,In_4090,In_2970);
nor U1376 (N_1376,In_2246,In_190);
or U1377 (N_1377,In_2797,In_560);
or U1378 (N_1378,In_1587,In_3390);
nor U1379 (N_1379,In_2389,In_293);
xnor U1380 (N_1380,In_723,In_3238);
and U1381 (N_1381,In_2889,In_2554);
nand U1382 (N_1382,In_3443,In_2823);
nand U1383 (N_1383,In_4146,In_542);
and U1384 (N_1384,In_2008,In_3466);
or U1385 (N_1385,In_642,In_429);
nor U1386 (N_1386,In_1776,In_375);
or U1387 (N_1387,In_1049,In_4534);
xor U1388 (N_1388,In_1846,In_1289);
nand U1389 (N_1389,In_3174,In_356);
and U1390 (N_1390,In_736,In_4023);
and U1391 (N_1391,In_3856,In_657);
and U1392 (N_1392,In_3564,In_4174);
xor U1393 (N_1393,In_721,In_944);
xnor U1394 (N_1394,In_441,In_2461);
or U1395 (N_1395,In_4305,In_882);
and U1396 (N_1396,In_2596,In_3221);
nand U1397 (N_1397,In_3143,In_4901);
nand U1398 (N_1398,In_1452,In_4845);
nor U1399 (N_1399,In_2785,In_1129);
nor U1400 (N_1400,In_242,In_4460);
xnor U1401 (N_1401,In_948,In_646);
nand U1402 (N_1402,In_3557,In_4586);
nor U1403 (N_1403,In_4740,In_867);
and U1404 (N_1404,In_1084,In_4821);
xnor U1405 (N_1405,In_4087,In_3099);
and U1406 (N_1406,In_2393,In_1333);
nand U1407 (N_1407,In_2266,In_1440);
xnor U1408 (N_1408,In_2345,In_4105);
and U1409 (N_1409,In_2126,In_3610);
nand U1410 (N_1410,In_2378,In_1366);
nand U1411 (N_1411,In_50,In_2996);
and U1412 (N_1412,In_266,In_4523);
xor U1413 (N_1413,In_4664,In_893);
nand U1414 (N_1414,In_3629,In_1298);
and U1415 (N_1415,In_3784,In_1163);
or U1416 (N_1416,In_42,In_4828);
nand U1417 (N_1417,In_887,In_746);
nand U1418 (N_1418,In_3735,In_2763);
or U1419 (N_1419,In_1438,In_3766);
or U1420 (N_1420,In_4414,In_2766);
xor U1421 (N_1421,In_4612,In_1978);
or U1422 (N_1422,In_2555,In_4530);
or U1423 (N_1423,In_397,In_4644);
xnor U1424 (N_1424,In_4323,In_320);
nand U1425 (N_1425,In_4922,In_1781);
xor U1426 (N_1426,In_1075,In_1796);
or U1427 (N_1427,In_3042,In_1778);
nor U1428 (N_1428,In_979,In_4362);
xor U1429 (N_1429,In_4129,In_4390);
xnor U1430 (N_1430,In_1950,In_1081);
and U1431 (N_1431,In_1990,In_3061);
or U1432 (N_1432,In_4539,In_1907);
nand U1433 (N_1433,In_2128,In_1854);
xor U1434 (N_1434,In_3192,In_1032);
nor U1435 (N_1435,In_4791,In_2247);
nor U1436 (N_1436,In_633,In_77);
and U1437 (N_1437,In_554,In_2864);
xor U1438 (N_1438,In_1370,In_2493);
nand U1439 (N_1439,In_798,In_96);
xor U1440 (N_1440,In_4170,In_1161);
or U1441 (N_1441,In_3633,In_518);
nor U1442 (N_1442,In_4679,In_3694);
xnor U1443 (N_1443,In_2144,In_1574);
xor U1444 (N_1444,In_4910,In_520);
or U1445 (N_1445,In_3199,In_740);
and U1446 (N_1446,In_4188,In_4952);
xor U1447 (N_1447,In_537,In_2925);
nand U1448 (N_1448,In_248,In_4367);
xor U1449 (N_1449,In_993,In_342);
nor U1450 (N_1450,In_4786,In_2947);
nand U1451 (N_1451,In_3434,In_3503);
and U1452 (N_1452,In_2819,In_3917);
xnor U1453 (N_1453,In_3927,In_3710);
nand U1454 (N_1454,In_2975,In_3100);
or U1455 (N_1455,In_1542,In_2792);
or U1456 (N_1456,In_3198,In_2278);
or U1457 (N_1457,In_84,In_3721);
and U1458 (N_1458,In_3558,In_151);
nand U1459 (N_1459,In_1121,In_654);
nand U1460 (N_1460,In_2363,In_1728);
nor U1461 (N_1461,In_1744,In_3681);
or U1462 (N_1462,In_519,In_1029);
nor U1463 (N_1463,In_3816,In_4719);
nand U1464 (N_1464,In_471,In_2077);
or U1465 (N_1465,In_2044,In_616);
nand U1466 (N_1466,In_795,In_3889);
and U1467 (N_1467,In_334,In_544);
or U1468 (N_1468,In_4816,In_3712);
xnor U1469 (N_1469,In_2808,In_2723);
nor U1470 (N_1470,In_4205,In_2599);
and U1471 (N_1471,In_1371,In_1719);
nor U1472 (N_1472,In_1556,In_1487);
and U1473 (N_1473,In_3071,In_3119);
and U1474 (N_1474,In_4044,In_3413);
xor U1475 (N_1475,In_2595,In_838);
and U1476 (N_1476,In_1418,In_1980);
nand U1477 (N_1477,In_1648,In_2488);
xnor U1478 (N_1478,In_2118,In_3597);
and U1479 (N_1479,In_3387,In_317);
or U1480 (N_1480,In_1866,In_1681);
or U1481 (N_1481,In_1762,In_3367);
nor U1482 (N_1482,In_1746,In_2629);
and U1483 (N_1483,In_3688,In_1352);
nor U1484 (N_1484,In_1410,In_2654);
or U1485 (N_1485,In_2106,In_3992);
and U1486 (N_1486,In_309,In_1529);
nor U1487 (N_1487,In_117,In_61);
or U1488 (N_1488,In_2038,In_659);
or U1489 (N_1489,In_1228,In_4633);
xor U1490 (N_1490,In_1954,In_4541);
xor U1491 (N_1491,In_3782,In_1953);
or U1492 (N_1492,In_4979,In_273);
nand U1493 (N_1493,In_3385,In_3883);
and U1494 (N_1494,In_2593,In_2614);
nand U1495 (N_1495,In_3834,In_3163);
nand U1496 (N_1496,In_4662,In_215);
xnor U1497 (N_1497,In_1292,In_2914);
and U1498 (N_1498,In_2799,In_1349);
nand U1499 (N_1499,In_3765,In_431);
nor U1500 (N_1500,In_4945,In_1984);
xor U1501 (N_1501,In_2115,In_2051);
or U1502 (N_1502,In_3475,In_961);
nor U1503 (N_1503,In_1601,In_3372);
or U1504 (N_1504,In_880,In_3960);
or U1505 (N_1505,In_4124,In_4685);
or U1506 (N_1506,In_4925,In_373);
or U1507 (N_1507,In_165,In_4582);
or U1508 (N_1508,In_592,In_2861);
nand U1509 (N_1509,In_922,In_166);
nand U1510 (N_1510,In_470,In_1201);
and U1511 (N_1511,In_796,In_4615);
nor U1512 (N_1512,In_3648,In_765);
or U1513 (N_1513,In_2567,In_2160);
nand U1514 (N_1514,In_4011,In_469);
nand U1515 (N_1515,In_4776,In_974);
nor U1516 (N_1516,In_329,In_896);
nand U1517 (N_1517,In_1651,In_3623);
xor U1518 (N_1518,In_26,In_3566);
xor U1519 (N_1519,In_4271,In_3222);
nor U1520 (N_1520,In_667,In_4521);
nor U1521 (N_1521,In_923,In_319);
xnor U1522 (N_1522,In_2632,In_1994);
nor U1523 (N_1523,In_1554,In_1754);
xor U1524 (N_1524,In_1881,In_3618);
or U1525 (N_1525,In_2907,In_4712);
xnor U1526 (N_1526,In_4997,In_920);
nand U1527 (N_1527,In_348,In_409);
and U1528 (N_1528,In_2374,In_2100);
and U1529 (N_1529,In_1304,In_1009);
xnor U1530 (N_1530,In_3997,In_1923);
nand U1531 (N_1531,In_473,In_863);
nand U1532 (N_1532,In_3957,In_2877);
nand U1533 (N_1533,In_696,In_883);
nor U1534 (N_1534,In_817,In_1564);
and U1535 (N_1535,In_3980,In_1178);
xor U1536 (N_1536,In_3371,In_2828);
nor U1537 (N_1537,In_406,In_1235);
nand U1538 (N_1538,In_4137,In_4295);
or U1539 (N_1539,In_4716,In_318);
xor U1540 (N_1540,In_3062,In_2377);
and U1541 (N_1541,In_527,In_994);
xor U1542 (N_1542,In_3005,In_3326);
nand U1543 (N_1543,In_603,In_971);
nor U1544 (N_1544,In_2605,In_1879);
and U1545 (N_1545,In_3705,In_4650);
nor U1546 (N_1546,In_4941,In_2026);
or U1547 (N_1547,In_4788,In_3035);
and U1548 (N_1548,In_4852,In_3871);
nor U1549 (N_1549,In_3295,In_3276);
and U1550 (N_1550,In_804,In_4632);
nor U1551 (N_1551,In_2254,In_4818);
xnor U1552 (N_1552,In_4091,In_4437);
nor U1553 (N_1553,In_4222,In_3958);
nand U1554 (N_1554,In_3474,In_2666);
nor U1555 (N_1555,In_3967,In_4286);
or U1556 (N_1556,In_186,In_1147);
or U1557 (N_1557,In_403,In_3435);
nand U1558 (N_1558,In_3235,In_3574);
xor U1559 (N_1559,In_4355,In_1701);
and U1560 (N_1560,In_4585,In_4476);
nand U1561 (N_1561,In_2707,In_2566);
nand U1562 (N_1562,In_1584,In_495);
and U1563 (N_1563,In_968,In_3089);
nand U1564 (N_1564,In_4532,In_1074);
xnor U1565 (N_1565,In_597,In_4611);
nand U1566 (N_1566,In_3286,In_229);
and U1567 (N_1567,In_1346,In_2286);
nor U1568 (N_1568,In_790,In_813);
or U1569 (N_1569,In_1813,In_4721);
xor U1570 (N_1570,In_1861,In_4370);
nand U1571 (N_1571,In_3278,In_3840);
and U1572 (N_1572,In_4686,In_4339);
nor U1573 (N_1573,In_2404,In_284);
and U1574 (N_1574,In_68,In_600);
and U1575 (N_1575,In_1412,In_2245);
nand U1576 (N_1576,In_253,In_1652);
nor U1577 (N_1577,In_1960,In_2138);
nand U1578 (N_1578,In_3934,In_1532);
and U1579 (N_1579,In_3901,In_4309);
nand U1580 (N_1580,In_388,In_1656);
xor U1581 (N_1581,In_4093,In_4207);
nor U1582 (N_1582,In_3977,In_1772);
nand U1583 (N_1583,In_1190,In_3890);
nand U1584 (N_1584,In_777,In_2177);
and U1585 (N_1585,In_3440,In_845);
nand U1586 (N_1586,In_3323,In_1551);
nand U1587 (N_1587,In_2276,In_3642);
nor U1588 (N_1588,In_497,In_2025);
or U1589 (N_1589,In_4084,In_917);
nor U1590 (N_1590,In_1996,In_4866);
nand U1591 (N_1591,In_2251,In_1481);
xor U1592 (N_1592,In_3338,In_750);
nor U1593 (N_1593,In_4318,In_2951);
xnor U1594 (N_1594,In_3939,In_3381);
nor U1595 (N_1595,In_1297,In_1491);
or U1596 (N_1596,In_2942,In_3459);
nor U1597 (N_1597,In_4288,In_4151);
xnor U1598 (N_1598,In_3116,In_4734);
nor U1599 (N_1599,In_2356,In_1218);
and U1600 (N_1600,In_2592,In_3098);
nor U1601 (N_1601,In_825,In_4485);
or U1602 (N_1602,In_1755,In_1697);
nand U1603 (N_1603,In_3131,In_1217);
and U1604 (N_1604,In_2796,In_4810);
xor U1605 (N_1605,In_311,In_2609);
nand U1606 (N_1606,In_1643,In_257);
xor U1607 (N_1607,In_154,In_1663);
nand U1608 (N_1608,In_3342,In_394);
or U1609 (N_1609,In_1672,In_1396);
and U1610 (N_1610,In_2146,In_3936);
nand U1611 (N_1611,In_3250,In_3024);
nor U1612 (N_1612,In_64,In_1069);
nand U1613 (N_1613,In_3464,In_2836);
xnor U1614 (N_1614,In_2618,In_4949);
or U1615 (N_1615,In_3245,In_853);
nand U1616 (N_1616,In_573,In_4076);
nor U1617 (N_1617,In_2441,In_124);
and U1618 (N_1618,In_2523,In_244);
xor U1619 (N_1619,In_3990,In_3055);
xnor U1620 (N_1620,In_3619,In_4990);
or U1621 (N_1621,In_4063,In_3768);
nand U1622 (N_1622,In_3302,In_4806);
or U1623 (N_1623,In_3339,In_756);
and U1624 (N_1624,In_4916,In_4012);
nor U1625 (N_1625,In_4032,In_3165);
xnor U1626 (N_1626,In_2424,In_2510);
and U1627 (N_1627,In_3513,In_4760);
nor U1628 (N_1628,In_719,In_224);
nand U1629 (N_1629,In_2668,In_536);
and U1630 (N_1630,In_3852,In_243);
nand U1631 (N_1631,In_6,In_2827);
xnor U1632 (N_1632,In_2862,In_299);
nor U1633 (N_1633,In_4496,In_1568);
nor U1634 (N_1634,In_4429,In_3410);
nor U1635 (N_1635,In_4846,In_3274);
and U1636 (N_1636,In_3660,In_2346);
and U1637 (N_1637,In_4191,In_4733);
nor U1638 (N_1638,In_1220,In_1896);
nand U1639 (N_1639,In_264,In_664);
nand U1640 (N_1640,In_2023,In_352);
nor U1641 (N_1641,In_1087,In_281);
or U1642 (N_1642,In_4535,In_2081);
or U1643 (N_1643,In_4658,In_2459);
and U1644 (N_1644,In_3029,In_4165);
xor U1645 (N_1645,In_3333,In_4921);
xnor U1646 (N_1646,In_608,In_351);
nand U1647 (N_1647,In_3357,In_4212);
nor U1648 (N_1648,In_4500,In_823);
xor U1649 (N_1649,In_4748,In_3573);
nand U1650 (N_1650,In_3288,In_4110);
nor U1651 (N_1651,In_3792,In_1489);
nor U1652 (N_1652,In_1699,In_4036);
nand U1653 (N_1653,In_980,In_672);
and U1654 (N_1654,In_3651,In_2570);
xor U1655 (N_1655,In_3407,In_3656);
xor U1656 (N_1656,In_1286,In_3081);
or U1657 (N_1657,In_3225,In_4825);
nand U1658 (N_1658,In_4113,In_324);
and U1659 (N_1659,In_3321,In_1505);
nand U1660 (N_1660,In_2422,In_3913);
xnor U1661 (N_1661,In_2744,In_645);
xnor U1662 (N_1662,In_1525,In_2059);
nand U1663 (N_1663,In_3114,In_1428);
and U1664 (N_1664,In_3719,In_3468);
or U1665 (N_1665,In_3726,In_78);
nor U1666 (N_1666,In_4176,In_4157);
xnor U1667 (N_1667,In_4516,In_500);
nand U1668 (N_1668,In_23,In_2367);
nand U1669 (N_1669,In_3264,In_2952);
and U1670 (N_1670,In_4718,In_1538);
and U1671 (N_1671,In_2486,In_3972);
nand U1672 (N_1672,In_1329,In_377);
and U1673 (N_1673,In_2644,In_692);
xor U1674 (N_1674,In_289,In_404);
or U1675 (N_1675,In_3334,In_4668);
or U1676 (N_1676,In_4617,In_4763);
nor U1677 (N_1677,In_4977,In_1018);
xor U1678 (N_1678,In_2826,In_108);
nor U1679 (N_1679,In_739,In_2487);
nor U1680 (N_1680,In_2444,In_4371);
and U1681 (N_1681,In_4795,In_157);
and U1682 (N_1682,In_4785,In_4031);
or U1683 (N_1683,In_3400,In_995);
xor U1684 (N_1684,In_1422,In_3058);
or U1685 (N_1685,In_5,In_3744);
xor U1686 (N_1686,In_2354,In_2845);
nand U1687 (N_1687,In_2625,In_2563);
and U1688 (N_1688,In_2615,In_1989);
nor U1689 (N_1689,In_1138,In_2760);
or U1690 (N_1690,In_1168,In_3038);
nand U1691 (N_1691,In_2878,In_4171);
xor U1692 (N_1692,In_3662,In_417);
xnor U1693 (N_1693,In_389,In_2758);
nand U1694 (N_1694,In_3788,In_3776);
nor U1695 (N_1695,In_3003,In_4104);
nand U1696 (N_1696,In_3849,In_3706);
or U1697 (N_1697,In_2980,In_4713);
nand U1698 (N_1698,In_1882,In_1785);
and U1699 (N_1699,In_2953,In_2740);
or U1700 (N_1700,In_162,In_4955);
and U1701 (N_1701,In_4262,In_682);
or U1702 (N_1702,In_2082,In_140);
and U1703 (N_1703,In_613,In_1034);
nor U1704 (N_1704,In_3877,In_802);
nand U1705 (N_1705,In_2831,In_1264);
xor U1706 (N_1706,In_3228,In_2518);
xnor U1707 (N_1707,In_1660,In_885);
xnor U1708 (N_1708,In_2141,In_1274);
nor U1709 (N_1709,In_4200,In_1000);
and U1710 (N_1710,In_2388,In_1197);
nor U1711 (N_1711,In_1599,In_2453);
nor U1712 (N_1712,In_2192,In_611);
nor U1713 (N_1713,In_4978,In_1206);
and U1714 (N_1714,In_591,In_3320);
nand U1715 (N_1715,In_3201,In_957);
xnor U1716 (N_1716,In_761,In_3577);
or U1717 (N_1717,In_4699,In_2516);
nor U1718 (N_1718,In_4039,In_3711);
xor U1719 (N_1719,In_3732,In_2950);
nor U1720 (N_1720,In_1294,In_454);
and U1721 (N_1721,In_3959,In_712);
or U1722 (N_1722,In_2052,In_118);
and U1723 (N_1723,In_3315,In_73);
xnor U1724 (N_1724,In_1504,In_2852);
or U1725 (N_1725,In_4871,In_385);
and U1726 (N_1726,In_4954,In_1267);
nor U1727 (N_1727,In_643,In_184);
and U1728 (N_1728,In_4669,In_1722);
or U1729 (N_1729,In_2743,In_4673);
xnor U1730 (N_1730,In_1209,In_1858);
nor U1731 (N_1731,In_4348,In_1044);
nor U1732 (N_1732,In_4005,In_4973);
and U1733 (N_1733,In_609,In_1827);
or U1734 (N_1734,In_1467,In_34);
nand U1735 (N_1735,In_3036,In_2170);
nand U1736 (N_1736,In_4918,In_2501);
or U1737 (N_1737,In_3820,In_2287);
and U1738 (N_1738,In_1447,In_1052);
or U1739 (N_1739,In_2841,In_2875);
nor U1740 (N_1740,In_212,In_1327);
nor U1741 (N_1741,In_3053,In_1341);
xnor U1742 (N_1742,In_4354,In_3998);
or U1743 (N_1743,In_1350,In_80);
and U1744 (N_1744,In_3246,In_4745);
or U1745 (N_1745,In_1745,In_1310);
and U1746 (N_1746,In_3000,In_2754);
xnor U1747 (N_1747,In_2791,In_1193);
or U1748 (N_1748,In_4882,In_809);
nor U1749 (N_1749,In_3895,In_2559);
nand U1750 (N_1750,In_1057,In_579);
nor U1751 (N_1751,In_2539,In_4817);
nor U1752 (N_1752,In_1938,In_799);
and U1753 (N_1753,In_2617,In_4133);
or U1754 (N_1754,In_4715,In_2373);
nand U1755 (N_1755,In_3587,In_1653);
nor U1756 (N_1756,In_2017,In_74);
and U1757 (N_1757,In_2460,In_2322);
and U1758 (N_1758,In_3445,In_2911);
and U1759 (N_1759,In_783,In_2124);
nand U1760 (N_1760,In_152,In_2189);
nand U1761 (N_1761,In_4394,In_4884);
nand U1762 (N_1762,In_1293,In_483);
nand U1763 (N_1763,In_2094,In_341);
and U1764 (N_1764,In_48,In_675);
or U1765 (N_1765,In_3065,In_1842);
and U1766 (N_1766,In_4028,In_4755);
xnor U1767 (N_1767,In_4839,In_370);
or U1768 (N_1768,In_3103,In_3754);
or U1769 (N_1769,In_4423,In_904);
or U1770 (N_1770,In_2640,In_2631);
nand U1771 (N_1771,In_4243,In_4221);
nor U1772 (N_1772,In_4303,In_2466);
or U1773 (N_1773,In_411,In_1696);
nor U1774 (N_1774,In_3077,In_2691);
xnor U1775 (N_1775,In_1809,In_4231);
xor U1776 (N_1776,In_3968,In_4620);
xnor U1777 (N_1777,In_182,In_4697);
and U1778 (N_1778,In_2020,In_1343);
nand U1779 (N_1779,In_4695,In_3447);
nor U1780 (N_1780,In_2281,In_2888);
and U1781 (N_1781,In_793,In_1915);
and U1782 (N_1782,In_1959,In_1473);
or U1783 (N_1783,In_4756,In_4930);
and U1784 (N_1784,In_962,In_1492);
nand U1785 (N_1785,In_3310,In_237);
xor U1786 (N_1786,In_4544,In_694);
nor U1787 (N_1787,In_4294,In_607);
xnor U1788 (N_1788,In_4626,In_4037);
and U1789 (N_1789,In_2337,In_2386);
xnor U1790 (N_1790,In_3585,In_2590);
xor U1791 (N_1791,In_2909,In_4405);
nor U1792 (N_1792,In_1271,In_1594);
and U1793 (N_1793,In_482,In_551);
nor U1794 (N_1794,In_1355,In_3316);
nand U1795 (N_1795,In_225,In_4879);
nand U1796 (N_1796,In_4635,In_1958);
and U1797 (N_1797,In_1066,In_977);
nand U1798 (N_1798,In_4928,In_3684);
nand U1799 (N_1799,In_2463,In_1512);
xnor U1800 (N_1800,In_2809,In_2517);
nand U1801 (N_1801,In_1887,In_3731);
xnor U1802 (N_1802,In_1369,In_3850);
nand U1803 (N_1803,In_3839,In_3509);
or U1804 (N_1804,In_2172,In_2964);
and U1805 (N_1805,In_51,In_1703);
or U1806 (N_1806,In_2333,In_2366);
nor U1807 (N_1807,In_3284,In_1462);
or U1808 (N_1808,In_4655,In_4445);
and U1809 (N_1809,In_2069,In_1205);
xnor U1810 (N_1810,In_129,In_3056);
or U1811 (N_1811,In_4366,In_2430);
or U1812 (N_1812,In_3908,In_233);
nand U1813 (N_1813,In_363,In_1674);
or U1814 (N_1814,In_2236,In_4943);
nand U1815 (N_1815,In_3742,In_1431);
and U1816 (N_1816,In_4993,In_3949);
and U1817 (N_1817,In_4483,In_2712);
nor U1818 (N_1818,In_2695,In_3601);
nor U1819 (N_1819,In_3500,In_2295);
nor U1820 (N_1820,In_1103,In_4466);
xnor U1821 (N_1821,In_4932,In_3737);
xor U1822 (N_1822,In_2832,In_1405);
nand U1823 (N_1823,In_870,In_1090);
or U1824 (N_1824,In_3027,In_612);
nand U1825 (N_1825,In_3515,In_2753);
and U1826 (N_1826,In_935,In_2770);
nand U1827 (N_1827,In_3843,In_786);
nor U1828 (N_1828,In_3202,In_3227);
nor U1829 (N_1829,In_4349,In_849);
xor U1830 (N_1830,In_2868,In_1654);
and U1831 (N_1831,In_3987,In_906);
or U1832 (N_1832,In_4351,In_2548);
xnor U1833 (N_1833,In_4484,In_2610);
nand U1834 (N_1834,In_1585,In_4446);
nor U1835 (N_1835,In_1445,In_2565);
xor U1836 (N_1836,In_2182,In_3093);
or U1837 (N_1837,In_1231,In_4403);
xnor U1838 (N_1838,In_1583,In_3287);
nor U1839 (N_1839,In_1884,In_1805);
and U1840 (N_1840,In_4489,In_1806);
xnor U1841 (N_1841,In_3146,In_1243);
or U1842 (N_1842,In_701,In_816);
nor U1843 (N_1843,In_2993,In_3394);
xnor U1844 (N_1844,In_945,In_727);
or U1845 (N_1845,In_1929,In_1682);
or U1846 (N_1846,In_3397,In_415);
xnor U1847 (N_1847,In_4661,In_4324);
xor U1848 (N_1848,In_4737,In_2371);
xnor U1849 (N_1849,In_2999,In_1510);
and U1850 (N_1850,In_4293,In_1761);
or U1851 (N_1851,In_3884,In_1638);
nor U1852 (N_1852,In_2148,In_179);
nand U1853 (N_1853,In_3299,In_623);
xor U1854 (N_1854,In_164,In_3389);
xnor U1855 (N_1855,In_4337,In_733);
nor U1856 (N_1856,In_2779,In_173);
nand U1857 (N_1857,In_2316,In_797);
nor U1858 (N_1858,In_3634,In_4159);
nor U1859 (N_1859,In_3576,In_2606);
nand U1860 (N_1860,In_1088,In_855);
or U1861 (N_1861,In_3140,In_1972);
nor U1862 (N_1862,In_766,In_1736);
xor U1863 (N_1863,In_4427,In_1631);
xnor U1864 (N_1864,In_2104,In_1839);
xnor U1865 (N_1865,In_4455,In_2314);
nor U1866 (N_1866,In_792,In_3489);
nand U1867 (N_1867,In_44,In_3008);
and U1868 (N_1868,In_4799,In_2270);
or U1869 (N_1869,In_911,In_4518);
xnor U1870 (N_1870,In_3073,In_4630);
or U1871 (N_1871,In_2,In_3398);
and U1872 (N_1872,In_1225,In_156);
nor U1873 (N_1873,In_976,In_1524);
and U1874 (N_1874,In_4602,In_2035);
xor U1875 (N_1875,In_847,In_1276);
or U1876 (N_1876,In_3693,In_4569);
or U1877 (N_1877,In_3860,In_1155);
and U1878 (N_1878,In_1295,In_2010);
or U1879 (N_1879,In_990,In_3516);
and U1880 (N_1880,In_3785,In_1775);
and U1881 (N_1881,In_3057,In_2540);
nor U1882 (N_1882,In_3230,In_620);
nor U1883 (N_1883,In_2600,In_3530);
nand U1884 (N_1884,In_4904,In_4344);
or U1885 (N_1885,In_1756,In_1425);
nand U1886 (N_1886,In_2419,In_3117);
nand U1887 (N_1887,In_1903,In_4717);
and U1888 (N_1888,In_350,In_3547);
and U1889 (N_1889,In_1300,In_3063);
or U1890 (N_1890,In_251,In_1157);
nand U1891 (N_1891,In_3563,In_1429);
nand U1892 (N_1892,In_2913,In_4422);
xor U1893 (N_1893,In_3525,In_4053);
nand U1894 (N_1894,In_942,In_2494);
nand U1895 (N_1895,In_3802,In_3191);
nor U1896 (N_1896,In_3875,In_3457);
nor U1897 (N_1897,In_4078,In_1680);
or U1898 (N_1898,In_938,In_1823);
and U1899 (N_1899,In_2698,In_3770);
nand U1900 (N_1900,In_4600,In_4002);
nor U1901 (N_1901,In_4714,In_4894);
nor U1902 (N_1902,In_2934,In_2893);
or U1903 (N_1903,In_3830,In_1064);
and U1904 (N_1904,In_4982,In_3049);
nand U1905 (N_1905,In_2525,In_1625);
xor U1906 (N_1906,In_3034,In_3954);
nand U1907 (N_1907,In_2854,In_4121);
nor U1908 (N_1908,In_4025,In_877);
xnor U1909 (N_1909,In_1312,In_2520);
and U1910 (N_1910,In_3079,In_3293);
or U1911 (N_1911,In_578,In_3125);
and U1912 (N_1912,In_2089,In_4359);
nand U1913 (N_1913,In_4209,In_1877);
or U1914 (N_1914,In_3519,In_3182);
nor U1915 (N_1915,In_840,In_2175);
and U1916 (N_1916,In_868,In_467);
nor U1917 (N_1917,In_1227,In_3155);
nand U1918 (N_1918,In_1718,In_3200);
or U1919 (N_1919,In_3178,In_3083);
xnor U1920 (N_1920,In_4327,In_686);
xnor U1921 (N_1921,In_4118,In_1931);
xor U1922 (N_1922,In_1127,In_1078);
xnor U1923 (N_1923,In_2768,In_4046);
nand U1924 (N_1924,In_4245,In_1486);
nand U1925 (N_1925,In_3031,In_2360);
nor U1926 (N_1926,In_3094,In_869);
nor U1927 (N_1927,In_2369,In_27);
nor U1928 (N_1928,In_1433,In_197);
nand U1929 (N_1929,In_1207,In_4469);
nand U1930 (N_1930,In_3666,In_3267);
nor U1931 (N_1931,In_2604,In_4096);
or U1932 (N_1932,In_2560,In_3017);
nor U1933 (N_1933,In_3216,In_2815);
nor U1934 (N_1934,In_3011,In_1572);
nor U1935 (N_1935,In_1480,In_1008);
or U1936 (N_1936,In_3544,In_3265);
or U1937 (N_1937,In_276,In_2532);
nor U1938 (N_1938,In_1125,In_2651);
xnor U1939 (N_1939,In_69,In_1768);
and U1940 (N_1940,In_3335,In_4055);
or U1941 (N_1941,In_1783,In_820);
nor U1942 (N_1942,In_4195,In_102);
nor U1943 (N_1943,In_3812,In_358);
and U1944 (N_1944,In_2817,In_3306);
or U1945 (N_1945,In_1098,In_3690);
nand U1946 (N_1946,In_3059,In_458);
nor U1947 (N_1947,In_3905,In_1124);
nand U1948 (N_1948,In_1715,In_2762);
or U1949 (N_1949,In_1598,In_4800);
nand U1950 (N_1950,In_4310,In_1434);
or U1951 (N_1951,In_4304,In_2390);
or U1952 (N_1952,In_581,In_2579);
nor U1953 (N_1953,In_1810,In_936);
xnor U1954 (N_1954,In_4154,In_4022);
nor U1955 (N_1955,In_2006,In_3976);
nand U1956 (N_1956,In_748,In_2880);
nor U1957 (N_1957,In_3676,In_3606);
nand U1958 (N_1958,In_4225,In_2690);
and U1959 (N_1959,In_526,In_1251);
xnor U1960 (N_1960,In_4919,In_3492);
nand U1961 (N_1961,In_2375,In_769);
and U1962 (N_1962,In_4027,In_3630);
and U1963 (N_1963,In_1256,In_3826);
and U1964 (N_1964,In_2856,In_4378);
nor U1965 (N_1965,In_3319,In_2634);
or U1966 (N_1966,In_848,In_277);
or U1967 (N_1967,In_4751,In_3141);
xor U1968 (N_1968,In_3305,In_2211);
nor U1969 (N_1969,In_2309,In_2674);
xnor U1970 (N_1970,In_4075,In_3798);
or U1971 (N_1971,In_307,In_2806);
nor U1972 (N_1972,In_3942,In_4856);
nand U1973 (N_1973,In_405,In_3416);
nor U1974 (N_1974,In_4316,In_1869);
and U1975 (N_1975,In_846,In_2883);
nand U1976 (N_1976,In_3904,In_2357);
and U1977 (N_1977,In_2490,In_4441);
and U1978 (N_1978,In_4313,In_3523);
xnor U1979 (N_1979,In_2063,In_1028);
nand U1980 (N_1980,In_4974,In_3897);
and U1981 (N_1981,In_1773,In_1458);
xor U1982 (N_1982,In_4030,In_924);
nor U1983 (N_1983,In_4073,In_2728);
or U1984 (N_1984,In_2923,In_4062);
nor U1985 (N_1985,In_99,In_4424);
nand U1986 (N_1986,In_3556,In_3115);
xnor U1987 (N_1987,In_3593,In_1615);
xor U1988 (N_1988,In_1610,In_3882);
nand U1989 (N_1989,In_523,In_3975);
xor U1990 (N_1990,In_779,In_2677);
nor U1991 (N_1991,In_3560,In_2102);
and U1992 (N_1992,In_3456,In_1273);
and U1993 (N_1993,In_2068,In_4522);
nor U1994 (N_1994,In_1769,In_563);
nor U1995 (N_1995,In_819,In_639);
and U1996 (N_1996,In_4988,In_2585);
xor U1997 (N_1997,In_1065,In_1685);
xor U1998 (N_1998,In_4905,In_2060);
nand U1999 (N_1999,In_2769,In_4765);
or U2000 (N_2000,In_209,In_2738);
nand U2001 (N_2001,In_1780,In_1150);
or U2002 (N_2002,In_512,In_2096);
nand U2003 (N_2003,In_4876,In_4089);
and U2004 (N_2004,In_1011,In_4768);
or U2005 (N_2005,In_3373,In_532);
nand U2006 (N_2006,In_3748,In_2262);
nand U2007 (N_2007,In_1374,In_4675);
nor U2008 (N_2008,In_4217,In_4067);
xnor U2009 (N_2009,In_1592,In_1751);
nor U2010 (N_2010,In_3864,In_3743);
xnor U2011 (N_2011,In_1726,In_207);
or U2012 (N_2012,In_3767,In_3602);
or U2013 (N_2013,In_1357,In_1305);
xor U2014 (N_2014,In_3906,In_2722);
xor U2015 (N_2015,In_1086,In_4834);
or U2016 (N_2016,In_180,In_3179);
and U2017 (N_2017,In_379,In_1816);
and U2018 (N_2018,In_1451,In_4560);
nor U2019 (N_2019,In_211,In_574);
or U2020 (N_2020,In_4196,In_3956);
nor U2021 (N_2021,In_4971,In_1763);
nor U2022 (N_2022,In_2937,In_2142);
xor U2023 (N_2023,In_661,In_4311);
xnor U2024 (N_2024,In_30,In_4481);
nor U2025 (N_2025,In_4723,In_2724);
nor U2026 (N_2026,In_1578,In_1245);
or U2027 (N_2027,In_1530,In_3947);
nor U2028 (N_2028,In_1880,In_2546);
nand U2029 (N_2029,In_767,In_839);
or U2030 (N_2030,In_3325,In_4453);
xnor U2031 (N_2031,In_3701,In_2101);
and U2032 (N_2032,In_172,In_693);
nor U2033 (N_2033,In_4578,In_4282);
and U2034 (N_2034,In_4761,In_4575);
xor U2035 (N_2035,In_1767,In_2264);
nor U2036 (N_2036,In_3272,In_3112);
and U2037 (N_2037,In_2005,In_568);
and U2038 (N_2038,In_2816,In_2508);
nand U2039 (N_2039,In_2212,In_3896);
xnor U2040 (N_2040,In_2303,In_11);
nand U2041 (N_2041,In_4681,In_3331);
and U2042 (N_2042,In_3022,In_4474);
nand U2043 (N_2043,In_2886,In_4428);
xor U2044 (N_2044,In_3582,In_133);
nor U2045 (N_2045,In_703,In_3714);
or U2046 (N_2046,In_1202,In_3858);
nand U2047 (N_2047,In_1181,In_1430);
and U2048 (N_2048,In_1782,In_3123);
nor U2049 (N_2049,In_4730,In_4649);
or U2050 (N_2050,In_4610,In_2932);
xnor U2051 (N_2051,In_1837,In_1116);
nor U2052 (N_2052,In_752,In_1162);
xnor U2053 (N_2053,In_1539,In_4343);
and U2054 (N_2054,In_1885,In_3615);
or U2055 (N_2055,In_1356,In_842);
xor U2056 (N_2056,In_1930,In_2848);
and U2057 (N_2057,In_624,In_4457);
or U2058 (N_2058,In_4203,In_4859);
nand U2059 (N_2059,In_4625,In_4891);
nand U2060 (N_2060,In_886,In_3391);
or U2061 (N_2061,In_301,In_768);
nor U2062 (N_2062,In_2990,In_1621);
and U2063 (N_2063,In_4128,In_584);
and U2064 (N_2064,In_4150,In_4319);
nor U2065 (N_2065,In_4461,In_1843);
nor U2066 (N_2066,In_1855,In_4660);
nand U2067 (N_2067,In_2894,In_2306);
nor U2068 (N_2068,In_3296,In_4214);
nor U2069 (N_2069,In_3794,In_1831);
or U2070 (N_2070,In_3769,In_4862);
xor U2071 (N_2071,In_2297,In_3236);
nand U2072 (N_2072,In_2218,In_2860);
nor U2073 (N_2073,In_119,In_1740);
nor U2074 (N_2074,In_2576,In_2865);
nand U2075 (N_2075,In_1570,In_2733);
nor U2076 (N_2076,In_295,In_2558);
and U2077 (N_2077,In_366,In_113);
xor U2078 (N_2078,In_1033,In_2240);
nor U2079 (N_2079,In_1688,In_3777);
nor U2080 (N_2080,In_4753,In_1894);
xnor U2081 (N_2081,In_4590,In_413);
nand U2082 (N_2082,In_4684,In_1446);
nor U2083 (N_2083,In_1019,In_3911);
and U2084 (N_2084,In_1092,In_3271);
and U2085 (N_2085,In_4588,In_2358);
and U2086 (N_2086,In_3156,In_3465);
and U2087 (N_2087,In_4462,In_4488);
nand U2088 (N_2088,In_1345,In_2134);
nand U2089 (N_2089,In_2061,In_4201);
xnor U2090 (N_2090,In_1145,In_4627);
nor U2091 (N_2091,In_1398,In_2057);
xor U2092 (N_2092,In_3080,In_4182);
and U2093 (N_2093,In_2415,In_4843);
nand U2094 (N_2094,In_1037,In_1095);
nor U2095 (N_2095,In_1046,In_803);
or U2096 (N_2096,In_2435,In_3032);
or U2097 (N_2097,In_625,In_1946);
xor U2098 (N_2098,In_3453,In_2135);
and U2099 (N_2099,In_2777,In_1200);
xnor U2100 (N_2100,In_1662,In_4898);
or U2101 (N_2101,In_4855,In_650);
and U2102 (N_2102,In_1272,In_2715);
or U2103 (N_2103,In_3951,In_4688);
and U2104 (N_2104,In_1945,In_2340);
xnor U2105 (N_2105,In_4693,In_1342);
and U2106 (N_2106,In_2153,In_2041);
xnor U2107 (N_2107,In_3847,In_3786);
and U2108 (N_2108,In_1322,In_2269);
and U2109 (N_2109,In_755,In_1362);
xor U2110 (N_2110,In_346,In_3184);
xor U2111 (N_2111,In_2470,In_3527);
xor U2112 (N_2112,In_4758,In_360);
nor U2113 (N_2113,In_4526,In_2083);
xor U2114 (N_2114,In_188,In_3118);
xnor U2115 (N_2115,In_136,In_3442);
nor U2116 (N_2116,In_3484,In_419);
and U2117 (N_2117,In_4777,In_1521);
or U2118 (N_2118,In_1468,In_572);
or U2119 (N_2119,In_4079,In_4415);
xor U2120 (N_2120,In_1130,In_4497);
or U2121 (N_2121,In_4198,In_2263);
nor U2122 (N_2122,In_3800,In_3589);
or U2123 (N_2123,In_220,In_2897);
nor U2124 (N_2124,In_4967,In_3745);
nand U2125 (N_2125,In_3971,In_2349);
nand U2126 (N_2126,In_3715,In_1828);
xnor U2127 (N_2127,In_3451,In_2641);
and U2128 (N_2128,In_1710,In_1632);
nor U2129 (N_2129,In_3680,In_399);
nand U2130 (N_2130,In_1199,In_1678);
and U2131 (N_2131,In_2741,In_3070);
nand U2132 (N_2132,In_3344,In_1913);
xor U2133 (N_2133,In_3455,In_2477);
xnor U2134 (N_2134,In_3350,In_3300);
nor U2135 (N_2135,In_2745,In_322);
or U2136 (N_2136,In_2842,In_2406);
or U2137 (N_2137,In_2623,In_1262);
nand U2138 (N_2138,In_228,In_4472);
or U2139 (N_2139,In_4594,In_1797);
nor U2140 (N_2140,In_3009,In_3845);
nand U2141 (N_2141,In_615,In_685);
and U2142 (N_2142,In_1914,In_638);
xnor U2143 (N_2143,In_1171,In_1977);
nor U2144 (N_2144,In_3823,In_3517);
or U2145 (N_2145,In_371,In_3824);
or U2146 (N_2146,In_3164,In_367);
xnor U2147 (N_2147,In_386,In_4246);
and U2148 (N_2148,In_2399,In_4368);
xnor U2149 (N_2149,In_770,In_3279);
nand U2150 (N_2150,In_1361,In_4145);
or U2151 (N_2151,In_3252,In_1698);
nor U2152 (N_2152,In_3471,In_1249);
nor U2153 (N_2153,In_2938,In_2229);
and U2154 (N_2154,In_4275,In_3810);
or U2155 (N_2155,In_4268,In_708);
nor U2156 (N_2156,In_1793,In_2611);
or U2157 (N_2157,In_2258,In_7);
or U2158 (N_2158,In_4914,In_788);
xor U2159 (N_2159,In_2658,In_1403);
nand U2160 (N_2160,In_865,In_2957);
xnor U2161 (N_2161,In_2859,In_39);
xor U2162 (N_2162,In_2046,In_3097);
xnor U2163 (N_2163,In_2157,In_3825);
xor U2164 (N_2164,In_2048,In_2418);
nand U2165 (N_2165,In_3449,In_3603);
nor U2166 (N_2166,In_3730,In_1758);
nand U2167 (N_2167,In_3653,In_2439);
and U2168 (N_2168,In_2042,In_4576);
nor U2169 (N_2169,In_1,In_4345);
nand U2170 (N_2170,In_4573,In_1857);
or U2171 (N_2171,In_4566,In_548);
nor U2172 (N_2172,In_2433,In_4279);
or U2173 (N_2173,In_440,In_605);
xnor U2174 (N_2174,In_20,In_3044);
nor U2175 (N_2175,In_2703,In_265);
and U2176 (N_2176,In_1511,In_4419);
xor U2177 (N_2177,In_4435,In_3001);
nor U2178 (N_2178,In_2529,In_812);
nand U2179 (N_2179,In_2255,In_3161);
xnor U2180 (N_2180,In_2001,In_567);
or U2181 (N_2181,In_1752,In_2066);
xnor U2182 (N_2182,In_2401,In_2140);
nor U2183 (N_2183,In_2412,In_3359);
and U2184 (N_2184,In_4584,In_3614);
nor U2185 (N_2185,In_4480,In_4647);
nor U2186 (N_2186,In_4652,In_67);
nor U2187 (N_2187,In_4562,In_569);
or U2188 (N_2188,In_4248,In_1847);
or U2189 (N_2189,In_4372,In_4155);
nor U2190 (N_2190,In_660,In_3257);
nand U2191 (N_2191,In_256,In_2203);
nor U2192 (N_2192,In_286,In_213);
and U2193 (N_2193,In_2922,In_1627);
xor U2194 (N_2194,In_3790,In_3944);
and U2195 (N_2195,In_407,In_988);
and U2196 (N_2196,In_2423,In_2293);
nand U2197 (N_2197,In_3599,In_4824);
and U2198 (N_2198,In_49,In_2542);
nor U2199 (N_2199,In_3086,In_1443);
xor U2200 (N_2200,In_1898,In_1727);
nor U2201 (N_2201,In_1817,In_2647);
nor U2202 (N_2202,In_203,In_4332);
and U2203 (N_2203,In_3356,In_4547);
or U2204 (N_2204,In_2503,In_1544);
and U2205 (N_2205,In_3665,In_1236);
xor U2206 (N_2206,In_451,In_3521);
nand U2207 (N_2207,In_1759,In_1192);
xor U2208 (N_2208,In_3322,In_4376);
and U2209 (N_2209,In_2926,In_1180);
nor U2210 (N_2210,In_3969,In_4387);
xor U2211 (N_2211,In_2571,In_4583);
nor U2212 (N_2212,In_3941,In_177);
xnor U2213 (N_2213,In_1455,In_763);
nand U2214 (N_2214,In_423,In_932);
nand U2215 (N_2215,In_4130,In_3072);
nand U2216 (N_2216,In_56,In_2335);
xnor U2217 (N_2217,In_3233,In_3808);
or U2218 (N_2218,In_456,In_4558);
xnor U2219 (N_2219,In_2299,In_4381);
xor U2220 (N_2220,In_4850,In_2997);
xnor U2221 (N_2221,In_673,In_1030);
and U2222 (N_2222,In_1799,In_3154);
and U2223 (N_2223,In_1874,In_4397);
xnor U2224 (N_2224,In_2178,In_3962);
xnor U2225 (N_2225,In_1634,In_637);
nand U2226 (N_2226,In_546,In_1905);
nor U2227 (N_2227,In_4870,In_4672);
nor U2228 (N_2228,In_3095,In_873);
nor U2229 (N_2229,In_1531,In_3429);
and U2230 (N_2230,In_1470,In_1247);
and U2231 (N_2231,In_1586,In_4671);
and U2232 (N_2232,In_2467,In_3106);
nor U2233 (N_2233,In_3148,In_1667);
nor U2234 (N_2234,In_2927,In_3571);
or U2235 (N_2235,In_3430,In_4487);
nor U2236 (N_2236,In_2330,In_1027);
nor U2237 (N_2237,In_2983,In_101);
nand U2238 (N_2238,In_1961,In_1717);
nor U2239 (N_2239,In_634,In_562);
and U2240 (N_2240,In_4557,In_2429);
and U2241 (N_2241,In_2765,In_2384);
and U2242 (N_2242,In_1275,In_4506);
or U2243 (N_2243,In_4135,In_4102);
or U2244 (N_2244,In_110,In_2323);
or U2245 (N_2245,In_268,In_4029);
and U2246 (N_2246,In_4909,In_444);
nand U2247 (N_2247,In_2223,In_683);
or U2248 (N_2248,In_398,In_2946);
and U2249 (N_2249,In_4454,In_4404);
nor U2250 (N_2250,In_1233,In_2221);
or U2251 (N_2251,In_3159,In_3176);
and U2252 (N_2252,In_1315,In_1031);
nor U2253 (N_2253,In_4651,In_2207);
nor U2254 (N_2254,In_4421,In_3575);
nand U2255 (N_2255,In_234,In_3285);
and U2256 (N_2256,In_3051,In_1395);
and U2257 (N_2257,In_2885,In_4881);
nand U2258 (N_2258,In_2252,In_14);
or U2259 (N_2259,In_1671,In_2235);
or U2260 (N_2260,In_4822,In_1035);
nand U2261 (N_2261,In_4451,In_4783);
nand U2262 (N_2262,In_1975,In_4543);
or U2263 (N_2263,In_2324,In_3313);
xor U2264 (N_2264,In_4985,In_2500);
or U2265 (N_2265,In_3144,In_4033);
and U2266 (N_2266,In_3716,In_4875);
xnor U2267 (N_2267,In_1055,In_3304);
xnor U2268 (N_2268,In_4350,In_1734);
and U2269 (N_2269,In_1724,In_2338);
xor U2270 (N_2270,In_3087,In_16);
xnor U2271 (N_2271,In_2108,In_4126);
nand U2272 (N_2272,In_4463,In_1875);
and U2273 (N_2273,In_202,In_1085);
and U2274 (N_2274,In_1499,In_1459);
or U2275 (N_2275,In_801,In_2103);
nor U2276 (N_2276,In_4,In_4285);
nand U2277 (N_2277,In_2473,In_3970);
nor U2278 (N_2278,In_4255,In_3678);
and U2279 (N_2279,In_4443,In_1819);
xnor U2280 (N_2280,In_1824,In_4770);
xnor U2281 (N_2281,In_814,In_2686);
and U2282 (N_2282,In_1795,In_2550);
xor U2283 (N_2283,In_3308,In_3846);
or U2284 (N_2284,In_1372,In_2935);
nand U2285 (N_2285,In_47,In_3865);
xnor U2286 (N_2286,In_2074,In_1692);
xor U2287 (N_2287,In_3774,In_1922);
nor U2288 (N_2288,In_543,In_1076);
and U2289 (N_2289,In_561,In_433);
or U2290 (N_2290,In_2033,In_4937);
and U2291 (N_2291,In_2867,In_3085);
xor U2292 (N_2292,In_2231,In_2637);
or U2293 (N_2293,In_2968,In_1388);
or U2294 (N_2294,In_3624,In_2462);
or U2295 (N_2295,In_718,In_2784);
xnor U2296 (N_2296,In_3431,In_339);
or U2297 (N_2297,In_3579,In_571);
or U2298 (N_2298,In_2727,In_2562);
and U2299 (N_2299,In_1417,In_3082);
nor U2300 (N_2300,In_4361,In_4657);
nor U2301 (N_2301,In_4619,In_4138);
and U2302 (N_2302,In_3835,In_2107);
nor U2303 (N_2303,In_4634,In_800);
or U2304 (N_2304,In_3497,In_3572);
nor U2305 (N_2305,In_1123,In_4147);
nor U2306 (N_2306,In_141,In_3142);
and U2307 (N_2307,In_1801,In_4807);
nand U2308 (N_2308,In_2482,In_4929);
nand U2309 (N_2309,In_25,In_4833);
xnor U2310 (N_2310,In_2960,In_1408);
or U2311 (N_2311,In_1777,In_1951);
and U2312 (N_2312,In_640,In_2085);
or U2313 (N_2313,In_3470,In_2191);
and U2314 (N_2314,In_1826,In_4103);
nor U2315 (N_2315,In_3266,In_3867);
nand U2316 (N_2316,In_3311,In_1479);
nand U2317 (N_2317,In_376,In_2119);
and U2318 (N_2318,In_1971,In_1254);
nor U2319 (N_2319,In_1943,In_1061);
nand U2320 (N_2320,In_3646,In_3483);
nand U2321 (N_2321,In_2168,In_474);
nand U2322 (N_2322,In_1640,In_2736);
xor U2323 (N_2323,In_263,In_109);
xor U2324 (N_2324,In_3487,In_2410);
nand U2325 (N_2325,In_2273,In_3345);
and U2326 (N_2326,In_446,In_4494);
or U2327 (N_2327,In_2133,In_946);
nand U2328 (N_2328,In_3717,In_4864);
nand U2329 (N_2329,In_2372,In_534);
xnor U2330 (N_2330,In_1187,In_4235);
nor U2331 (N_2331,In_2731,In_2661);
nand U2332 (N_2332,In_325,In_4220);
xor U2333 (N_2333,In_1265,In_3401);
nand U2334 (N_2334,In_59,In_3508);
or U2335 (N_2335,In_4426,In_1332);
xnor U2336 (N_2336,In_2380,In_3592);
or U2337 (N_2337,In_1172,In_2709);
xor U2338 (N_2338,In_4065,In_3912);
xnor U2339 (N_2339,In_3747,In_3995);
nand U2340 (N_2340,In_3439,In_123);
or U2341 (N_2341,In_462,In_138);
nor U2342 (N_2342,In_2846,In_1482);
nor U2343 (N_2343,In_2032,In_1003);
nor U2344 (N_2344,In_291,In_1102);
nor U2345 (N_2345,In_1498,In_4329);
and U2346 (N_2346,In_2446,In_2573);
nor U2347 (N_2347,In_2931,In_4885);
nor U2348 (N_2348,In_3403,In_826);
nand U2349 (N_2349,In_1659,In_1956);
xor U2350 (N_2350,In_4616,In_3763);
and U2351 (N_2351,In_691,In_1365);
or U2352 (N_2352,In_262,In_4292);
nand U2353 (N_2353,In_296,In_4732);
nor U2354 (N_2354,In_3595,In_4659);
nor U2355 (N_2355,In_4781,In_2627);
nor U2356 (N_2356,In_4607,In_178);
and U2357 (N_2357,In_789,In_3691);
nand U2358 (N_2358,In_3925,In_2013);
xnor U2359 (N_2359,In_1270,In_3107);
nor U2360 (N_2360,In_2398,In_3441);
or U2361 (N_2361,In_463,In_372);
or U2362 (N_2362,In_775,In_442);
or U2363 (N_2363,In_4744,In_751);
or U2364 (N_2364,In_1784,In_2166);
xnor U2365 (N_2365,In_1416,In_144);
xor U2366 (N_2366,In_4410,In_2718);
xor U2367 (N_2367,In_4889,In_4187);
nand U2368 (N_2368,In_3533,In_1414);
xnor U2369 (N_2369,In_391,In_418);
xor U2370 (N_2370,In_4470,In_1463);
nand U2371 (N_2371,In_1708,In_17);
nor U2372 (N_2372,In_1604,In_1947);
or U2373 (N_2373,In_2277,In_2022);
xnor U2374 (N_2374,In_4449,In_4141);
nor U2375 (N_2375,In_1261,In_618);
and U2376 (N_2376,In_1284,In_949);
xor U2377 (N_2377,In_1567,In_15);
nor U2378 (N_2378,In_176,In_4767);
and U2379 (N_2379,In_4724,In_3183);
xor U2380 (N_2380,In_4623,In_535);
or U2381 (N_2381,In_3251,In_4142);
nor U2382 (N_2382,In_552,In_4491);
and U2383 (N_2383,In_1104,In_2431);
xnor U2384 (N_2384,In_3126,In_4006);
or U2385 (N_2385,In_3880,In_808);
or U2386 (N_2386,In_3374,In_4106);
and U2387 (N_2387,In_4477,In_2551);
nand U2388 (N_2388,In_3787,In_3419);
xnor U2389 (N_2389,In_3713,In_3020);
and U2390 (N_2390,In_3552,In_3781);
nor U2391 (N_2391,In_4549,In_3703);
xor U2392 (N_2392,In_1432,In_4389);
nor U2393 (N_2393,In_2161,In_2930);
or U2394 (N_2394,In_1005,In_717);
xor U2395 (N_2395,In_4194,In_3738);
and U2396 (N_2396,In_4867,In_1203);
nor U2397 (N_2397,In_2259,In_4700);
nor U2398 (N_2398,In_2243,In_43);
nor U2399 (N_2399,In_3428,In_206);
and U2400 (N_2400,In_997,In_2012);
or U2401 (N_2401,In_1115,In_4676);
and U2402 (N_2402,In_2283,In_851);
or U2403 (N_2403,In_582,In_1204);
or U2404 (N_2404,In_2998,In_1888);
or U2405 (N_2405,In_1266,In_4490);
nor U2406 (N_2406,In_4897,In_3695);
or U2407 (N_2407,In_2737,In_1732);
xor U2408 (N_2408,In_1609,In_3659);
nand U2409 (N_2409,In_4694,In_2055);
and U2410 (N_2410,In_1788,In_3999);
or U2411 (N_2411,In_4960,In_65);
or U2412 (N_2412,In_4068,In_2989);
nand U2413 (N_2413,In_2261,In_4264);
nand U2414 (N_2414,In_498,In_1891);
nor U2415 (N_2415,In_4912,In_2489);
nand U2416 (N_2416,In_4074,In_871);
nor U2417 (N_2417,In_3076,In_1800);
nor U2418 (N_2418,In_1017,In_4007);
and U2419 (N_2419,In_2855,In_3196);
nand U2420 (N_2420,In_1378,In_4436);
and U2421 (N_2421,In_4551,In_90);
and U2422 (N_2422,In_517,In_4307);
or U2423 (N_2423,In_3938,In_4924);
and U2424 (N_2424,In_4479,In_2219);
and U2425 (N_2425,In_3640,In_4857);
nand U2426 (N_2426,In_2409,In_4432);
nand U2427 (N_2427,In_2588,In_4581);
or U2428 (N_2428,In_1794,In_4408);
nor U2429 (N_2429,In_1965,In_4570);
nand U2430 (N_2430,In_3277,In_3273);
or U2431 (N_2431,In_1949,In_2291);
or U2432 (N_2432,In_3379,In_2476);
xnor U2433 (N_2433,In_3128,In_3420);
nand U2434 (N_2434,In_1981,In_2795);
nor U2435 (N_2435,In_3303,In_1670);
nand U2436 (N_2436,In_4771,In_678);
nor U2437 (N_2437,In_908,In_1421);
and U2438 (N_2438,In_3255,In_4531);
or U2439 (N_2439,In_3979,In_915);
and U2440 (N_2440,In_3751,In_2233);
and U2441 (N_2441,In_3358,In_1450);
xnor U2442 (N_2442,In_1006,In_200);
and U2443 (N_2443,In_1863,In_983);
or U2444 (N_2444,In_2176,In_4347);
and U2445 (N_2445,In_4308,In_3607);
nor U2446 (N_2446,In_671,In_2578);
nand U2447 (N_2447,In_1522,In_589);
xor U2448 (N_2448,In_1731,In_189);
or U2449 (N_2449,In_2484,In_449);
or U2450 (N_2450,In_1835,In_35);
and U2451 (N_2451,In_3755,In_1993);
or U2452 (N_2452,In_580,In_555);
xor U2453 (N_2453,In_854,In_861);
nor U2454 (N_2454,In_716,In_1496);
or U2455 (N_2455,In_4070,In_3376);
nor U2456 (N_2456,In_1559,In_1684);
nand U2457 (N_2457,In_3291,In_1258);
nor U2458 (N_2458,In_3669,In_4230);
and U2459 (N_2459,In_425,In_85);
xor U2460 (N_2460,In_859,In_4809);
nand U2461 (N_2461,In_3189,In_684);
and U2462 (N_2462,In_747,In_1851);
nor U2463 (N_2463,In_1690,In_2643);
and U2464 (N_2464,In_1807,In_3628);
nand U2465 (N_2465,In_2079,In_3611);
nand U2466 (N_2466,In_1402,In_1375);
xnor U2467 (N_2467,In_3078,In_137);
or U2468 (N_2468,In_1170,In_4273);
xor U2469 (N_2469,In_2699,In_2910);
xnor U2470 (N_2470,In_1211,In_1691);
xnor U2471 (N_2471,In_2851,In_287);
nand U2472 (N_2472,In_3383,In_1655);
xor U2473 (N_2473,In_2692,In_3740);
or U2474 (N_2474,In_2581,In_1808);
xor U2475 (N_2475,In_3170,In_486);
nor U2476 (N_2476,In_2663,In_4204);
nor U2477 (N_2477,In_1094,In_1893);
xnor U2478 (N_2478,In_1401,In_196);
nor U2479 (N_2479,In_1883,In_3369);
or U2480 (N_2480,In_2416,In_3568);
nand U2481 (N_2481,In_2365,In_1336);
xnor U2482 (N_2482,In_695,In_918);
and U2483 (N_2483,In_1523,In_1392);
nand U2484 (N_2484,In_3919,In_3479);
xnor U2485 (N_2485,In_1739,In_3671);
or U2486 (N_2486,In_2171,In_2547);
nor U2487 (N_2487,In_1789,In_3702);
nand U2488 (N_2488,In_344,In_2534);
and U2489 (N_2489,In_4747,In_3495);
or U2490 (N_2490,In_975,In_2788);
or U2491 (N_2491,In_4179,In_2099);
and U2492 (N_2492,In_773,In_3213);
xor U2493 (N_2493,In_255,In_1133);
nor U2494 (N_2494,In_575,In_2933);
or U2495 (N_2495,In_688,In_2665);
and U2496 (N_2496,In_2195,In_221);
xor U2497 (N_2497,In_3145,In_4792);
nor U2498 (N_2498,In_28,In_3425);
nand U2499 (N_2499,In_950,In_46);
xnor U2500 (N_2500,In_216,In_3767);
or U2501 (N_2501,In_825,In_3565);
nand U2502 (N_2502,In_2503,In_2625);
nor U2503 (N_2503,In_4077,In_2912);
nand U2504 (N_2504,In_993,In_187);
nand U2505 (N_2505,In_2688,In_1943);
nor U2506 (N_2506,In_3268,In_905);
xnor U2507 (N_2507,In_1148,In_4351);
or U2508 (N_2508,In_1979,In_1472);
xor U2509 (N_2509,In_1249,In_567);
or U2510 (N_2510,In_2643,In_3902);
nor U2511 (N_2511,In_2219,In_1012);
xor U2512 (N_2512,In_2784,In_2719);
nand U2513 (N_2513,In_1012,In_720);
xor U2514 (N_2514,In_4,In_3011);
nor U2515 (N_2515,In_2894,In_537);
or U2516 (N_2516,In_4388,In_4423);
nor U2517 (N_2517,In_742,In_4508);
and U2518 (N_2518,In_2819,In_3131);
nor U2519 (N_2519,In_1391,In_4084);
xnor U2520 (N_2520,In_2943,In_761);
nand U2521 (N_2521,In_270,In_97);
and U2522 (N_2522,In_2348,In_4430);
xor U2523 (N_2523,In_4174,In_635);
or U2524 (N_2524,In_462,In_2277);
and U2525 (N_2525,In_2746,In_2619);
nor U2526 (N_2526,In_1571,In_720);
xnor U2527 (N_2527,In_3387,In_1028);
and U2528 (N_2528,In_4441,In_2304);
and U2529 (N_2529,In_4906,In_3383);
nor U2530 (N_2530,In_210,In_3908);
or U2531 (N_2531,In_4776,In_539);
nor U2532 (N_2532,In_3773,In_1421);
xnor U2533 (N_2533,In_4857,In_1976);
and U2534 (N_2534,In_2067,In_428);
and U2535 (N_2535,In_4962,In_2763);
xor U2536 (N_2536,In_3071,In_2522);
nor U2537 (N_2537,In_999,In_1312);
or U2538 (N_2538,In_2113,In_2538);
xor U2539 (N_2539,In_4545,In_925);
nand U2540 (N_2540,In_2691,In_1945);
nor U2541 (N_2541,In_1869,In_3199);
xor U2542 (N_2542,In_2194,In_2418);
nand U2543 (N_2543,In_4151,In_4415);
nand U2544 (N_2544,In_4836,In_3420);
or U2545 (N_2545,In_981,In_3407);
nand U2546 (N_2546,In_238,In_4505);
and U2547 (N_2547,In_1350,In_3857);
nor U2548 (N_2548,In_3629,In_1582);
xor U2549 (N_2549,In_1633,In_4773);
nand U2550 (N_2550,In_3466,In_4186);
xor U2551 (N_2551,In_1265,In_1559);
xnor U2552 (N_2552,In_4705,In_557);
or U2553 (N_2553,In_321,In_1928);
nand U2554 (N_2554,In_942,In_1814);
or U2555 (N_2555,In_2142,In_3640);
nor U2556 (N_2556,In_104,In_3463);
nor U2557 (N_2557,In_10,In_1913);
xor U2558 (N_2558,In_3960,In_4117);
or U2559 (N_2559,In_148,In_4997);
nor U2560 (N_2560,In_4905,In_72);
or U2561 (N_2561,In_2873,In_4747);
or U2562 (N_2562,In_425,In_576);
nor U2563 (N_2563,In_4570,In_3810);
or U2564 (N_2564,In_4994,In_1397);
xnor U2565 (N_2565,In_2782,In_3174);
or U2566 (N_2566,In_2087,In_1971);
nand U2567 (N_2567,In_1276,In_4535);
or U2568 (N_2568,In_3795,In_4209);
and U2569 (N_2569,In_3360,In_4031);
nand U2570 (N_2570,In_4477,In_4777);
xor U2571 (N_2571,In_4923,In_1250);
and U2572 (N_2572,In_1663,In_4541);
nor U2573 (N_2573,In_3707,In_3887);
xor U2574 (N_2574,In_3329,In_808);
and U2575 (N_2575,In_1608,In_4313);
nor U2576 (N_2576,In_2173,In_2153);
or U2577 (N_2577,In_1943,In_4637);
nor U2578 (N_2578,In_451,In_2208);
nand U2579 (N_2579,In_3062,In_3486);
or U2580 (N_2580,In_1498,In_2493);
xnor U2581 (N_2581,In_1382,In_3784);
or U2582 (N_2582,In_62,In_4227);
or U2583 (N_2583,In_1791,In_3974);
nand U2584 (N_2584,In_2428,In_1657);
xor U2585 (N_2585,In_4786,In_4358);
nand U2586 (N_2586,In_3248,In_1704);
xor U2587 (N_2587,In_996,In_1752);
or U2588 (N_2588,In_2386,In_4102);
xnor U2589 (N_2589,In_3444,In_932);
and U2590 (N_2590,In_4223,In_302);
nor U2591 (N_2591,In_862,In_1578);
or U2592 (N_2592,In_380,In_4005);
and U2593 (N_2593,In_4583,In_2878);
nor U2594 (N_2594,In_1255,In_2575);
nand U2595 (N_2595,In_858,In_305);
nor U2596 (N_2596,In_2940,In_2655);
or U2597 (N_2597,In_1489,In_1776);
or U2598 (N_2598,In_443,In_3661);
nand U2599 (N_2599,In_3659,In_721);
and U2600 (N_2600,In_3748,In_3773);
nand U2601 (N_2601,In_893,In_583);
or U2602 (N_2602,In_4079,In_1384);
xor U2603 (N_2603,In_2313,In_2716);
xor U2604 (N_2604,In_4889,In_3009);
nor U2605 (N_2605,In_481,In_3756);
and U2606 (N_2606,In_3093,In_3872);
or U2607 (N_2607,In_4681,In_2230);
or U2608 (N_2608,In_327,In_4981);
nor U2609 (N_2609,In_1191,In_2382);
or U2610 (N_2610,In_4549,In_4771);
nor U2611 (N_2611,In_2756,In_3630);
xor U2612 (N_2612,In_1610,In_4018);
nand U2613 (N_2613,In_2018,In_2306);
and U2614 (N_2614,In_3675,In_875);
or U2615 (N_2615,In_3433,In_4742);
nand U2616 (N_2616,In_4371,In_4031);
nor U2617 (N_2617,In_4590,In_1081);
nand U2618 (N_2618,In_955,In_3260);
or U2619 (N_2619,In_3289,In_986);
nor U2620 (N_2620,In_1947,In_435);
nand U2621 (N_2621,In_1429,In_1040);
nand U2622 (N_2622,In_3091,In_3256);
or U2623 (N_2623,In_105,In_2719);
nor U2624 (N_2624,In_3446,In_823);
nand U2625 (N_2625,In_3006,In_2082);
nand U2626 (N_2626,In_2635,In_2710);
and U2627 (N_2627,In_4802,In_904);
or U2628 (N_2628,In_1390,In_2499);
nand U2629 (N_2629,In_3321,In_3516);
nor U2630 (N_2630,In_2079,In_2479);
or U2631 (N_2631,In_3324,In_3515);
xnor U2632 (N_2632,In_1146,In_3653);
nand U2633 (N_2633,In_3053,In_625);
nor U2634 (N_2634,In_2293,In_3016);
or U2635 (N_2635,In_2923,In_1346);
nor U2636 (N_2636,In_248,In_2697);
or U2637 (N_2637,In_334,In_4597);
xnor U2638 (N_2638,In_2811,In_1826);
xnor U2639 (N_2639,In_4711,In_4807);
nand U2640 (N_2640,In_921,In_244);
xnor U2641 (N_2641,In_4706,In_1141);
and U2642 (N_2642,In_448,In_583);
nand U2643 (N_2643,In_1223,In_2553);
and U2644 (N_2644,In_2470,In_4851);
nand U2645 (N_2645,In_4915,In_1654);
and U2646 (N_2646,In_1357,In_1791);
and U2647 (N_2647,In_1127,In_1695);
xnor U2648 (N_2648,In_1385,In_4469);
nor U2649 (N_2649,In_2391,In_1760);
or U2650 (N_2650,In_2323,In_1763);
and U2651 (N_2651,In_1468,In_2304);
xor U2652 (N_2652,In_716,In_4581);
or U2653 (N_2653,In_963,In_694);
or U2654 (N_2654,In_78,In_249);
and U2655 (N_2655,In_2292,In_4083);
nor U2656 (N_2656,In_309,In_4289);
nand U2657 (N_2657,In_4218,In_3587);
xnor U2658 (N_2658,In_912,In_2801);
and U2659 (N_2659,In_4514,In_3964);
nand U2660 (N_2660,In_3711,In_4688);
or U2661 (N_2661,In_3284,In_420);
nand U2662 (N_2662,In_1523,In_3968);
nand U2663 (N_2663,In_909,In_2207);
nor U2664 (N_2664,In_4391,In_1006);
and U2665 (N_2665,In_776,In_3595);
xnor U2666 (N_2666,In_2493,In_3910);
and U2667 (N_2667,In_1867,In_4523);
nand U2668 (N_2668,In_4409,In_1583);
nor U2669 (N_2669,In_3701,In_2446);
or U2670 (N_2670,In_87,In_1701);
or U2671 (N_2671,In_4545,In_2851);
and U2672 (N_2672,In_2079,In_2413);
and U2673 (N_2673,In_4762,In_4026);
xor U2674 (N_2674,In_1042,In_3237);
nand U2675 (N_2675,In_2552,In_2977);
xnor U2676 (N_2676,In_2145,In_1236);
or U2677 (N_2677,In_4026,In_2330);
and U2678 (N_2678,In_2637,In_494);
nor U2679 (N_2679,In_354,In_1166);
nor U2680 (N_2680,In_4138,In_2304);
nor U2681 (N_2681,In_3491,In_700);
nor U2682 (N_2682,In_2798,In_2216);
xnor U2683 (N_2683,In_2795,In_1438);
nor U2684 (N_2684,In_331,In_3791);
and U2685 (N_2685,In_2557,In_1110);
or U2686 (N_2686,In_2337,In_1539);
xor U2687 (N_2687,In_498,In_3379);
nor U2688 (N_2688,In_215,In_3787);
or U2689 (N_2689,In_1583,In_1773);
xnor U2690 (N_2690,In_4993,In_3264);
or U2691 (N_2691,In_2204,In_2094);
xor U2692 (N_2692,In_3019,In_2075);
and U2693 (N_2693,In_2478,In_1105);
and U2694 (N_2694,In_4516,In_410);
nor U2695 (N_2695,In_548,In_299);
or U2696 (N_2696,In_110,In_3181);
or U2697 (N_2697,In_4292,In_3690);
and U2698 (N_2698,In_352,In_2914);
xor U2699 (N_2699,In_1531,In_482);
nor U2700 (N_2700,In_4474,In_3770);
or U2701 (N_2701,In_2409,In_116);
or U2702 (N_2702,In_621,In_3381);
xnor U2703 (N_2703,In_3415,In_4685);
nor U2704 (N_2704,In_4428,In_4946);
xnor U2705 (N_2705,In_3725,In_194);
and U2706 (N_2706,In_3898,In_3817);
or U2707 (N_2707,In_3329,In_2008);
xor U2708 (N_2708,In_4144,In_1878);
nand U2709 (N_2709,In_4253,In_3761);
xor U2710 (N_2710,In_1476,In_2232);
nand U2711 (N_2711,In_2365,In_1098);
or U2712 (N_2712,In_1481,In_1444);
and U2713 (N_2713,In_3076,In_929);
nor U2714 (N_2714,In_3612,In_890);
nand U2715 (N_2715,In_2299,In_1511);
nor U2716 (N_2716,In_3964,In_4033);
and U2717 (N_2717,In_4372,In_1814);
and U2718 (N_2718,In_4804,In_1967);
and U2719 (N_2719,In_1576,In_1312);
nor U2720 (N_2720,In_4338,In_3985);
xor U2721 (N_2721,In_2598,In_3199);
xnor U2722 (N_2722,In_2841,In_4361);
xnor U2723 (N_2723,In_591,In_3611);
nand U2724 (N_2724,In_2079,In_4166);
or U2725 (N_2725,In_407,In_3519);
nand U2726 (N_2726,In_3618,In_3532);
nand U2727 (N_2727,In_823,In_3690);
and U2728 (N_2728,In_124,In_975);
nand U2729 (N_2729,In_2986,In_1489);
and U2730 (N_2730,In_855,In_964);
nor U2731 (N_2731,In_2615,In_4459);
xor U2732 (N_2732,In_2943,In_4412);
nor U2733 (N_2733,In_2417,In_2226);
nand U2734 (N_2734,In_2102,In_2458);
xnor U2735 (N_2735,In_2373,In_4786);
nor U2736 (N_2736,In_2001,In_3421);
xor U2737 (N_2737,In_1786,In_3884);
and U2738 (N_2738,In_2095,In_2241);
nor U2739 (N_2739,In_4826,In_648);
and U2740 (N_2740,In_2588,In_1405);
nand U2741 (N_2741,In_118,In_1312);
xor U2742 (N_2742,In_3271,In_4125);
nor U2743 (N_2743,In_2885,In_2563);
nand U2744 (N_2744,In_1961,In_3844);
nor U2745 (N_2745,In_1091,In_4726);
nand U2746 (N_2746,In_2209,In_4511);
or U2747 (N_2747,In_503,In_40);
and U2748 (N_2748,In_189,In_4038);
and U2749 (N_2749,In_1312,In_3276);
nor U2750 (N_2750,In_2023,In_3721);
and U2751 (N_2751,In_3233,In_1791);
nand U2752 (N_2752,In_2515,In_3773);
nand U2753 (N_2753,In_1873,In_3377);
and U2754 (N_2754,In_1582,In_1240);
xnor U2755 (N_2755,In_1153,In_3045);
xor U2756 (N_2756,In_4190,In_2629);
nor U2757 (N_2757,In_3544,In_3759);
xnor U2758 (N_2758,In_1162,In_1518);
or U2759 (N_2759,In_320,In_137);
or U2760 (N_2760,In_2902,In_205);
and U2761 (N_2761,In_3594,In_4059);
nand U2762 (N_2762,In_3142,In_1227);
nor U2763 (N_2763,In_1688,In_3267);
nand U2764 (N_2764,In_953,In_4991);
and U2765 (N_2765,In_4370,In_3879);
or U2766 (N_2766,In_1951,In_4888);
nand U2767 (N_2767,In_56,In_791);
nand U2768 (N_2768,In_4877,In_98);
and U2769 (N_2769,In_2621,In_4728);
nand U2770 (N_2770,In_1639,In_2442);
nor U2771 (N_2771,In_1305,In_61);
nand U2772 (N_2772,In_4133,In_1393);
nor U2773 (N_2773,In_4012,In_3353);
and U2774 (N_2774,In_3202,In_2494);
or U2775 (N_2775,In_3512,In_2928);
nand U2776 (N_2776,In_2349,In_2709);
or U2777 (N_2777,In_2176,In_2458);
or U2778 (N_2778,In_113,In_803);
and U2779 (N_2779,In_2962,In_1545);
or U2780 (N_2780,In_920,In_4487);
nor U2781 (N_2781,In_3040,In_1309);
and U2782 (N_2782,In_1673,In_3941);
xor U2783 (N_2783,In_781,In_3614);
or U2784 (N_2784,In_2434,In_587);
and U2785 (N_2785,In_3609,In_2771);
nand U2786 (N_2786,In_1187,In_1751);
and U2787 (N_2787,In_3267,In_4053);
nand U2788 (N_2788,In_1837,In_4585);
nand U2789 (N_2789,In_4337,In_1138);
and U2790 (N_2790,In_2738,In_3120);
and U2791 (N_2791,In_1924,In_1304);
and U2792 (N_2792,In_1529,In_3248);
and U2793 (N_2793,In_3771,In_3674);
xor U2794 (N_2794,In_2524,In_473);
and U2795 (N_2795,In_1547,In_3334);
and U2796 (N_2796,In_1344,In_3021);
and U2797 (N_2797,In_2090,In_2307);
or U2798 (N_2798,In_497,In_2141);
and U2799 (N_2799,In_254,In_3289);
nand U2800 (N_2800,In_3557,In_227);
nor U2801 (N_2801,In_3794,In_1877);
and U2802 (N_2802,In_160,In_641);
nor U2803 (N_2803,In_4023,In_4167);
and U2804 (N_2804,In_1001,In_3579);
and U2805 (N_2805,In_4519,In_2675);
or U2806 (N_2806,In_1769,In_1415);
nand U2807 (N_2807,In_2060,In_873);
xnor U2808 (N_2808,In_1880,In_4676);
nand U2809 (N_2809,In_3568,In_1102);
or U2810 (N_2810,In_4938,In_1366);
nor U2811 (N_2811,In_3612,In_3140);
xor U2812 (N_2812,In_1317,In_2496);
nor U2813 (N_2813,In_3375,In_2429);
and U2814 (N_2814,In_511,In_2307);
xnor U2815 (N_2815,In_3001,In_443);
or U2816 (N_2816,In_72,In_3146);
and U2817 (N_2817,In_2455,In_2110);
nand U2818 (N_2818,In_2920,In_4048);
nor U2819 (N_2819,In_1516,In_2265);
xor U2820 (N_2820,In_3919,In_3468);
nand U2821 (N_2821,In_3854,In_3136);
xor U2822 (N_2822,In_4482,In_555);
nand U2823 (N_2823,In_2263,In_4611);
or U2824 (N_2824,In_4547,In_4878);
nor U2825 (N_2825,In_4155,In_3184);
and U2826 (N_2826,In_2433,In_4470);
xnor U2827 (N_2827,In_4388,In_2884);
or U2828 (N_2828,In_2934,In_3934);
and U2829 (N_2829,In_3341,In_1222);
or U2830 (N_2830,In_4436,In_4100);
and U2831 (N_2831,In_3689,In_2942);
nor U2832 (N_2832,In_993,In_2203);
xor U2833 (N_2833,In_3606,In_1072);
nor U2834 (N_2834,In_3236,In_3194);
nand U2835 (N_2835,In_4649,In_4772);
nor U2836 (N_2836,In_2213,In_3575);
nand U2837 (N_2837,In_3699,In_2625);
nor U2838 (N_2838,In_260,In_4814);
nand U2839 (N_2839,In_1634,In_3872);
nor U2840 (N_2840,In_3051,In_4991);
xor U2841 (N_2841,In_982,In_795);
nand U2842 (N_2842,In_1526,In_2329);
nand U2843 (N_2843,In_3962,In_4939);
xor U2844 (N_2844,In_3052,In_1656);
or U2845 (N_2845,In_486,In_4625);
nor U2846 (N_2846,In_39,In_4552);
and U2847 (N_2847,In_834,In_4026);
nand U2848 (N_2848,In_3594,In_4693);
nand U2849 (N_2849,In_4598,In_4731);
nor U2850 (N_2850,In_1239,In_2749);
nor U2851 (N_2851,In_4198,In_3876);
xnor U2852 (N_2852,In_2182,In_4789);
nor U2853 (N_2853,In_2891,In_4874);
and U2854 (N_2854,In_299,In_1130);
and U2855 (N_2855,In_3306,In_1170);
nand U2856 (N_2856,In_3993,In_262);
and U2857 (N_2857,In_1187,In_3506);
xor U2858 (N_2858,In_2186,In_903);
or U2859 (N_2859,In_4129,In_512);
nand U2860 (N_2860,In_2310,In_2783);
or U2861 (N_2861,In_2239,In_1773);
nor U2862 (N_2862,In_3599,In_4671);
and U2863 (N_2863,In_2640,In_4146);
or U2864 (N_2864,In_3222,In_278);
or U2865 (N_2865,In_1879,In_4132);
nand U2866 (N_2866,In_2551,In_2817);
nand U2867 (N_2867,In_939,In_2901);
xnor U2868 (N_2868,In_4073,In_1224);
xnor U2869 (N_2869,In_3379,In_3855);
or U2870 (N_2870,In_4889,In_1667);
nand U2871 (N_2871,In_2094,In_3102);
or U2872 (N_2872,In_1172,In_3684);
or U2873 (N_2873,In_3173,In_2311);
nand U2874 (N_2874,In_4754,In_238);
and U2875 (N_2875,In_2906,In_2448);
nand U2876 (N_2876,In_2530,In_2727);
xnor U2877 (N_2877,In_574,In_657);
xor U2878 (N_2878,In_4520,In_949);
or U2879 (N_2879,In_855,In_1425);
and U2880 (N_2880,In_1217,In_1121);
or U2881 (N_2881,In_641,In_2025);
or U2882 (N_2882,In_2444,In_4264);
xor U2883 (N_2883,In_1367,In_2008);
nand U2884 (N_2884,In_4528,In_3865);
nand U2885 (N_2885,In_420,In_2989);
or U2886 (N_2886,In_1624,In_1819);
nand U2887 (N_2887,In_2561,In_1055);
and U2888 (N_2888,In_2688,In_3039);
xnor U2889 (N_2889,In_296,In_3291);
nor U2890 (N_2890,In_948,In_3292);
and U2891 (N_2891,In_2208,In_4367);
and U2892 (N_2892,In_1323,In_409);
or U2893 (N_2893,In_1623,In_2098);
and U2894 (N_2894,In_2565,In_4661);
or U2895 (N_2895,In_4313,In_1605);
xor U2896 (N_2896,In_4989,In_1580);
or U2897 (N_2897,In_1017,In_4032);
nor U2898 (N_2898,In_1127,In_2720);
xor U2899 (N_2899,In_1,In_4770);
and U2900 (N_2900,In_1133,In_2658);
and U2901 (N_2901,In_626,In_1931);
or U2902 (N_2902,In_4166,In_290);
and U2903 (N_2903,In_2849,In_3191);
xor U2904 (N_2904,In_3227,In_1708);
xor U2905 (N_2905,In_3869,In_4399);
or U2906 (N_2906,In_590,In_3726);
xor U2907 (N_2907,In_2292,In_335);
xnor U2908 (N_2908,In_2085,In_3784);
nand U2909 (N_2909,In_1540,In_4863);
nor U2910 (N_2910,In_2326,In_3681);
and U2911 (N_2911,In_1128,In_4221);
nand U2912 (N_2912,In_704,In_512);
nand U2913 (N_2913,In_26,In_1241);
or U2914 (N_2914,In_1831,In_2070);
nor U2915 (N_2915,In_384,In_658);
or U2916 (N_2916,In_4973,In_4645);
nor U2917 (N_2917,In_542,In_4185);
nand U2918 (N_2918,In_211,In_1381);
xor U2919 (N_2919,In_801,In_3109);
xnor U2920 (N_2920,In_380,In_2855);
and U2921 (N_2921,In_4044,In_4701);
and U2922 (N_2922,In_2850,In_4633);
or U2923 (N_2923,In_2028,In_3034);
nand U2924 (N_2924,In_92,In_4099);
nor U2925 (N_2925,In_3944,In_4325);
and U2926 (N_2926,In_598,In_2255);
xnor U2927 (N_2927,In_4455,In_4162);
nand U2928 (N_2928,In_4049,In_915);
xnor U2929 (N_2929,In_772,In_4845);
or U2930 (N_2930,In_2750,In_710);
or U2931 (N_2931,In_237,In_944);
xnor U2932 (N_2932,In_2109,In_3487);
xor U2933 (N_2933,In_3389,In_963);
xor U2934 (N_2934,In_199,In_1450);
nand U2935 (N_2935,In_2730,In_1606);
xor U2936 (N_2936,In_2609,In_3277);
and U2937 (N_2937,In_641,In_3935);
or U2938 (N_2938,In_864,In_3300);
nor U2939 (N_2939,In_3317,In_3816);
nand U2940 (N_2940,In_2186,In_1548);
nand U2941 (N_2941,In_2007,In_3843);
xor U2942 (N_2942,In_4177,In_2752);
or U2943 (N_2943,In_1566,In_4649);
nor U2944 (N_2944,In_2855,In_987);
nor U2945 (N_2945,In_9,In_4464);
and U2946 (N_2946,In_1116,In_3136);
xor U2947 (N_2947,In_2227,In_2134);
or U2948 (N_2948,In_3427,In_2230);
and U2949 (N_2949,In_2907,In_2783);
nor U2950 (N_2950,In_2747,In_3065);
xor U2951 (N_2951,In_1879,In_2426);
nand U2952 (N_2952,In_1610,In_2413);
xnor U2953 (N_2953,In_4285,In_3283);
nor U2954 (N_2954,In_3506,In_1464);
nor U2955 (N_2955,In_696,In_2920);
xor U2956 (N_2956,In_4346,In_2832);
nor U2957 (N_2957,In_3911,In_4203);
xor U2958 (N_2958,In_47,In_1663);
nor U2959 (N_2959,In_246,In_354);
nand U2960 (N_2960,In_3476,In_2851);
or U2961 (N_2961,In_4314,In_580);
nor U2962 (N_2962,In_4677,In_119);
and U2963 (N_2963,In_2012,In_3315);
and U2964 (N_2964,In_599,In_3177);
nor U2965 (N_2965,In_3235,In_504);
or U2966 (N_2966,In_707,In_4561);
xor U2967 (N_2967,In_3318,In_4576);
nor U2968 (N_2968,In_40,In_2924);
xor U2969 (N_2969,In_4618,In_2996);
or U2970 (N_2970,In_1534,In_1078);
nand U2971 (N_2971,In_1269,In_152);
xor U2972 (N_2972,In_2719,In_4939);
xnor U2973 (N_2973,In_1083,In_482);
nor U2974 (N_2974,In_4683,In_527);
nand U2975 (N_2975,In_2871,In_2015);
nand U2976 (N_2976,In_4752,In_3445);
or U2977 (N_2977,In_4573,In_4131);
or U2978 (N_2978,In_3761,In_714);
nor U2979 (N_2979,In_25,In_3030);
or U2980 (N_2980,In_1759,In_4487);
nand U2981 (N_2981,In_2989,In_1907);
nand U2982 (N_2982,In_3366,In_674);
nor U2983 (N_2983,In_4654,In_4111);
nor U2984 (N_2984,In_4926,In_3146);
xor U2985 (N_2985,In_3666,In_4438);
nand U2986 (N_2986,In_2938,In_660);
nor U2987 (N_2987,In_1639,In_2731);
or U2988 (N_2988,In_4250,In_4599);
xnor U2989 (N_2989,In_2081,In_4729);
and U2990 (N_2990,In_4229,In_2126);
or U2991 (N_2991,In_1013,In_2733);
or U2992 (N_2992,In_3753,In_789);
xor U2993 (N_2993,In_1053,In_2192);
and U2994 (N_2994,In_531,In_133);
nand U2995 (N_2995,In_3578,In_4184);
nor U2996 (N_2996,In_1392,In_2801);
nand U2997 (N_2997,In_3552,In_2297);
or U2998 (N_2998,In_3075,In_1575);
nor U2999 (N_2999,In_304,In_2660);
xor U3000 (N_3000,In_2253,In_1180);
or U3001 (N_3001,In_2918,In_1185);
xnor U3002 (N_3002,In_2831,In_3495);
and U3003 (N_3003,In_4128,In_355);
nand U3004 (N_3004,In_4254,In_2715);
and U3005 (N_3005,In_3826,In_3134);
nand U3006 (N_3006,In_351,In_4413);
xor U3007 (N_3007,In_4309,In_2144);
and U3008 (N_3008,In_3382,In_2421);
or U3009 (N_3009,In_1057,In_2281);
and U3010 (N_3010,In_647,In_82);
and U3011 (N_3011,In_96,In_2030);
xnor U3012 (N_3012,In_685,In_2479);
or U3013 (N_3013,In_4516,In_4149);
nand U3014 (N_3014,In_1209,In_3689);
nand U3015 (N_3015,In_1268,In_3287);
xor U3016 (N_3016,In_4807,In_2448);
xnor U3017 (N_3017,In_4317,In_3389);
xnor U3018 (N_3018,In_746,In_4549);
xnor U3019 (N_3019,In_34,In_4130);
and U3020 (N_3020,In_2658,In_1095);
or U3021 (N_3021,In_92,In_832);
and U3022 (N_3022,In_3025,In_405);
or U3023 (N_3023,In_2069,In_2941);
xor U3024 (N_3024,In_3614,In_484);
and U3025 (N_3025,In_644,In_660);
or U3026 (N_3026,In_1684,In_652);
xnor U3027 (N_3027,In_4148,In_1172);
nand U3028 (N_3028,In_1964,In_2144);
or U3029 (N_3029,In_245,In_4921);
xnor U3030 (N_3030,In_1610,In_2227);
nor U3031 (N_3031,In_645,In_4485);
nor U3032 (N_3032,In_458,In_365);
or U3033 (N_3033,In_2010,In_598);
or U3034 (N_3034,In_954,In_156);
or U3035 (N_3035,In_3974,In_297);
or U3036 (N_3036,In_1766,In_4537);
nor U3037 (N_3037,In_1376,In_1667);
xnor U3038 (N_3038,In_3808,In_3860);
nand U3039 (N_3039,In_772,In_259);
or U3040 (N_3040,In_1179,In_1869);
or U3041 (N_3041,In_3402,In_3335);
nand U3042 (N_3042,In_3738,In_4321);
and U3043 (N_3043,In_1845,In_309);
or U3044 (N_3044,In_309,In_4192);
and U3045 (N_3045,In_1924,In_4720);
nor U3046 (N_3046,In_2451,In_3695);
nor U3047 (N_3047,In_529,In_1327);
or U3048 (N_3048,In_4697,In_2316);
and U3049 (N_3049,In_986,In_3269);
nand U3050 (N_3050,In_2139,In_1822);
nand U3051 (N_3051,In_1620,In_4346);
nor U3052 (N_3052,In_3527,In_1241);
and U3053 (N_3053,In_391,In_1284);
nor U3054 (N_3054,In_3604,In_2925);
or U3055 (N_3055,In_4524,In_4441);
and U3056 (N_3056,In_4165,In_2309);
and U3057 (N_3057,In_1159,In_2897);
and U3058 (N_3058,In_1730,In_2114);
nor U3059 (N_3059,In_4255,In_244);
nand U3060 (N_3060,In_3704,In_1430);
xnor U3061 (N_3061,In_2610,In_670);
or U3062 (N_3062,In_2472,In_2371);
nand U3063 (N_3063,In_629,In_886);
nor U3064 (N_3064,In_3024,In_264);
nand U3065 (N_3065,In_209,In_4740);
or U3066 (N_3066,In_2543,In_1739);
xor U3067 (N_3067,In_4013,In_4276);
xnor U3068 (N_3068,In_1217,In_1167);
nand U3069 (N_3069,In_607,In_2052);
nor U3070 (N_3070,In_2535,In_1661);
nor U3071 (N_3071,In_3682,In_476);
and U3072 (N_3072,In_3084,In_4691);
nand U3073 (N_3073,In_1399,In_4654);
xor U3074 (N_3074,In_656,In_4787);
nor U3075 (N_3075,In_2916,In_3817);
and U3076 (N_3076,In_2817,In_634);
xor U3077 (N_3077,In_2013,In_2427);
and U3078 (N_3078,In_3830,In_1582);
xnor U3079 (N_3079,In_1861,In_1462);
and U3080 (N_3080,In_693,In_1);
nor U3081 (N_3081,In_4410,In_2662);
and U3082 (N_3082,In_4855,In_80);
xor U3083 (N_3083,In_588,In_2198);
nor U3084 (N_3084,In_4937,In_2699);
and U3085 (N_3085,In_1342,In_1909);
nor U3086 (N_3086,In_1990,In_3552);
and U3087 (N_3087,In_2128,In_4245);
and U3088 (N_3088,In_1950,In_3520);
nor U3089 (N_3089,In_4406,In_915);
xor U3090 (N_3090,In_3376,In_3163);
or U3091 (N_3091,In_4865,In_4630);
or U3092 (N_3092,In_2662,In_1776);
or U3093 (N_3093,In_3590,In_597);
nor U3094 (N_3094,In_4442,In_2302);
xnor U3095 (N_3095,In_4257,In_2852);
nand U3096 (N_3096,In_776,In_1130);
xor U3097 (N_3097,In_1659,In_4094);
xor U3098 (N_3098,In_4004,In_214);
and U3099 (N_3099,In_1040,In_3672);
xor U3100 (N_3100,In_1931,In_223);
nand U3101 (N_3101,In_3696,In_421);
xor U3102 (N_3102,In_4165,In_556);
nand U3103 (N_3103,In_769,In_1460);
or U3104 (N_3104,In_312,In_3679);
xnor U3105 (N_3105,In_1574,In_1825);
and U3106 (N_3106,In_4204,In_1710);
or U3107 (N_3107,In_148,In_3066);
nand U3108 (N_3108,In_1996,In_211);
nand U3109 (N_3109,In_4879,In_747);
xor U3110 (N_3110,In_4365,In_1101);
and U3111 (N_3111,In_4256,In_3576);
and U3112 (N_3112,In_1159,In_3755);
nand U3113 (N_3113,In_4130,In_1068);
nor U3114 (N_3114,In_3347,In_4182);
xnor U3115 (N_3115,In_1967,In_4950);
nand U3116 (N_3116,In_3405,In_2609);
xnor U3117 (N_3117,In_2483,In_547);
and U3118 (N_3118,In_926,In_1993);
nand U3119 (N_3119,In_1137,In_4533);
nor U3120 (N_3120,In_3720,In_1904);
nand U3121 (N_3121,In_1997,In_4670);
xor U3122 (N_3122,In_3964,In_298);
and U3123 (N_3123,In_980,In_1570);
nand U3124 (N_3124,In_2394,In_547);
and U3125 (N_3125,In_2200,In_4821);
nor U3126 (N_3126,In_2555,In_3388);
xnor U3127 (N_3127,In_1199,In_4949);
or U3128 (N_3128,In_885,In_2029);
nor U3129 (N_3129,In_4494,In_3295);
and U3130 (N_3130,In_2758,In_396);
and U3131 (N_3131,In_1207,In_634);
nand U3132 (N_3132,In_4247,In_2927);
xor U3133 (N_3133,In_359,In_809);
nand U3134 (N_3134,In_3939,In_3217);
xnor U3135 (N_3135,In_2157,In_4133);
and U3136 (N_3136,In_708,In_732);
and U3137 (N_3137,In_429,In_3202);
and U3138 (N_3138,In_3264,In_2226);
and U3139 (N_3139,In_3434,In_2264);
xor U3140 (N_3140,In_15,In_2541);
nand U3141 (N_3141,In_2374,In_2842);
xnor U3142 (N_3142,In_2131,In_3676);
nor U3143 (N_3143,In_1316,In_3879);
nand U3144 (N_3144,In_3813,In_3280);
nor U3145 (N_3145,In_488,In_1375);
xor U3146 (N_3146,In_2672,In_3269);
nor U3147 (N_3147,In_4536,In_3276);
or U3148 (N_3148,In_4611,In_4661);
nor U3149 (N_3149,In_3816,In_2582);
nor U3150 (N_3150,In_1452,In_3433);
or U3151 (N_3151,In_3614,In_2760);
and U3152 (N_3152,In_3035,In_539);
and U3153 (N_3153,In_1990,In_3074);
nor U3154 (N_3154,In_746,In_3550);
and U3155 (N_3155,In_696,In_2880);
and U3156 (N_3156,In_3769,In_2887);
xnor U3157 (N_3157,In_31,In_2944);
xor U3158 (N_3158,In_4444,In_1596);
and U3159 (N_3159,In_4652,In_1274);
nor U3160 (N_3160,In_2656,In_2998);
or U3161 (N_3161,In_3901,In_2397);
xor U3162 (N_3162,In_4491,In_3026);
nor U3163 (N_3163,In_3676,In_4010);
xnor U3164 (N_3164,In_4053,In_3762);
xnor U3165 (N_3165,In_2153,In_574);
nand U3166 (N_3166,In_3737,In_267);
xnor U3167 (N_3167,In_4509,In_2213);
nor U3168 (N_3168,In_115,In_394);
nor U3169 (N_3169,In_598,In_3419);
xor U3170 (N_3170,In_3965,In_2231);
and U3171 (N_3171,In_4144,In_4864);
nor U3172 (N_3172,In_3456,In_2705);
nand U3173 (N_3173,In_2988,In_413);
or U3174 (N_3174,In_3571,In_4424);
xor U3175 (N_3175,In_947,In_104);
or U3176 (N_3176,In_2941,In_674);
nor U3177 (N_3177,In_3561,In_4378);
xnor U3178 (N_3178,In_1753,In_1206);
nand U3179 (N_3179,In_3846,In_3532);
nand U3180 (N_3180,In_1646,In_2100);
nor U3181 (N_3181,In_2526,In_1676);
xor U3182 (N_3182,In_3076,In_670);
nand U3183 (N_3183,In_4732,In_1307);
nor U3184 (N_3184,In_3072,In_4812);
or U3185 (N_3185,In_1815,In_43);
nand U3186 (N_3186,In_3067,In_2515);
nand U3187 (N_3187,In_2611,In_3693);
nand U3188 (N_3188,In_113,In_2781);
nand U3189 (N_3189,In_1070,In_515);
xor U3190 (N_3190,In_1804,In_1151);
nand U3191 (N_3191,In_4969,In_4274);
and U3192 (N_3192,In_350,In_2418);
nor U3193 (N_3193,In_4531,In_1941);
nor U3194 (N_3194,In_2963,In_3187);
xor U3195 (N_3195,In_1987,In_3756);
xnor U3196 (N_3196,In_594,In_4599);
or U3197 (N_3197,In_1229,In_2609);
xor U3198 (N_3198,In_2917,In_989);
nor U3199 (N_3199,In_1550,In_460);
xnor U3200 (N_3200,In_4034,In_1894);
nand U3201 (N_3201,In_2398,In_4727);
and U3202 (N_3202,In_1161,In_1535);
xnor U3203 (N_3203,In_2844,In_3464);
nand U3204 (N_3204,In_1314,In_1272);
nor U3205 (N_3205,In_1794,In_4478);
nand U3206 (N_3206,In_2747,In_3040);
nand U3207 (N_3207,In_2477,In_853);
nand U3208 (N_3208,In_4620,In_3226);
and U3209 (N_3209,In_791,In_4789);
nand U3210 (N_3210,In_2468,In_4191);
nor U3211 (N_3211,In_2603,In_3569);
xor U3212 (N_3212,In_455,In_6);
nor U3213 (N_3213,In_3782,In_3125);
nand U3214 (N_3214,In_2773,In_2671);
nor U3215 (N_3215,In_722,In_554);
nor U3216 (N_3216,In_3131,In_1732);
xor U3217 (N_3217,In_3056,In_59);
xnor U3218 (N_3218,In_129,In_3117);
xor U3219 (N_3219,In_1963,In_3635);
or U3220 (N_3220,In_2929,In_1443);
nor U3221 (N_3221,In_3476,In_437);
xor U3222 (N_3222,In_2071,In_232);
xnor U3223 (N_3223,In_265,In_1805);
and U3224 (N_3224,In_2034,In_3247);
nand U3225 (N_3225,In_2883,In_1643);
nor U3226 (N_3226,In_3754,In_4117);
and U3227 (N_3227,In_2014,In_3501);
nor U3228 (N_3228,In_2848,In_4611);
xnor U3229 (N_3229,In_4216,In_2954);
and U3230 (N_3230,In_1216,In_3195);
xor U3231 (N_3231,In_2112,In_343);
or U3232 (N_3232,In_2108,In_3448);
or U3233 (N_3233,In_290,In_1805);
nand U3234 (N_3234,In_4481,In_758);
nand U3235 (N_3235,In_4359,In_1621);
and U3236 (N_3236,In_4368,In_1873);
or U3237 (N_3237,In_4872,In_1565);
nand U3238 (N_3238,In_1452,In_4544);
or U3239 (N_3239,In_2934,In_4213);
and U3240 (N_3240,In_4957,In_2898);
nor U3241 (N_3241,In_3607,In_2215);
nor U3242 (N_3242,In_4939,In_2653);
or U3243 (N_3243,In_3047,In_30);
nor U3244 (N_3244,In_4188,In_598);
xor U3245 (N_3245,In_4077,In_4994);
or U3246 (N_3246,In_640,In_4837);
or U3247 (N_3247,In_3853,In_61);
and U3248 (N_3248,In_4535,In_229);
xor U3249 (N_3249,In_592,In_2392);
nand U3250 (N_3250,In_4973,In_1917);
nor U3251 (N_3251,In_3655,In_680);
nor U3252 (N_3252,In_4968,In_4563);
or U3253 (N_3253,In_3645,In_2236);
xnor U3254 (N_3254,In_1345,In_4897);
nor U3255 (N_3255,In_303,In_598);
nand U3256 (N_3256,In_4313,In_142);
and U3257 (N_3257,In_3416,In_2299);
xnor U3258 (N_3258,In_4550,In_2561);
nor U3259 (N_3259,In_1245,In_1511);
xnor U3260 (N_3260,In_651,In_4364);
and U3261 (N_3261,In_3321,In_4460);
and U3262 (N_3262,In_855,In_1012);
xor U3263 (N_3263,In_2145,In_20);
or U3264 (N_3264,In_238,In_4630);
and U3265 (N_3265,In_1731,In_1171);
and U3266 (N_3266,In_3176,In_450);
nand U3267 (N_3267,In_1593,In_1381);
or U3268 (N_3268,In_4448,In_2760);
xnor U3269 (N_3269,In_4304,In_4448);
and U3270 (N_3270,In_3883,In_3779);
nor U3271 (N_3271,In_925,In_3760);
and U3272 (N_3272,In_2695,In_3910);
xnor U3273 (N_3273,In_2278,In_610);
nand U3274 (N_3274,In_2294,In_2231);
nor U3275 (N_3275,In_708,In_3658);
and U3276 (N_3276,In_2306,In_1913);
nand U3277 (N_3277,In_2282,In_4146);
nand U3278 (N_3278,In_3184,In_2841);
xnor U3279 (N_3279,In_732,In_1045);
xor U3280 (N_3280,In_680,In_2958);
nor U3281 (N_3281,In_279,In_320);
nand U3282 (N_3282,In_3128,In_1378);
and U3283 (N_3283,In_799,In_968);
or U3284 (N_3284,In_1133,In_4877);
xnor U3285 (N_3285,In_1317,In_1006);
xor U3286 (N_3286,In_622,In_26);
nor U3287 (N_3287,In_2432,In_4832);
or U3288 (N_3288,In_1216,In_2143);
xnor U3289 (N_3289,In_2531,In_2292);
and U3290 (N_3290,In_389,In_3273);
nor U3291 (N_3291,In_817,In_3547);
xnor U3292 (N_3292,In_3722,In_4551);
and U3293 (N_3293,In_4485,In_2606);
nor U3294 (N_3294,In_3557,In_4809);
or U3295 (N_3295,In_4243,In_1478);
or U3296 (N_3296,In_4089,In_1104);
and U3297 (N_3297,In_1476,In_541);
and U3298 (N_3298,In_343,In_3678);
xnor U3299 (N_3299,In_2648,In_2728);
or U3300 (N_3300,In_3492,In_4748);
nand U3301 (N_3301,In_1133,In_4969);
nor U3302 (N_3302,In_3616,In_1248);
nor U3303 (N_3303,In_4176,In_3562);
xor U3304 (N_3304,In_1938,In_982);
nor U3305 (N_3305,In_3909,In_3960);
xor U3306 (N_3306,In_2329,In_747);
nand U3307 (N_3307,In_2011,In_1952);
xor U3308 (N_3308,In_3643,In_3511);
nor U3309 (N_3309,In_3540,In_846);
xor U3310 (N_3310,In_3662,In_59);
xor U3311 (N_3311,In_3229,In_210);
or U3312 (N_3312,In_1206,In_3943);
nor U3313 (N_3313,In_2097,In_2639);
nor U3314 (N_3314,In_92,In_61);
nand U3315 (N_3315,In_4493,In_2416);
nor U3316 (N_3316,In_4216,In_231);
and U3317 (N_3317,In_37,In_2395);
nor U3318 (N_3318,In_4794,In_953);
and U3319 (N_3319,In_1954,In_2249);
and U3320 (N_3320,In_1493,In_663);
nor U3321 (N_3321,In_2973,In_1243);
or U3322 (N_3322,In_2411,In_2636);
and U3323 (N_3323,In_2716,In_3462);
nor U3324 (N_3324,In_252,In_1758);
and U3325 (N_3325,In_1198,In_4896);
xor U3326 (N_3326,In_1830,In_549);
nor U3327 (N_3327,In_4818,In_4869);
or U3328 (N_3328,In_4040,In_44);
or U3329 (N_3329,In_3424,In_4925);
or U3330 (N_3330,In_1176,In_2674);
and U3331 (N_3331,In_2812,In_211);
nor U3332 (N_3332,In_294,In_3533);
nor U3333 (N_3333,In_4122,In_4918);
nor U3334 (N_3334,In_2083,In_1631);
xor U3335 (N_3335,In_1545,In_4720);
nor U3336 (N_3336,In_3197,In_697);
and U3337 (N_3337,In_3494,In_4014);
and U3338 (N_3338,In_3331,In_1636);
nand U3339 (N_3339,In_1119,In_1207);
nor U3340 (N_3340,In_1203,In_287);
nor U3341 (N_3341,In_763,In_3967);
or U3342 (N_3342,In_1313,In_345);
nor U3343 (N_3343,In_1790,In_4457);
nor U3344 (N_3344,In_1105,In_3048);
nor U3345 (N_3345,In_2230,In_1777);
and U3346 (N_3346,In_853,In_4081);
nor U3347 (N_3347,In_1468,In_2890);
xor U3348 (N_3348,In_4817,In_603);
and U3349 (N_3349,In_3460,In_1202);
and U3350 (N_3350,In_87,In_2115);
xnor U3351 (N_3351,In_1457,In_4861);
nor U3352 (N_3352,In_1327,In_693);
xor U3353 (N_3353,In_2735,In_1003);
xor U3354 (N_3354,In_2244,In_775);
or U3355 (N_3355,In_1100,In_4721);
and U3356 (N_3356,In_4782,In_924);
xnor U3357 (N_3357,In_1562,In_1351);
and U3358 (N_3358,In_3112,In_1095);
nand U3359 (N_3359,In_2455,In_704);
nand U3360 (N_3360,In_2648,In_1571);
nor U3361 (N_3361,In_4268,In_1558);
xnor U3362 (N_3362,In_3820,In_4500);
nand U3363 (N_3363,In_1746,In_1597);
nor U3364 (N_3364,In_3966,In_3532);
nand U3365 (N_3365,In_3084,In_1599);
xnor U3366 (N_3366,In_1203,In_1311);
xor U3367 (N_3367,In_2671,In_3660);
xnor U3368 (N_3368,In_3706,In_175);
or U3369 (N_3369,In_4544,In_3401);
xor U3370 (N_3370,In_336,In_2969);
nor U3371 (N_3371,In_864,In_726);
nand U3372 (N_3372,In_1067,In_3615);
xor U3373 (N_3373,In_1864,In_4349);
and U3374 (N_3374,In_2483,In_537);
xor U3375 (N_3375,In_2773,In_3738);
nor U3376 (N_3376,In_525,In_2694);
nand U3377 (N_3377,In_1828,In_4547);
xor U3378 (N_3378,In_2795,In_4218);
or U3379 (N_3379,In_90,In_3338);
or U3380 (N_3380,In_3627,In_759);
and U3381 (N_3381,In_3620,In_3978);
and U3382 (N_3382,In_1350,In_2403);
nor U3383 (N_3383,In_1500,In_1505);
or U3384 (N_3384,In_4982,In_2787);
xor U3385 (N_3385,In_4398,In_4232);
and U3386 (N_3386,In_2376,In_1355);
nor U3387 (N_3387,In_2579,In_291);
nor U3388 (N_3388,In_1447,In_1015);
nand U3389 (N_3389,In_1341,In_1206);
nor U3390 (N_3390,In_3,In_3914);
nand U3391 (N_3391,In_4306,In_3396);
and U3392 (N_3392,In_3585,In_2398);
xnor U3393 (N_3393,In_398,In_63);
nor U3394 (N_3394,In_1516,In_3731);
xnor U3395 (N_3395,In_4196,In_547);
nand U3396 (N_3396,In_4809,In_1042);
nor U3397 (N_3397,In_4727,In_986);
nand U3398 (N_3398,In_2341,In_4033);
nand U3399 (N_3399,In_1623,In_728);
nand U3400 (N_3400,In_1241,In_2779);
xnor U3401 (N_3401,In_3590,In_2371);
nand U3402 (N_3402,In_3396,In_1585);
or U3403 (N_3403,In_1956,In_1745);
nand U3404 (N_3404,In_1863,In_3660);
or U3405 (N_3405,In_3503,In_3487);
nor U3406 (N_3406,In_3101,In_4929);
nand U3407 (N_3407,In_3087,In_1627);
nand U3408 (N_3408,In_2212,In_1138);
nand U3409 (N_3409,In_1990,In_3320);
or U3410 (N_3410,In_1342,In_2366);
nor U3411 (N_3411,In_1165,In_2807);
nand U3412 (N_3412,In_1697,In_2126);
nand U3413 (N_3413,In_596,In_4838);
xnor U3414 (N_3414,In_1330,In_2290);
xor U3415 (N_3415,In_3751,In_512);
nand U3416 (N_3416,In_502,In_4912);
and U3417 (N_3417,In_4153,In_1598);
and U3418 (N_3418,In_4453,In_4602);
xor U3419 (N_3419,In_4651,In_159);
nand U3420 (N_3420,In_3218,In_4329);
and U3421 (N_3421,In_1008,In_1736);
or U3422 (N_3422,In_1812,In_2389);
and U3423 (N_3423,In_3815,In_4521);
and U3424 (N_3424,In_1662,In_1335);
xor U3425 (N_3425,In_4146,In_2731);
nand U3426 (N_3426,In_3189,In_4194);
and U3427 (N_3427,In_2889,In_764);
and U3428 (N_3428,In_329,In_4196);
xor U3429 (N_3429,In_522,In_958);
xnor U3430 (N_3430,In_3275,In_3286);
and U3431 (N_3431,In_4881,In_3654);
or U3432 (N_3432,In_4623,In_2357);
or U3433 (N_3433,In_4193,In_1052);
nand U3434 (N_3434,In_4033,In_4254);
or U3435 (N_3435,In_2725,In_2332);
and U3436 (N_3436,In_3256,In_2655);
nor U3437 (N_3437,In_2778,In_1452);
nor U3438 (N_3438,In_679,In_2993);
nand U3439 (N_3439,In_2567,In_280);
xnor U3440 (N_3440,In_3965,In_3409);
xnor U3441 (N_3441,In_3695,In_647);
xor U3442 (N_3442,In_4645,In_1078);
xor U3443 (N_3443,In_4587,In_2751);
and U3444 (N_3444,In_1597,In_2307);
xor U3445 (N_3445,In_4553,In_258);
nand U3446 (N_3446,In_4343,In_2417);
nand U3447 (N_3447,In_3485,In_2581);
and U3448 (N_3448,In_1583,In_137);
xor U3449 (N_3449,In_2330,In_538);
xnor U3450 (N_3450,In_4334,In_2732);
or U3451 (N_3451,In_4443,In_3281);
xnor U3452 (N_3452,In_3775,In_4200);
nand U3453 (N_3453,In_2972,In_2289);
and U3454 (N_3454,In_326,In_3480);
xnor U3455 (N_3455,In_1693,In_4280);
nand U3456 (N_3456,In_3570,In_2572);
or U3457 (N_3457,In_4622,In_793);
xor U3458 (N_3458,In_4779,In_667);
nor U3459 (N_3459,In_2557,In_2313);
or U3460 (N_3460,In_1478,In_4872);
and U3461 (N_3461,In_3284,In_1854);
or U3462 (N_3462,In_4653,In_493);
nand U3463 (N_3463,In_4058,In_643);
or U3464 (N_3464,In_1027,In_3101);
nor U3465 (N_3465,In_3117,In_2741);
and U3466 (N_3466,In_77,In_1722);
nor U3467 (N_3467,In_1683,In_1604);
nor U3468 (N_3468,In_765,In_3465);
xor U3469 (N_3469,In_2822,In_1432);
xnor U3470 (N_3470,In_829,In_1470);
nand U3471 (N_3471,In_3132,In_1484);
and U3472 (N_3472,In_2183,In_2942);
and U3473 (N_3473,In_177,In_2845);
nor U3474 (N_3474,In_3920,In_1547);
and U3475 (N_3475,In_4647,In_4366);
nor U3476 (N_3476,In_214,In_1414);
nor U3477 (N_3477,In_1085,In_1486);
nand U3478 (N_3478,In_2087,In_3092);
nand U3479 (N_3479,In_145,In_4983);
or U3480 (N_3480,In_4428,In_574);
or U3481 (N_3481,In_522,In_1546);
xnor U3482 (N_3482,In_3895,In_4730);
xor U3483 (N_3483,In_2244,In_4323);
xnor U3484 (N_3484,In_4318,In_1497);
nor U3485 (N_3485,In_1679,In_3554);
xnor U3486 (N_3486,In_4498,In_1015);
or U3487 (N_3487,In_4721,In_82);
xnor U3488 (N_3488,In_3796,In_226);
nor U3489 (N_3489,In_3220,In_2631);
xor U3490 (N_3490,In_2640,In_1667);
or U3491 (N_3491,In_3922,In_4850);
or U3492 (N_3492,In_2962,In_238);
nand U3493 (N_3493,In_3423,In_4914);
nor U3494 (N_3494,In_1709,In_4481);
nor U3495 (N_3495,In_4608,In_4892);
or U3496 (N_3496,In_1617,In_2966);
or U3497 (N_3497,In_1879,In_1493);
and U3498 (N_3498,In_4082,In_3068);
xor U3499 (N_3499,In_2439,In_1121);
xnor U3500 (N_3500,In_1744,In_3033);
and U3501 (N_3501,In_283,In_4306);
xnor U3502 (N_3502,In_2152,In_2255);
nand U3503 (N_3503,In_644,In_4413);
nand U3504 (N_3504,In_288,In_2439);
nor U3505 (N_3505,In_4212,In_3522);
xnor U3506 (N_3506,In_950,In_634);
and U3507 (N_3507,In_3002,In_3679);
and U3508 (N_3508,In_2308,In_4421);
or U3509 (N_3509,In_2306,In_3374);
or U3510 (N_3510,In_1672,In_236);
xnor U3511 (N_3511,In_1420,In_3185);
and U3512 (N_3512,In_872,In_2006);
and U3513 (N_3513,In_3206,In_2363);
nor U3514 (N_3514,In_858,In_2734);
xnor U3515 (N_3515,In_2268,In_3827);
nor U3516 (N_3516,In_4167,In_2061);
xnor U3517 (N_3517,In_4982,In_4069);
or U3518 (N_3518,In_1538,In_4112);
or U3519 (N_3519,In_1186,In_2488);
and U3520 (N_3520,In_4250,In_4029);
or U3521 (N_3521,In_708,In_2676);
nand U3522 (N_3522,In_4455,In_3941);
or U3523 (N_3523,In_2786,In_3548);
or U3524 (N_3524,In_3099,In_1844);
and U3525 (N_3525,In_2712,In_3195);
xor U3526 (N_3526,In_2866,In_360);
or U3527 (N_3527,In_4615,In_739);
nor U3528 (N_3528,In_2668,In_4963);
and U3529 (N_3529,In_4347,In_3288);
or U3530 (N_3530,In_1669,In_1789);
xor U3531 (N_3531,In_2729,In_4432);
nand U3532 (N_3532,In_4614,In_4061);
xnor U3533 (N_3533,In_2478,In_1601);
xor U3534 (N_3534,In_1814,In_1725);
nand U3535 (N_3535,In_1376,In_2185);
xnor U3536 (N_3536,In_1982,In_3846);
nand U3537 (N_3537,In_4045,In_3381);
nor U3538 (N_3538,In_369,In_1409);
xnor U3539 (N_3539,In_3597,In_1531);
xnor U3540 (N_3540,In_3160,In_2688);
nor U3541 (N_3541,In_3186,In_3);
xor U3542 (N_3542,In_2059,In_800);
and U3543 (N_3543,In_3144,In_3749);
xor U3544 (N_3544,In_3220,In_2288);
or U3545 (N_3545,In_561,In_493);
xor U3546 (N_3546,In_3963,In_1281);
xnor U3547 (N_3547,In_1579,In_2465);
nand U3548 (N_3548,In_3565,In_3402);
nand U3549 (N_3549,In_2408,In_4231);
xor U3550 (N_3550,In_4591,In_2951);
xnor U3551 (N_3551,In_1302,In_331);
nand U3552 (N_3552,In_3609,In_1338);
and U3553 (N_3553,In_3184,In_1820);
nand U3554 (N_3554,In_1547,In_119);
nor U3555 (N_3555,In_3617,In_2086);
nor U3556 (N_3556,In_3745,In_2122);
or U3557 (N_3557,In_2672,In_469);
xor U3558 (N_3558,In_2638,In_1071);
nor U3559 (N_3559,In_3070,In_4884);
or U3560 (N_3560,In_4300,In_3428);
nand U3561 (N_3561,In_4781,In_587);
nand U3562 (N_3562,In_2415,In_533);
and U3563 (N_3563,In_2800,In_4595);
nand U3564 (N_3564,In_2350,In_2463);
nor U3565 (N_3565,In_2561,In_1404);
and U3566 (N_3566,In_3616,In_2428);
nand U3567 (N_3567,In_1384,In_4210);
and U3568 (N_3568,In_1150,In_3723);
nand U3569 (N_3569,In_4431,In_3733);
nor U3570 (N_3570,In_3246,In_652);
nand U3571 (N_3571,In_3575,In_4315);
nand U3572 (N_3572,In_4350,In_2260);
nand U3573 (N_3573,In_3290,In_3308);
or U3574 (N_3574,In_3504,In_3010);
nor U3575 (N_3575,In_4131,In_1273);
xnor U3576 (N_3576,In_4446,In_2674);
or U3577 (N_3577,In_2925,In_71);
and U3578 (N_3578,In_1557,In_3549);
and U3579 (N_3579,In_2940,In_4417);
nand U3580 (N_3580,In_4539,In_3460);
and U3581 (N_3581,In_2759,In_3891);
xnor U3582 (N_3582,In_1188,In_3913);
or U3583 (N_3583,In_301,In_2745);
or U3584 (N_3584,In_3890,In_53);
xnor U3585 (N_3585,In_3090,In_1851);
xnor U3586 (N_3586,In_1797,In_1794);
and U3587 (N_3587,In_103,In_4448);
or U3588 (N_3588,In_1216,In_4155);
and U3589 (N_3589,In_3655,In_222);
xor U3590 (N_3590,In_3930,In_1816);
xnor U3591 (N_3591,In_462,In_1653);
nand U3592 (N_3592,In_4264,In_3604);
and U3593 (N_3593,In_4760,In_3482);
xnor U3594 (N_3594,In_527,In_4018);
nand U3595 (N_3595,In_4697,In_2212);
nand U3596 (N_3596,In_2682,In_2479);
or U3597 (N_3597,In_2523,In_3895);
or U3598 (N_3598,In_3515,In_1304);
nor U3599 (N_3599,In_2079,In_1553);
and U3600 (N_3600,In_2792,In_4981);
or U3601 (N_3601,In_2644,In_4875);
and U3602 (N_3602,In_997,In_3775);
or U3603 (N_3603,In_2060,In_1163);
nand U3604 (N_3604,In_3822,In_4091);
nand U3605 (N_3605,In_2108,In_1884);
nand U3606 (N_3606,In_1611,In_3414);
and U3607 (N_3607,In_4717,In_1518);
and U3608 (N_3608,In_482,In_1367);
or U3609 (N_3609,In_807,In_4779);
or U3610 (N_3610,In_1157,In_3613);
and U3611 (N_3611,In_3749,In_913);
xnor U3612 (N_3612,In_2952,In_4283);
nor U3613 (N_3613,In_1864,In_4564);
nand U3614 (N_3614,In_2220,In_4740);
and U3615 (N_3615,In_1125,In_4144);
nand U3616 (N_3616,In_2912,In_1361);
nor U3617 (N_3617,In_3940,In_945);
and U3618 (N_3618,In_1244,In_905);
nor U3619 (N_3619,In_2658,In_3640);
nor U3620 (N_3620,In_3472,In_4333);
or U3621 (N_3621,In_568,In_668);
nand U3622 (N_3622,In_1613,In_644);
and U3623 (N_3623,In_4774,In_4617);
xor U3624 (N_3624,In_139,In_3682);
xnor U3625 (N_3625,In_4816,In_3441);
or U3626 (N_3626,In_4668,In_2735);
nor U3627 (N_3627,In_1517,In_3886);
xor U3628 (N_3628,In_658,In_4544);
and U3629 (N_3629,In_4727,In_883);
nand U3630 (N_3630,In_4229,In_4759);
or U3631 (N_3631,In_657,In_665);
and U3632 (N_3632,In_4711,In_1539);
nor U3633 (N_3633,In_4084,In_1287);
xnor U3634 (N_3634,In_1218,In_3255);
nor U3635 (N_3635,In_2760,In_1972);
and U3636 (N_3636,In_4787,In_490);
and U3637 (N_3637,In_190,In_4699);
xnor U3638 (N_3638,In_1523,In_2360);
or U3639 (N_3639,In_4854,In_965);
nand U3640 (N_3640,In_2734,In_1225);
nor U3641 (N_3641,In_2048,In_2796);
xnor U3642 (N_3642,In_2159,In_231);
nor U3643 (N_3643,In_1395,In_87);
nand U3644 (N_3644,In_2408,In_3714);
nor U3645 (N_3645,In_3768,In_4344);
or U3646 (N_3646,In_776,In_1950);
and U3647 (N_3647,In_3889,In_1527);
nand U3648 (N_3648,In_1772,In_3381);
or U3649 (N_3649,In_4355,In_3603);
xor U3650 (N_3650,In_3095,In_3060);
and U3651 (N_3651,In_1999,In_2726);
and U3652 (N_3652,In_451,In_1296);
xor U3653 (N_3653,In_1894,In_2943);
nor U3654 (N_3654,In_1544,In_3789);
xor U3655 (N_3655,In_1548,In_2938);
or U3656 (N_3656,In_963,In_580);
or U3657 (N_3657,In_797,In_4227);
or U3658 (N_3658,In_432,In_4994);
xnor U3659 (N_3659,In_4536,In_1215);
nand U3660 (N_3660,In_1839,In_3997);
nor U3661 (N_3661,In_3186,In_2637);
nand U3662 (N_3662,In_845,In_2883);
xnor U3663 (N_3663,In_3221,In_4874);
or U3664 (N_3664,In_1725,In_4102);
nor U3665 (N_3665,In_904,In_713);
nor U3666 (N_3666,In_629,In_4622);
and U3667 (N_3667,In_2913,In_2648);
nor U3668 (N_3668,In_1585,In_1301);
nand U3669 (N_3669,In_2216,In_2555);
and U3670 (N_3670,In_931,In_453);
nor U3671 (N_3671,In_2317,In_3846);
nand U3672 (N_3672,In_1363,In_410);
and U3673 (N_3673,In_4860,In_3534);
xor U3674 (N_3674,In_1121,In_4748);
nor U3675 (N_3675,In_866,In_4782);
and U3676 (N_3676,In_792,In_2298);
or U3677 (N_3677,In_2311,In_1331);
and U3678 (N_3678,In_865,In_3381);
xnor U3679 (N_3679,In_2359,In_614);
nor U3680 (N_3680,In_1995,In_4902);
nand U3681 (N_3681,In_4596,In_862);
or U3682 (N_3682,In_3316,In_932);
or U3683 (N_3683,In_4143,In_1556);
nand U3684 (N_3684,In_4932,In_1373);
nand U3685 (N_3685,In_2355,In_1405);
and U3686 (N_3686,In_2824,In_3432);
nor U3687 (N_3687,In_3542,In_2058);
and U3688 (N_3688,In_2125,In_3945);
and U3689 (N_3689,In_3815,In_4035);
nand U3690 (N_3690,In_1596,In_1570);
or U3691 (N_3691,In_3111,In_4992);
xnor U3692 (N_3692,In_22,In_1064);
nor U3693 (N_3693,In_4853,In_3856);
or U3694 (N_3694,In_349,In_457);
nor U3695 (N_3695,In_1134,In_4137);
xnor U3696 (N_3696,In_154,In_3662);
or U3697 (N_3697,In_2990,In_327);
xor U3698 (N_3698,In_3118,In_2254);
and U3699 (N_3699,In_2671,In_227);
nand U3700 (N_3700,In_2686,In_1376);
nand U3701 (N_3701,In_771,In_3231);
or U3702 (N_3702,In_3816,In_117);
nand U3703 (N_3703,In_1806,In_2953);
nor U3704 (N_3704,In_1062,In_2067);
nor U3705 (N_3705,In_2815,In_162);
or U3706 (N_3706,In_2154,In_1487);
and U3707 (N_3707,In_4137,In_3890);
xnor U3708 (N_3708,In_3430,In_2874);
nor U3709 (N_3709,In_3474,In_1695);
nand U3710 (N_3710,In_543,In_4548);
nor U3711 (N_3711,In_1990,In_2787);
nor U3712 (N_3712,In_1575,In_1659);
xor U3713 (N_3713,In_4887,In_2778);
and U3714 (N_3714,In_947,In_3507);
or U3715 (N_3715,In_4257,In_1376);
and U3716 (N_3716,In_1737,In_3672);
nand U3717 (N_3717,In_4098,In_2259);
and U3718 (N_3718,In_409,In_875);
nand U3719 (N_3719,In_4253,In_4972);
or U3720 (N_3720,In_3873,In_707);
nand U3721 (N_3721,In_1706,In_3339);
nand U3722 (N_3722,In_4393,In_2819);
xnor U3723 (N_3723,In_2545,In_540);
nand U3724 (N_3724,In_1120,In_2964);
and U3725 (N_3725,In_944,In_4771);
xor U3726 (N_3726,In_2766,In_2784);
and U3727 (N_3727,In_3171,In_4073);
nand U3728 (N_3728,In_984,In_1836);
or U3729 (N_3729,In_4619,In_706);
xnor U3730 (N_3730,In_4584,In_1055);
and U3731 (N_3731,In_1699,In_4920);
and U3732 (N_3732,In_1099,In_2705);
or U3733 (N_3733,In_1212,In_987);
and U3734 (N_3734,In_147,In_4507);
and U3735 (N_3735,In_2396,In_2155);
or U3736 (N_3736,In_912,In_3066);
or U3737 (N_3737,In_1167,In_1976);
xor U3738 (N_3738,In_3158,In_4454);
nand U3739 (N_3739,In_3007,In_518);
and U3740 (N_3740,In_4713,In_1956);
xor U3741 (N_3741,In_3396,In_1932);
and U3742 (N_3742,In_2186,In_1364);
and U3743 (N_3743,In_1282,In_1001);
nand U3744 (N_3744,In_1380,In_1140);
or U3745 (N_3745,In_521,In_1625);
and U3746 (N_3746,In_4303,In_4350);
and U3747 (N_3747,In_4076,In_3952);
and U3748 (N_3748,In_1944,In_583);
xor U3749 (N_3749,In_1530,In_6);
nor U3750 (N_3750,In_3405,In_69);
xnor U3751 (N_3751,In_1760,In_1366);
or U3752 (N_3752,In_2563,In_4390);
xor U3753 (N_3753,In_4895,In_1531);
and U3754 (N_3754,In_2739,In_3928);
or U3755 (N_3755,In_171,In_1206);
and U3756 (N_3756,In_3825,In_2131);
or U3757 (N_3757,In_2638,In_2823);
and U3758 (N_3758,In_4093,In_4862);
nand U3759 (N_3759,In_4240,In_2433);
or U3760 (N_3760,In_205,In_2409);
or U3761 (N_3761,In_3455,In_2606);
nor U3762 (N_3762,In_819,In_2126);
and U3763 (N_3763,In_2395,In_3006);
and U3764 (N_3764,In_87,In_1424);
nand U3765 (N_3765,In_2957,In_903);
and U3766 (N_3766,In_2409,In_2178);
nand U3767 (N_3767,In_3192,In_2748);
nand U3768 (N_3768,In_2198,In_4619);
xor U3769 (N_3769,In_3453,In_1655);
xnor U3770 (N_3770,In_310,In_4485);
nor U3771 (N_3771,In_4499,In_1730);
nor U3772 (N_3772,In_2963,In_3760);
nand U3773 (N_3773,In_1759,In_440);
and U3774 (N_3774,In_670,In_2964);
nand U3775 (N_3775,In_4948,In_4463);
nand U3776 (N_3776,In_2103,In_2784);
nand U3777 (N_3777,In_238,In_1481);
nand U3778 (N_3778,In_3226,In_1702);
and U3779 (N_3779,In_1599,In_1301);
or U3780 (N_3780,In_40,In_4891);
xnor U3781 (N_3781,In_975,In_4528);
or U3782 (N_3782,In_2940,In_4904);
nand U3783 (N_3783,In_2233,In_1197);
and U3784 (N_3784,In_4189,In_4557);
nor U3785 (N_3785,In_2641,In_4637);
nand U3786 (N_3786,In_4077,In_1310);
nor U3787 (N_3787,In_461,In_740);
nor U3788 (N_3788,In_4980,In_4541);
or U3789 (N_3789,In_3796,In_2780);
or U3790 (N_3790,In_2506,In_4459);
or U3791 (N_3791,In_3676,In_3203);
nand U3792 (N_3792,In_167,In_2041);
and U3793 (N_3793,In_2431,In_1567);
nor U3794 (N_3794,In_1548,In_346);
or U3795 (N_3795,In_697,In_2988);
or U3796 (N_3796,In_2444,In_4276);
or U3797 (N_3797,In_942,In_2014);
and U3798 (N_3798,In_1327,In_4612);
xnor U3799 (N_3799,In_1848,In_2587);
nand U3800 (N_3800,In_3043,In_2661);
xor U3801 (N_3801,In_1460,In_3705);
or U3802 (N_3802,In_3390,In_1717);
xor U3803 (N_3803,In_542,In_4974);
or U3804 (N_3804,In_3482,In_2397);
or U3805 (N_3805,In_2476,In_1040);
nand U3806 (N_3806,In_2362,In_1504);
and U3807 (N_3807,In_4101,In_812);
nand U3808 (N_3808,In_1531,In_621);
and U3809 (N_3809,In_446,In_4579);
xnor U3810 (N_3810,In_3178,In_419);
nand U3811 (N_3811,In_2865,In_1794);
and U3812 (N_3812,In_52,In_2181);
or U3813 (N_3813,In_472,In_1715);
nand U3814 (N_3814,In_1397,In_2930);
or U3815 (N_3815,In_2900,In_4909);
or U3816 (N_3816,In_2379,In_2783);
or U3817 (N_3817,In_1455,In_3630);
and U3818 (N_3818,In_1138,In_718);
or U3819 (N_3819,In_1029,In_3163);
xnor U3820 (N_3820,In_1808,In_531);
and U3821 (N_3821,In_2025,In_294);
or U3822 (N_3822,In_1894,In_2973);
nor U3823 (N_3823,In_2082,In_3337);
or U3824 (N_3824,In_2950,In_1452);
nor U3825 (N_3825,In_578,In_3923);
nor U3826 (N_3826,In_935,In_4417);
nor U3827 (N_3827,In_2793,In_765);
and U3828 (N_3828,In_4954,In_4351);
and U3829 (N_3829,In_3195,In_4732);
nand U3830 (N_3830,In_943,In_3884);
xor U3831 (N_3831,In_3863,In_1423);
nand U3832 (N_3832,In_3433,In_4175);
and U3833 (N_3833,In_4143,In_1836);
or U3834 (N_3834,In_1160,In_2213);
and U3835 (N_3835,In_3815,In_3081);
nor U3836 (N_3836,In_35,In_2577);
and U3837 (N_3837,In_3089,In_3156);
nor U3838 (N_3838,In_2324,In_2756);
nor U3839 (N_3839,In_3549,In_3704);
or U3840 (N_3840,In_3677,In_4947);
or U3841 (N_3841,In_544,In_4519);
nand U3842 (N_3842,In_2800,In_2289);
or U3843 (N_3843,In_1030,In_4610);
and U3844 (N_3844,In_2583,In_4021);
xor U3845 (N_3845,In_3180,In_1295);
or U3846 (N_3846,In_4784,In_3906);
xnor U3847 (N_3847,In_2417,In_4201);
or U3848 (N_3848,In_1485,In_1757);
and U3849 (N_3849,In_4071,In_3959);
or U3850 (N_3850,In_3943,In_1081);
and U3851 (N_3851,In_2255,In_858);
or U3852 (N_3852,In_1676,In_230);
xnor U3853 (N_3853,In_1942,In_2922);
nor U3854 (N_3854,In_2219,In_475);
or U3855 (N_3855,In_2013,In_2678);
xor U3856 (N_3856,In_2433,In_2990);
xor U3857 (N_3857,In_2839,In_3150);
nand U3858 (N_3858,In_4928,In_1869);
nand U3859 (N_3859,In_3276,In_2336);
and U3860 (N_3860,In_2839,In_1306);
and U3861 (N_3861,In_2637,In_1775);
nand U3862 (N_3862,In_4136,In_3330);
xnor U3863 (N_3863,In_508,In_1564);
or U3864 (N_3864,In_671,In_4438);
or U3865 (N_3865,In_3263,In_569);
and U3866 (N_3866,In_1747,In_4754);
nand U3867 (N_3867,In_3972,In_3339);
xnor U3868 (N_3868,In_2687,In_3108);
nor U3869 (N_3869,In_21,In_218);
xor U3870 (N_3870,In_752,In_3852);
xnor U3871 (N_3871,In_1024,In_1784);
nand U3872 (N_3872,In_4009,In_901);
or U3873 (N_3873,In_3947,In_1072);
nand U3874 (N_3874,In_1235,In_2418);
or U3875 (N_3875,In_1762,In_641);
xnor U3876 (N_3876,In_3485,In_1083);
and U3877 (N_3877,In_2604,In_294);
nand U3878 (N_3878,In_1410,In_3827);
nand U3879 (N_3879,In_2988,In_494);
xnor U3880 (N_3880,In_1592,In_4301);
xor U3881 (N_3881,In_542,In_2841);
xor U3882 (N_3882,In_765,In_2053);
nor U3883 (N_3883,In_2040,In_2752);
nand U3884 (N_3884,In_15,In_4130);
nand U3885 (N_3885,In_2250,In_3440);
nor U3886 (N_3886,In_1250,In_2687);
xor U3887 (N_3887,In_4345,In_2980);
or U3888 (N_3888,In_2251,In_3914);
nand U3889 (N_3889,In_991,In_4553);
xnor U3890 (N_3890,In_4844,In_970);
nor U3891 (N_3891,In_123,In_1913);
xor U3892 (N_3892,In_1651,In_3620);
nor U3893 (N_3893,In_2241,In_9);
or U3894 (N_3894,In_4444,In_4073);
and U3895 (N_3895,In_4969,In_3176);
or U3896 (N_3896,In_911,In_2678);
and U3897 (N_3897,In_4720,In_3466);
nand U3898 (N_3898,In_2675,In_750);
or U3899 (N_3899,In_2546,In_4130);
and U3900 (N_3900,In_1303,In_3445);
xor U3901 (N_3901,In_2927,In_1708);
nand U3902 (N_3902,In_3906,In_3126);
or U3903 (N_3903,In_4372,In_893);
or U3904 (N_3904,In_4807,In_4856);
and U3905 (N_3905,In_2033,In_209);
xor U3906 (N_3906,In_2376,In_4398);
and U3907 (N_3907,In_4188,In_2922);
xnor U3908 (N_3908,In_245,In_234);
and U3909 (N_3909,In_609,In_4421);
nand U3910 (N_3910,In_3200,In_4799);
and U3911 (N_3911,In_3455,In_1216);
or U3912 (N_3912,In_2527,In_4882);
nor U3913 (N_3913,In_1252,In_4663);
nor U3914 (N_3914,In_397,In_1277);
nand U3915 (N_3915,In_3810,In_4068);
or U3916 (N_3916,In_33,In_3816);
xor U3917 (N_3917,In_1666,In_2222);
and U3918 (N_3918,In_591,In_4979);
nor U3919 (N_3919,In_4897,In_2894);
nand U3920 (N_3920,In_3807,In_3382);
nor U3921 (N_3921,In_1034,In_3705);
nor U3922 (N_3922,In_2341,In_120);
xnor U3923 (N_3923,In_1952,In_1867);
nand U3924 (N_3924,In_2486,In_3684);
or U3925 (N_3925,In_4911,In_3802);
or U3926 (N_3926,In_3530,In_1468);
and U3927 (N_3927,In_1576,In_4989);
or U3928 (N_3928,In_1267,In_2411);
or U3929 (N_3929,In_1938,In_2488);
nand U3930 (N_3930,In_3918,In_686);
nor U3931 (N_3931,In_2889,In_769);
and U3932 (N_3932,In_54,In_2909);
nor U3933 (N_3933,In_4824,In_826);
nand U3934 (N_3934,In_1849,In_4758);
nand U3935 (N_3935,In_4673,In_79);
and U3936 (N_3936,In_487,In_723);
nor U3937 (N_3937,In_3773,In_4963);
xnor U3938 (N_3938,In_73,In_1899);
nor U3939 (N_3939,In_1280,In_1691);
xnor U3940 (N_3940,In_2701,In_3267);
xor U3941 (N_3941,In_837,In_1343);
xor U3942 (N_3942,In_873,In_2657);
or U3943 (N_3943,In_1029,In_2480);
or U3944 (N_3944,In_1650,In_1901);
xnor U3945 (N_3945,In_31,In_2780);
or U3946 (N_3946,In_876,In_2317);
xnor U3947 (N_3947,In_4180,In_1481);
xnor U3948 (N_3948,In_2865,In_3418);
and U3949 (N_3949,In_3070,In_3748);
nand U3950 (N_3950,In_1602,In_1054);
or U3951 (N_3951,In_2890,In_3993);
nor U3952 (N_3952,In_3848,In_789);
or U3953 (N_3953,In_402,In_2177);
or U3954 (N_3954,In_4548,In_564);
and U3955 (N_3955,In_1852,In_3009);
and U3956 (N_3956,In_207,In_553);
and U3957 (N_3957,In_179,In_1679);
or U3958 (N_3958,In_495,In_2134);
nor U3959 (N_3959,In_1732,In_1421);
nor U3960 (N_3960,In_24,In_4534);
nand U3961 (N_3961,In_1107,In_2332);
xor U3962 (N_3962,In_1121,In_4337);
nand U3963 (N_3963,In_3671,In_3943);
xor U3964 (N_3964,In_3337,In_2684);
xor U3965 (N_3965,In_4202,In_3325);
nand U3966 (N_3966,In_3965,In_3238);
nand U3967 (N_3967,In_3351,In_701);
nor U3968 (N_3968,In_2720,In_1845);
xnor U3969 (N_3969,In_2648,In_2447);
nand U3970 (N_3970,In_751,In_2648);
or U3971 (N_3971,In_4888,In_4367);
xor U3972 (N_3972,In_4054,In_1172);
nor U3973 (N_3973,In_4833,In_20);
xor U3974 (N_3974,In_207,In_1731);
nor U3975 (N_3975,In_3890,In_2988);
nor U3976 (N_3976,In_451,In_3450);
nand U3977 (N_3977,In_3811,In_3796);
xor U3978 (N_3978,In_4520,In_2818);
or U3979 (N_3979,In_3866,In_3317);
nor U3980 (N_3980,In_528,In_1860);
xor U3981 (N_3981,In_2004,In_2999);
nor U3982 (N_3982,In_4649,In_4419);
nand U3983 (N_3983,In_474,In_989);
nor U3984 (N_3984,In_855,In_470);
nor U3985 (N_3985,In_3843,In_2506);
xor U3986 (N_3986,In_1285,In_1197);
or U3987 (N_3987,In_2023,In_3954);
nor U3988 (N_3988,In_3987,In_1090);
and U3989 (N_3989,In_2044,In_187);
nor U3990 (N_3990,In_29,In_4128);
or U3991 (N_3991,In_4775,In_3323);
and U3992 (N_3992,In_3290,In_3118);
nor U3993 (N_3993,In_1925,In_2911);
xor U3994 (N_3994,In_3246,In_3236);
nand U3995 (N_3995,In_3028,In_3854);
nand U3996 (N_3996,In_2533,In_3320);
nor U3997 (N_3997,In_2890,In_4961);
or U3998 (N_3998,In_2459,In_2864);
xor U3999 (N_3999,In_2991,In_2865);
and U4000 (N_4000,In_54,In_4999);
and U4001 (N_4001,In_2489,In_3867);
nand U4002 (N_4002,In_1615,In_2423);
or U4003 (N_4003,In_4265,In_3352);
or U4004 (N_4004,In_4612,In_4754);
and U4005 (N_4005,In_4076,In_3699);
or U4006 (N_4006,In_268,In_1450);
or U4007 (N_4007,In_1482,In_1628);
or U4008 (N_4008,In_4512,In_3919);
xnor U4009 (N_4009,In_4965,In_2897);
nor U4010 (N_4010,In_388,In_3522);
and U4011 (N_4011,In_1507,In_718);
xor U4012 (N_4012,In_3444,In_2080);
xnor U4013 (N_4013,In_3648,In_4568);
nand U4014 (N_4014,In_1192,In_4557);
nand U4015 (N_4015,In_3608,In_4842);
xor U4016 (N_4016,In_1480,In_1275);
nor U4017 (N_4017,In_3861,In_632);
and U4018 (N_4018,In_772,In_3035);
xor U4019 (N_4019,In_3010,In_2360);
and U4020 (N_4020,In_1863,In_3380);
and U4021 (N_4021,In_616,In_1557);
or U4022 (N_4022,In_900,In_882);
and U4023 (N_4023,In_3140,In_2327);
and U4024 (N_4024,In_1127,In_4118);
xnor U4025 (N_4025,In_4849,In_2325);
nand U4026 (N_4026,In_4722,In_4310);
and U4027 (N_4027,In_4231,In_2117);
and U4028 (N_4028,In_4105,In_813);
nor U4029 (N_4029,In_4473,In_4925);
xor U4030 (N_4030,In_2146,In_565);
or U4031 (N_4031,In_4144,In_397);
nor U4032 (N_4032,In_471,In_962);
nor U4033 (N_4033,In_4266,In_4664);
and U4034 (N_4034,In_4942,In_2976);
nor U4035 (N_4035,In_4928,In_2218);
nor U4036 (N_4036,In_4500,In_1716);
xor U4037 (N_4037,In_4930,In_2863);
and U4038 (N_4038,In_766,In_1221);
and U4039 (N_4039,In_3234,In_1662);
xor U4040 (N_4040,In_4682,In_3050);
nand U4041 (N_4041,In_623,In_4309);
or U4042 (N_4042,In_1362,In_1753);
and U4043 (N_4043,In_317,In_4688);
xor U4044 (N_4044,In_3400,In_2664);
nor U4045 (N_4045,In_1051,In_512);
or U4046 (N_4046,In_108,In_4757);
or U4047 (N_4047,In_2595,In_4281);
or U4048 (N_4048,In_1065,In_4872);
xnor U4049 (N_4049,In_1878,In_4046);
nor U4050 (N_4050,In_500,In_621);
nand U4051 (N_4051,In_3551,In_4189);
nor U4052 (N_4052,In_4901,In_4669);
nand U4053 (N_4053,In_4263,In_4113);
or U4054 (N_4054,In_4737,In_4843);
or U4055 (N_4055,In_3606,In_1639);
and U4056 (N_4056,In_3172,In_4755);
or U4057 (N_4057,In_187,In_312);
nand U4058 (N_4058,In_1037,In_4361);
nand U4059 (N_4059,In_1278,In_1585);
xnor U4060 (N_4060,In_4415,In_3949);
and U4061 (N_4061,In_2494,In_4497);
xnor U4062 (N_4062,In_1248,In_2079);
nand U4063 (N_4063,In_2434,In_536);
and U4064 (N_4064,In_2508,In_1803);
nand U4065 (N_4065,In_2787,In_3635);
nor U4066 (N_4066,In_2540,In_2058);
nand U4067 (N_4067,In_382,In_65);
nand U4068 (N_4068,In_1454,In_2162);
or U4069 (N_4069,In_1457,In_1208);
and U4070 (N_4070,In_2044,In_4578);
nand U4071 (N_4071,In_4598,In_4793);
or U4072 (N_4072,In_3726,In_255);
and U4073 (N_4073,In_1937,In_2599);
or U4074 (N_4074,In_1312,In_2013);
nor U4075 (N_4075,In_4448,In_2915);
xnor U4076 (N_4076,In_628,In_4805);
and U4077 (N_4077,In_3365,In_4678);
nor U4078 (N_4078,In_685,In_3377);
xnor U4079 (N_4079,In_2114,In_4229);
xor U4080 (N_4080,In_189,In_4895);
nand U4081 (N_4081,In_1759,In_4185);
xor U4082 (N_4082,In_3862,In_1429);
xor U4083 (N_4083,In_1609,In_229);
nand U4084 (N_4084,In_1672,In_1465);
nand U4085 (N_4085,In_117,In_4159);
nand U4086 (N_4086,In_971,In_1844);
nor U4087 (N_4087,In_2281,In_2768);
and U4088 (N_4088,In_3035,In_2382);
and U4089 (N_4089,In_1902,In_3896);
nor U4090 (N_4090,In_1355,In_1633);
or U4091 (N_4091,In_717,In_3336);
nor U4092 (N_4092,In_2094,In_1429);
or U4093 (N_4093,In_2863,In_4276);
nor U4094 (N_4094,In_782,In_2201);
and U4095 (N_4095,In_2062,In_2060);
xnor U4096 (N_4096,In_2838,In_1807);
nor U4097 (N_4097,In_1804,In_1593);
nand U4098 (N_4098,In_3870,In_649);
xor U4099 (N_4099,In_1659,In_973);
nor U4100 (N_4100,In_32,In_852);
nor U4101 (N_4101,In_4960,In_4408);
nand U4102 (N_4102,In_4572,In_1513);
nor U4103 (N_4103,In_1140,In_1730);
nor U4104 (N_4104,In_3721,In_2085);
nand U4105 (N_4105,In_3219,In_1043);
nand U4106 (N_4106,In_1577,In_1146);
xnor U4107 (N_4107,In_1839,In_4023);
nand U4108 (N_4108,In_4713,In_522);
nor U4109 (N_4109,In_3025,In_2965);
xor U4110 (N_4110,In_170,In_2838);
xor U4111 (N_4111,In_2110,In_3044);
xnor U4112 (N_4112,In_3368,In_3010);
and U4113 (N_4113,In_705,In_3287);
nor U4114 (N_4114,In_4075,In_1179);
nor U4115 (N_4115,In_4273,In_4439);
or U4116 (N_4116,In_2320,In_3845);
xnor U4117 (N_4117,In_4428,In_3820);
xnor U4118 (N_4118,In_2210,In_4595);
or U4119 (N_4119,In_4170,In_1857);
xnor U4120 (N_4120,In_1456,In_1679);
nor U4121 (N_4121,In_2835,In_838);
or U4122 (N_4122,In_973,In_1117);
or U4123 (N_4123,In_4134,In_2871);
or U4124 (N_4124,In_2942,In_3313);
nor U4125 (N_4125,In_3122,In_4688);
nand U4126 (N_4126,In_2134,In_2401);
and U4127 (N_4127,In_2672,In_271);
nor U4128 (N_4128,In_1850,In_294);
nand U4129 (N_4129,In_2313,In_1964);
nor U4130 (N_4130,In_1960,In_218);
and U4131 (N_4131,In_4942,In_2606);
and U4132 (N_4132,In_1402,In_2336);
nor U4133 (N_4133,In_478,In_3516);
and U4134 (N_4134,In_1456,In_2283);
and U4135 (N_4135,In_2764,In_2382);
nand U4136 (N_4136,In_3568,In_1048);
xnor U4137 (N_4137,In_3584,In_1686);
and U4138 (N_4138,In_4384,In_4961);
nor U4139 (N_4139,In_2915,In_2971);
nor U4140 (N_4140,In_642,In_938);
nor U4141 (N_4141,In_1554,In_718);
nand U4142 (N_4142,In_1450,In_328);
xor U4143 (N_4143,In_2250,In_2871);
or U4144 (N_4144,In_1444,In_4656);
or U4145 (N_4145,In_4343,In_2886);
or U4146 (N_4146,In_1540,In_3519);
xnor U4147 (N_4147,In_64,In_3942);
xnor U4148 (N_4148,In_603,In_3981);
or U4149 (N_4149,In_307,In_409);
xnor U4150 (N_4150,In_1604,In_1583);
and U4151 (N_4151,In_1387,In_2120);
or U4152 (N_4152,In_3979,In_3992);
nand U4153 (N_4153,In_3157,In_4618);
nand U4154 (N_4154,In_4710,In_3727);
xnor U4155 (N_4155,In_1579,In_9);
or U4156 (N_4156,In_2240,In_2426);
xnor U4157 (N_4157,In_526,In_380);
and U4158 (N_4158,In_4253,In_2477);
nor U4159 (N_4159,In_2040,In_718);
nand U4160 (N_4160,In_949,In_4007);
nor U4161 (N_4161,In_1745,In_4160);
or U4162 (N_4162,In_1475,In_4665);
xor U4163 (N_4163,In_3245,In_2005);
and U4164 (N_4164,In_1585,In_4792);
and U4165 (N_4165,In_2763,In_3783);
nor U4166 (N_4166,In_1481,In_2268);
nand U4167 (N_4167,In_1654,In_823);
nor U4168 (N_4168,In_1293,In_3885);
nor U4169 (N_4169,In_4993,In_2642);
xor U4170 (N_4170,In_2380,In_3933);
or U4171 (N_4171,In_567,In_714);
nand U4172 (N_4172,In_3229,In_4998);
nand U4173 (N_4173,In_902,In_1589);
and U4174 (N_4174,In_4536,In_4286);
and U4175 (N_4175,In_3092,In_1973);
and U4176 (N_4176,In_1036,In_3324);
and U4177 (N_4177,In_1188,In_3949);
xnor U4178 (N_4178,In_3103,In_1972);
nor U4179 (N_4179,In_2180,In_2911);
xor U4180 (N_4180,In_3442,In_3886);
or U4181 (N_4181,In_4903,In_3926);
nand U4182 (N_4182,In_3814,In_3200);
nor U4183 (N_4183,In_2291,In_283);
nand U4184 (N_4184,In_4397,In_2170);
nand U4185 (N_4185,In_114,In_4864);
or U4186 (N_4186,In_719,In_867);
nand U4187 (N_4187,In_1175,In_971);
or U4188 (N_4188,In_635,In_2879);
nand U4189 (N_4189,In_2069,In_26);
xor U4190 (N_4190,In_3630,In_68);
or U4191 (N_4191,In_631,In_1745);
and U4192 (N_4192,In_3320,In_1790);
or U4193 (N_4193,In_3304,In_4447);
or U4194 (N_4194,In_1159,In_3952);
and U4195 (N_4195,In_3737,In_4612);
or U4196 (N_4196,In_2872,In_1884);
and U4197 (N_4197,In_1112,In_1278);
or U4198 (N_4198,In_4878,In_46);
xor U4199 (N_4199,In_1528,In_969);
and U4200 (N_4200,In_3580,In_3833);
nor U4201 (N_4201,In_2537,In_2428);
or U4202 (N_4202,In_542,In_4547);
nor U4203 (N_4203,In_588,In_907);
nor U4204 (N_4204,In_2388,In_4404);
xnor U4205 (N_4205,In_3824,In_1204);
nor U4206 (N_4206,In_1178,In_1960);
and U4207 (N_4207,In_559,In_3958);
nor U4208 (N_4208,In_2996,In_2790);
nand U4209 (N_4209,In_667,In_4118);
xor U4210 (N_4210,In_4035,In_421);
and U4211 (N_4211,In_4582,In_754);
nor U4212 (N_4212,In_4808,In_1063);
xnor U4213 (N_4213,In_1068,In_195);
nor U4214 (N_4214,In_306,In_2278);
and U4215 (N_4215,In_2324,In_3116);
xor U4216 (N_4216,In_1727,In_4161);
and U4217 (N_4217,In_1988,In_2891);
and U4218 (N_4218,In_1720,In_2490);
nand U4219 (N_4219,In_1272,In_3341);
or U4220 (N_4220,In_4889,In_2161);
xnor U4221 (N_4221,In_544,In_2024);
xor U4222 (N_4222,In_1630,In_4291);
nor U4223 (N_4223,In_191,In_1650);
nand U4224 (N_4224,In_3678,In_3320);
nand U4225 (N_4225,In_349,In_649);
xor U4226 (N_4226,In_4253,In_4145);
nor U4227 (N_4227,In_2523,In_3516);
nand U4228 (N_4228,In_2502,In_3195);
nand U4229 (N_4229,In_2323,In_4115);
nand U4230 (N_4230,In_2167,In_3115);
xor U4231 (N_4231,In_1624,In_1050);
and U4232 (N_4232,In_4222,In_2343);
nor U4233 (N_4233,In_3083,In_4286);
nor U4234 (N_4234,In_1169,In_508);
nor U4235 (N_4235,In_2553,In_1771);
and U4236 (N_4236,In_4816,In_1956);
or U4237 (N_4237,In_1729,In_2403);
xor U4238 (N_4238,In_2299,In_683);
xnor U4239 (N_4239,In_1859,In_3209);
xnor U4240 (N_4240,In_236,In_2095);
nor U4241 (N_4241,In_3503,In_4716);
xor U4242 (N_4242,In_3245,In_3978);
or U4243 (N_4243,In_3467,In_1253);
or U4244 (N_4244,In_1447,In_1300);
nand U4245 (N_4245,In_2086,In_586);
nor U4246 (N_4246,In_3830,In_976);
xor U4247 (N_4247,In_615,In_4899);
nand U4248 (N_4248,In_1867,In_4024);
or U4249 (N_4249,In_2044,In_4176);
or U4250 (N_4250,In_1306,In_2541);
xor U4251 (N_4251,In_579,In_996);
nor U4252 (N_4252,In_4877,In_1627);
nand U4253 (N_4253,In_498,In_1512);
nor U4254 (N_4254,In_2772,In_849);
nor U4255 (N_4255,In_2431,In_3088);
and U4256 (N_4256,In_1296,In_2044);
xor U4257 (N_4257,In_3814,In_4276);
and U4258 (N_4258,In_1684,In_560);
or U4259 (N_4259,In_4674,In_2361);
or U4260 (N_4260,In_2427,In_3850);
or U4261 (N_4261,In_1401,In_3849);
xor U4262 (N_4262,In_2836,In_1313);
and U4263 (N_4263,In_3148,In_4020);
nand U4264 (N_4264,In_3036,In_1152);
or U4265 (N_4265,In_1118,In_4871);
and U4266 (N_4266,In_2242,In_3100);
nor U4267 (N_4267,In_1375,In_3313);
and U4268 (N_4268,In_3060,In_420);
or U4269 (N_4269,In_3761,In_1676);
xor U4270 (N_4270,In_1018,In_2672);
xnor U4271 (N_4271,In_716,In_1305);
nor U4272 (N_4272,In_1319,In_658);
xor U4273 (N_4273,In_3375,In_4906);
or U4274 (N_4274,In_3836,In_4846);
nand U4275 (N_4275,In_4786,In_2304);
or U4276 (N_4276,In_926,In_1520);
or U4277 (N_4277,In_800,In_1771);
and U4278 (N_4278,In_3375,In_327);
xor U4279 (N_4279,In_218,In_2987);
or U4280 (N_4280,In_2709,In_1281);
or U4281 (N_4281,In_1360,In_3749);
xor U4282 (N_4282,In_1291,In_1408);
or U4283 (N_4283,In_344,In_4083);
and U4284 (N_4284,In_4013,In_3587);
xnor U4285 (N_4285,In_3933,In_1970);
nor U4286 (N_4286,In_2928,In_514);
nor U4287 (N_4287,In_2951,In_2944);
nor U4288 (N_4288,In_3807,In_4426);
nand U4289 (N_4289,In_1437,In_2451);
nand U4290 (N_4290,In_398,In_107);
xnor U4291 (N_4291,In_3520,In_3628);
and U4292 (N_4292,In_1119,In_3077);
or U4293 (N_4293,In_592,In_4902);
and U4294 (N_4294,In_1992,In_1090);
or U4295 (N_4295,In_3875,In_646);
nand U4296 (N_4296,In_2965,In_4338);
and U4297 (N_4297,In_2446,In_405);
and U4298 (N_4298,In_4627,In_1661);
nand U4299 (N_4299,In_128,In_1233);
nor U4300 (N_4300,In_1430,In_331);
or U4301 (N_4301,In_3534,In_4311);
xnor U4302 (N_4302,In_2273,In_3281);
xnor U4303 (N_4303,In_1840,In_2757);
or U4304 (N_4304,In_4935,In_4412);
nor U4305 (N_4305,In_4702,In_3368);
nand U4306 (N_4306,In_4030,In_838);
and U4307 (N_4307,In_2582,In_3691);
nand U4308 (N_4308,In_4943,In_694);
xnor U4309 (N_4309,In_563,In_4415);
or U4310 (N_4310,In_3945,In_4872);
and U4311 (N_4311,In_1221,In_4907);
nor U4312 (N_4312,In_855,In_543);
xnor U4313 (N_4313,In_1621,In_3494);
nand U4314 (N_4314,In_1760,In_211);
and U4315 (N_4315,In_2430,In_3484);
xor U4316 (N_4316,In_512,In_1981);
or U4317 (N_4317,In_2333,In_4474);
nor U4318 (N_4318,In_548,In_1899);
or U4319 (N_4319,In_2701,In_961);
or U4320 (N_4320,In_892,In_2620);
nor U4321 (N_4321,In_4253,In_397);
nor U4322 (N_4322,In_3961,In_2315);
and U4323 (N_4323,In_531,In_603);
nor U4324 (N_4324,In_4841,In_4813);
nand U4325 (N_4325,In_1451,In_4942);
or U4326 (N_4326,In_4958,In_2418);
xor U4327 (N_4327,In_1266,In_738);
nor U4328 (N_4328,In_3554,In_4250);
xnor U4329 (N_4329,In_674,In_1975);
or U4330 (N_4330,In_3145,In_4954);
nand U4331 (N_4331,In_717,In_4916);
nor U4332 (N_4332,In_4138,In_3276);
and U4333 (N_4333,In_3543,In_4139);
xnor U4334 (N_4334,In_2,In_3262);
xnor U4335 (N_4335,In_988,In_1840);
xnor U4336 (N_4336,In_167,In_3226);
xnor U4337 (N_4337,In_4171,In_1116);
nor U4338 (N_4338,In_1315,In_4927);
and U4339 (N_4339,In_1834,In_1965);
or U4340 (N_4340,In_239,In_756);
and U4341 (N_4341,In_1386,In_421);
or U4342 (N_4342,In_894,In_4917);
nor U4343 (N_4343,In_3328,In_2270);
nor U4344 (N_4344,In_4238,In_4446);
nand U4345 (N_4345,In_1143,In_2144);
xor U4346 (N_4346,In_2151,In_1410);
nand U4347 (N_4347,In_1071,In_3997);
and U4348 (N_4348,In_542,In_1326);
and U4349 (N_4349,In_1169,In_3807);
nor U4350 (N_4350,In_794,In_2653);
or U4351 (N_4351,In_833,In_275);
xnor U4352 (N_4352,In_1280,In_1519);
or U4353 (N_4353,In_1561,In_3118);
nor U4354 (N_4354,In_3278,In_2651);
or U4355 (N_4355,In_48,In_274);
or U4356 (N_4356,In_395,In_4760);
nand U4357 (N_4357,In_4927,In_1375);
nor U4358 (N_4358,In_1679,In_1452);
or U4359 (N_4359,In_1834,In_1550);
nor U4360 (N_4360,In_3150,In_4086);
and U4361 (N_4361,In_3597,In_68);
nand U4362 (N_4362,In_1465,In_1035);
or U4363 (N_4363,In_1225,In_849);
nand U4364 (N_4364,In_1785,In_1772);
xnor U4365 (N_4365,In_3310,In_3933);
nor U4366 (N_4366,In_3976,In_4424);
nor U4367 (N_4367,In_3048,In_2895);
and U4368 (N_4368,In_2564,In_237);
and U4369 (N_4369,In_3461,In_3463);
xor U4370 (N_4370,In_4747,In_4318);
nor U4371 (N_4371,In_3449,In_4786);
nand U4372 (N_4372,In_1080,In_2090);
and U4373 (N_4373,In_3582,In_1226);
and U4374 (N_4374,In_2349,In_3131);
or U4375 (N_4375,In_981,In_2904);
xnor U4376 (N_4376,In_4676,In_2846);
and U4377 (N_4377,In_3648,In_78);
nor U4378 (N_4378,In_714,In_814);
nor U4379 (N_4379,In_3893,In_638);
xor U4380 (N_4380,In_3411,In_4974);
or U4381 (N_4381,In_245,In_2031);
and U4382 (N_4382,In_2737,In_4783);
or U4383 (N_4383,In_4979,In_3096);
or U4384 (N_4384,In_2210,In_2186);
xnor U4385 (N_4385,In_2681,In_4292);
and U4386 (N_4386,In_1619,In_2534);
nor U4387 (N_4387,In_1673,In_4206);
nand U4388 (N_4388,In_3580,In_4668);
xnor U4389 (N_4389,In_2154,In_4860);
or U4390 (N_4390,In_3073,In_1447);
xnor U4391 (N_4391,In_97,In_1718);
and U4392 (N_4392,In_2955,In_4719);
xor U4393 (N_4393,In_2869,In_4897);
nand U4394 (N_4394,In_3384,In_319);
xor U4395 (N_4395,In_936,In_4779);
or U4396 (N_4396,In_1225,In_4285);
xor U4397 (N_4397,In_1581,In_2976);
or U4398 (N_4398,In_3720,In_1435);
nand U4399 (N_4399,In_4539,In_3554);
nor U4400 (N_4400,In_168,In_3597);
and U4401 (N_4401,In_2240,In_1673);
xnor U4402 (N_4402,In_1095,In_3224);
or U4403 (N_4403,In_4371,In_2230);
xor U4404 (N_4404,In_492,In_1044);
and U4405 (N_4405,In_4260,In_2798);
xor U4406 (N_4406,In_661,In_3313);
xor U4407 (N_4407,In_2570,In_4177);
or U4408 (N_4408,In_230,In_2519);
and U4409 (N_4409,In_4939,In_2294);
or U4410 (N_4410,In_1247,In_673);
and U4411 (N_4411,In_1367,In_2853);
or U4412 (N_4412,In_4113,In_2052);
nand U4413 (N_4413,In_4357,In_2927);
and U4414 (N_4414,In_3818,In_1556);
and U4415 (N_4415,In_1532,In_4389);
and U4416 (N_4416,In_2772,In_3177);
xnor U4417 (N_4417,In_2815,In_401);
and U4418 (N_4418,In_3281,In_1995);
xnor U4419 (N_4419,In_3393,In_2257);
xnor U4420 (N_4420,In_3041,In_1138);
nand U4421 (N_4421,In_110,In_1451);
nand U4422 (N_4422,In_4121,In_1088);
and U4423 (N_4423,In_2409,In_2441);
or U4424 (N_4424,In_312,In_300);
nand U4425 (N_4425,In_2017,In_1797);
or U4426 (N_4426,In_1431,In_1827);
or U4427 (N_4427,In_2635,In_3549);
and U4428 (N_4428,In_3024,In_3961);
nand U4429 (N_4429,In_4330,In_4780);
or U4430 (N_4430,In_4182,In_67);
or U4431 (N_4431,In_4255,In_3038);
xor U4432 (N_4432,In_1414,In_1435);
nand U4433 (N_4433,In_786,In_2405);
or U4434 (N_4434,In_3748,In_283);
or U4435 (N_4435,In_2550,In_4552);
xnor U4436 (N_4436,In_1376,In_3097);
nand U4437 (N_4437,In_4247,In_1434);
nor U4438 (N_4438,In_4927,In_3248);
or U4439 (N_4439,In_2079,In_2339);
or U4440 (N_4440,In_327,In_4555);
and U4441 (N_4441,In_303,In_23);
and U4442 (N_4442,In_2087,In_2625);
or U4443 (N_4443,In_478,In_3186);
and U4444 (N_4444,In_348,In_1290);
nor U4445 (N_4445,In_145,In_3309);
and U4446 (N_4446,In_4188,In_344);
nor U4447 (N_4447,In_3068,In_2391);
and U4448 (N_4448,In_4908,In_1183);
and U4449 (N_4449,In_1459,In_1054);
and U4450 (N_4450,In_4914,In_3919);
or U4451 (N_4451,In_3382,In_240);
nor U4452 (N_4452,In_3737,In_2046);
xnor U4453 (N_4453,In_2824,In_2967);
xor U4454 (N_4454,In_723,In_2632);
nand U4455 (N_4455,In_4455,In_331);
nand U4456 (N_4456,In_4945,In_1998);
xnor U4457 (N_4457,In_3901,In_1033);
nand U4458 (N_4458,In_1233,In_4405);
nand U4459 (N_4459,In_4437,In_481);
nand U4460 (N_4460,In_3516,In_2732);
nor U4461 (N_4461,In_907,In_4073);
nor U4462 (N_4462,In_1255,In_2464);
xnor U4463 (N_4463,In_591,In_4278);
nor U4464 (N_4464,In_4583,In_2874);
and U4465 (N_4465,In_1814,In_462);
xnor U4466 (N_4466,In_2378,In_267);
or U4467 (N_4467,In_3546,In_2263);
nand U4468 (N_4468,In_2991,In_2176);
nor U4469 (N_4469,In_159,In_2272);
or U4470 (N_4470,In_3708,In_4635);
or U4471 (N_4471,In_2873,In_8);
or U4472 (N_4472,In_1584,In_1804);
xnor U4473 (N_4473,In_1698,In_4244);
or U4474 (N_4474,In_245,In_4154);
nor U4475 (N_4475,In_4179,In_4616);
and U4476 (N_4476,In_4244,In_685);
xnor U4477 (N_4477,In_1412,In_3869);
nand U4478 (N_4478,In_2644,In_4487);
and U4479 (N_4479,In_132,In_1076);
nor U4480 (N_4480,In_1725,In_2372);
or U4481 (N_4481,In_2722,In_4486);
nor U4482 (N_4482,In_1291,In_1701);
and U4483 (N_4483,In_2157,In_681);
xor U4484 (N_4484,In_3590,In_1568);
nand U4485 (N_4485,In_1884,In_4320);
and U4486 (N_4486,In_2558,In_3523);
nor U4487 (N_4487,In_3288,In_4690);
and U4488 (N_4488,In_2588,In_4824);
nor U4489 (N_4489,In_2204,In_162);
nor U4490 (N_4490,In_80,In_3238);
xnor U4491 (N_4491,In_2790,In_1746);
and U4492 (N_4492,In_1506,In_1539);
and U4493 (N_4493,In_1844,In_382);
nor U4494 (N_4494,In_4011,In_3370);
or U4495 (N_4495,In_4902,In_2539);
or U4496 (N_4496,In_4437,In_3355);
xnor U4497 (N_4497,In_4306,In_3999);
xnor U4498 (N_4498,In_3783,In_4061);
nand U4499 (N_4499,In_2586,In_4354);
nor U4500 (N_4500,In_4797,In_3091);
and U4501 (N_4501,In_1779,In_4224);
nor U4502 (N_4502,In_239,In_3135);
and U4503 (N_4503,In_3946,In_2212);
or U4504 (N_4504,In_2525,In_1979);
xor U4505 (N_4505,In_1269,In_256);
nor U4506 (N_4506,In_1842,In_2046);
and U4507 (N_4507,In_1182,In_3470);
xnor U4508 (N_4508,In_3591,In_4351);
and U4509 (N_4509,In_4670,In_3482);
and U4510 (N_4510,In_1756,In_4912);
and U4511 (N_4511,In_4889,In_4912);
and U4512 (N_4512,In_1302,In_3389);
nor U4513 (N_4513,In_1682,In_4757);
and U4514 (N_4514,In_2699,In_1138);
or U4515 (N_4515,In_1135,In_4856);
nor U4516 (N_4516,In_3661,In_212);
nand U4517 (N_4517,In_1771,In_4112);
xnor U4518 (N_4518,In_1372,In_2189);
and U4519 (N_4519,In_4246,In_4137);
nor U4520 (N_4520,In_1831,In_3589);
xor U4521 (N_4521,In_347,In_4336);
nand U4522 (N_4522,In_774,In_3220);
xnor U4523 (N_4523,In_2054,In_1326);
xor U4524 (N_4524,In_3666,In_260);
and U4525 (N_4525,In_346,In_3094);
nor U4526 (N_4526,In_915,In_1999);
xnor U4527 (N_4527,In_3510,In_1584);
or U4528 (N_4528,In_1965,In_1939);
nor U4529 (N_4529,In_850,In_3790);
or U4530 (N_4530,In_20,In_228);
nor U4531 (N_4531,In_3832,In_4051);
or U4532 (N_4532,In_2787,In_393);
nand U4533 (N_4533,In_2403,In_3581);
and U4534 (N_4534,In_1358,In_4202);
and U4535 (N_4535,In_3329,In_3647);
nor U4536 (N_4536,In_3736,In_161);
nor U4537 (N_4537,In_2715,In_4240);
or U4538 (N_4538,In_3289,In_2067);
nand U4539 (N_4539,In_2967,In_4301);
nor U4540 (N_4540,In_1721,In_3097);
nand U4541 (N_4541,In_4455,In_2496);
xor U4542 (N_4542,In_1350,In_743);
and U4543 (N_4543,In_4253,In_1505);
nand U4544 (N_4544,In_2363,In_2650);
xor U4545 (N_4545,In_3145,In_1515);
nand U4546 (N_4546,In_2392,In_29);
xor U4547 (N_4547,In_3187,In_2086);
nor U4548 (N_4548,In_432,In_2914);
or U4549 (N_4549,In_2567,In_1559);
nor U4550 (N_4550,In_2993,In_642);
xnor U4551 (N_4551,In_3581,In_1412);
and U4552 (N_4552,In_3187,In_1848);
xnor U4553 (N_4553,In_375,In_1423);
nor U4554 (N_4554,In_1604,In_804);
xnor U4555 (N_4555,In_4479,In_1579);
and U4556 (N_4556,In_4119,In_3175);
or U4557 (N_4557,In_4704,In_1903);
or U4558 (N_4558,In_270,In_3158);
xnor U4559 (N_4559,In_11,In_2823);
xor U4560 (N_4560,In_805,In_3837);
and U4561 (N_4561,In_2385,In_2680);
or U4562 (N_4562,In_4665,In_1415);
and U4563 (N_4563,In_1378,In_3069);
nand U4564 (N_4564,In_1163,In_1020);
nand U4565 (N_4565,In_2915,In_2680);
and U4566 (N_4566,In_4824,In_3400);
xnor U4567 (N_4567,In_1632,In_4628);
or U4568 (N_4568,In_1708,In_2197);
nand U4569 (N_4569,In_2366,In_4468);
xor U4570 (N_4570,In_1756,In_2614);
nor U4571 (N_4571,In_1280,In_3235);
and U4572 (N_4572,In_2235,In_4339);
or U4573 (N_4573,In_3394,In_2153);
and U4574 (N_4574,In_2156,In_1026);
and U4575 (N_4575,In_2924,In_4118);
nor U4576 (N_4576,In_3795,In_1815);
or U4577 (N_4577,In_4637,In_1432);
nor U4578 (N_4578,In_1084,In_861);
nor U4579 (N_4579,In_4690,In_3568);
nand U4580 (N_4580,In_1833,In_3945);
xor U4581 (N_4581,In_2022,In_3875);
nand U4582 (N_4582,In_1608,In_2164);
or U4583 (N_4583,In_816,In_4099);
nand U4584 (N_4584,In_4346,In_4320);
or U4585 (N_4585,In_2647,In_1515);
and U4586 (N_4586,In_1481,In_3845);
xor U4587 (N_4587,In_3886,In_1300);
and U4588 (N_4588,In_4816,In_1211);
nor U4589 (N_4589,In_466,In_478);
and U4590 (N_4590,In_2392,In_4635);
nor U4591 (N_4591,In_2196,In_1968);
nor U4592 (N_4592,In_229,In_3416);
and U4593 (N_4593,In_4462,In_1832);
and U4594 (N_4594,In_3014,In_3549);
nor U4595 (N_4595,In_4816,In_911);
nand U4596 (N_4596,In_2501,In_70);
or U4597 (N_4597,In_3340,In_446);
nor U4598 (N_4598,In_1655,In_4549);
nor U4599 (N_4599,In_767,In_2169);
xnor U4600 (N_4600,In_3214,In_1277);
xnor U4601 (N_4601,In_1930,In_2849);
nor U4602 (N_4602,In_1296,In_1231);
nor U4603 (N_4603,In_3687,In_1007);
and U4604 (N_4604,In_1675,In_1337);
nand U4605 (N_4605,In_1784,In_846);
nand U4606 (N_4606,In_2078,In_4103);
xnor U4607 (N_4607,In_4744,In_2719);
nor U4608 (N_4608,In_3253,In_996);
nand U4609 (N_4609,In_4052,In_1609);
nand U4610 (N_4610,In_4894,In_88);
or U4611 (N_4611,In_4211,In_3694);
nor U4612 (N_4612,In_2983,In_4726);
xnor U4613 (N_4613,In_2739,In_1574);
nand U4614 (N_4614,In_3431,In_963);
and U4615 (N_4615,In_1799,In_2200);
nand U4616 (N_4616,In_4769,In_1482);
xor U4617 (N_4617,In_4503,In_4788);
nand U4618 (N_4618,In_2394,In_1757);
nor U4619 (N_4619,In_4904,In_3896);
and U4620 (N_4620,In_2637,In_1960);
nand U4621 (N_4621,In_3259,In_2976);
and U4622 (N_4622,In_1124,In_4104);
or U4623 (N_4623,In_420,In_4314);
nor U4624 (N_4624,In_1251,In_3181);
nand U4625 (N_4625,In_4725,In_2608);
xor U4626 (N_4626,In_1135,In_4760);
nor U4627 (N_4627,In_2644,In_3338);
or U4628 (N_4628,In_1040,In_3673);
nor U4629 (N_4629,In_3415,In_728);
nand U4630 (N_4630,In_1174,In_1730);
or U4631 (N_4631,In_4512,In_1886);
nor U4632 (N_4632,In_2245,In_1666);
xor U4633 (N_4633,In_2941,In_2788);
or U4634 (N_4634,In_4063,In_110);
and U4635 (N_4635,In_360,In_3052);
xnor U4636 (N_4636,In_4493,In_3821);
or U4637 (N_4637,In_4733,In_3151);
xor U4638 (N_4638,In_4068,In_1743);
nand U4639 (N_4639,In_4070,In_1609);
nor U4640 (N_4640,In_3241,In_3833);
nand U4641 (N_4641,In_3774,In_823);
xor U4642 (N_4642,In_485,In_2847);
xnor U4643 (N_4643,In_1563,In_631);
xor U4644 (N_4644,In_4403,In_4366);
and U4645 (N_4645,In_3869,In_54);
and U4646 (N_4646,In_2764,In_3946);
or U4647 (N_4647,In_3649,In_2269);
or U4648 (N_4648,In_3168,In_1272);
or U4649 (N_4649,In_4538,In_1854);
xnor U4650 (N_4650,In_4301,In_2481);
nor U4651 (N_4651,In_4644,In_1077);
nor U4652 (N_4652,In_4794,In_4774);
xnor U4653 (N_4653,In_3827,In_4439);
nand U4654 (N_4654,In_2816,In_4653);
or U4655 (N_4655,In_2280,In_4911);
nor U4656 (N_4656,In_1007,In_352);
xnor U4657 (N_4657,In_1153,In_2663);
and U4658 (N_4658,In_781,In_4521);
nand U4659 (N_4659,In_3659,In_6);
nor U4660 (N_4660,In_816,In_442);
nand U4661 (N_4661,In_635,In_1901);
nor U4662 (N_4662,In_1547,In_282);
nand U4663 (N_4663,In_938,In_803);
nand U4664 (N_4664,In_2824,In_894);
or U4665 (N_4665,In_746,In_3687);
nor U4666 (N_4666,In_2905,In_1031);
nand U4667 (N_4667,In_4518,In_1413);
xnor U4668 (N_4668,In_1327,In_4148);
nand U4669 (N_4669,In_3245,In_653);
or U4670 (N_4670,In_2831,In_3254);
and U4671 (N_4671,In_1514,In_1264);
and U4672 (N_4672,In_2206,In_2593);
or U4673 (N_4673,In_1472,In_4690);
nor U4674 (N_4674,In_4545,In_514);
nor U4675 (N_4675,In_4841,In_2470);
nor U4676 (N_4676,In_4798,In_2902);
xnor U4677 (N_4677,In_4014,In_4937);
or U4678 (N_4678,In_4335,In_4958);
and U4679 (N_4679,In_2838,In_2977);
or U4680 (N_4680,In_860,In_4332);
xor U4681 (N_4681,In_2553,In_4352);
nand U4682 (N_4682,In_1094,In_1712);
nand U4683 (N_4683,In_2572,In_1072);
or U4684 (N_4684,In_1685,In_2152);
nor U4685 (N_4685,In_1455,In_3012);
nand U4686 (N_4686,In_3910,In_2930);
xor U4687 (N_4687,In_2398,In_2222);
or U4688 (N_4688,In_3866,In_172);
or U4689 (N_4689,In_1338,In_1114);
nor U4690 (N_4690,In_3005,In_598);
nor U4691 (N_4691,In_2614,In_3170);
and U4692 (N_4692,In_4455,In_1611);
xor U4693 (N_4693,In_4037,In_3514);
nand U4694 (N_4694,In_3722,In_2509);
nor U4695 (N_4695,In_1928,In_807);
nor U4696 (N_4696,In_3355,In_2048);
nor U4697 (N_4697,In_1513,In_2516);
xor U4698 (N_4698,In_612,In_1597);
and U4699 (N_4699,In_3697,In_1240);
xnor U4700 (N_4700,In_775,In_2325);
xnor U4701 (N_4701,In_2973,In_2584);
and U4702 (N_4702,In_3741,In_353);
nor U4703 (N_4703,In_3812,In_2390);
or U4704 (N_4704,In_3951,In_1932);
xnor U4705 (N_4705,In_1726,In_4673);
nand U4706 (N_4706,In_4567,In_2233);
and U4707 (N_4707,In_893,In_2119);
nand U4708 (N_4708,In_3281,In_2386);
nor U4709 (N_4709,In_1775,In_3388);
xor U4710 (N_4710,In_2520,In_1074);
xnor U4711 (N_4711,In_3841,In_2996);
xor U4712 (N_4712,In_2520,In_2653);
xor U4713 (N_4713,In_4983,In_4294);
nand U4714 (N_4714,In_1254,In_2284);
nand U4715 (N_4715,In_2487,In_3634);
or U4716 (N_4716,In_155,In_2356);
or U4717 (N_4717,In_2323,In_2223);
nand U4718 (N_4718,In_1473,In_4050);
nor U4719 (N_4719,In_4907,In_4706);
xnor U4720 (N_4720,In_1480,In_1593);
xnor U4721 (N_4721,In_3496,In_3959);
nor U4722 (N_4722,In_3004,In_4463);
nand U4723 (N_4723,In_4965,In_2743);
and U4724 (N_4724,In_1465,In_2712);
or U4725 (N_4725,In_2943,In_4948);
and U4726 (N_4726,In_1886,In_1312);
and U4727 (N_4727,In_2379,In_2891);
nand U4728 (N_4728,In_4556,In_3886);
and U4729 (N_4729,In_4405,In_1031);
nor U4730 (N_4730,In_782,In_2188);
nor U4731 (N_4731,In_401,In_3744);
xnor U4732 (N_4732,In_1640,In_2271);
or U4733 (N_4733,In_3049,In_3804);
and U4734 (N_4734,In_1885,In_3212);
nor U4735 (N_4735,In_3105,In_3346);
nand U4736 (N_4736,In_185,In_1369);
and U4737 (N_4737,In_2013,In_1000);
or U4738 (N_4738,In_2864,In_4135);
nor U4739 (N_4739,In_4053,In_4563);
and U4740 (N_4740,In_4539,In_381);
xnor U4741 (N_4741,In_3120,In_3923);
and U4742 (N_4742,In_4431,In_334);
or U4743 (N_4743,In_3038,In_2048);
and U4744 (N_4744,In_1297,In_2696);
nor U4745 (N_4745,In_1253,In_4543);
nor U4746 (N_4746,In_3526,In_2272);
xor U4747 (N_4747,In_2260,In_751);
or U4748 (N_4748,In_875,In_3278);
and U4749 (N_4749,In_1152,In_1941);
nor U4750 (N_4750,In_3788,In_4697);
nor U4751 (N_4751,In_1562,In_2304);
or U4752 (N_4752,In_3342,In_1899);
or U4753 (N_4753,In_1119,In_475);
or U4754 (N_4754,In_4921,In_2062);
nor U4755 (N_4755,In_4606,In_4156);
and U4756 (N_4756,In_2495,In_2291);
or U4757 (N_4757,In_3489,In_2656);
xor U4758 (N_4758,In_4109,In_379);
xor U4759 (N_4759,In_3086,In_2324);
and U4760 (N_4760,In_3395,In_25);
or U4761 (N_4761,In_1297,In_924);
nor U4762 (N_4762,In_4037,In_3871);
nor U4763 (N_4763,In_1379,In_150);
xor U4764 (N_4764,In_844,In_2454);
nor U4765 (N_4765,In_2470,In_4700);
xor U4766 (N_4766,In_927,In_112);
or U4767 (N_4767,In_4380,In_2772);
nor U4768 (N_4768,In_2324,In_1702);
and U4769 (N_4769,In_4659,In_2239);
nor U4770 (N_4770,In_290,In_4894);
or U4771 (N_4771,In_4194,In_3412);
nor U4772 (N_4772,In_1411,In_1002);
and U4773 (N_4773,In_2946,In_2420);
xor U4774 (N_4774,In_2646,In_22);
nor U4775 (N_4775,In_527,In_4412);
and U4776 (N_4776,In_3801,In_3419);
xnor U4777 (N_4777,In_4124,In_1656);
and U4778 (N_4778,In_213,In_4498);
and U4779 (N_4779,In_459,In_4413);
or U4780 (N_4780,In_755,In_840);
or U4781 (N_4781,In_1029,In_1580);
xor U4782 (N_4782,In_1076,In_280);
and U4783 (N_4783,In_4340,In_2368);
nand U4784 (N_4784,In_597,In_4268);
or U4785 (N_4785,In_4280,In_978);
nor U4786 (N_4786,In_3066,In_1448);
and U4787 (N_4787,In_763,In_2912);
nor U4788 (N_4788,In_3962,In_748);
or U4789 (N_4789,In_539,In_684);
nor U4790 (N_4790,In_2438,In_1440);
or U4791 (N_4791,In_3247,In_2486);
nand U4792 (N_4792,In_1819,In_3132);
or U4793 (N_4793,In_714,In_4229);
and U4794 (N_4794,In_1186,In_2203);
nor U4795 (N_4795,In_525,In_3515);
and U4796 (N_4796,In_4818,In_3485);
nand U4797 (N_4797,In_3048,In_3683);
or U4798 (N_4798,In_1674,In_2261);
nor U4799 (N_4799,In_2464,In_1360);
nand U4800 (N_4800,In_1273,In_2547);
xnor U4801 (N_4801,In_2933,In_141);
nor U4802 (N_4802,In_2061,In_1092);
and U4803 (N_4803,In_19,In_2463);
xor U4804 (N_4804,In_4881,In_3244);
xnor U4805 (N_4805,In_30,In_2093);
nand U4806 (N_4806,In_416,In_229);
nor U4807 (N_4807,In_4753,In_4491);
and U4808 (N_4808,In_1227,In_3902);
nand U4809 (N_4809,In_197,In_847);
and U4810 (N_4810,In_43,In_4589);
and U4811 (N_4811,In_255,In_1884);
xor U4812 (N_4812,In_4018,In_3186);
xnor U4813 (N_4813,In_777,In_3431);
and U4814 (N_4814,In_3740,In_1766);
or U4815 (N_4815,In_1192,In_2521);
xnor U4816 (N_4816,In_1907,In_4056);
or U4817 (N_4817,In_1325,In_3248);
or U4818 (N_4818,In_1757,In_4654);
and U4819 (N_4819,In_3135,In_1219);
nor U4820 (N_4820,In_4160,In_1015);
xnor U4821 (N_4821,In_3902,In_596);
and U4822 (N_4822,In_3663,In_1631);
nor U4823 (N_4823,In_4392,In_4079);
and U4824 (N_4824,In_1204,In_3371);
nor U4825 (N_4825,In_2456,In_368);
nand U4826 (N_4826,In_4097,In_4807);
and U4827 (N_4827,In_3973,In_3722);
and U4828 (N_4828,In_2458,In_373);
and U4829 (N_4829,In_216,In_4206);
and U4830 (N_4830,In_1279,In_2705);
xnor U4831 (N_4831,In_852,In_3069);
xor U4832 (N_4832,In_8,In_732);
xnor U4833 (N_4833,In_3064,In_1525);
nand U4834 (N_4834,In_2889,In_4742);
or U4835 (N_4835,In_1132,In_103);
xnor U4836 (N_4836,In_1749,In_3188);
nand U4837 (N_4837,In_2934,In_4840);
nand U4838 (N_4838,In_1584,In_4902);
nand U4839 (N_4839,In_2970,In_265);
nand U4840 (N_4840,In_2995,In_741);
and U4841 (N_4841,In_4412,In_4498);
or U4842 (N_4842,In_4191,In_892);
and U4843 (N_4843,In_3934,In_79);
nor U4844 (N_4844,In_4977,In_2259);
and U4845 (N_4845,In_3015,In_4949);
nor U4846 (N_4846,In_2612,In_4027);
nor U4847 (N_4847,In_4993,In_3640);
xor U4848 (N_4848,In_4868,In_952);
and U4849 (N_4849,In_4552,In_3698);
and U4850 (N_4850,In_1471,In_126);
nand U4851 (N_4851,In_4074,In_2336);
nor U4852 (N_4852,In_4889,In_2092);
and U4853 (N_4853,In_1372,In_2945);
xnor U4854 (N_4854,In_3001,In_23);
xnor U4855 (N_4855,In_3845,In_691);
nor U4856 (N_4856,In_2096,In_3809);
xor U4857 (N_4857,In_3547,In_2646);
nand U4858 (N_4858,In_3035,In_2831);
and U4859 (N_4859,In_4900,In_4057);
nand U4860 (N_4860,In_1889,In_3114);
xor U4861 (N_4861,In_4035,In_335);
xor U4862 (N_4862,In_3737,In_3097);
nand U4863 (N_4863,In_492,In_834);
or U4864 (N_4864,In_1299,In_2670);
xor U4865 (N_4865,In_852,In_1309);
or U4866 (N_4866,In_1076,In_1756);
nor U4867 (N_4867,In_4972,In_1692);
xnor U4868 (N_4868,In_658,In_2390);
and U4869 (N_4869,In_4208,In_709);
nor U4870 (N_4870,In_1749,In_1188);
xor U4871 (N_4871,In_471,In_3190);
xor U4872 (N_4872,In_1985,In_2689);
and U4873 (N_4873,In_529,In_3023);
or U4874 (N_4874,In_3181,In_1250);
or U4875 (N_4875,In_4405,In_3655);
nand U4876 (N_4876,In_3774,In_470);
xnor U4877 (N_4877,In_3420,In_4416);
nand U4878 (N_4878,In_2342,In_2288);
nand U4879 (N_4879,In_305,In_31);
or U4880 (N_4880,In_842,In_760);
xnor U4881 (N_4881,In_4389,In_129);
xor U4882 (N_4882,In_1539,In_2926);
and U4883 (N_4883,In_4012,In_2675);
xnor U4884 (N_4884,In_3312,In_2070);
nor U4885 (N_4885,In_2269,In_3482);
or U4886 (N_4886,In_4382,In_4759);
nor U4887 (N_4887,In_350,In_1696);
and U4888 (N_4888,In_2554,In_4032);
or U4889 (N_4889,In_914,In_2703);
or U4890 (N_4890,In_121,In_3128);
nor U4891 (N_4891,In_1525,In_3741);
xor U4892 (N_4892,In_248,In_1772);
nor U4893 (N_4893,In_1194,In_3305);
nand U4894 (N_4894,In_3847,In_3848);
nand U4895 (N_4895,In_3312,In_3219);
or U4896 (N_4896,In_1840,In_1535);
or U4897 (N_4897,In_4947,In_3801);
nor U4898 (N_4898,In_290,In_525);
and U4899 (N_4899,In_3335,In_4376);
xor U4900 (N_4900,In_3668,In_4764);
xnor U4901 (N_4901,In_3082,In_3285);
or U4902 (N_4902,In_510,In_4018);
nor U4903 (N_4903,In_1608,In_322);
nand U4904 (N_4904,In_3755,In_4432);
xnor U4905 (N_4905,In_1567,In_405);
or U4906 (N_4906,In_4806,In_3785);
and U4907 (N_4907,In_187,In_3126);
xor U4908 (N_4908,In_3427,In_1919);
xnor U4909 (N_4909,In_1829,In_2322);
nor U4910 (N_4910,In_3366,In_3735);
and U4911 (N_4911,In_3458,In_3363);
and U4912 (N_4912,In_4460,In_794);
xnor U4913 (N_4913,In_322,In_4421);
nor U4914 (N_4914,In_4925,In_2562);
and U4915 (N_4915,In_4921,In_2582);
xor U4916 (N_4916,In_1857,In_630);
or U4917 (N_4917,In_3432,In_3078);
or U4918 (N_4918,In_458,In_4552);
xnor U4919 (N_4919,In_4284,In_2089);
nor U4920 (N_4920,In_1227,In_4602);
or U4921 (N_4921,In_4758,In_4539);
and U4922 (N_4922,In_2811,In_645);
or U4923 (N_4923,In_4394,In_908);
or U4924 (N_4924,In_4096,In_417);
nand U4925 (N_4925,In_1858,In_4956);
xnor U4926 (N_4926,In_3111,In_736);
xor U4927 (N_4927,In_1066,In_3405);
and U4928 (N_4928,In_4869,In_3261);
nor U4929 (N_4929,In_3189,In_4759);
nor U4930 (N_4930,In_2792,In_3415);
nor U4931 (N_4931,In_1160,In_2104);
and U4932 (N_4932,In_1879,In_4361);
and U4933 (N_4933,In_3972,In_2655);
nor U4934 (N_4934,In_4468,In_4455);
or U4935 (N_4935,In_225,In_3252);
nor U4936 (N_4936,In_3747,In_460);
nand U4937 (N_4937,In_3935,In_3002);
or U4938 (N_4938,In_4257,In_3153);
xnor U4939 (N_4939,In_2252,In_571);
and U4940 (N_4940,In_1860,In_1493);
nand U4941 (N_4941,In_835,In_3978);
nand U4942 (N_4942,In_695,In_2020);
or U4943 (N_4943,In_39,In_4377);
nand U4944 (N_4944,In_4542,In_760);
and U4945 (N_4945,In_1937,In_1547);
and U4946 (N_4946,In_4790,In_250);
xor U4947 (N_4947,In_4715,In_1533);
and U4948 (N_4948,In_2912,In_3544);
nor U4949 (N_4949,In_500,In_539);
nand U4950 (N_4950,In_4155,In_605);
or U4951 (N_4951,In_3412,In_4705);
nand U4952 (N_4952,In_4487,In_1207);
and U4953 (N_4953,In_2166,In_1062);
nand U4954 (N_4954,In_2459,In_3537);
or U4955 (N_4955,In_4483,In_4133);
or U4956 (N_4956,In_4444,In_1875);
and U4957 (N_4957,In_500,In_327);
nor U4958 (N_4958,In_2355,In_2288);
and U4959 (N_4959,In_1260,In_463);
xnor U4960 (N_4960,In_945,In_3287);
and U4961 (N_4961,In_4626,In_831);
or U4962 (N_4962,In_1809,In_4285);
or U4963 (N_4963,In_1871,In_3301);
or U4964 (N_4964,In_2324,In_3177);
nor U4965 (N_4965,In_2226,In_824);
xor U4966 (N_4966,In_3062,In_439);
nand U4967 (N_4967,In_3056,In_127);
and U4968 (N_4968,In_4417,In_1467);
and U4969 (N_4969,In_899,In_296);
nor U4970 (N_4970,In_1471,In_2181);
nand U4971 (N_4971,In_4990,In_4729);
nand U4972 (N_4972,In_333,In_2529);
nand U4973 (N_4973,In_3225,In_2119);
nand U4974 (N_4974,In_2477,In_635);
and U4975 (N_4975,In_3973,In_683);
nor U4976 (N_4976,In_1261,In_310);
nor U4977 (N_4977,In_3859,In_880);
and U4978 (N_4978,In_726,In_3162);
and U4979 (N_4979,In_1992,In_1094);
xnor U4980 (N_4980,In_1411,In_2313);
nand U4981 (N_4981,In_1654,In_537);
and U4982 (N_4982,In_2317,In_1618);
nand U4983 (N_4983,In_2159,In_1066);
and U4984 (N_4984,In_492,In_3776);
nand U4985 (N_4985,In_1751,In_101);
or U4986 (N_4986,In_2702,In_1991);
xor U4987 (N_4987,In_3506,In_2338);
xnor U4988 (N_4988,In_2339,In_3455);
and U4989 (N_4989,In_4372,In_2765);
xor U4990 (N_4990,In_387,In_4384);
or U4991 (N_4991,In_1959,In_1453);
nor U4992 (N_4992,In_2392,In_1853);
or U4993 (N_4993,In_2033,In_945);
xnor U4994 (N_4994,In_1654,In_124);
or U4995 (N_4995,In_1447,In_3678);
nor U4996 (N_4996,In_2399,In_1204);
or U4997 (N_4997,In_3208,In_4934);
nand U4998 (N_4998,In_3629,In_3393);
or U4999 (N_4999,In_3619,In_3820);
and U5000 (N_5000,N_1771,N_3919);
xnor U5001 (N_5001,N_875,N_188);
nor U5002 (N_5002,N_2422,N_4370);
and U5003 (N_5003,N_991,N_4088);
xnor U5004 (N_5004,N_1298,N_3097);
nand U5005 (N_5005,N_229,N_4933);
or U5006 (N_5006,N_1330,N_3020);
xnor U5007 (N_5007,N_909,N_2418);
nor U5008 (N_5008,N_1648,N_778);
nor U5009 (N_5009,N_3987,N_3714);
or U5010 (N_5010,N_2297,N_3180);
and U5011 (N_5011,N_418,N_4753);
and U5012 (N_5012,N_4608,N_4747);
and U5013 (N_5013,N_9,N_2638);
nor U5014 (N_5014,N_1905,N_3659);
nand U5015 (N_5015,N_3776,N_956);
nand U5016 (N_5016,N_3536,N_2936);
nand U5017 (N_5017,N_1015,N_1937);
nand U5018 (N_5018,N_2487,N_3938);
nand U5019 (N_5019,N_2261,N_819);
nor U5020 (N_5020,N_444,N_466);
nor U5021 (N_5021,N_628,N_1312);
or U5022 (N_5022,N_4401,N_103);
nand U5023 (N_5023,N_1918,N_1406);
and U5024 (N_5024,N_1521,N_929);
and U5025 (N_5025,N_1802,N_234);
or U5026 (N_5026,N_3770,N_3062);
or U5027 (N_5027,N_1269,N_2636);
and U5028 (N_5028,N_36,N_893);
xnor U5029 (N_5029,N_4552,N_2732);
nor U5030 (N_5030,N_1014,N_205);
nand U5031 (N_5031,N_3881,N_1026);
nand U5032 (N_5032,N_1795,N_1819);
or U5033 (N_5033,N_3174,N_2416);
nand U5034 (N_5034,N_2104,N_3578);
nand U5035 (N_5035,N_2408,N_3069);
or U5036 (N_5036,N_3668,N_4635);
or U5037 (N_5037,N_4331,N_3329);
nand U5038 (N_5038,N_2207,N_4882);
xnor U5039 (N_5039,N_517,N_2913);
xnor U5040 (N_5040,N_4542,N_1793);
nand U5041 (N_5041,N_3205,N_2459);
and U5042 (N_5042,N_2172,N_2330);
or U5043 (N_5043,N_3417,N_4839);
nand U5044 (N_5044,N_2637,N_4354);
and U5045 (N_5045,N_1071,N_3311);
nor U5046 (N_5046,N_3043,N_242);
xor U5047 (N_5047,N_3628,N_1168);
nand U5048 (N_5048,N_2568,N_2042);
nand U5049 (N_5049,N_691,N_195);
nand U5050 (N_5050,N_2316,N_2489);
and U5051 (N_5051,N_2883,N_368);
xnor U5052 (N_5052,N_1579,N_2824);
nor U5053 (N_5053,N_4550,N_855);
nor U5054 (N_5054,N_2731,N_4588);
xor U5055 (N_5055,N_2255,N_808);
or U5056 (N_5056,N_2246,N_3806);
nor U5057 (N_5057,N_112,N_4132);
xnor U5058 (N_5058,N_2524,N_3240);
xor U5059 (N_5059,N_1753,N_3051);
or U5060 (N_5060,N_3252,N_4150);
nor U5061 (N_5061,N_2492,N_2988);
or U5062 (N_5062,N_2480,N_1779);
nand U5063 (N_5063,N_1765,N_4901);
nand U5064 (N_5064,N_1293,N_52);
or U5065 (N_5065,N_3980,N_4572);
or U5066 (N_5066,N_3907,N_3200);
nor U5067 (N_5067,N_3842,N_1173);
xnor U5068 (N_5068,N_212,N_178);
nor U5069 (N_5069,N_1083,N_1124);
xor U5070 (N_5070,N_3281,N_2598);
xnor U5071 (N_5071,N_1759,N_3670);
nand U5072 (N_5072,N_4907,N_256);
or U5073 (N_5073,N_4970,N_3528);
nor U5074 (N_5074,N_115,N_1136);
nand U5075 (N_5075,N_568,N_1824);
or U5076 (N_5076,N_3272,N_1361);
xor U5077 (N_5077,N_3588,N_4272);
and U5078 (N_5078,N_2143,N_3331);
or U5079 (N_5079,N_4186,N_4081);
and U5080 (N_5080,N_4028,N_1678);
or U5081 (N_5081,N_3944,N_1376);
xor U5082 (N_5082,N_454,N_796);
and U5083 (N_5083,N_4214,N_4064);
nand U5084 (N_5084,N_2135,N_4738);
nand U5085 (N_5085,N_4978,N_398);
nor U5086 (N_5086,N_1481,N_1319);
or U5087 (N_5087,N_251,N_2682);
and U5088 (N_5088,N_233,N_4265);
and U5089 (N_5089,N_3832,N_1776);
xnor U5090 (N_5090,N_3928,N_385);
nor U5091 (N_5091,N_1559,N_4743);
or U5092 (N_5092,N_19,N_138);
xor U5093 (N_5093,N_2550,N_1955);
nand U5094 (N_5094,N_1531,N_4498);
nor U5095 (N_5095,N_4180,N_3756);
xnor U5096 (N_5096,N_270,N_4380);
nand U5097 (N_5097,N_2192,N_1954);
and U5098 (N_5098,N_709,N_1249);
nor U5099 (N_5099,N_3170,N_2890);
or U5100 (N_5100,N_4304,N_4042);
or U5101 (N_5101,N_349,N_2663);
and U5102 (N_5102,N_63,N_2496);
nor U5103 (N_5103,N_4590,N_2968);
or U5104 (N_5104,N_4493,N_3204);
nor U5105 (N_5105,N_4917,N_1630);
nor U5106 (N_5106,N_2806,N_3103);
xnor U5107 (N_5107,N_2558,N_4709);
nand U5108 (N_5108,N_3593,N_551);
xor U5109 (N_5109,N_3385,N_2937);
nor U5110 (N_5110,N_2884,N_872);
and U5111 (N_5111,N_2033,N_4696);
or U5112 (N_5112,N_4843,N_4564);
xor U5113 (N_5113,N_2364,N_213);
xnor U5114 (N_5114,N_2193,N_2784);
or U5115 (N_5115,N_23,N_2775);
and U5116 (N_5116,N_4545,N_3924);
xnor U5117 (N_5117,N_4622,N_859);
nand U5118 (N_5118,N_1898,N_4189);
xnor U5119 (N_5119,N_2363,N_4688);
and U5120 (N_5120,N_155,N_4016);
and U5121 (N_5121,N_1513,N_4101);
xnor U5122 (N_5122,N_3219,N_2191);
xnor U5123 (N_5123,N_2914,N_3558);
nor U5124 (N_5124,N_140,N_3638);
nor U5125 (N_5125,N_743,N_2012);
and U5126 (N_5126,N_146,N_1394);
or U5127 (N_5127,N_76,N_1030);
nor U5128 (N_5128,N_3175,N_1257);
nand U5129 (N_5129,N_4321,N_2082);
nand U5130 (N_5130,N_2978,N_4513);
xnor U5131 (N_5131,N_1138,N_1037);
xor U5132 (N_5132,N_3126,N_1960);
nand U5133 (N_5133,N_2702,N_3468);
nand U5134 (N_5134,N_3306,N_3683);
and U5135 (N_5135,N_4202,N_2867);
nand U5136 (N_5136,N_489,N_3887);
nand U5137 (N_5137,N_3786,N_457);
nor U5138 (N_5138,N_2287,N_1265);
xnor U5139 (N_5139,N_3132,N_4068);
xnor U5140 (N_5140,N_2462,N_4296);
nand U5141 (N_5141,N_3393,N_3239);
xnor U5142 (N_5142,N_373,N_4115);
nor U5143 (N_5143,N_2960,N_2752);
xor U5144 (N_5144,N_4934,N_2774);
xor U5145 (N_5145,N_4117,N_1963);
or U5146 (N_5146,N_3816,N_32);
xor U5147 (N_5147,N_3811,N_3474);
or U5148 (N_5148,N_2751,N_1130);
nand U5149 (N_5149,N_2923,N_1000);
nor U5150 (N_5150,N_2281,N_235);
nor U5151 (N_5151,N_1214,N_3493);
nand U5152 (N_5152,N_4636,N_4899);
xor U5153 (N_5153,N_1402,N_2705);
nand U5154 (N_5154,N_571,N_2121);
nor U5155 (N_5155,N_2861,N_2763);
xnor U5156 (N_5156,N_4480,N_3241);
and U5157 (N_5157,N_3696,N_815);
nand U5158 (N_5158,N_3686,N_3420);
nand U5159 (N_5159,N_399,N_4277);
nor U5160 (N_5160,N_1268,N_2669);
nand U5161 (N_5161,N_2668,N_2372);
nand U5162 (N_5162,N_2974,N_1749);
nand U5163 (N_5163,N_4430,N_1989);
nand U5164 (N_5164,N_1271,N_608);
nand U5165 (N_5165,N_3015,N_210);
nor U5166 (N_5166,N_3692,N_3017);
nand U5167 (N_5167,N_4518,N_2110);
xor U5168 (N_5168,N_3632,N_4848);
or U5169 (N_5169,N_3287,N_1877);
or U5170 (N_5170,N_4928,N_3922);
and U5171 (N_5171,N_972,N_1238);
nor U5172 (N_5172,N_3517,N_1606);
nand U5173 (N_5173,N_2595,N_1456);
or U5174 (N_5174,N_2223,N_2176);
or U5175 (N_5175,N_4908,N_1573);
nor U5176 (N_5176,N_4144,N_1430);
nand U5177 (N_5177,N_166,N_1808);
nor U5178 (N_5178,N_4911,N_2684);
nor U5179 (N_5179,N_2235,N_4662);
or U5180 (N_5180,N_1529,N_2106);
or U5181 (N_5181,N_1517,N_4558);
nor U5182 (N_5182,N_1099,N_1964);
or U5183 (N_5183,N_2819,N_3809);
and U5184 (N_5184,N_3934,N_72);
nand U5185 (N_5185,N_3551,N_354);
and U5186 (N_5186,N_4192,N_591);
nor U5187 (N_5187,N_326,N_2551);
and U5188 (N_5188,N_3077,N_1499);
nor U5189 (N_5189,N_330,N_684);
nor U5190 (N_5190,N_2917,N_3253);
or U5191 (N_5191,N_3815,N_537);
or U5192 (N_5192,N_2412,N_1936);
xnor U5193 (N_5193,N_4685,N_1328);
and U5194 (N_5194,N_4773,N_423);
xnor U5195 (N_5195,N_1869,N_4121);
xor U5196 (N_5196,N_1763,N_3102);
and U5197 (N_5197,N_2066,N_3572);
nor U5198 (N_5198,N_2383,N_3118);
or U5199 (N_5199,N_3926,N_254);
or U5200 (N_5200,N_1151,N_107);
xnor U5201 (N_5201,N_1798,N_1429);
xor U5202 (N_5202,N_1073,N_3391);
xnor U5203 (N_5203,N_2538,N_4829);
xnor U5204 (N_5204,N_4656,N_4168);
and U5205 (N_5205,N_891,N_4169);
nor U5206 (N_5206,N_2304,N_4642);
and U5207 (N_5207,N_4789,N_1595);
or U5208 (N_5208,N_3633,N_455);
nor U5209 (N_5209,N_4898,N_669);
or U5210 (N_5210,N_586,N_2864);
xnor U5211 (N_5211,N_400,N_4626);
and U5212 (N_5212,N_87,N_3247);
or U5213 (N_5213,N_3750,N_3500);
nor U5214 (N_5214,N_1641,N_4505);
nor U5215 (N_5215,N_2366,N_4851);
nor U5216 (N_5216,N_2660,N_3554);
nor U5217 (N_5217,N_2655,N_3024);
nand U5218 (N_5218,N_3847,N_805);
or U5219 (N_5219,N_1618,N_4867);
and U5220 (N_5220,N_827,N_3257);
and U5221 (N_5221,N_2738,N_4066);
xor U5222 (N_5222,N_2132,N_3605);
and U5223 (N_5223,N_777,N_3462);
nand U5224 (N_5224,N_1666,N_2181);
xor U5225 (N_5225,N_4262,N_3469);
nand U5226 (N_5226,N_1993,N_4301);
or U5227 (N_5227,N_1598,N_3758);
nand U5228 (N_5228,N_3330,N_1346);
or U5229 (N_5229,N_3580,N_4473);
nand U5230 (N_5230,N_696,N_2471);
nor U5231 (N_5231,N_2685,N_1719);
and U5232 (N_5232,N_2486,N_4963);
nand U5233 (N_5233,N_4457,N_3206);
xnor U5234 (N_5234,N_1305,N_3216);
or U5235 (N_5235,N_611,N_1734);
and U5236 (N_5236,N_1029,N_1275);
nand U5237 (N_5237,N_3761,N_262);
nor U5238 (N_5238,N_1290,N_2482);
and U5239 (N_5239,N_550,N_468);
xor U5240 (N_5240,N_1196,N_4417);
and U5241 (N_5241,N_2761,N_1075);
or U5242 (N_5242,N_1100,N_2163);
nor U5243 (N_5243,N_2177,N_981);
nand U5244 (N_5244,N_1757,N_1823);
nand U5245 (N_5245,N_1875,N_4669);
xor U5246 (N_5246,N_862,N_480);
and U5247 (N_5247,N_3989,N_4313);
nor U5248 (N_5248,N_2182,N_222);
nand U5249 (N_5249,N_887,N_297);
nor U5250 (N_5250,N_4159,N_3261);
or U5251 (N_5251,N_1803,N_1581);
nand U5252 (N_5252,N_534,N_2530);
nand U5253 (N_5253,N_3590,N_3121);
and U5254 (N_5254,N_1236,N_3155);
and U5255 (N_5255,N_4534,N_157);
nor U5256 (N_5256,N_1737,N_3752);
nor U5257 (N_5257,N_4004,N_4008);
nand U5258 (N_5258,N_4673,N_3600);
nand U5259 (N_5259,N_1863,N_4061);
nand U5260 (N_5260,N_704,N_1609);
xor U5261 (N_5261,N_3160,N_4694);
xor U5262 (N_5262,N_1174,N_720);
or U5263 (N_5263,N_4295,N_3757);
and U5264 (N_5264,N_3158,N_1644);
nand U5265 (N_5265,N_976,N_4665);
xnor U5266 (N_5266,N_477,N_4187);
xor U5267 (N_5267,N_1384,N_3697);
nor U5268 (N_5268,N_3250,N_4085);
and U5269 (N_5269,N_2903,N_375);
xor U5270 (N_5270,N_3603,N_3728);
nand U5271 (N_5271,N_2696,N_3610);
nor U5272 (N_5272,N_4631,N_1280);
xnor U5273 (N_5273,N_2034,N_4952);
or U5274 (N_5274,N_3969,N_4616);
and U5275 (N_5275,N_869,N_2577);
xnor U5276 (N_5276,N_177,N_3125);
nand U5277 (N_5277,N_4757,N_1629);
nand U5278 (N_5278,N_3315,N_4543);
or U5279 (N_5279,N_800,N_2724);
nor U5280 (N_5280,N_1398,N_4739);
or U5281 (N_5281,N_2814,N_3111);
nand U5282 (N_5282,N_3716,N_782);
nand U5283 (N_5283,N_2590,N_3258);
or U5284 (N_5284,N_3585,N_4357);
xnor U5285 (N_5285,N_857,N_2718);
or U5286 (N_5286,N_3013,N_1575);
xnor U5287 (N_5287,N_1811,N_207);
nand U5288 (N_5288,N_3695,N_3361);
xor U5289 (N_5289,N_2678,N_126);
xor U5290 (N_5290,N_3073,N_3357);
nand U5291 (N_5291,N_1334,N_3779);
and U5292 (N_5292,N_4499,N_1534);
nor U5293 (N_5293,N_1544,N_106);
nor U5294 (N_5294,N_2020,N_657);
or U5295 (N_5295,N_2885,N_2714);
and U5296 (N_5296,N_3983,N_2527);
nor U5297 (N_5297,N_4352,N_4976);
xor U5298 (N_5298,N_2664,N_2274);
or U5299 (N_5299,N_498,N_4387);
or U5300 (N_5300,N_2057,N_593);
or U5301 (N_5301,N_2321,N_2510);
or U5302 (N_5302,N_749,N_1580);
xnor U5303 (N_5303,N_2679,N_201);
or U5304 (N_5304,N_578,N_3727);
and U5305 (N_5305,N_1087,N_1885);
or U5306 (N_5306,N_163,N_273);
nor U5307 (N_5307,N_930,N_836);
nor U5308 (N_5308,N_1184,N_728);
or U5309 (N_5309,N_2634,N_2841);
nor U5310 (N_5310,N_4926,N_3165);
and U5311 (N_5311,N_695,N_1682);
and U5312 (N_5312,N_4078,N_4177);
or U5313 (N_5313,N_3228,N_727);
nand U5314 (N_5314,N_2945,N_2098);
nand U5315 (N_5315,N_1395,N_1343);
nor U5316 (N_5316,N_2107,N_459);
nor U5317 (N_5317,N_4835,N_3507);
xnor U5318 (N_5318,N_3461,N_1426);
and U5319 (N_5319,N_48,N_4200);
and U5320 (N_5320,N_4120,N_2357);
nand U5321 (N_5321,N_1274,N_2210);
nand U5322 (N_5322,N_2313,N_4967);
nor U5323 (N_5323,N_573,N_221);
nor U5324 (N_5324,N_154,N_3355);
or U5325 (N_5325,N_948,N_773);
xnor U5326 (N_5326,N_760,N_1929);
xor U5327 (N_5327,N_2961,N_4392);
nand U5328 (N_5328,N_4778,N_34);
nor U5329 (N_5329,N_676,N_171);
nand U5330 (N_5330,N_452,N_492);
xor U5331 (N_5331,N_4951,N_785);
xnor U5332 (N_5332,N_253,N_3340);
and U5333 (N_5333,N_3095,N_3753);
and U5334 (N_5334,N_3854,N_4174);
and U5335 (N_5335,N_3196,N_2564);
and U5336 (N_5336,N_89,N_3034);
nand U5337 (N_5337,N_2847,N_886);
or U5338 (N_5338,N_464,N_2710);
nor U5339 (N_5339,N_1225,N_70);
xnor U5340 (N_5340,N_1552,N_1654);
and U5341 (N_5341,N_44,N_2445);
nand U5342 (N_5342,N_2686,N_3777);
or U5343 (N_5343,N_2365,N_4808);
or U5344 (N_5344,N_1339,N_3530);
nor U5345 (N_5345,N_4344,N_864);
or U5346 (N_5346,N_1267,N_2320);
or U5347 (N_5347,N_129,N_3504);
nand U5348 (N_5348,N_342,N_4259);
or U5349 (N_5349,N_580,N_309);
nor U5350 (N_5350,N_2153,N_3424);
xnor U5351 (N_5351,N_4010,N_791);
or U5352 (N_5352,N_4707,N_4258);
nand U5353 (N_5353,N_3181,N_223);
or U5354 (N_5354,N_1953,N_376);
and U5355 (N_5355,N_4030,N_3434);
or U5356 (N_5356,N_833,N_1461);
nand U5357 (N_5357,N_2131,N_1047);
xor U5358 (N_5358,N_1323,N_3033);
nand U5359 (N_5359,N_2901,N_2629);
or U5360 (N_5360,N_3794,N_69);
xnor U5361 (N_5361,N_481,N_2973);
xnor U5362 (N_5362,N_2232,N_3268);
xnor U5363 (N_5363,N_609,N_4591);
nor U5364 (N_5364,N_1601,N_1787);
nand U5365 (N_5365,N_595,N_4675);
and U5366 (N_5366,N_2800,N_2815);
nor U5367 (N_5367,N_2859,N_2842);
or U5368 (N_5368,N_4684,N_1002);
xnor U5369 (N_5369,N_3943,N_4939);
xor U5370 (N_5370,N_3769,N_3350);
nor U5371 (N_5371,N_4825,N_1414);
xor U5372 (N_5372,N_4724,N_130);
and U5373 (N_5373,N_4514,N_4651);
xor U5374 (N_5374,N_3429,N_2954);
nor U5375 (N_5375,N_2713,N_3341);
xor U5376 (N_5376,N_2370,N_3245);
xor U5377 (N_5377,N_2866,N_3886);
nor U5378 (N_5378,N_1012,N_3259);
nor U5379 (N_5379,N_3706,N_2582);
nand U5380 (N_5380,N_671,N_2644);
or U5381 (N_5381,N_3319,N_1976);
xnor U5382 (N_5382,N_1605,N_190);
nand U5383 (N_5383,N_3273,N_732);
or U5384 (N_5384,N_3722,N_473);
or U5385 (N_5385,N_2312,N_964);
nor U5386 (N_5386,N_1519,N_3318);
or U5387 (N_5387,N_4810,N_1175);
and U5388 (N_5388,N_3356,N_3168);
xor U5389 (N_5389,N_2144,N_4657);
xnor U5390 (N_5390,N_364,N_4379);
nor U5391 (N_5391,N_96,N_4198);
xnor U5392 (N_5392,N_4962,N_41);
and U5393 (N_5393,N_3230,N_4912);
nand U5394 (N_5394,N_1696,N_3667);
and U5395 (N_5395,N_4361,N_1566);
xor U5396 (N_5396,N_4220,N_3260);
or U5397 (N_5397,N_420,N_2349);
xnor U5398 (N_5398,N_2491,N_4680);
nand U5399 (N_5399,N_3140,N_4371);
nand U5400 (N_5400,N_4623,N_3251);
or U5401 (N_5401,N_91,N_1471);
xor U5402 (N_5402,N_750,N_3295);
xor U5403 (N_5403,N_2015,N_2028);
or U5404 (N_5404,N_2501,N_2241);
nor U5405 (N_5405,N_2778,N_3263);
and U5406 (N_5406,N_323,N_2848);
nand U5407 (N_5407,N_4408,N_1279);
nor U5408 (N_5408,N_1235,N_54);
xnor U5409 (N_5409,N_2301,N_3618);
nand U5410 (N_5410,N_2173,N_3332);
xnor U5411 (N_5411,N_3211,N_4815);
and U5412 (N_5412,N_4666,N_2151);
xor U5413 (N_5413,N_2683,N_1388);
and U5414 (N_5414,N_892,N_3787);
or U5415 (N_5415,N_1739,N_1549);
nand U5416 (N_5416,N_652,N_3105);
nand U5417 (N_5417,N_3370,N_831);
or U5418 (N_5418,N_1736,N_2230);
xor U5419 (N_5419,N_2100,N_822);
or U5420 (N_5420,N_1234,N_3972);
xor U5421 (N_5421,N_3209,N_474);
and U5422 (N_5422,N_4698,N_1986);
nor U5423 (N_5423,N_2242,N_799);
nor U5424 (N_5424,N_61,N_2058);
and U5425 (N_5425,N_2803,N_896);
nand U5426 (N_5426,N_4640,N_81);
nor U5427 (N_5427,N_2935,N_4178);
xor U5428 (N_5428,N_1464,N_4960);
nor U5429 (N_5429,N_2873,N_1747);
nand U5430 (N_5430,N_4628,N_4625);
xor U5431 (N_5431,N_110,N_1935);
or U5432 (N_5432,N_3369,N_3129);
xor U5433 (N_5433,N_2495,N_2675);
or U5434 (N_5434,N_3030,N_4569);
nand U5435 (N_5435,N_2839,N_2105);
and U5436 (N_5436,N_532,N_2265);
and U5437 (N_5437,N_963,N_3120);
xnor U5438 (N_5438,N_1387,N_1418);
nor U5439 (N_5439,N_172,N_2055);
and U5440 (N_5440,N_4025,N_2017);
nand U5441 (N_5441,N_2562,N_2161);
nor U5442 (N_5442,N_1326,N_4598);
nand U5443 (N_5443,N_411,N_2025);
or U5444 (N_5444,N_1299,N_2236);
and U5445 (N_5445,N_248,N_3741);
and U5446 (N_5446,N_2248,N_456);
nand U5447 (N_5447,N_638,N_3755);
and U5448 (N_5448,N_2478,N_4799);
xor U5449 (N_5449,N_3547,N_4054);
nand U5450 (N_5450,N_4497,N_3669);
xnor U5451 (N_5451,N_4268,N_2249);
and U5452 (N_5452,N_4209,N_2918);
nor U5453 (N_5453,N_3560,N_3465);
nor U5454 (N_5454,N_4643,N_3231);
xnor U5455 (N_5455,N_2203,N_4393);
xnor U5456 (N_5456,N_3471,N_28);
and U5457 (N_5457,N_1220,N_3297);
and U5458 (N_5458,N_2219,N_1347);
nand U5459 (N_5459,N_3436,N_4073);
xnor U5460 (N_5460,N_565,N_1480);
and U5461 (N_5461,N_243,N_581);
nor U5462 (N_5462,N_1389,N_94);
nor U5463 (N_5463,N_49,N_445);
xor U5464 (N_5464,N_1622,N_3836);
nor U5465 (N_5465,N_852,N_3657);
nand U5466 (N_5466,N_3541,N_4780);
and U5467 (N_5467,N_1061,N_4982);
nand U5468 (N_5468,N_2838,N_1427);
nand U5469 (N_5469,N_2267,N_1159);
xor U5470 (N_5470,N_215,N_525);
or U5471 (N_5471,N_4440,N_4583);
and U5472 (N_5472,N_4148,N_4172);
xnor U5473 (N_5473,N_3454,N_78);
or U5474 (N_5474,N_1616,N_4489);
nand U5475 (N_5475,N_3409,N_3171);
and U5476 (N_5476,N_3278,N_3437);
and U5477 (N_5477,N_3133,N_632);
and U5478 (N_5478,N_479,N_3195);
or U5479 (N_5479,N_3110,N_1673);
nor U5480 (N_5480,N_574,N_4332);
xor U5481 (N_5481,N_4728,N_1192);
and U5482 (N_5482,N_4965,N_3872);
or U5483 (N_5483,N_3719,N_1836);
nor U5484 (N_5484,N_2650,N_3040);
nor U5485 (N_5485,N_1610,N_1643);
or U5486 (N_5486,N_4119,N_3921);
xor U5487 (N_5487,N_3704,N_3920);
and U5488 (N_5488,N_3303,N_3049);
xnor U5489 (N_5489,N_3635,N_125);
and U5490 (N_5490,N_2342,N_564);
or U5491 (N_5491,N_3905,N_167);
and U5492 (N_5492,N_3394,N_2581);
and U5493 (N_5493,N_3068,N_2456);
nand U5494 (N_5494,N_4394,N_4968);
nor U5495 (N_5495,N_4525,N_2437);
or U5496 (N_5496,N_1,N_2289);
nor U5497 (N_5497,N_4095,N_1158);
nand U5498 (N_5498,N_4069,N_4745);
and U5499 (N_5499,N_2962,N_3372);
nor U5500 (N_5500,N_3518,N_3720);
nand U5501 (N_5501,N_2658,N_4244);
or U5502 (N_5502,N_1215,N_3364);
nand U5503 (N_5503,N_3799,N_1864);
nand U5504 (N_5504,N_2114,N_4058);
nor U5505 (N_5505,N_3984,N_4208);
nand U5506 (N_5506,N_4985,N_1469);
xor U5507 (N_5507,N_3499,N_1526);
xor U5508 (N_5508,N_3028,N_2288);
nor U5509 (N_5509,N_1442,N_282);
nor U5510 (N_5510,N_4281,N_1243);
and U5511 (N_5511,N_2570,N_1490);
nor U5512 (N_5512,N_1498,N_3337);
nand U5513 (N_5513,N_798,N_1072);
or U5514 (N_5514,N_2215,N_320);
or U5515 (N_5515,N_3660,N_3896);
and U5516 (N_5516,N_2130,N_1909);
and U5517 (N_5517,N_4864,N_1946);
or U5518 (N_5518,N_1096,N_4043);
or U5519 (N_5519,N_4914,N_4524);
or U5520 (N_5520,N_362,N_2880);
xor U5521 (N_5521,N_3127,N_790);
nor U5522 (N_5522,N_1313,N_3875);
nand U5523 (N_5523,N_1171,N_1665);
and U5524 (N_5524,N_4326,N_2833);
xnor U5525 (N_5525,N_1185,N_511);
xnor U5526 (N_5526,N_4872,N_4718);
or U5527 (N_5527,N_2943,N_2958);
and U5528 (N_5528,N_2295,N_3060);
nor U5529 (N_5529,N_1169,N_165);
nor U5530 (N_5530,N_1239,N_1664);
xor U5531 (N_5531,N_3869,N_3721);
nor U5532 (N_5532,N_355,N_804);
and U5533 (N_5533,N_2258,N_2387);
nand U5534 (N_5534,N_4317,N_3059);
nand U5535 (N_5535,N_3177,N_915);
xnor U5536 (N_5536,N_1651,N_100);
xor U5537 (N_5537,N_3452,N_2208);
nand U5538 (N_5538,N_4731,N_3128);
nor U5539 (N_5539,N_4467,N_3785);
xnor U5540 (N_5540,N_4182,N_2979);
nand U5541 (N_5541,N_1781,N_634);
nor U5542 (N_5542,N_3843,N_2196);
nand U5543 (N_5543,N_4536,N_942);
xor U5544 (N_5544,N_507,N_2701);
or U5545 (N_5545,N_3149,N_4045);
nor U5546 (N_5546,N_2910,N_1038);
xnor U5547 (N_5547,N_899,N_3407);
xnor U5548 (N_5548,N_2212,N_4248);
or U5549 (N_5549,N_4097,N_2292);
and U5550 (N_5550,N_2218,N_555);
xor U5551 (N_5551,N_1633,N_203);
nand U5552 (N_5552,N_850,N_3626);
or U5553 (N_5553,N_4110,N_1143);
nor U5554 (N_5554,N_2073,N_741);
and U5555 (N_5555,N_1379,N_768);
or U5556 (N_5556,N_4155,N_3651);
or U5557 (N_5557,N_3225,N_3100);
xnor U5558 (N_5558,N_2608,N_3803);
and U5559 (N_5559,N_2475,N_3478);
xnor U5560 (N_5560,N_2790,N_504);
and U5561 (N_5561,N_1942,N_4959);
nand U5562 (N_5562,N_521,N_3388);
xnor U5563 (N_5563,N_1021,N_4170);
or U5564 (N_5564,N_353,N_1358);
or U5565 (N_5565,N_4719,N_4779);
xor U5566 (N_5566,N_3783,N_1721);
nor U5567 (N_5567,N_316,N_2730);
and U5568 (N_5568,N_4659,N_2715);
nand U5569 (N_5569,N_1908,N_1216);
nor U5570 (N_5570,N_2499,N_1971);
or U5571 (N_5571,N_1483,N_1679);
xnor U5572 (N_5572,N_2504,N_2755);
nor U5573 (N_5573,N_367,N_1163);
or U5574 (N_5574,N_1539,N_2128);
nor U5575 (N_5575,N_3362,N_3673);
nor U5576 (N_5576,N_2152,N_3201);
or U5577 (N_5577,N_4411,N_617);
xnor U5578 (N_5578,N_2381,N_3583);
nand U5579 (N_5579,N_3718,N_3269);
and U5580 (N_5580,N_3487,N_3130);
nor U5581 (N_5581,N_1359,N_2200);
and U5582 (N_5582,N_3192,N_1300);
nor U5583 (N_5583,N_1463,N_3495);
nand U5584 (N_5584,N_1125,N_3932);
and U5585 (N_5585,N_516,N_3930);
or U5586 (N_5586,N_1367,N_384);
nand U5587 (N_5587,N_1371,N_56);
nor U5588 (N_5588,N_2785,N_3965);
nor U5589 (N_5589,N_3035,N_2594);
or U5590 (N_5590,N_2506,N_2627);
and U5591 (N_5591,N_700,N_422);
xor U5592 (N_5592,N_3690,N_3613);
or U5593 (N_5593,N_4213,N_1981);
nor U5594 (N_5594,N_1915,N_1608);
nor U5595 (N_5595,N_2989,N_2977);
or U5596 (N_5596,N_1887,N_969);
nand U5597 (N_5597,N_1102,N_4544);
or U5598 (N_5598,N_1540,N_1292);
nor U5599 (N_5599,N_3691,N_4141);
xnor U5600 (N_5600,N_4979,N_118);
and U5601 (N_5601,N_390,N_1548);
nor U5602 (N_5602,N_3022,N_350);
or U5603 (N_5603,N_3446,N_2079);
xnor U5604 (N_5604,N_3851,N_4462);
nand U5605 (N_5605,N_4384,N_1470);
xor U5606 (N_5606,N_1467,N_1045);
or U5607 (N_5607,N_4935,N_762);
nand U5608 (N_5608,N_3870,N_2578);
or U5609 (N_5609,N_623,N_2007);
or U5610 (N_5610,N_1341,N_435);
xor U5611 (N_5611,N_182,N_4775);
nor U5612 (N_5612,N_4305,N_3898);
nand U5613 (N_5613,N_2836,N_2165);
or U5614 (N_5614,N_1767,N_3492);
or U5615 (N_5615,N_3453,N_4002);
nor U5616 (N_5616,N_4887,N_841);
nor U5617 (N_5617,N_4236,N_4548);
nand U5618 (N_5618,N_1401,N_1888);
nand U5619 (N_5619,N_1327,N_629);
nand U5620 (N_5620,N_2334,N_3814);
nor U5621 (N_5621,N_965,N_1592);
nor U5622 (N_5622,N_2314,N_3929);
xor U5623 (N_5623,N_4785,N_547);
nand U5624 (N_5624,N_4059,N_3652);
or U5625 (N_5625,N_3455,N_2041);
nand U5626 (N_5626,N_3701,N_1166);
xnor U5627 (N_5627,N_2704,N_2975);
or U5628 (N_5628,N_3857,N_2070);
nand U5629 (N_5629,N_4336,N_3218);
or U5630 (N_5630,N_1801,N_1127);
and U5631 (N_5631,N_1843,N_38);
nand U5632 (N_5632,N_3484,N_3116);
and U5633 (N_5633,N_4190,N_1766);
xor U5634 (N_5634,N_686,N_1625);
nor U5635 (N_5635,N_4927,N_4961);
nand U5636 (N_5636,N_1403,N_1692);
nor U5637 (N_5637,N_1497,N_2169);
xnor U5638 (N_5638,N_102,N_4712);
and U5639 (N_5639,N_4230,N_4644);
or U5640 (N_5640,N_494,N_3354);
or U5641 (N_5641,N_1761,N_216);
nor U5642 (N_5642,N_2623,N_1956);
and U5643 (N_5643,N_4014,N_1662);
nand U5644 (N_5644,N_1276,N_4369);
or U5645 (N_5645,N_1631,N_3169);
nand U5646 (N_5646,N_735,N_1537);
nand U5647 (N_5647,N_4287,N_425);
xor U5648 (N_5648,N_2460,N_369);
and U5649 (N_5649,N_4140,N_101);
or U5650 (N_5650,N_3038,N_1287);
and U5651 (N_5651,N_959,N_12);
xnor U5652 (N_5652,N_446,N_2111);
and U5653 (N_5653,N_1478,N_4019);
nand U5654 (N_5654,N_4271,N_2092);
nor U5655 (N_5655,N_2532,N_1348);
nand U5656 (N_5656,N_757,N_2619);
or U5657 (N_5657,N_2693,N_1382);
nor U5658 (N_5658,N_2938,N_17);
nand U5659 (N_5659,N_1035,N_4116);
nand U5660 (N_5660,N_4368,N_4565);
xor U5661 (N_5661,N_2950,N_3699);
or U5662 (N_5662,N_2722,N_677);
and U5663 (N_5663,N_3732,N_2119);
and U5664 (N_5664,N_1465,N_4026);
and U5665 (N_5665,N_4511,N_2014);
nor U5666 (N_5666,N_43,N_3190);
xor U5667 (N_5667,N_3075,N_2244);
nor U5668 (N_5668,N_1799,N_2605);
xnor U5669 (N_5669,N_3525,N_1951);
nand U5670 (N_5670,N_2272,N_88);
nand U5671 (N_5671,N_645,N_85);
nand U5672 (N_5672,N_230,N_3210);
or U5673 (N_5673,N_71,N_1515);
or U5674 (N_5674,N_4693,N_1285);
or U5675 (N_5675,N_3185,N_2138);
or U5676 (N_5676,N_3672,N_1370);
nor U5677 (N_5677,N_2240,N_4479);
or U5678 (N_5678,N_3009,N_1212);
or U5679 (N_5679,N_4400,N_4905);
nor U5680 (N_5680,N_1448,N_3604);
nand U5681 (N_5681,N_2514,N_3607);
or U5682 (N_5682,N_1289,N_4996);
and U5683 (N_5683,N_4431,N_3894);
nor U5684 (N_5684,N_57,N_1068);
nand U5685 (N_5685,N_4356,N_1003);
or U5686 (N_5686,N_4717,N_3426);
and U5687 (N_5687,N_1646,N_1782);
nor U5688 (N_5688,N_1057,N_1070);
xnor U5689 (N_5689,N_1372,N_1294);
or U5690 (N_5690,N_1254,N_2455);
nand U5691 (N_5691,N_2857,N_1871);
nor U5692 (N_5692,N_627,N_610);
nor U5693 (N_5693,N_3144,N_1975);
nor U5694 (N_5694,N_4319,N_1504);
nand U5695 (N_5695,N_3602,N_966);
xor U5696 (N_5696,N_642,N_2736);
nand U5697 (N_5697,N_2344,N_1904);
nor U5698 (N_5698,N_397,N_2812);
or U5699 (N_5699,N_3226,N_2952);
nor U5700 (N_5700,N_4920,N_4435);
and U5701 (N_5701,N_2198,N_3113);
nor U5702 (N_5702,N_2967,N_2561);
nand U5703 (N_5703,N_4991,N_1482);
and U5704 (N_5704,N_4330,N_589);
and U5705 (N_5705,N_2624,N_4247);
xor U5706 (N_5706,N_1695,N_3654);
and U5707 (N_5707,N_541,N_888);
and U5708 (N_5708,N_3900,N_3645);
or U5709 (N_5709,N_1556,N_2270);
xor U5710 (N_5710,N_4218,N_2502);
and U5711 (N_5711,N_2882,N_4274);
xnor U5712 (N_5712,N_3056,N_4476);
and U5713 (N_5713,N_2046,N_134);
nor U5714 (N_5714,N_2436,N_4089);
nand U5715 (N_5715,N_1880,N_2593);
or U5716 (N_5716,N_1231,N_4827);
nor U5717 (N_5717,N_136,N_1706);
and U5718 (N_5718,N_4458,N_388);
nand U5719 (N_5719,N_4535,N_2569);
nor U5720 (N_5720,N_802,N_2659);
or U5721 (N_5721,N_2733,N_3865);
or U5722 (N_5722,N_345,N_693);
nand U5723 (N_5723,N_3003,N_2779);
and U5724 (N_5724,N_2516,N_889);
or U5725 (N_5725,N_2987,N_1959);
nand U5726 (N_5726,N_4832,N_3957);
nand U5727 (N_5727,N_502,N_1210);
nor U5728 (N_5728,N_2703,N_845);
nor U5729 (N_5729,N_890,N_1594);
or U5730 (N_5730,N_92,N_731);
nand U5731 (N_5731,N_1455,N_1369);
or U5732 (N_5732,N_2711,N_4945);
and U5733 (N_5733,N_2505,N_1431);
nor U5734 (N_5734,N_4065,N_2764);
or U5735 (N_5735,N_245,N_3788);
and U5736 (N_5736,N_2285,N_3797);
and U5737 (N_5737,N_4612,N_2394);
xnor U5738 (N_5738,N_4954,N_3951);
xnor U5739 (N_5739,N_2720,N_2692);
or U5740 (N_5740,N_4423,N_1085);
nand U5741 (N_5741,N_2672,N_3153);
or U5742 (N_5742,N_854,N_2002);
nor U5743 (N_5743,N_3490,N_3846);
nor U5744 (N_5744,N_1411,N_2458);
nand U5745 (N_5745,N_1345,N_868);
nand U5746 (N_5746,N_2222,N_3912);
or U5747 (N_5747,N_324,N_2003);
nand U5748 (N_5748,N_912,N_4809);
or U5749 (N_5749,N_493,N_2399);
or U5750 (N_5750,N_1322,N_391);
nand U5751 (N_5751,N_4152,N_2126);
nand U5752 (N_5752,N_291,N_543);
xor U5753 (N_5753,N_4957,N_1825);
or U5754 (N_5754,N_4242,N_3978);
nor U5755 (N_5755,N_941,N_3419);
nand U5756 (N_5756,N_2202,N_5);
nand U5757 (N_5757,N_1775,N_1701);
xor U5758 (N_5758,N_2472,N_4009);
nor U5759 (N_5759,N_2547,N_3104);
nor U5760 (N_5760,N_1487,N_2645);
nor U5761 (N_5761,N_2996,N_2583);
nor U5762 (N_5762,N_1031,N_3675);
or U5763 (N_5763,N_3284,N_2415);
or U5764 (N_5764,N_281,N_16);
and U5765 (N_5765,N_873,N_680);
or U5766 (N_5766,N_1363,N_2539);
nand U5767 (N_5767,N_842,N_1067);
or U5768 (N_5768,N_3743,N_2463);
or U5769 (N_5769,N_1224,N_3342);
nand U5770 (N_5770,N_3023,N_3966);
nor U5771 (N_5771,N_1383,N_4072);
nor U5772 (N_5772,N_2450,N_2101);
nand U5773 (N_5773,N_1137,N_3693);
nand U5774 (N_5774,N_2753,N_4406);
and U5775 (N_5775,N_3106,N_962);
nor U5776 (N_5776,N_4617,N_4681);
or U5777 (N_5777,N_4063,N_3304);
or U5778 (N_5778,N_4486,N_79);
or U5779 (N_5779,N_2116,N_347);
xnor U5780 (N_5780,N_2868,N_4263);
nor U5781 (N_5781,N_1690,N_4495);
xor U5782 (N_5782,N_1010,N_3988);
and U5783 (N_5783,N_4610,N_51);
nor U5784 (N_5784,N_4818,N_2448);
nand U5785 (N_5785,N_4714,N_4364);
nor U5786 (N_5786,N_3335,N_447);
xor U5787 (N_5787,N_93,N_2929);
or U5788 (N_5788,N_74,N_1560);
and U5789 (N_5789,N_3054,N_4878);
or U5790 (N_5790,N_1660,N_220);
or U5791 (N_5791,N_3745,N_3595);
nor U5792 (N_5792,N_3546,N_1994);
xor U5793 (N_5793,N_272,N_393);
or U5794 (N_5794,N_4701,N_2770);
nand U5795 (N_5795,N_856,N_1441);
and U5796 (N_5796,N_4160,N_204);
xnor U5797 (N_5797,N_557,N_4556);
and U5798 (N_5798,N_988,N_840);
and U5799 (N_5799,N_1302,N_1028);
nand U5800 (N_5800,N_2051,N_488);
and U5801 (N_5801,N_1738,N_1740);
xor U5802 (N_5802,N_219,N_358);
xor U5803 (N_5803,N_1318,N_4754);
xnor U5804 (N_5804,N_4075,N_4080);
and U5805 (N_5805,N_1848,N_3399);
xor U5806 (N_5806,N_458,N_4201);
nand U5807 (N_5807,N_4436,N_2481);
nand U5808 (N_5808,N_3435,N_1997);
and U5809 (N_5809,N_2117,N_404);
nor U5810 (N_5810,N_2296,N_936);
nand U5811 (N_5811,N_3387,N_3868);
or U5812 (N_5812,N_3942,N_1098);
nor U5813 (N_5813,N_1505,N_189);
xor U5814 (N_5814,N_1723,N_1172);
nor U5815 (N_5815,N_4269,N_4568);
xor U5816 (N_5816,N_4679,N_158);
or U5817 (N_5817,N_4158,N_4704);
nor U5818 (N_5818,N_1796,N_655);
or U5819 (N_5819,N_3556,N_2617);
xor U5820 (N_5820,N_67,N_834);
or U5821 (N_5821,N_185,N_3917);
nor U5822 (N_5822,N_1051,N_3682);
and U5823 (N_5823,N_979,N_2064);
and U5824 (N_5824,N_4594,N_1245);
nand U5825 (N_5825,N_3433,N_596);
and U5826 (N_5826,N_1851,N_2559);
nand U5827 (N_5827,N_3415,N_3101);
nand U5828 (N_5828,N_2099,N_1378);
or U5829 (N_5829,N_3973,N_2435);
and U5830 (N_5830,N_460,N_3176);
nor U5831 (N_5831,N_3991,N_3711);
nand U5832 (N_5832,N_3486,N_882);
nand U5833 (N_5833,N_3457,N_2758);
nor U5834 (N_5834,N_3935,N_4418);
nor U5835 (N_5835,N_2369,N_674);
and U5836 (N_5836,N_1281,N_1111);
nand U5837 (N_5837,N_4171,N_4297);
and U5838 (N_5838,N_202,N_3947);
or U5839 (N_5839,N_4454,N_1855);
and U5840 (N_5840,N_2479,N_2681);
nor U5841 (N_5841,N_4216,N_2677);
or U5842 (N_5842,N_3143,N_2500);
nand U5843 (N_5843,N_542,N_2498);
and U5844 (N_5844,N_1742,N_4940);
and U5845 (N_5845,N_2123,N_4532);
or U5846 (N_5846,N_1019,N_3601);
xor U5847 (N_5847,N_2453,N_2310);
nor U5848 (N_5848,N_2091,N_4537);
or U5849 (N_5849,N_2094,N_2810);
or U5850 (N_5850,N_3380,N_3405);
nor U5851 (N_5851,N_470,N_1355);
or U5852 (N_5852,N_2837,N_4634);
nor U5853 (N_5853,N_3606,N_3189);
and U5854 (N_5854,N_4231,N_3901);
nor U5855 (N_5855,N_4938,N_1545);
and U5856 (N_5856,N_1685,N_6);
and U5857 (N_5857,N_2286,N_274);
or U5858 (N_5858,N_4875,N_4749);
nor U5859 (N_5859,N_1921,N_4285);
or U5860 (N_5860,N_4800,N_2413);
and U5861 (N_5861,N_4660,N_4254);
and U5862 (N_5862,N_3863,N_619);
nor U5863 (N_5863,N_884,N_1479);
xor U5864 (N_5864,N_2333,N_3611);
nor U5865 (N_5865,N_1221,N_2010);
and U5866 (N_5866,N_3724,N_794);
nor U5867 (N_5867,N_2719,N_4871);
and U5868 (N_5868,N_1812,N_1511);
or U5869 (N_5869,N_4191,N_3964);
xor U5870 (N_5870,N_4756,N_4397);
and U5871 (N_5871,N_4385,N_3810);
xor U5872 (N_5872,N_4035,N_3581);
xnor U5873 (N_5873,N_2951,N_2656);
nand U5874 (N_5874,N_4539,N_797);
nand U5875 (N_5875,N_4700,N_692);
and U5876 (N_5876,N_1046,N_1854);
xnor U5877 (N_5877,N_3198,N_4139);
and U5878 (N_5878,N_4267,N_4836);
and U5879 (N_5879,N_1180,N_2368);
and U5880 (N_5880,N_4000,N_2024);
xnor U5881 (N_5881,N_4238,N_371);
nor U5882 (N_5882,N_2970,N_2980);
or U5883 (N_5883,N_2016,N_4921);
nand U5884 (N_5884,N_4894,N_3873);
and U5885 (N_5885,N_4207,N_4705);
nor U5886 (N_5886,N_1984,N_2377);
nor U5887 (N_5887,N_1947,N_2120);
or U5888 (N_5888,N_3025,N_4001);
or U5889 (N_5889,N_3496,N_1613);
or U5890 (N_5890,N_2955,N_2553);
or U5891 (N_5891,N_4715,N_4234);
and U5892 (N_5892,N_4620,N_4212);
xor U5893 (N_5893,N_1827,N_3447);
nand U5894 (N_5894,N_4695,N_440);
and U5895 (N_5895,N_3879,N_2186);
nor U5896 (N_5896,N_4215,N_913);
xnor U5897 (N_5897,N_4339,N_1004);
nor U5898 (N_5898,N_2807,N_861);
xnor U5899 (N_5899,N_4444,N_3569);
nand U5900 (N_5900,N_3463,N_1416);
nand U5901 (N_5901,N_847,N_4797);
or U5902 (N_5902,N_3418,N_978);
nor U5903 (N_5903,N_3074,N_4087);
nand U5904 (N_5904,N_2351,N_723);
nand U5905 (N_5905,N_4146,N_4530);
xor U5906 (N_5906,N_927,N_4570);
and U5907 (N_5907,N_1494,N_2519);
nand U5908 (N_5908,N_226,N_3117);
nand U5909 (N_5909,N_3223,N_900);
or U5910 (N_5910,N_2205,N_2157);
nor U5911 (N_5911,N_4855,N_863);
xor U5912 (N_5912,N_651,N_1809);
nor U5913 (N_5913,N_552,N_2739);
or U5914 (N_5914,N_4455,N_615);
nor U5915 (N_5915,N_2133,N_3456);
xnor U5916 (N_5916,N_2888,N_4029);
and U5917 (N_5917,N_2080,N_3725);
or U5918 (N_5918,N_3520,N_3124);
xor U5919 (N_5919,N_1218,N_3639);
nor U5920 (N_5920,N_1049,N_2273);
xor U5921 (N_5921,N_4241,N_3325);
or U5922 (N_5922,N_4475,N_4973);
nor U5923 (N_5923,N_2944,N_2322);
nor U5924 (N_5924,N_305,N_1768);
xnor U5925 (N_5925,N_2630,N_1698);
nand U5926 (N_5926,N_10,N_786);
or U5927 (N_5927,N_3006,N_1110);
xor U5928 (N_5928,N_3977,N_1007);
and U5929 (N_5929,N_2670,N_2474);
xor U5930 (N_5930,N_381,N_3359);
or U5931 (N_5931,N_4036,N_4204);
xnor U5932 (N_5932,N_3173,N_897);
nor U5933 (N_5933,N_3609,N_697);
xor U5934 (N_5934,N_989,N_169);
and U5935 (N_5935,N_4892,N_2926);
xor U5936 (N_5936,N_3402,N_2367);
nand U5937 (N_5937,N_2325,N_4733);
nor U5938 (N_5938,N_4930,N_1600);
or U5939 (N_5939,N_1912,N_3772);
xnor U5940 (N_5940,N_2136,N_4856);
nor U5941 (N_5941,N_1440,N_1861);
or U5942 (N_5942,N_643,N_1650);
or U5943 (N_5943,N_472,N_1876);
nand U5944 (N_5944,N_4349,N_2688);
nor U5945 (N_5945,N_1060,N_14);
nor U5946 (N_5946,N_2697,N_2793);
and U5947 (N_5947,N_55,N_4947);
nor U5948 (N_5948,N_4834,N_1452);
xor U5949 (N_5949,N_501,N_4599);
xnor U5950 (N_5950,N_1444,N_1638);
xnor U5951 (N_5951,N_1086,N_2062);
xor U5952 (N_5952,N_2823,N_649);
nor U5953 (N_5953,N_284,N_83);
xor U5954 (N_5954,N_1817,N_4410);
nor U5955 (N_5955,N_1055,N_4691);
or U5956 (N_5956,N_3537,N_1602);
nand U5957 (N_5957,N_4858,N_1807);
and U5958 (N_5958,N_4318,N_2610);
and U5959 (N_5959,N_1324,N_1568);
or U5960 (N_5960,N_2335,N_111);
and U5961 (N_5961,N_4184,N_2346);
nor U5962 (N_5962,N_4661,N_1399);
or U5963 (N_5963,N_3575,N_2328);
xnor U5964 (N_5964,N_2147,N_1129);
and U5965 (N_5965,N_4402,N_848);
and U5966 (N_5966,N_3213,N_1170);
nor U5967 (N_5967,N_584,N_902);
nor U5968 (N_5968,N_3333,N_2609);
or U5969 (N_5969,N_1939,N_1380);
nand U5970 (N_5970,N_3826,N_340);
or U5971 (N_5971,N_2197,N_1162);
xor U5972 (N_5972,N_4197,N_3663);
nand U5973 (N_5973,N_3032,N_3637);
nand U5974 (N_5974,N_3191,N_1746);
and U5975 (N_5975,N_2411,N_1684);
nand U5976 (N_5976,N_616,N_439);
xor U5977 (N_5977,N_1726,N_2433);
or U5978 (N_5978,N_1157,N_4706);
and U5979 (N_5979,N_236,N_3277);
and U5980 (N_5980,N_3238,N_4750);
or U5981 (N_5981,N_1572,N_238);
nand U5982 (N_5982,N_4723,N_4578);
nor U5983 (N_5983,N_1998,N_742);
or U5984 (N_5984,N_3515,N_225);
nor U5985 (N_5985,N_1190,N_3087);
nor U5986 (N_5986,N_1495,N_2820);
xnor U5987 (N_5987,N_2699,N_1336);
or U5988 (N_5988,N_4805,N_3442);
or U5989 (N_5989,N_4515,N_1304);
or U5990 (N_5990,N_4811,N_4157);
xor U5991 (N_5991,N_1134,N_4219);
and U5992 (N_5992,N_4761,N_2187);
and U5993 (N_5993,N_267,N_4381);
nand U5994 (N_5994,N_197,N_2671);
and U5995 (N_5995,N_1838,N_2308);
and U5996 (N_5996,N_2440,N_2468);
nor U5997 (N_5997,N_476,N_4774);
or U5998 (N_5998,N_2757,N_3910);
nor U5999 (N_5999,N_1458,N_4438);
xor U6000 (N_6000,N_1900,N_4857);
nand U6001 (N_6001,N_3373,N_4290);
nand U6002 (N_6002,N_2231,N_2744);
xnor U6003 (N_6003,N_211,N_66);
xnor U6004 (N_6004,N_3353,N_3048);
xnor U6005 (N_6005,N_2378,N_2054);
and U6006 (N_6006,N_3443,N_3384);
or U6007 (N_6007,N_1390,N_3685);
nand U6008 (N_6008,N_4039,N_299);
or U6009 (N_6009,N_592,N_179);
xor U6010 (N_6010,N_3915,N_3768);
nor U6011 (N_6011,N_3365,N_1351);
or U6012 (N_6012,N_2545,N_1818);
nor U6013 (N_6013,N_3571,N_719);
xnor U6014 (N_6014,N_4528,N_2898);
nand U6015 (N_6015,N_1846,N_3784);
or U6016 (N_6016,N_3574,N_2687);
and U6017 (N_6017,N_2560,N_3828);
or U6018 (N_6018,N_3773,N_4686);
and U6019 (N_6019,N_4549,N_601);
nand U6020 (N_6020,N_2984,N_622);
or U6021 (N_6021,N_3861,N_3244);
or U6022 (N_6022,N_2257,N_2149);
nand U6023 (N_6023,N_926,N_1597);
and U6024 (N_6024,N_752,N_147);
nand U6025 (N_6025,N_4324,N_3466);
xor U6026 (N_6026,N_302,N_4390);
xor U6027 (N_6027,N_405,N_4958);
nor U6028 (N_6028,N_1459,N_145);
nor U6029 (N_6029,N_175,N_407);
xnor U6030 (N_6030,N_4512,N_934);
nor U6031 (N_6031,N_1264,N_973);
and U6032 (N_6032,N_2194,N_3813);
xor U6033 (N_6033,N_4441,N_4040);
nand U6034 (N_6034,N_2188,N_2621);
xor U6035 (N_6035,N_2523,N_2090);
xor U6036 (N_6036,N_4546,N_1538);
or U6037 (N_6037,N_4108,N_753);
xor U6038 (N_6038,N_660,N_1357);
nand U6039 (N_6039,N_1069,N_2362);
xor U6040 (N_6040,N_2373,N_3314);
and U6041 (N_6041,N_3093,N_4279);
and U6042 (N_6042,N_2741,N_4605);
nand U6043 (N_6043,N_3516,N_687);
xor U6044 (N_6044,N_3091,N_290);
and U6045 (N_6045,N_572,N_3731);
or U6046 (N_6046,N_4273,N_951);
nand U6047 (N_6047,N_2737,N_1604);
and U6048 (N_6048,N_4300,N_2184);
nor U6049 (N_6049,N_4022,N_2507);
nand U6050 (N_6050,N_2393,N_1420);
nand U6051 (N_6051,N_3631,N_1637);
and U6052 (N_6052,N_3945,N_506);
or U6053 (N_6053,N_2488,N_3292);
nor U6054 (N_6054,N_2904,N_1123);
nand U6055 (N_6055,N_4725,N_1438);
nand U6056 (N_6056,N_4409,N_3963);
xnor U6057 (N_6057,N_2444,N_3052);
or U6058 (N_6058,N_2781,N_3748);
nor U6059 (N_6059,N_1536,N_2886);
nand U6060 (N_6060,N_1714,N_3464);
or U6061 (N_6061,N_2374,N_4702);
and U6062 (N_6062,N_513,N_2410);
or U6063 (N_6063,N_1916,N_3055);
nand U6064 (N_6064,N_3931,N_661);
nand U6065 (N_6065,N_1132,N_825);
xor U6066 (N_6066,N_1509,N_4067);
nand U6067 (N_6067,N_3286,N_1820);
and U6068 (N_6068,N_641,N_1693);
or U6069 (N_6069,N_2084,N_232);
or U6070 (N_6070,N_967,N_3482);
and U6071 (N_6071,N_1835,N_1732);
nand U6072 (N_6072,N_2611,N_3004);
xor U6073 (N_6073,N_3058,N_2596);
or U6074 (N_6074,N_1530,N_1962);
and U6075 (N_6075,N_1349,N_1034);
nand U6076 (N_6076,N_4424,N_3308);
nor U6077 (N_6077,N_2398,N_40);
nand U6078 (N_6078,N_3893,N_1607);
nor U6079 (N_6079,N_715,N_3999);
nor U6080 (N_6080,N_917,N_1585);
and U6081 (N_6081,N_1451,N_3563);
and U6082 (N_6082,N_183,N_1404);
xnor U6083 (N_6083,N_4826,N_1553);
and U6084 (N_6084,N_1522,N_1547);
and U6085 (N_6085,N_3584,N_4720);
and U6086 (N_6086,N_2804,N_4837);
nor U6087 (N_6087,N_3985,N_4652);
or U6088 (N_6088,N_679,N_3298);
and U6089 (N_6089,N_4496,N_285);
xnor U6090 (N_6090,N_209,N_4162);
or U6091 (N_6091,N_3994,N_1596);
nand U6092 (N_6092,N_3265,N_3640);
or U6093 (N_6093,N_4682,N_4275);
xor U6094 (N_6094,N_4151,N_4886);
nand U6095 (N_6095,N_4255,N_99);
nor U6096 (N_6096,N_2306,N_1058);
nor U6097 (N_6097,N_4697,N_4577);
xor U6098 (N_6098,N_3123,N_3064);
and U6099 (N_6099,N_1619,N_1800);
nand U6100 (N_6100,N_3299,N_2250);
and U6101 (N_6101,N_2380,N_2895);
nand U6102 (N_6102,N_3946,N_3367);
nor U6103 (N_6103,N_975,N_2986);
xnor U6104 (N_6104,N_4027,N_705);
or U6105 (N_6105,N_4093,N_1152);
and U6106 (N_6106,N_1790,N_2788);
nand U6107 (N_6107,N_1506,N_787);
and U6108 (N_6108,N_1496,N_2359);
and U6109 (N_6109,N_1308,N_2916);
and U6110 (N_6110,N_2840,N_3392);
and U6111 (N_6111,N_3916,N_2591);
nor U6112 (N_6112,N_1017,N_3646);
nand U6113 (N_6113,N_4193,N_1972);
or U6114 (N_6114,N_2081,N_1436);
nand U6115 (N_6115,N_4752,N_160);
xnor U6116 (N_6116,N_450,N_1114);
nand U6117 (N_6117,N_3021,N_604);
nor U6118 (N_6118,N_682,N_4597);
xnor U6119 (N_6119,N_761,N_820);
nand U6120 (N_6120,N_1131,N_3830);
nand U6121 (N_6121,N_2443,N_775);
nor U6122 (N_6122,N_3831,N_870);
xor U6123 (N_6123,N_1186,N_1832);
and U6124 (N_6124,N_3853,N_1805);
nand U6125 (N_6125,N_945,N_3962);
xnor U6126 (N_6126,N_153,N_4689);
or U6127 (N_6127,N_4226,N_441);
nor U6128 (N_6128,N_1773,N_4541);
nor U6129 (N_6129,N_4413,N_462);
xnor U6130 (N_6130,N_3953,N_4386);
and U6131 (N_6131,N_4547,N_4919);
or U6132 (N_6132,N_4237,N_277);
or U6133 (N_6133,N_3624,N_1725);
and U6134 (N_6134,N_1342,N_4948);
or U6135 (N_6135,N_874,N_999);
nor U6136 (N_6136,N_3523,N_920);
xnor U6137 (N_6137,N_2324,N_4488);
nand U6138 (N_6138,N_1472,N_1155);
and U6139 (N_6139,N_789,N_1025);
nor U6140 (N_6140,N_1457,N_1840);
and U6141 (N_6141,N_3242,N_3057);
or U6142 (N_6142,N_261,N_4051);
or U6143 (N_6143,N_1940,N_3078);
or U6144 (N_6144,N_1780,N_871);
and U6145 (N_6145,N_1542,N_3970);
nand U6146 (N_6146,N_2827,N_2981);
nand U6147 (N_6147,N_3576,N_4249);
xor U6148 (N_6148,N_3289,N_3012);
nor U6149 (N_6149,N_4964,N_4429);
and U6150 (N_6150,N_2580,N_1146);
xnor U6151 (N_6151,N_3542,N_3911);
and U6152 (N_6152,N_894,N_1577);
xor U6153 (N_6153,N_2323,N_725);
and U6154 (N_6154,N_2964,N_18);
nand U6155 (N_6155,N_2228,N_2771);
xnor U6156 (N_6156,N_4342,N_475);
and U6157 (N_6157,N_1217,N_2816);
and U6158 (N_6158,N_1866,N_2392);
xor U6159 (N_6159,N_4195,N_3636);
and U6160 (N_6160,N_4082,N_389);
nor U6161 (N_6161,N_1407,N_2211);
or U6162 (N_6162,N_4123,N_1423);
or U6163 (N_6163,N_336,N_4203);
or U6164 (N_6164,N_289,N_132);
and U6165 (N_6165,N_1016,N_803);
nand U6166 (N_6166,N_137,N_64);
or U6167 (N_6167,N_3889,N_774);
nor U6168 (N_6168,N_1273,N_2676);
and U6169 (N_6169,N_148,N_566);
nand U6170 (N_6170,N_3996,N_1751);
and U6171 (N_6171,N_4942,N_2858);
nor U6172 (N_6172,N_3641,N_1278);
nand U6173 (N_6173,N_983,N_613);
nand U6174 (N_6174,N_1493,N_4823);
nand U6175 (N_6175,N_1042,N_2728);
nand U6176 (N_6176,N_3085,N_1392);
xor U6177 (N_6177,N_357,N_3617);
xor U6178 (N_6178,N_1990,N_4145);
nor U6179 (N_6179,N_4619,N_736);
xor U6180 (N_6180,N_2798,N_4323);
and U6181 (N_6181,N_718,N_1325);
and U6182 (N_6182,N_4288,N_409);
or U6183 (N_6183,N_4980,N_1284);
nand U6184 (N_6184,N_1240,N_1623);
nand U6185 (N_6185,N_3876,N_1211);
or U6186 (N_6186,N_2434,N_1867);
and U6187 (N_6187,N_602,N_2805);
and U6188 (N_6188,N_1052,N_3063);
xnor U6189 (N_6189,N_4880,N_2854);
or U6190 (N_6190,N_2745,N_4099);
or U6191 (N_6191,N_3421,N_1421);
nand U6192 (N_6192,N_2808,N_2794);
xnor U6193 (N_6193,N_333,N_3428);
xor U6194 (N_6194,N_4795,N_918);
and U6195 (N_6195,N_1938,N_2828);
or U6196 (N_6196,N_4106,N_553);
nor U6197 (N_6197,N_0,N_490);
nor U6198 (N_6198,N_3448,N_1033);
nor U6199 (N_6199,N_1657,N_901);
and U6200 (N_6200,N_2932,N_1872);
nand U6201 (N_6201,N_461,N_1764);
or U6202 (N_6202,N_2311,N_3771);
xnor U6203 (N_6203,N_3795,N_4425);
nor U6204 (N_6204,N_97,N_1847);
nor U6205 (N_6205,N_878,N_4478);
nand U6206 (N_6206,N_2224,N_2872);
nor U6207 (N_6207,N_4031,N_4671);
xor U6208 (N_6208,N_1862,N_4931);
nand U6209 (N_6209,N_4156,N_161);
nand U6210 (N_6210,N_635,N_3703);
and U6211 (N_6211,N_3227,N_1145);
xor U6212 (N_6212,N_1941,N_4109);
xor U6213 (N_6213,N_2616,N_4373);
and U6214 (N_6214,N_1147,N_2432);
nand U6215 (N_6215,N_569,N_3164);
or U6216 (N_6216,N_283,N_3855);
or U6217 (N_6217,N_1518,N_437);
nor U6218 (N_6218,N_3122,N_1772);
nor U6219 (N_6219,N_952,N_3766);
and U6220 (N_6220,N_255,N_4494);
and U6221 (N_6221,N_4849,N_4741);
nand U6222 (N_6222,N_767,N_2576);
xor U6223 (N_6223,N_2327,N_374);
or U6224 (N_6224,N_442,N_2993);
or U6225 (N_6225,N_372,N_3790);
or U6226 (N_6226,N_4969,N_1743);
or U6227 (N_6227,N_3858,N_4637);
or U6228 (N_6228,N_1460,N_4365);
and U6229 (N_6229,N_1354,N_2855);
nor U6230 (N_6230,N_3754,N_4760);
and U6231 (N_6231,N_2013,N_2293);
and U6232 (N_6232,N_2001,N_3291);
nor U6233 (N_6233,N_3561,N_2949);
nor U6234 (N_6234,N_4860,N_3532);
and U6235 (N_6235,N_1844,N_2300);
xnor U6236 (N_6236,N_4699,N_4046);
or U6237 (N_6237,N_3958,N_793);
nor U6238 (N_6238,N_3172,N_1391);
or U6239 (N_6239,N_570,N_730);
and U6240 (N_6240,N_828,N_4989);
or U6241 (N_6241,N_240,N_4710);
and U6242 (N_6242,N_4863,N_2765);
or U6243 (N_6243,N_3707,N_2927);
or U6244 (N_6244,N_2030,N_2832);
xnor U6245 (N_6245,N_483,N_426);
nand U6246 (N_6246,N_4276,N_2768);
xor U6247 (N_6247,N_4250,N_62);
and U6248 (N_6248,N_77,N_2009);
xor U6249 (N_6249,N_1520,N_1331);
or U6250 (N_6250,N_1934,N_3061);
and U6251 (N_6251,N_540,N_1859);
and U6252 (N_6252,N_4734,N_4481);
or U6253 (N_6253,N_548,N_84);
nand U6254 (N_6254,N_4521,N_722);
nor U6255 (N_6255,N_1617,N_3000);
and U6256 (N_6256,N_2939,N_128);
or U6257 (N_6257,N_998,N_1717);
nor U6258 (N_6258,N_4477,N_3655);
nor U6259 (N_6259,N_2183,N_3334);
xnor U6260 (N_6260,N_3016,N_772);
nor U6261 (N_6261,N_1627,N_4859);
or U6262 (N_6262,N_4302,N_4674);
nor U6263 (N_6263,N_2206,N_2018);
xnor U6264 (N_6264,N_382,N_3254);
nor U6265 (N_6265,N_2543,N_1229);
and U6266 (N_6266,N_518,N_1612);
or U6267 (N_6267,N_699,N_3840);
nor U6268 (N_6268,N_2204,N_1919);
nand U6269 (N_6269,N_266,N_3839);
nand U6270 (N_6270,N_879,N_4314);
nor U6271 (N_6271,N_3156,N_3390);
nand U6272 (N_6272,N_1062,N_3310);
and U6273 (N_6273,N_4769,N_3891);
nand U6274 (N_6274,N_4310,N_2613);
nor U6275 (N_6275,N_162,N_4037);
nand U6276 (N_6276,N_3562,N_3146);
xor U6277 (N_6277,N_614,N_3248);
nand U6278 (N_6278,N_467,N_3026);
nand U6279 (N_6279,N_1797,N_4796);
xnor U6280 (N_6280,N_2522,N_2137);
nand U6281 (N_6281,N_463,N_3363);
xnor U6282 (N_6282,N_2019,N_2512);
nor U6283 (N_6283,N_681,N_3232);
xor U6284 (N_6284,N_4663,N_843);
or U6285 (N_6285,N_3680,N_4790);
or U6286 (N_6286,N_944,N_1816);
nand U6287 (N_6287,N_4175,N_365);
nand U6288 (N_6288,N_1857,N_3859);
and U6289 (N_6289,N_4690,N_1365);
and U6290 (N_6290,N_4639,N_2946);
nor U6291 (N_6291,N_2379,N_4916);
or U6292 (N_6292,N_2298,N_3162);
or U6293 (N_6293,N_1965,N_545);
xnor U6294 (N_6294,N_3202,N_308);
and U6295 (N_6295,N_4194,N_4451);
and U6296 (N_6296,N_2740,N_3347);
xor U6297 (N_6297,N_585,N_263);
or U6298 (N_6298,N_1445,N_1550);
or U6299 (N_6299,N_3612,N_567);
nand U6300 (N_6300,N_47,N_421);
nor U6301 (N_6301,N_4050,N_1571);
nand U6302 (N_6302,N_4997,N_1473);
and U6303 (N_6303,N_3877,N_3979);
xor U6304 (N_6304,N_2573,N_4211);
nand U6305 (N_6305,N_1561,N_2280);
nor U6306 (N_6306,N_2124,N_2004);
nand U6307 (N_6307,N_2642,N_2649);
or U6308 (N_6308,N_1412,N_4090);
nand U6309 (N_6309,N_3031,N_1507);
nor U6310 (N_6310,N_3997,N_3187);
xnor U6311 (N_6311,N_3011,N_4645);
or U6312 (N_6312,N_2747,N_1907);
xor U6313 (N_6313,N_2877,N_788);
nand U6314 (N_6314,N_268,N_438);
nor U6315 (N_6315,N_4338,N_2085);
or U6316 (N_6316,N_1178,N_1024);
nand U6317 (N_6317,N_3650,N_2584);
nor U6318 (N_6318,N_526,N_2167);
nor U6319 (N_6319,N_763,N_3623);
xor U6320 (N_6320,N_626,N_2405);
and U6321 (N_6321,N_338,N_2102);
and U6322 (N_6322,N_3119,N_3586);
or U6323 (N_6323,N_3163,N_744);
or U6324 (N_6324,N_1202,N_3892);
nor U6325 (N_6325,N_2743,N_4446);
nor U6326 (N_6326,N_3642,N_1118);
nand U6327 (N_6327,N_1059,N_3076);
nand U6328 (N_6328,N_2725,N_3166);
nor U6329 (N_6329,N_4333,N_3401);
or U6330 (N_6330,N_2040,N_2451);
nor U6331 (N_6331,N_1828,N_1669);
or U6332 (N_6332,N_4877,N_26);
xnor U6333 (N_6333,N_2260,N_4383);
and U6334 (N_6334,N_1054,N_2168);
xor U6335 (N_6335,N_806,N_1670);
xor U6336 (N_6336,N_4261,N_3109);
or U6337 (N_6337,N_2227,N_4199);
nand U6338 (N_6338,N_4910,N_2587);
nand U6339 (N_6339,N_3108,N_2307);
nor U6340 (N_6340,N_4563,N_606);
and U6341 (N_6341,N_3092,N_3408);
or U6342 (N_6342,N_1842,N_4589);
nor U6343 (N_6343,N_4466,N_60);
nor U6344 (N_6344,N_3856,N_780);
and U6345 (N_6345,N_4553,N_3378);
and U6346 (N_6346,N_2424,N_1671);
nand U6347 (N_6347,N_1791,N_946);
and U6348 (N_6348,N_4506,N_2180);
and U6349 (N_6349,N_3759,N_2160);
nor U6350 (N_6350,N_1865,N_4367);
nor U6351 (N_6351,N_1428,N_2643);
and U6352 (N_6352,N_2179,N_1228);
or U6353 (N_6353,N_3472,N_293);
nor U6354 (N_6354,N_4726,N_3557);
nor U6355 (N_6355,N_2900,N_883);
or U6356 (N_6356,N_156,N_2461);
and U6357 (N_6357,N_4447,N_2389);
or U6358 (N_6358,N_1194,N_4167);
xor U6359 (N_6359,N_1933,N_1653);
xnor U6360 (N_6360,N_4526,N_3084);
or U6361 (N_6361,N_2529,N_4841);
xor U6362 (N_6362,N_2271,N_4667);
and U6363 (N_6363,N_560,N_1044);
nor U6364 (N_6364,N_7,N_2069);
xnor U6365 (N_6365,N_2830,N_2390);
or U6366 (N_6366,N_4469,N_748);
xnor U6367 (N_6367,N_4266,N_1957);
xnor U6368 (N_6368,N_4044,N_1716);
nor U6369 (N_6369,N_1923,N_2254);
or U6370 (N_6370,N_2909,N_3533);
or U6371 (N_6371,N_4879,N_554);
xnor U6372 (N_6372,N_3072,N_765);
or U6373 (N_6373,N_2011,N_1462);
and U6374 (N_6374,N_3522,N_3674);
xor U6375 (N_6375,N_4842,N_1593);
nand U6376 (N_6376,N_3591,N_1663);
nor U6377 (N_6377,N_672,N_3559);
nand U6378 (N_6378,N_4432,N_3526);
or U6379 (N_6379,N_1756,N_3577);
xnor U6380 (N_6380,N_3666,N_2089);
nand U6381 (N_6381,N_3616,N_4098);
xor U6382 (N_6382,N_590,N_427);
xor U6383 (N_6383,N_2641,N_348);
or U6384 (N_6384,N_1774,N_770);
nor U6385 (N_6385,N_453,N_3824);
nand U6386 (N_6386,N_15,N_683);
xnor U6387 (N_6387,N_2735,N_11);
nand U6388 (N_6388,N_471,N_3339);
nand U6389 (N_6389,N_327,N_4389);
nand U6390 (N_6390,N_3993,N_3598);
or U6391 (N_6391,N_4164,N_1116);
and U6392 (N_6392,N_2164,N_3377);
nor U6393 (N_6393,N_1978,N_4802);
nand U6394 (N_6394,N_3927,N_241);
nand U6395 (N_6395,N_82,N_702);
or U6396 (N_6396,N_3096,N_497);
nand U6397 (N_6397,N_295,N_3656);
xnor U6398 (N_6398,N_3643,N_2825);
nor U6399 (N_6399,N_2667,N_4551);
nor U6400 (N_6400,N_4020,N_2976);
xnor U6401 (N_6401,N_4580,N_758);
or U6402 (N_6402,N_4134,N_287);
nand U6403 (N_6403,N_527,N_1090);
xor U6404 (N_6404,N_2284,N_3760);
nor U6405 (N_6405,N_3647,N_4355);
nor U6406 (N_6406,N_310,N_2072);
and U6407 (N_6407,N_1164,N_4683);
or U6408 (N_6408,N_1645,N_3488);
xor U6409 (N_6409,N_3221,N_2113);
and U6410 (N_6410,N_1804,N_2843);
or U6411 (N_6411,N_2493,N_3792);
or U6412 (N_6412,N_4852,N_4721);
nand U6413 (N_6413,N_1973,N_4742);
or U6414 (N_6414,N_510,N_4103);
xnor U6415 (N_6415,N_3804,N_3403);
nor U6416 (N_6416,N_3416,N_2620);
nand U6417 (N_6417,N_620,N_1020);
xor U6418 (N_6418,N_237,N_378);
and U6419 (N_6419,N_1718,N_950);
nand U6420 (N_6420,N_3345,N_4981);
nand U6421 (N_6421,N_2465,N_1516);
nand U6422 (N_6422,N_4092,N_4813);
xor U6423 (N_6423,N_1574,N_881);
nor U6424 (N_6424,N_4308,N_2575);
xnor U6425 (N_6425,N_2956,N_4377);
nor U6426 (N_6426,N_2467,N_4845);
and U6427 (N_6427,N_690,N_3614);
xor U6428 (N_6428,N_1668,N_265);
or U6429 (N_6429,N_335,N_1419);
nor U6430 (N_6430,N_1434,N_960);
nand U6431 (N_6431,N_4374,N_2347);
or U6432 (N_6432,N_940,N_1722);
and U6433 (N_6433,N_4471,N_2606);
nand U6434 (N_6434,N_3212,N_4830);
nand U6435 (N_6435,N_3135,N_3094);
or U6436 (N_6436,N_380,N_1591);
nor U6437 (N_6437,N_135,N_1266);
nor U6438 (N_6438,N_4133,N_1242);
xnor U6439 (N_6439,N_4320,N_4744);
xor U6440 (N_6440,N_694,N_180);
or U6441 (N_6441,N_4399,N_2509);
nor U6442 (N_6442,N_1813,N_4654);
nor U6443 (N_6443,N_1634,N_4388);
nor U6444 (N_6444,N_2027,N_3800);
or U6445 (N_6445,N_4507,N_2604);
or U6446 (N_6446,N_4461,N_4456);
nand U6447 (N_6447,N_1091,N_664);
xnor U6448 (N_6448,N_1165,N_1729);
and U6449 (N_6449,N_663,N_633);
and U6450 (N_6450,N_1586,N_2759);
or U6451 (N_6451,N_2863,N_3596);
xor U6452 (N_6452,N_164,N_4988);
xor U6453 (N_6453,N_703,N_1967);
xnor U6454 (N_6454,N_181,N_2464);
or U6455 (N_6455,N_710,N_239);
nand U6456 (N_6456,N_3313,N_346);
xor U6457 (N_6457,N_4870,N_2657);
and U6458 (N_6458,N_2966,N_3702);
and U6459 (N_6459,N_1400,N_3282);
or U6460 (N_6460,N_3737,N_1676);
or U6461 (N_6461,N_3713,N_2348);
xor U6462 (N_6462,N_2994,N_3511);
nand U6463 (N_6463,N_4819,N_830);
nor U6464 (N_6464,N_2972,N_2908);
nor U6465 (N_6465,N_644,N_531);
xnor U6466 (N_6466,N_3107,N_3485);
and U6467 (N_6467,N_3936,N_1283);
or U6468 (N_6468,N_1582,N_279);
and U6469 (N_6469,N_4472,N_3902);
nand U6470 (N_6470,N_1375,N_575);
nand U6471 (N_6471,N_2648,N_515);
nand U6472 (N_6472,N_3627,N_1296);
nand U6473 (N_6473,N_4223,N_4376);
and U6474 (N_6474,N_2844,N_4581);
xor U6475 (N_6475,N_4024,N_2263);
or U6476 (N_6476,N_3751,N_318);
xnor U6477 (N_6477,N_4329,N_1177);
or U6478 (N_6478,N_4284,N_2071);
nor U6479 (N_6479,N_2925,N_1128);
or U6480 (N_6480,N_2552,N_312);
nand U6481 (N_6481,N_2597,N_3908);
xnor U6482 (N_6482,N_1611,N_4055);
or U6483 (N_6483,N_4487,N_4618);
xor U6484 (N_6484,N_2382,N_2315);
and U6485 (N_6485,N_496,N_2039);
and U6486 (N_6486,N_3782,N_997);
xnor U6487 (N_6487,N_2356,N_4771);
xor U6488 (N_6488,N_2229,N_3083);
or U6489 (N_6489,N_818,N_1697);
or U6490 (N_6490,N_1689,N_1894);
and U6491 (N_6491,N_1262,N_4233);
nand U6492 (N_6492,N_3328,N_1373);
and U6493 (N_6493,N_2385,N_751);
or U6494 (N_6494,N_3406,N_95);
nand U6495 (N_6495,N_2050,N_2896);
nor U6496 (N_6496,N_13,N_1839);
nor U6497 (N_6497,N_4792,N_2541);
or U6498 (N_6498,N_4762,N_1329);
and U6499 (N_6499,N_3450,N_2933);
nor U6500 (N_6500,N_667,N_3005);
nor U6501 (N_6501,N_152,N_764);
xor U6502 (N_6502,N_1896,N_3709);
nor U6503 (N_6503,N_1892,N_1150);
xnor U6504 (N_6504,N_2490,N_4240);
or U6505 (N_6505,N_3662,N_2291);
xor U6506 (N_6506,N_1076,N_3193);
nor U6507 (N_6507,N_1040,N_414);
and U6508 (N_6508,N_3137,N_1491);
xor U6509 (N_6509,N_535,N_4221);
and U6510 (N_6510,N_1204,N_3599);
xor U6511 (N_6511,N_4658,N_4923);
nand U6512 (N_6512,N_3573,N_4345);
xnor U6513 (N_6513,N_2140,N_2777);
and U6514 (N_6514,N_668,N_2792);
nor U6515 (N_6515,N_3270,N_1066);
or U6516 (N_6516,N_4509,N_996);
xor U6517 (N_6517,N_2338,N_935);
xor U6518 (N_6518,N_2652,N_2817);
and U6519 (N_6519,N_3266,N_206);
xor U6520 (N_6520,N_4866,N_1476);
nand U6521 (N_6521,N_2673,N_328);
or U6522 (N_6522,N_1952,N_2195);
or U6523 (N_6523,N_3352,N_3506);
xor U6524 (N_6524,N_4362,N_1564);
xor U6525 (N_6525,N_3344,N_3157);
nand U6526 (N_6526,N_2221,N_3047);
nor U6527 (N_6527,N_4776,N_947);
xor U6528 (N_6528,N_247,N_3955);
and U6529 (N_6529,N_837,N_3545);
nand U6530 (N_6530,N_2905,N_698);
or U6531 (N_6531,N_2332,N_2717);
nand U6532 (N_6532,N_4803,N_4517);
nor U6533 (N_6533,N_2589,N_659);
xor U6534 (N_6534,N_4113,N_3730);
and U6535 (N_6535,N_587,N_3044);
nor U6536 (N_6536,N_1758,N_3838);
nor U6537 (N_6537,N_1297,N_4540);
xnor U6538 (N_6538,N_1167,N_2086);
nor U6539 (N_6539,N_2665,N_1652);
xnor U6540 (N_6540,N_4895,N_4687);
nand U6541 (N_6541,N_1786,N_68);
nand U6542 (N_6542,N_4574,N_2277);
and U6543 (N_6543,N_4915,N_4070);
and U6544 (N_6544,N_1039,N_4414);
xnor U6545 (N_6545,N_3351,N_2694);
xor U6546 (N_6546,N_523,N_4299);
nor U6547 (N_6547,N_2115,N_4516);
and U6548 (N_6548,N_3949,N_3400);
or U6549 (N_6549,N_4452,N_2076);
or U6550 (N_6550,N_3615,N_603);
nand U6551 (N_6551,N_939,N_2442);
nor U6552 (N_6552,N_325,N_3414);
nand U6553 (N_6553,N_4291,N_4614);
or U6554 (N_6554,N_2401,N_2691);
nand U6555 (N_6555,N_1360,N_1362);
and U6556 (N_6556,N_665,N_113);
or U6557 (N_6557,N_1056,N_1858);
or U6558 (N_6558,N_2238,N_227);
xor U6559 (N_6559,N_4584,N_3582);
or U6560 (N_6560,N_3852,N_280);
and U6561 (N_6561,N_528,N_3712);
nor U6562 (N_6562,N_1187,N_1733);
and U6563 (N_6563,N_3317,N_3735);
xor U6564 (N_6564,N_1316,N_298);
nor U6565 (N_6565,N_4758,N_921);
or U6566 (N_6566,N_3552,N_108);
nand U6567 (N_6567,N_176,N_533);
xor U6568 (N_6568,N_1853,N_1945);
xnor U6569 (N_6569,N_2403,N_3544);
xor U6570 (N_6570,N_2899,N_1583);
xor U6571 (N_6571,N_3874,N_4737);
xor U6572 (N_6572,N_2125,N_3802);
nor U6573 (N_6573,N_636,N_1063);
or U6574 (N_6574,N_4994,N_2870);
xnor U6575 (N_6575,N_2407,N_2892);
nor U6576 (N_6576,N_59,N_2339);
nand U6577 (N_6577,N_1160,N_599);
xnor U6578 (N_6578,N_4084,N_194);
nand U6579 (N_6579,N_579,N_3801);
nor U6580 (N_6580,N_4966,N_4503);
nand U6581 (N_6581,N_717,N_1636);
nor U6582 (N_6582,N_1141,N_1486);
xor U6583 (N_6583,N_3723,N_485);
and U6584 (N_6584,N_4971,N_1562);
or U6585 (N_6585,N_4586,N_4522);
and U6586 (N_6586,N_2159,N_4794);
or U6587 (N_6587,N_2112,N_1850);
and U6588 (N_6588,N_1944,N_3184);
nand U6589 (N_6589,N_199,N_1528);
or U6590 (N_6590,N_4334,N_4071);
xor U6591 (N_6591,N_4868,N_1112);
and U6592 (N_6592,N_413,N_1510);
nand U6593 (N_6593,N_3749,N_1422);
nand U6594 (N_6594,N_2096,N_3262);
and U6595 (N_6595,N_3236,N_4889);
xnor U6596 (N_6596,N_3734,N_1208);
nor U6597 (N_6597,N_2484,N_4766);
or U6598 (N_6598,N_4122,N_1985);
or U6599 (N_6599,N_2542,N_3444);
or U6600 (N_6600,N_2998,N_1792);
and U6601 (N_6601,N_4153,N_1153);
nor U6602 (N_6602,N_1966,N_1149);
and U6603 (N_6603,N_708,N_3882);
and U6604 (N_6604,N_3327,N_495);
or U6605 (N_6605,N_1193,N_3671);
nor U6606 (N_6606,N_4840,N_3549);
or U6607 (N_6607,N_987,N_1344);
or U6608 (N_6608,N_3089,N_1250);
nand U6609 (N_6609,N_1980,N_4990);
or U6610 (N_6610,N_3740,N_1181);
and U6611 (N_6611,N_1277,N_142);
nand U6612 (N_6612,N_2309,N_1097);
or U6613 (N_6613,N_2826,N_4897);
nor U6614 (N_6614,N_1333,N_3620);
nor U6615 (N_6615,N_4023,N_1206);
or U6616 (N_6616,N_4510,N_3531);
nor U6617 (N_6617,N_2707,N_4445);
xnor U6618 (N_6618,N_839,N_1705);
and U6619 (N_6619,N_2129,N_3148);
nor U6620 (N_6620,N_781,N_3825);
or U6621 (N_6621,N_3812,N_2602);
xnor U6622 (N_6622,N_2999,N_1891);
or U6623 (N_6623,N_482,N_4944);
nand U6624 (N_6624,N_4592,N_4913);
or U6625 (N_6625,N_4812,N_4074);
xnor U6626 (N_6626,N_1286,N_2108);
and U6627 (N_6627,N_307,N_4788);
and U6628 (N_6628,N_4245,N_524);
xor U6629 (N_6629,N_2148,N_1001);
nand U6630 (N_6630,N_4736,N_2360);
or U6631 (N_6631,N_3336,N_4328);
or U6632 (N_6632,N_3475,N_3717);
and U6633 (N_6633,N_1563,N_706);
and U6634 (N_6634,N_3974,N_1911);
nand U6635 (N_6635,N_1077,N_428);
nand U6636 (N_6636,N_2689,N_1248);
xor U6637 (N_6637,N_810,N_1821);
or U6638 (N_6638,N_3220,N_2156);
nor U6639 (N_6639,N_3041,N_2517);
xor U6640 (N_6640,N_4573,N_1332);
and U6641 (N_6641,N_2566,N_3296);
or U6642 (N_6642,N_1992,N_3480);
or U6643 (N_6643,N_512,N_1272);
and U6644 (N_6644,N_4833,N_3161);
or U6645 (N_6645,N_2216,N_4232);
nor U6646 (N_6646,N_4210,N_2483);
xnor U6647 (N_6647,N_2341,N_1079);
nor U6648 (N_6648,N_4943,N_2045);
nand U6649 (N_6649,N_4251,N_1683);
or U6650 (N_6650,N_2799,N_4984);
and U6651 (N_6651,N_4079,N_4034);
and U6652 (N_6652,N_4846,N_1532);
nor U6653 (N_6653,N_631,N_1320);
or U6654 (N_6654,N_2698,N_86);
and U6655 (N_6655,N_3767,N_876);
nand U6656 (N_6656,N_1105,N_402);
xor U6657 (N_6657,N_424,N_2661);
xnor U6658 (N_6658,N_1201,N_2441);
nand U6659 (N_6659,N_4282,N_1450);
nor U6660 (N_6660,N_3397,N_1702);
nand U6661 (N_6661,N_877,N_2329);
nor U6662 (N_6662,N_3422,N_2940);
and U6663 (N_6663,N_184,N_3217);
nor U6664 (N_6664,N_168,N_4427);
xnor U6665 (N_6665,N_278,N_2760);
nor U6666 (N_6666,N_2600,N_933);
xor U6667 (N_6667,N_4624,N_3738);
nand U6668 (N_6668,N_974,N_2247);
xor U6669 (N_6669,N_1080,N_258);
or U6670 (N_6670,N_2850,N_361);
nand U6671 (N_6671,N_925,N_2941);
nor U6672 (N_6672,N_4311,N_1263);
xor U6673 (N_6673,N_4293,N_916);
and U6674 (N_6674,N_3502,N_3019);
nand U6675 (N_6675,N_4936,N_3845);
xor U6676 (N_6676,N_2397,N_3565);
and U6677 (N_6677,N_2503,N_612);
nand U6678 (N_6678,N_4127,N_4278);
xnor U6679 (N_6679,N_4995,N_65);
xor U6680 (N_6680,N_2068,N_2252);
or U6681 (N_6681,N_1991,N_1309);
or U6682 (N_6682,N_3899,N_1443);
nand U6683 (N_6683,N_3837,N_3243);
nor U6684 (N_6684,N_1213,N_2022);
nor U6685 (N_6685,N_3071,N_4366);
xor U6686 (N_6686,N_4853,N_1140);
nand U6687 (N_6687,N_1485,N_4751);
nor U6688 (N_6688,N_1914,N_4003);
xor U6689 (N_6689,N_675,N_2544);
and U6690 (N_6690,N_1890,N_478);
nand U6691 (N_6691,N_3543,N_2533);
xnor U6692 (N_6692,N_3008,N_3);
and U6693 (N_6693,N_4847,N_1258);
and U6694 (N_6694,N_2881,N_2388);
or U6695 (N_6695,N_961,N_3383);
and U6696 (N_6696,N_3679,N_394);
and U6697 (N_6697,N_196,N_2603);
nor U6698 (N_6698,N_3018,N_844);
xor U6699 (N_6699,N_3358,N_1447);
and U6700 (N_6700,N_747,N_3224);
xnor U6701 (N_6701,N_1845,N_3246);
nor U6702 (N_6702,N_1849,N_3070);
xnor U6703 (N_6703,N_4460,N_2639);
or U6704 (N_6704,N_3410,N_1084);
nand U6705 (N_6705,N_1970,N_2035);
xor U6706 (N_6706,N_1661,N_4638);
or U6707 (N_6707,N_2995,N_605);
or U6708 (N_6708,N_984,N_2985);
or U6709 (N_6709,N_1179,N_3629);
or U6710 (N_6710,N_2879,N_2948);
or U6711 (N_6711,N_4005,N_1261);
nand U6712 (N_6712,N_1599,N_4312);
xor U6713 (N_6713,N_4206,N_3940);
xnor U6714 (N_6714,N_24,N_430);
nor U6715 (N_6715,N_2762,N_2199);
nor U6716 (N_6716,N_1270,N_2521);
xor U6717 (N_6717,N_738,N_3625);
and U6718 (N_6718,N_3411,N_1437);
nor U6719 (N_6719,N_914,N_2556);
or U6720 (N_6720,N_3152,N_3954);
xnor U6721 (N_6721,N_294,N_3512);
and U6722 (N_6722,N_505,N_45);
nor U6723 (N_6723,N_4727,N_1009);
or U6724 (N_6724,N_257,N_3283);
and U6725 (N_6725,N_3587,N_1710);
or U6726 (N_6726,N_322,N_816);
or U6727 (N_6727,N_4420,N_1658);
and U6728 (N_6728,N_4306,N_4977);
nor U6729 (N_6729,N_1148,N_1374);
xor U6730 (N_6730,N_25,N_217);
or U6731 (N_6731,N_795,N_4765);
nor U6732 (N_6732,N_4538,N_2586);
nor U6733 (N_6733,N_360,N_2942);
nor U6734 (N_6734,N_4711,N_3255);
or U6735 (N_6735,N_500,N_1681);
nand U6736 (N_6736,N_4138,N_4820);
xor U6737 (N_6737,N_334,N_1656);
nand U6738 (N_6738,N_2813,N_3139);
and U6739 (N_6739,N_4746,N_4824);
nor U6740 (N_6740,N_4196,N_938);
and U6741 (N_6741,N_4464,N_2449);
nand U6742 (N_6742,N_122,N_1209);
or U6743 (N_6743,N_1107,N_127);
or U6744 (N_6744,N_4576,N_1897);
xor U6745 (N_6745,N_1686,N_104);
and U6746 (N_6746,N_724,N_3677);
xnor U6747 (N_6747,N_4217,N_3498);
nand U6748 (N_6748,N_4925,N_4405);
and U6749 (N_6749,N_2384,N_3941);
or U6750 (N_6750,N_1925,N_1961);
xnor U6751 (N_6751,N_264,N_2983);
nand U6752 (N_6752,N_4391,N_1901);
or U6753 (N_6753,N_2225,N_2742);
xnor U6754 (N_6754,N_838,N_3001);
and U6755 (N_6755,N_3320,N_1314);
or U6756 (N_6756,N_2511,N_4953);
nor U6757 (N_6757,N_3067,N_712);
xor U6758 (N_6758,N_3658,N_3449);
xnor U6759 (N_6759,N_994,N_1006);
and U6760 (N_6760,N_1569,N_919);
or U6761 (N_6761,N_1834,N_3817);
xnor U6762 (N_6762,N_3798,N_2438);
nand U6763 (N_6763,N_4422,N_2818);
and U6764 (N_6764,N_249,N_4956);
or U6765 (N_6765,N_1108,N_3293);
or U6766 (N_6766,N_3884,N_1903);
and U6767 (N_6767,N_2766,N_835);
or U6768 (N_6768,N_865,N_4949);
nand U6769 (N_6769,N_3301,N_2534);
nand U6770 (N_6770,N_713,N_2162);
and U6771 (N_6771,N_1829,N_3850);
or U6772 (N_6772,N_2931,N_2894);
nand U6773 (N_6773,N_662,N_4378);
or U6774 (N_6774,N_1222,N_4316);
xor U6775 (N_6775,N_370,N_3494);
nand U6776 (N_6776,N_3866,N_1413);
nor U6777 (N_6777,N_1711,N_3271);
nor U6778 (N_6778,N_4280,N_434);
or U6779 (N_6779,N_1088,N_4554);
nand U6780 (N_6780,N_1101,N_4582);
nor U6781 (N_6781,N_4575,N_2723);
and U6782 (N_6782,N_544,N_3042);
and U6783 (N_6783,N_1769,N_3214);
nor U6784 (N_6784,N_1924,N_716);
nor U6785 (N_6785,N_3396,N_4235);
or U6786 (N_6786,N_4854,N_2787);
xor U6787 (N_6787,N_2134,N_1785);
xnor U6788 (N_6788,N_2243,N_1674);
and U6789 (N_6789,N_754,N_3939);
xnor U6790 (N_6790,N_1755,N_3744);
nor U6791 (N_6791,N_4613,N_678);
nand U6792 (N_6792,N_4083,N_1253);
xor U6793 (N_6793,N_658,N_3275);
or U6794 (N_6794,N_2647,N_3395);
nor U6795 (N_6795,N_688,N_2361);
or U6796 (N_6796,N_771,N_4501);
nor U6797 (N_6797,N_1439,N_2494);
and U6798 (N_6798,N_4587,N_1356);
nand U6799 (N_6799,N_451,N_1082);
and U6800 (N_6800,N_4861,N_4057);
nand U6801 (N_6801,N_3425,N_1353);
nand U6802 (N_6802,N_499,N_4434);
nor U6803 (N_6803,N_4713,N_1874);
and U6804 (N_6804,N_1899,N_4606);
or U6805 (N_6805,N_1754,N_3971);
or U6806 (N_6806,N_1008,N_4692);
nor U6807 (N_6807,N_3871,N_562);
nand U6808 (N_6808,N_4786,N_3307);
nor U6809 (N_6809,N_2947,N_2185);
xnor U6810 (N_6810,N_4716,N_1712);
nand U6811 (N_6811,N_1488,N_4468);
nor U6812 (N_6812,N_4844,N_2141);
nor U6813 (N_6813,N_1425,N_2773);
nor U6814 (N_6814,N_3808,N_2654);
nor U6815 (N_6815,N_4062,N_4428);
xnor U6816 (N_6816,N_3115,N_4449);
nor U6817 (N_6817,N_2802,N_4018);
and U6818 (N_6818,N_860,N_311);
nor U6819 (N_6819,N_2266,N_1512);
or U6820 (N_6820,N_1133,N_288);
xor U6821 (N_6821,N_3082,N_1788);
nand U6822 (N_6822,N_3906,N_670);
nor U6823 (N_6823,N_1237,N_2834);
or U6824 (N_6824,N_356,N_1022);
nand U6825 (N_6825,N_4228,N_4941);
or U6826 (N_6826,N_943,N_186);
nor U6827 (N_6827,N_1317,N_2337);
xor U6828 (N_6828,N_4375,N_4975);
or U6829 (N_6829,N_2632,N_1831);
nor U6830 (N_6830,N_275,N_3053);
xor U6831 (N_6831,N_351,N_2414);
or U6832 (N_6832,N_4918,N_1078);
nand U6833 (N_6833,N_3764,N_2614);
xnor U6834 (N_6834,N_2915,N_1368);
xnor U6835 (N_6835,N_1043,N_1103);
xor U6836 (N_6836,N_2727,N_784);
nand U6837 (N_6837,N_1655,N_2345);
nor U6838 (N_6838,N_2796,N_3780);
xnor U6839 (N_6839,N_539,N_846);
nor U6840 (N_6840,N_1700,N_2749);
nor U6841 (N_6841,N_3497,N_1565);
xor U6842 (N_6842,N_529,N_2919);
nor U6843 (N_6843,N_3235,N_853);
xnor U6844 (N_6844,N_924,N_4482);
and U6845 (N_6845,N_2856,N_2906);
nand U6846 (N_6846,N_546,N_2);
nand U6847 (N_6847,N_42,N_2897);
or U6848 (N_6848,N_4303,N_559);
and U6849 (N_6849,N_911,N_2355);
and U6850 (N_6850,N_1223,N_2574);
or U6851 (N_6851,N_746,N_1640);
nor U6852 (N_6852,N_3256,N_1311);
nor U6853 (N_6853,N_2750,N_3821);
nor U6854 (N_6854,N_2571,N_2326);
xnor U6855 (N_6855,N_352,N_1906);
or U6856 (N_6856,N_1806,N_558);
and U6857 (N_6857,N_1870,N_2145);
or U6858 (N_6858,N_949,N_1337);
and U6859 (N_6859,N_2318,N_1856);
and U6860 (N_6860,N_1879,N_2282);
xnor U6861 (N_6861,N_4358,N_630);
xnor U6862 (N_6862,N_4755,N_3178);
xnor U6863 (N_6863,N_3807,N_1433);
and U6864 (N_6864,N_1183,N_3346);
and U6865 (N_6865,N_4561,N_4729);
and U6866 (N_6866,N_4615,N_4520);
nor U6867 (N_6867,N_3470,N_2259);
and U6868 (N_6868,N_3398,N_1748);
nand U6869 (N_6869,N_2400,N_2166);
and U6870 (N_6870,N_27,N_4347);
and U6871 (N_6871,N_2845,N_556);
nand U6872 (N_6872,N_2922,N_8);
xor U6873 (N_6873,N_880,N_733);
nand U6874 (N_6874,N_1303,N_2567);
xor U6875 (N_6875,N_2220,N_3079);
nor U6876 (N_6876,N_4102,N_2336);
or U6877 (N_6877,N_904,N_1735);
xor U6878 (N_6878,N_4653,N_4396);
nor U6879 (N_6879,N_2852,N_1410);
or U6880 (N_6880,N_1672,N_359);
xor U6881 (N_6881,N_2457,N_3312);
nor U6882 (N_6882,N_2821,N_2426);
xnor U6883 (N_6883,N_1282,N_4791);
xnor U6884 (N_6884,N_2969,N_3705);
or U6885 (N_6885,N_3326,N_2417);
nor U6886 (N_6886,N_3918,N_582);
and U6887 (N_6887,N_2299,N_1156);
or U6888 (N_6888,N_1624,N_813);
nand U6889 (N_6889,N_809,N_3199);
nor U6890 (N_6890,N_3147,N_141);
and U6891 (N_6891,N_3739,N_4629);
nor U6892 (N_6892,N_3142,N_4294);
nand U6893 (N_6893,N_2425,N_3438);
nand U6894 (N_6894,N_3366,N_2549);
or U6895 (N_6895,N_4633,N_1524);
or U6896 (N_6896,N_3796,N_2920);
xnor U6897 (N_6897,N_1930,N_2849);
xor U6898 (N_6898,N_625,N_1523);
nor U6899 (N_6899,N_2043,N_1041);
or U6900 (N_6900,N_2588,N_4600);
and U6901 (N_6901,N_392,N_2721);
or U6902 (N_6902,N_990,N_187);
nand U6903 (N_6903,N_3793,N_2083);
nor U6904 (N_6904,N_3249,N_1053);
or U6905 (N_6905,N_321,N_2103);
xnor U6906 (N_6906,N_2756,N_832);
nor U6907 (N_6907,N_1815,N_538);
and U6908 (N_6908,N_429,N_3451);
nor U6909 (N_6909,N_2563,N_1200);
xnor U6910 (N_6910,N_673,N_4529);
nand U6911 (N_6911,N_598,N_4126);
or U6912 (N_6912,N_3267,N_4904);
nor U6913 (N_6913,N_4896,N_339);
xnor U6914 (N_6914,N_3237,N_4289);
xnor U6915 (N_6915,N_2139,N_4421);
nand U6916 (N_6916,N_4053,N_4086);
nor U6917 (N_6917,N_4531,N_4993);
or U6918 (N_6918,N_1036,N_4185);
and U6919 (N_6919,N_1139,N_1115);
or U6920 (N_6920,N_4348,N_4781);
nor U6921 (N_6921,N_4453,N_4124);
nand U6922 (N_6922,N_3321,N_296);
nand U6923 (N_6923,N_4593,N_3805);
or U6924 (N_6924,N_1741,N_4601);
xnor U6925 (N_6925,N_4048,N_2865);
xnor U6926 (N_6926,N_4650,N_2666);
xnor U6927 (N_6927,N_954,N_2036);
or U6928 (N_6928,N_3948,N_3822);
and U6929 (N_6929,N_2477,N_898);
or U6930 (N_6930,N_4909,N_3503);
and U6931 (N_6931,N_4850,N_2518);
and U6932 (N_6932,N_4013,N_1197);
or U6933 (N_6933,N_2662,N_379);
or U6934 (N_6934,N_2427,N_4322);
nand U6935 (N_6935,N_2065,N_1724);
xor U6936 (N_6936,N_259,N_1873);
and U6937 (N_6937,N_2680,N_807);
nor U6938 (N_6938,N_1620,N_208);
or U6939 (N_6939,N_2026,N_4502);
and U6940 (N_6940,N_1927,N_4100);
or U6941 (N_6941,N_1381,N_35);
nor U6942 (N_6942,N_2269,N_4270);
or U6943 (N_6943,N_4315,N_3539);
and U6944 (N_6944,N_1922,N_3099);
or U6945 (N_6945,N_1950,N_4433);
nand U6946 (N_6946,N_214,N_3145);
and U6947 (N_6947,N_4804,N_600);
nand U6948 (N_6948,N_3234,N_3914);
and U6949 (N_6949,N_2256,N_2226);
nand U6950 (N_6950,N_1011,N_3183);
nand U6951 (N_6951,N_304,N_3774);
and U6952 (N_6952,N_4360,N_1065);
and U6953 (N_6953,N_1589,N_3844);
or U6954 (N_6954,N_4395,N_1409);
or U6955 (N_6955,N_3039,N_776);
nand U6956 (N_6956,N_2536,N_759);
nand U6957 (N_6957,N_811,N_1833);
nand U6958 (N_6958,N_3540,N_417);
nor U6959 (N_6959,N_2087,N_2572);
and U6960 (N_6960,N_3897,N_4974);
xnor U6961 (N_6961,N_1948,N_2283);
nand U6962 (N_6962,N_2928,N_1744);
xnor U6963 (N_6963,N_3775,N_2635);
nor U6964 (N_6964,N_3046,N_465);
nor U6965 (N_6965,N_4999,N_198);
or U6966 (N_6966,N_583,N_1715);
nor U6967 (N_6967,N_1182,N_955);
nor U6968 (N_6968,N_922,N_4566);
xnor U6969 (N_6969,N_2540,N_618);
and U6970 (N_6970,N_4337,N_3374);
and U6971 (N_6971,N_1968,N_2053);
nand U6972 (N_6972,N_3098,N_2395);
and U6973 (N_6973,N_2038,N_2546);
nor U6974 (N_6974,N_2772,N_4049);
nand U6975 (N_6975,N_4740,N_729);
nand U6976 (N_6976,N_2585,N_433);
or U6977 (N_6977,N_1081,N_740);
nor U6978 (N_6978,N_3483,N_4166);
xnor U6979 (N_6979,N_53,N_3222);
and U6980 (N_6980,N_4041,N_2930);
and U6981 (N_6981,N_982,N_1567);
and U6982 (N_6982,N_2555,N_3848);
nor U6983 (N_6983,N_3982,N_4777);
nand U6984 (N_6984,N_4677,N_2525);
nor U6985 (N_6985,N_2251,N_2789);
nand U6986 (N_6986,N_3644,N_3508);
xnor U6987 (N_6987,N_4372,N_151);
and U6988 (N_6988,N_4125,N_3736);
nand U6989 (N_6989,N_4655,N_2189);
nand U6990 (N_6990,N_75,N_4419);
nor U6991 (N_6991,N_2175,N_4555);
or U6992 (N_6992,N_931,N_2420);
xor U6993 (N_6993,N_4708,N_1810);
or U6994 (N_6994,N_1590,N_3029);
or U6995 (N_6995,N_4225,N_4782);
nand U6996 (N_6996,N_4609,N_4224);
or U6997 (N_6997,N_3888,N_2893);
and U6998 (N_6998,N_2150,N_1449);
or U6999 (N_6999,N_1659,N_1621);
nand U7000 (N_7000,N_231,N_487);
and U7001 (N_7001,N_3883,N_315);
nor U7002 (N_7002,N_3207,N_2404);
and U7003 (N_7003,N_549,N_2878);
nand U7004 (N_7004,N_2640,N_1475);
and U7005 (N_7005,N_1154,N_2353);
xnor U7006 (N_7006,N_3763,N_1195);
and U7007 (N_7007,N_1255,N_173);
nor U7008 (N_7008,N_2982,N_4627);
xor U7009 (N_7009,N_2047,N_4179);
or U7010 (N_7010,N_2376,N_4873);
and U7011 (N_7011,N_1048,N_1578);
or U7012 (N_7012,N_4950,N_1094);
nand U7013 (N_7013,N_1256,N_50);
nand U7014 (N_7014,N_4937,N_594);
nand U7015 (N_7015,N_707,N_514);
or U7016 (N_7016,N_3661,N_1260);
xor U7017 (N_7017,N_3867,N_2748);
and U7018 (N_7018,N_4283,N_2419);
xor U7019 (N_7019,N_3458,N_4732);
or U7020 (N_7020,N_2520,N_4286);
nor U7021 (N_7021,N_1306,N_2631);
nand U7022 (N_7022,N_4527,N_1188);
nor U7023 (N_7023,N_3513,N_3676);
or U7024 (N_7024,N_4415,N_3687);
and U7025 (N_7025,N_2209,N_408);
or U7026 (N_7026,N_3829,N_2317);
and U7027 (N_7027,N_3710,N_953);
nand U7028 (N_7028,N_2776,N_4448);
nor U7029 (N_7029,N_646,N_1352);
nand U7030 (N_7030,N_3925,N_4011);
or U7031 (N_7031,N_2971,N_3505);
nand U7032 (N_7032,N_3781,N_4253);
and U7033 (N_7033,N_1032,N_4678);
or U7034 (N_7034,N_3570,N_4443);
nor U7035 (N_7035,N_1527,N_858);
or U7036 (N_7036,N_3937,N_1335);
or U7037 (N_7037,N_2871,N_2466);
nor U7038 (N_7038,N_1691,N_1503);
or U7039 (N_7039,N_484,N_739);
xnor U7040 (N_7040,N_3208,N_37);
xnor U7041 (N_7041,N_2473,N_116);
nand U7042 (N_7042,N_123,N_2122);
xnor U7043 (N_7043,N_4630,N_1988);
nor U7044 (N_7044,N_4730,N_2371);
nor U7045 (N_7045,N_1106,N_701);
and U7046 (N_7046,N_377,N_3622);
and U7047 (N_7047,N_826,N_2358);
nand U7048 (N_7048,N_1315,N_4307);
xnor U7049 (N_7049,N_3045,N_1694);
xnor U7050 (N_7050,N_1018,N_637);
nor U7051 (N_7051,N_1246,N_4264);
or U7052 (N_7052,N_3529,N_2319);
nor U7053 (N_7053,N_2712,N_1233);
xnor U7054 (N_7054,N_2579,N_3880);
and U7055 (N_7055,N_3371,N_387);
nor U7056 (N_7056,N_1555,N_3960);
xor U7057 (N_7057,N_4112,N_3589);
nand U7058 (N_7058,N_1910,N_4647);
and U7059 (N_7059,N_2331,N_2234);
xor U7060 (N_7060,N_783,N_2869);
nand U7061 (N_7061,N_503,N_4163);
nor U7062 (N_7062,N_3375,N_193);
xor U7063 (N_7063,N_1708,N_1762);
or U7064 (N_7064,N_98,N_3182);
and U7065 (N_7065,N_3233,N_133);
nand U7066 (N_7066,N_4890,N_4104);
or U7067 (N_7067,N_2048,N_689);
nor U7068 (N_7068,N_3534,N_1704);
xnor U7069 (N_7069,N_448,N_2754);
nor U7070 (N_7070,N_4883,N_1259);
nand U7071 (N_7071,N_1639,N_755);
xnor U7072 (N_7072,N_4664,N_867);
and U7073 (N_7073,N_4862,N_121);
xnor U7074 (N_7074,N_1543,N_653);
nand U7075 (N_7075,N_319,N_4972);
and U7076 (N_7076,N_4903,N_1752);
nor U7077 (N_7077,N_509,N_2513);
and U7078 (N_7078,N_1113,N_4893);
xnor U7079 (N_7079,N_3368,N_1350);
or U7080 (N_7080,N_3923,N_745);
and U7081 (N_7081,N_4135,N_2391);
xor U7082 (N_7082,N_1680,N_1191);
and U7083 (N_7083,N_1943,N_292);
xor U7084 (N_7084,N_3981,N_1432);
and U7085 (N_7085,N_1244,N_3086);
xnor U7086 (N_7086,N_2991,N_4350);
or U7087 (N_7087,N_4885,N_1535);
nand U7088 (N_7088,N_2213,N_3376);
nor U7089 (N_7089,N_563,N_131);
nor U7090 (N_7090,N_2851,N_228);
xor U7091 (N_7091,N_756,N_170);
xor U7092 (N_7092,N_3597,N_2716);
xor U7093 (N_7093,N_1699,N_1886);
xor U7094 (N_7094,N_980,N_2924);
nor U7095 (N_7095,N_1987,N_1466);
and U7096 (N_7096,N_3309,N_4607);
and U7097 (N_7097,N_486,N_3305);
and U7098 (N_7098,N_4806,N_1730);
xor U7099 (N_7099,N_3649,N_114);
or U7100 (N_7100,N_1688,N_2889);
and U7101 (N_7101,N_1628,N_3648);
nand U7102 (N_7102,N_332,N_3389);
nand U7103 (N_7103,N_2797,N_1321);
or U7104 (N_7104,N_331,N_191);
nor U7105 (N_7105,N_2526,N_3264);
xor U7106 (N_7106,N_3007,N_4353);
xnor U7107 (N_7107,N_4021,N_3909);
nor U7108 (N_7108,N_3665,N_4351);
nor U7109 (N_7109,N_1778,N_4567);
xnor U7110 (N_7110,N_2239,N_4012);
and U7111 (N_7111,N_337,N_3746);
nor U7112 (N_7112,N_1247,N_2278);
nand U7113 (N_7113,N_1558,N_2439);
or U7114 (N_7114,N_4881,N_1241);
nor U7115 (N_7115,N_1881,N_3404);
nor U7116 (N_7116,N_2430,N_986);
or U7117 (N_7117,N_4557,N_58);
nand U7118 (N_7118,N_383,N_4426);
nand U7119 (N_7119,N_3412,N_1074);
or U7120 (N_7120,N_1176,N_2997);
or U7121 (N_7121,N_3476,N_817);
nand U7122 (N_7122,N_4801,N_1525);
nor U7123 (N_7123,N_4137,N_4748);
or U7124 (N_7124,N_3860,N_3322);
or U7125 (N_7125,N_3290,N_4735);
xor U7126 (N_7126,N_218,N_2783);
nand U7127 (N_7127,N_814,N_4621);
xor U7128 (N_7128,N_1603,N_1205);
nand U7129 (N_7129,N_3302,N_4047);
nor U7130 (N_7130,N_329,N_2874);
or U7131 (N_7131,N_2109,N_4929);
xnor U7132 (N_7132,N_2887,N_2853);
nand U7133 (N_7133,N_4143,N_1789);
nand U7134 (N_7134,N_3081,N_4983);
or U7135 (N_7135,N_2262,N_4770);
nor U7136 (N_7136,N_2452,N_588);
and U7137 (N_7137,N_3564,N_4955);
xnor U7138 (N_7138,N_3967,N_2653);
nor U7139 (N_7139,N_1920,N_1830);
nand U7140 (N_7140,N_2862,N_46);
nand U7141 (N_7141,N_2423,N_2734);
and U7142 (N_7142,N_2052,N_1584);
and U7143 (N_7143,N_2032,N_1826);
and U7144 (N_7144,N_1977,N_2005);
and U7145 (N_7145,N_3010,N_449);
nand U7146 (N_7146,N_4884,N_1454);
or U7147 (N_7147,N_415,N_1713);
nor U7148 (N_7148,N_4341,N_1626);
nand U7149 (N_7149,N_3594,N_597);
or U7150 (N_7150,N_992,N_685);
and U7151 (N_7151,N_1889,N_314);
xor U7152 (N_7152,N_4161,N_2963);
and U7153 (N_7153,N_3150,N_1750);
nand U7154 (N_7154,N_1667,N_1005);
xnor U7155 (N_7155,N_224,N_4822);
nor U7156 (N_7156,N_4602,N_4052);
xnor U7157 (N_7157,N_2170,N_1227);
nor U7158 (N_7158,N_3167,N_993);
or U7159 (N_7159,N_4900,N_1397);
and U7160 (N_7160,N_1982,N_4946);
nand U7161 (N_7161,N_1784,N_1415);
nand U7162 (N_7162,N_2409,N_958);
or U7163 (N_7163,N_2245,N_3765);
and U7164 (N_7164,N_200,N_1251);
and U7165 (N_7165,N_1484,N_343);
nor U7166 (N_7166,N_2835,N_3527);
and U7167 (N_7167,N_2822,N_3439);
and U7168 (N_7168,N_419,N_3968);
nor U7169 (N_7169,N_3348,N_410);
xor U7170 (N_7170,N_119,N_4131);
or U7171 (N_7171,N_4798,N_1703);
xor U7172 (N_7172,N_779,N_2290);
nor U7173 (N_7173,N_3834,N_3151);
nand U7174 (N_7174,N_3833,N_4111);
nor U7175 (N_7175,N_3460,N_2446);
or U7176 (N_7176,N_4105,N_1514);
or U7177 (N_7177,N_3413,N_2396);
xor U7178 (N_7178,N_1393,N_734);
and U7179 (N_7179,N_4986,N_3491);
or U7180 (N_7180,N_2078,N_1408);
nand U7181 (N_7181,N_3050,N_3014);
or U7182 (N_7182,N_4828,N_647);
and U7183 (N_7183,N_3519,N_1983);
nor U7184 (N_7184,N_4922,N_2352);
xnor U7185 (N_7185,N_3215,N_2029);
xor U7186 (N_7186,N_4641,N_2769);
and U7187 (N_7187,N_1219,N_2515);
or U7188 (N_7188,N_4821,N_3514);
and U7189 (N_7189,N_4229,N_3913);
xor U7190 (N_7190,N_1468,N_2934);
nand U7191 (N_7191,N_4227,N_4924);
or U7192 (N_7192,N_124,N_812);
and U7193 (N_7193,N_866,N_968);
xnor U7194 (N_7194,N_301,N_640);
nand U7195 (N_7195,N_3956,N_2907);
and U7196 (N_7196,N_2607,N_977);
and U7197 (N_7197,N_3473,N_823);
and U7198 (N_7198,N_4450,N_2276);
xnor U7199 (N_7199,N_4107,N_1508);
and U7200 (N_7200,N_396,N_4437);
and U7201 (N_7201,N_2891,N_2343);
nand U7202 (N_7202,N_1104,N_4814);
nand U7203 (N_7203,N_491,N_2074);
nand U7204 (N_7204,N_1446,N_4309);
nand U7205 (N_7205,N_2008,N_3878);
and U7206 (N_7206,N_4442,N_2782);
and U7207 (N_7207,N_2706,N_303);
nor U7208 (N_7208,N_80,N_3698);
nor U7209 (N_7209,N_4783,N_1198);
and U7210 (N_7210,N_3608,N_300);
xor U7211 (N_7211,N_3995,N_3592);
nor U7212 (N_7212,N_766,N_3700);
nor U7213 (N_7213,N_4772,N_3630);
nor U7214 (N_7214,N_3904,N_1501);
or U7215 (N_7215,N_344,N_508);
nand U7216 (N_7216,N_3159,N_4154);
nand U7217 (N_7217,N_2497,N_3194);
and U7218 (N_7218,N_2811,N_1675);
nor U7219 (N_7219,N_2155,N_1949);
and U7220 (N_7220,N_3653,N_432);
and U7221 (N_7221,N_824,N_3179);
nand U7222 (N_7222,N_4404,N_1417);
xnor U7223 (N_7223,N_2077,N_1588);
or U7224 (N_7224,N_4603,N_3681);
xor U7225 (N_7225,N_3538,N_1969);
and U7226 (N_7226,N_431,N_1092);
and U7227 (N_7227,N_3386,N_150);
nor U7228 (N_7228,N_21,N_3501);
xor U7229 (N_7229,N_4038,N_2429);
xor U7230 (N_7230,N_250,N_3862);
or U7231 (N_7231,N_1777,N_4571);
xor U7232 (N_7232,N_711,N_907);
xor U7233 (N_7233,N_1301,N_4403);
nor U7234 (N_7234,N_1064,N_1117);
xor U7235 (N_7235,N_2528,N_2000);
or U7236 (N_7236,N_985,N_3694);
or U7237 (N_7237,N_4,N_1377);
or U7238 (N_7238,N_851,N_306);
nor U7239 (N_7239,N_401,N_4523);
and U7240 (N_7240,N_3285,N_821);
nand U7241 (N_7241,N_3890,N_654);
and U7242 (N_7242,N_4335,N_4759);
nand U7243 (N_7243,N_721,N_3131);
or U7244 (N_7244,N_932,N_3818);
nor U7245 (N_7245,N_2088,N_2279);
and U7246 (N_7246,N_576,N_4340);
nor U7247 (N_7247,N_3990,N_1477);
or U7248 (N_7248,N_2253,N_4056);
nor U7249 (N_7249,N_4060,N_4987);
nand U7250 (N_7250,N_1291,N_2470);
nor U7251 (N_7251,N_1013,N_3708);
and U7252 (N_7252,N_906,N_639);
and U7253 (N_7253,N_3431,N_2911);
xnor U7254 (N_7254,N_29,N_3550);
xor U7255 (N_7255,N_3567,N_4533);
or U7256 (N_7256,N_2791,N_2217);
nor U7257 (N_7257,N_1649,N_3027);
and U7258 (N_7258,N_4147,N_1307);
xnor U7259 (N_7259,N_1541,N_3791);
xor U7260 (N_7260,N_4205,N_3381);
and U7261 (N_7261,N_1841,N_3279);
nand U7262 (N_7262,N_3992,N_2031);
nor U7263 (N_7263,N_1860,N_1868);
nand U7264 (N_7264,N_4483,N_3535);
and U7265 (N_7265,N_366,N_416);
and U7266 (N_7266,N_2708,N_624);
or U7267 (N_7267,N_4519,N_4722);
nand U7268 (N_7268,N_3090,N_3789);
xnor U7269 (N_7269,N_2846,N_4017);
and U7270 (N_7270,N_3684,N_2875);
or U7271 (N_7271,N_3036,N_443);
and U7272 (N_7272,N_1089,N_4585);
nand U7273 (N_7273,N_4767,N_928);
and U7274 (N_7274,N_2190,N_2142);
xnor U7275 (N_7275,N_2214,N_4559);
or U7276 (N_7276,N_4676,N_2601);
or U7277 (N_7277,N_4784,N_3524);
xnor U7278 (N_7278,N_4646,N_4398);
nor U7279 (N_7279,N_403,N_3747);
xor U7280 (N_7280,N_2628,N_2801);
or U7281 (N_7281,N_4474,N_3197);
nor U7282 (N_7282,N_3762,N_4188);
xnor U7283 (N_7283,N_1928,N_2060);
and U7284 (N_7284,N_1554,N_3112);
or U7285 (N_7285,N_1727,N_1500);
xnor U7286 (N_7286,N_1587,N_648);
or U7287 (N_7287,N_1995,N_4470);
nand U7288 (N_7288,N_4579,N_3619);
xnor U7289 (N_7289,N_1557,N_3864);
nor U7290 (N_7290,N_4128,N_1878);
nor U7291 (N_7291,N_1794,N_3689);
and U7292 (N_7292,N_4343,N_1917);
nor U7293 (N_7293,N_1288,N_4504);
and U7294 (N_7294,N_908,N_1546);
xnor U7295 (N_7295,N_4560,N_1893);
nand U7296 (N_7296,N_2831,N_2746);
xnor U7297 (N_7297,N_3568,N_3688);
nand U7298 (N_7298,N_341,N_1707);
or U7299 (N_7299,N_4703,N_4292);
or U7300 (N_7300,N_246,N_3664);
and U7301 (N_7301,N_39,N_3280);
and U7302 (N_7302,N_3489,N_1632);
nor U7303 (N_7303,N_3959,N_3088);
nor U7304 (N_7304,N_363,N_2537);
or U7305 (N_7305,N_2006,N_895);
and U7306 (N_7306,N_4865,N_317);
nand U7307 (N_7307,N_4768,N_4485);
and U7308 (N_7308,N_1120,N_3835);
and U7309 (N_7309,N_2075,N_2625);
nand U7310 (N_7310,N_903,N_4298);
nand U7311 (N_7311,N_3441,N_3430);
nand U7312 (N_7312,N_3841,N_2729);
nand U7313 (N_7313,N_4668,N_937);
nor U7314 (N_7314,N_412,N_4932);
nor U7315 (N_7315,N_2375,N_2992);
or U7316 (N_7316,N_1979,N_3138);
nand U7317 (N_7317,N_2548,N_1109);
or U7318 (N_7318,N_2795,N_1135);
and U7319 (N_7319,N_905,N_3445);
nor U7320 (N_7320,N_143,N_2860);
nor U7321 (N_7321,N_4500,N_4596);
and U7322 (N_7322,N_957,N_2726);
xnor U7323 (N_7323,N_1884,N_4902);
and U7324 (N_7324,N_22,N_4672);
and U7325 (N_7325,N_1882,N_2990);
and U7326 (N_7326,N_3379,N_3065);
xor U7327 (N_7327,N_4764,N_3427);
and U7328 (N_7328,N_2095,N_4891);
and U7329 (N_7329,N_395,N_3778);
or U7330 (N_7330,N_3229,N_4181);
xnor U7331 (N_7331,N_2959,N_3324);
xor U7332 (N_7332,N_1687,N_436);
or U7333 (N_7333,N_3555,N_4670);
and U7334 (N_7334,N_33,N_1958);
or U7335 (N_7335,N_4327,N_2340);
or U7336 (N_7336,N_1050,N_1386);
nand U7337 (N_7337,N_2953,N_849);
or U7338 (N_7338,N_3002,N_2615);
nor U7339 (N_7339,N_3300,N_1207);
nand U7340 (N_7340,N_4032,N_3733);
nor U7341 (N_7341,N_2469,N_120);
or U7342 (N_7342,N_3276,N_1385);
and U7343 (N_7343,N_4077,N_4091);
or U7344 (N_7344,N_2695,N_4611);
and U7345 (N_7345,N_1489,N_4998);
and U7346 (N_7346,N_3885,N_1926);
and U7347 (N_7347,N_3998,N_4007);
nand U7348 (N_7348,N_1203,N_1647);
and U7349 (N_7349,N_2633,N_4165);
or U7350 (N_7350,N_1126,N_1822);
nand U7351 (N_7351,N_252,N_1677);
xor U7352 (N_7352,N_2700,N_3986);
and U7353 (N_7353,N_3742,N_3188);
or U7354 (N_7354,N_885,N_3952);
and U7355 (N_7355,N_1931,N_3477);
nand U7356 (N_7356,N_4252,N_3186);
and U7357 (N_7357,N_3316,N_4491);
nor U7358 (N_7358,N_4129,N_2709);
xor U7359 (N_7359,N_561,N_3440);
xnor U7360 (N_7360,N_1533,N_117);
and U7361 (N_7361,N_2618,N_2044);
or U7362 (N_7362,N_801,N_3360);
or U7363 (N_7363,N_3715,N_4363);
or U7364 (N_7364,N_3136,N_3114);
and U7365 (N_7365,N_4359,N_522);
xnor U7366 (N_7366,N_4015,N_3634);
and U7367 (N_7367,N_3343,N_3154);
nor U7368 (N_7368,N_1027,N_4508);
or U7369 (N_7369,N_3903,N_2535);
or U7370 (N_7370,N_519,N_4604);
nand U7371 (N_7371,N_2651,N_2626);
nand U7372 (N_7372,N_4632,N_1492);
nor U7373 (N_7373,N_1095,N_2174);
nand U7374 (N_7374,N_1453,N_1913);
or U7375 (N_7375,N_4006,N_4817);
or U7376 (N_7376,N_1837,N_4256);
nor U7377 (N_7377,N_2599,N_923);
and U7378 (N_7378,N_3481,N_2531);
xor U7379 (N_7379,N_192,N_2037);
xor U7380 (N_7380,N_3294,N_536);
and U7381 (N_7381,N_4114,N_2063);
nand U7382 (N_7382,N_2021,N_2622);
nand U7383 (N_7383,N_1720,N_3510);
xnor U7384 (N_7384,N_1189,N_174);
or U7385 (N_7385,N_2557,N_4183);
xnor U7386 (N_7386,N_3819,N_4243);
and U7387 (N_7387,N_1199,N_3849);
nor U7388 (N_7388,N_1161,N_469);
and U7389 (N_7389,N_2118,N_3423);
nand U7390 (N_7390,N_269,N_1122);
nor U7391 (N_7391,N_3467,N_3459);
nor U7392 (N_7392,N_2476,N_2485);
and U7393 (N_7393,N_1709,N_4906);
nand U7394 (N_7394,N_1783,N_2093);
and U7395 (N_7395,N_276,N_1396);
and U7396 (N_7396,N_4831,N_4325);
nor U7397 (N_7397,N_4648,N_4490);
nand U7398 (N_7398,N_149,N_4118);
and U7399 (N_7399,N_4257,N_3338);
nor U7400 (N_7400,N_3432,N_31);
and U7401 (N_7401,N_4649,N_2178);
and U7402 (N_7402,N_2386,N_244);
or U7403 (N_7403,N_4763,N_1226);
and U7404 (N_7404,N_2097,N_1230);
nor U7405 (N_7405,N_2154,N_2690);
xor U7406 (N_7406,N_2674,N_4033);
xor U7407 (N_7407,N_3729,N_4874);
xor U7408 (N_7408,N_2061,N_4463);
nand U7409 (N_7409,N_3509,N_271);
nor U7410 (N_7410,N_2059,N_4492);
xnor U7411 (N_7411,N_1551,N_4465);
xor U7412 (N_7412,N_4246,N_4992);
nand U7413 (N_7413,N_1474,N_1642);
nand U7414 (N_7414,N_530,N_3976);
xnor U7415 (N_7415,N_4787,N_607);
and U7416 (N_7416,N_1023,N_1424);
nor U7417 (N_7417,N_3134,N_4888);
nand U7418 (N_7418,N_1974,N_2158);
xor U7419 (N_7419,N_4096,N_90);
nor U7420 (N_7420,N_2350,N_3349);
nand U7421 (N_7421,N_4346,N_621);
nand U7422 (N_7422,N_3823,N_2421);
or U7423 (N_7423,N_4222,N_3553);
or U7424 (N_7424,N_2431,N_1760);
or U7425 (N_7425,N_4136,N_3080);
nand U7426 (N_7426,N_4260,N_577);
or U7427 (N_7427,N_2780,N_3141);
xor U7428 (N_7428,N_2876,N_4869);
nor U7429 (N_7429,N_1902,N_3827);
nand U7430 (N_7430,N_4142,N_73);
or U7431 (N_7431,N_2264,N_2275);
and U7432 (N_7432,N_520,N_995);
nand U7433 (N_7433,N_3950,N_1366);
xor U7434 (N_7434,N_3933,N_4382);
nor U7435 (N_7435,N_406,N_2067);
xnor U7436 (N_7436,N_2023,N_1093);
nor U7437 (N_7437,N_1814,N_386);
xor U7438 (N_7438,N_2592,N_2565);
xor U7439 (N_7439,N_2201,N_4562);
nand U7440 (N_7440,N_666,N_2612);
nand U7441 (N_7441,N_1576,N_1502);
and U7442 (N_7442,N_3895,N_1364);
or U7443 (N_7443,N_1883,N_313);
nand U7444 (N_7444,N_4094,N_2354);
nor U7445 (N_7445,N_2237,N_3274);
xor U7446 (N_7446,N_3203,N_3288);
nand U7447 (N_7447,N_4173,N_1142);
or U7448 (N_7448,N_159,N_1635);
or U7449 (N_7449,N_1144,N_4416);
xor U7450 (N_7450,N_656,N_4816);
or U7451 (N_7451,N_3726,N_1852);
xnor U7452 (N_7452,N_971,N_2146);
xnor U7453 (N_7453,N_2454,N_3566);
xor U7454 (N_7454,N_3479,N_3678);
or U7455 (N_7455,N_1119,N_4149);
and U7456 (N_7456,N_1731,N_726);
nor U7457 (N_7457,N_20,N_105);
nand U7458 (N_7458,N_3037,N_3066);
and U7459 (N_7459,N_910,N_1338);
or U7460 (N_7460,N_1728,N_2049);
and U7461 (N_7461,N_1999,N_1745);
xnor U7462 (N_7462,N_1405,N_4412);
and U7463 (N_7463,N_4876,N_4239);
or U7464 (N_7464,N_2809,N_4838);
nand U7465 (N_7465,N_714,N_1121);
xor U7466 (N_7466,N_1996,N_3975);
nand U7467 (N_7467,N_260,N_4176);
and U7468 (N_7468,N_1340,N_3382);
or U7469 (N_7469,N_1614,N_4484);
nor U7470 (N_7470,N_2294,N_3961);
nor U7471 (N_7471,N_650,N_3548);
nand U7472 (N_7472,N_4439,N_1615);
nor U7473 (N_7473,N_792,N_30);
xor U7474 (N_7474,N_1932,N_737);
nand U7475 (N_7475,N_109,N_1310);
xnor U7476 (N_7476,N_2786,N_1232);
xnor U7477 (N_7477,N_3521,N_2127);
or U7478 (N_7478,N_4130,N_2965);
or U7479 (N_7479,N_2646,N_2447);
or U7480 (N_7480,N_2305,N_970);
xor U7481 (N_7481,N_1252,N_2268);
xor U7482 (N_7482,N_2056,N_4407);
and U7483 (N_7483,N_286,N_4595);
nand U7484 (N_7484,N_1295,N_3323);
nand U7485 (N_7485,N_4076,N_2302);
and U7486 (N_7486,N_3820,N_1435);
or U7487 (N_7487,N_2554,N_3621);
nor U7488 (N_7488,N_1770,N_4459);
or U7489 (N_7489,N_2428,N_4807);
nor U7490 (N_7490,N_829,N_2921);
xnor U7491 (N_7491,N_2233,N_139);
or U7492 (N_7492,N_3579,N_144);
nor U7493 (N_7493,N_2303,N_2912);
and U7494 (N_7494,N_2406,N_2767);
xor U7495 (N_7495,N_769,N_2402);
xor U7496 (N_7496,N_1570,N_2957);
or U7497 (N_7497,N_2171,N_2902);
nor U7498 (N_7498,N_4793,N_1895);
nand U7499 (N_7499,N_2829,N_2508);
nand U7500 (N_7500,N_4045,N_3683);
or U7501 (N_7501,N_4360,N_3411);
xor U7502 (N_7502,N_803,N_2548);
or U7503 (N_7503,N_1188,N_3656);
and U7504 (N_7504,N_3871,N_556);
and U7505 (N_7505,N_1999,N_3531);
or U7506 (N_7506,N_797,N_4132);
nand U7507 (N_7507,N_1219,N_3082);
xor U7508 (N_7508,N_167,N_2768);
nand U7509 (N_7509,N_2762,N_4416);
nand U7510 (N_7510,N_2163,N_4042);
xor U7511 (N_7511,N_963,N_1108);
or U7512 (N_7512,N_4652,N_3888);
and U7513 (N_7513,N_3767,N_2123);
or U7514 (N_7514,N_2655,N_351);
nand U7515 (N_7515,N_3100,N_4255);
and U7516 (N_7516,N_3972,N_3408);
nand U7517 (N_7517,N_2559,N_1973);
nor U7518 (N_7518,N_4699,N_2950);
nor U7519 (N_7519,N_3092,N_232);
xor U7520 (N_7520,N_2440,N_3564);
nand U7521 (N_7521,N_1162,N_3473);
xor U7522 (N_7522,N_1780,N_2284);
xnor U7523 (N_7523,N_1376,N_4506);
or U7524 (N_7524,N_1890,N_692);
and U7525 (N_7525,N_618,N_2997);
xor U7526 (N_7526,N_2201,N_195);
and U7527 (N_7527,N_1852,N_4439);
and U7528 (N_7528,N_309,N_1506);
xor U7529 (N_7529,N_1814,N_2934);
xnor U7530 (N_7530,N_205,N_906);
or U7531 (N_7531,N_1721,N_214);
xnor U7532 (N_7532,N_1479,N_178);
nand U7533 (N_7533,N_2680,N_3944);
nand U7534 (N_7534,N_1662,N_2010);
and U7535 (N_7535,N_4574,N_1095);
and U7536 (N_7536,N_2749,N_3978);
nor U7537 (N_7537,N_4370,N_476);
or U7538 (N_7538,N_2404,N_961);
xnor U7539 (N_7539,N_1677,N_1418);
or U7540 (N_7540,N_3294,N_3891);
nor U7541 (N_7541,N_4591,N_837);
xnor U7542 (N_7542,N_1046,N_1830);
or U7543 (N_7543,N_909,N_4398);
nand U7544 (N_7544,N_2803,N_603);
xor U7545 (N_7545,N_214,N_1984);
or U7546 (N_7546,N_126,N_608);
xnor U7547 (N_7547,N_720,N_4506);
nand U7548 (N_7548,N_2111,N_4588);
nor U7549 (N_7549,N_1173,N_4644);
xnor U7550 (N_7550,N_4296,N_4679);
nor U7551 (N_7551,N_1861,N_3699);
or U7552 (N_7552,N_1460,N_173);
and U7553 (N_7553,N_476,N_665);
nor U7554 (N_7554,N_3444,N_3884);
xnor U7555 (N_7555,N_2672,N_1259);
nor U7556 (N_7556,N_590,N_1590);
xnor U7557 (N_7557,N_2756,N_1238);
or U7558 (N_7558,N_2868,N_1383);
and U7559 (N_7559,N_4799,N_3487);
and U7560 (N_7560,N_4152,N_140);
nand U7561 (N_7561,N_3808,N_658);
and U7562 (N_7562,N_3953,N_3132);
nand U7563 (N_7563,N_4030,N_2731);
or U7564 (N_7564,N_4,N_4143);
xor U7565 (N_7565,N_3957,N_1568);
nand U7566 (N_7566,N_3903,N_4836);
or U7567 (N_7567,N_286,N_924);
xor U7568 (N_7568,N_4256,N_3985);
or U7569 (N_7569,N_2134,N_1408);
or U7570 (N_7570,N_1988,N_3780);
or U7571 (N_7571,N_51,N_1777);
nor U7572 (N_7572,N_4200,N_2068);
xnor U7573 (N_7573,N_4895,N_3047);
xor U7574 (N_7574,N_2673,N_2730);
nand U7575 (N_7575,N_2147,N_2007);
nand U7576 (N_7576,N_245,N_2101);
nor U7577 (N_7577,N_717,N_1966);
nor U7578 (N_7578,N_3603,N_2832);
xnor U7579 (N_7579,N_1206,N_1860);
xnor U7580 (N_7580,N_2289,N_2363);
xnor U7581 (N_7581,N_3032,N_948);
and U7582 (N_7582,N_4596,N_1792);
xnor U7583 (N_7583,N_1784,N_1917);
nand U7584 (N_7584,N_1485,N_4386);
and U7585 (N_7585,N_4423,N_4957);
or U7586 (N_7586,N_560,N_938);
nor U7587 (N_7587,N_1049,N_1255);
xnor U7588 (N_7588,N_3277,N_3808);
xnor U7589 (N_7589,N_4853,N_104);
and U7590 (N_7590,N_2915,N_1378);
nand U7591 (N_7591,N_4537,N_2145);
and U7592 (N_7592,N_3158,N_2585);
and U7593 (N_7593,N_4738,N_3274);
or U7594 (N_7594,N_4750,N_608);
nor U7595 (N_7595,N_956,N_4370);
nand U7596 (N_7596,N_3308,N_3759);
or U7597 (N_7597,N_3323,N_3910);
nor U7598 (N_7598,N_1779,N_2490);
xnor U7599 (N_7599,N_3346,N_4758);
xnor U7600 (N_7600,N_4618,N_1531);
or U7601 (N_7601,N_1823,N_1434);
xor U7602 (N_7602,N_3422,N_773);
nand U7603 (N_7603,N_1305,N_557);
nor U7604 (N_7604,N_1771,N_2276);
and U7605 (N_7605,N_1799,N_3554);
and U7606 (N_7606,N_353,N_1940);
nand U7607 (N_7607,N_3463,N_4212);
xor U7608 (N_7608,N_4654,N_720);
xnor U7609 (N_7609,N_2305,N_1881);
xor U7610 (N_7610,N_4875,N_1835);
nor U7611 (N_7611,N_1746,N_4292);
nor U7612 (N_7612,N_400,N_5);
or U7613 (N_7613,N_2923,N_3109);
and U7614 (N_7614,N_554,N_4136);
xor U7615 (N_7615,N_2798,N_4216);
or U7616 (N_7616,N_4320,N_1131);
or U7617 (N_7617,N_2976,N_3636);
and U7618 (N_7618,N_441,N_1294);
xor U7619 (N_7619,N_2938,N_2696);
xor U7620 (N_7620,N_1676,N_3919);
nor U7621 (N_7621,N_1156,N_3284);
nor U7622 (N_7622,N_297,N_3110);
or U7623 (N_7623,N_763,N_2412);
nand U7624 (N_7624,N_3612,N_2385);
and U7625 (N_7625,N_1287,N_2992);
nand U7626 (N_7626,N_4388,N_1860);
nor U7627 (N_7627,N_3318,N_2551);
nand U7628 (N_7628,N_1332,N_3862);
or U7629 (N_7629,N_4092,N_775);
nor U7630 (N_7630,N_1346,N_4224);
nand U7631 (N_7631,N_2983,N_4847);
nor U7632 (N_7632,N_2567,N_1807);
and U7633 (N_7633,N_1366,N_4876);
and U7634 (N_7634,N_4244,N_3917);
nor U7635 (N_7635,N_740,N_4767);
nand U7636 (N_7636,N_2093,N_2090);
nor U7637 (N_7637,N_1182,N_2737);
or U7638 (N_7638,N_3055,N_3616);
nand U7639 (N_7639,N_3937,N_51);
xor U7640 (N_7640,N_130,N_27);
or U7641 (N_7641,N_2063,N_1872);
nor U7642 (N_7642,N_1562,N_3865);
and U7643 (N_7643,N_3099,N_1066);
xor U7644 (N_7644,N_2110,N_1928);
xor U7645 (N_7645,N_1453,N_2843);
nand U7646 (N_7646,N_2332,N_1718);
or U7647 (N_7647,N_1707,N_2106);
xor U7648 (N_7648,N_4234,N_642);
or U7649 (N_7649,N_1046,N_4961);
and U7650 (N_7650,N_3135,N_128);
xor U7651 (N_7651,N_517,N_543);
nor U7652 (N_7652,N_3306,N_3190);
nor U7653 (N_7653,N_1280,N_707);
or U7654 (N_7654,N_1839,N_3762);
and U7655 (N_7655,N_4289,N_1012);
and U7656 (N_7656,N_3521,N_1237);
or U7657 (N_7657,N_1218,N_2069);
nand U7658 (N_7658,N_1323,N_3978);
nor U7659 (N_7659,N_4242,N_4362);
nand U7660 (N_7660,N_463,N_3908);
nor U7661 (N_7661,N_2463,N_2146);
nor U7662 (N_7662,N_3103,N_4269);
xor U7663 (N_7663,N_2710,N_4405);
nand U7664 (N_7664,N_3370,N_3948);
or U7665 (N_7665,N_3492,N_3634);
nand U7666 (N_7666,N_287,N_1934);
and U7667 (N_7667,N_2005,N_238);
xor U7668 (N_7668,N_2101,N_687);
or U7669 (N_7669,N_1692,N_4869);
nor U7670 (N_7670,N_1114,N_4077);
or U7671 (N_7671,N_1538,N_1466);
or U7672 (N_7672,N_1707,N_3518);
nand U7673 (N_7673,N_1071,N_3255);
and U7674 (N_7674,N_2196,N_2748);
nand U7675 (N_7675,N_471,N_3514);
nor U7676 (N_7676,N_332,N_1564);
nand U7677 (N_7677,N_3098,N_4133);
or U7678 (N_7678,N_4321,N_2322);
nand U7679 (N_7679,N_3004,N_857);
xnor U7680 (N_7680,N_658,N_2257);
or U7681 (N_7681,N_3030,N_123);
nor U7682 (N_7682,N_3462,N_3792);
and U7683 (N_7683,N_3030,N_4114);
or U7684 (N_7684,N_1010,N_674);
xor U7685 (N_7685,N_4572,N_2949);
xnor U7686 (N_7686,N_3333,N_4924);
and U7687 (N_7687,N_3785,N_4268);
or U7688 (N_7688,N_4608,N_1086);
or U7689 (N_7689,N_3887,N_4942);
or U7690 (N_7690,N_2476,N_5);
or U7691 (N_7691,N_1236,N_2667);
nor U7692 (N_7692,N_2568,N_1493);
nor U7693 (N_7693,N_3154,N_3553);
nand U7694 (N_7694,N_2542,N_4792);
xnor U7695 (N_7695,N_1850,N_4841);
and U7696 (N_7696,N_4123,N_1635);
and U7697 (N_7697,N_1033,N_1605);
nand U7698 (N_7698,N_4317,N_86);
nor U7699 (N_7699,N_4133,N_2562);
or U7700 (N_7700,N_3875,N_4613);
nor U7701 (N_7701,N_342,N_1136);
nor U7702 (N_7702,N_157,N_3088);
nand U7703 (N_7703,N_1292,N_494);
nor U7704 (N_7704,N_3465,N_1048);
or U7705 (N_7705,N_1393,N_4244);
nand U7706 (N_7706,N_4294,N_468);
nand U7707 (N_7707,N_3883,N_573);
xnor U7708 (N_7708,N_4406,N_561);
or U7709 (N_7709,N_3033,N_33);
xnor U7710 (N_7710,N_1118,N_2189);
nand U7711 (N_7711,N_3255,N_2812);
and U7712 (N_7712,N_4248,N_4975);
and U7713 (N_7713,N_4449,N_3596);
nor U7714 (N_7714,N_99,N_4964);
nand U7715 (N_7715,N_1588,N_3696);
and U7716 (N_7716,N_2579,N_2560);
nor U7717 (N_7717,N_2044,N_1692);
or U7718 (N_7718,N_3092,N_1530);
or U7719 (N_7719,N_1830,N_1592);
or U7720 (N_7720,N_284,N_437);
nor U7721 (N_7721,N_4181,N_1955);
or U7722 (N_7722,N_2884,N_772);
xor U7723 (N_7723,N_1994,N_3459);
and U7724 (N_7724,N_4226,N_2572);
nand U7725 (N_7725,N_199,N_372);
nor U7726 (N_7726,N_95,N_4180);
nand U7727 (N_7727,N_4762,N_4576);
and U7728 (N_7728,N_1593,N_2549);
or U7729 (N_7729,N_1081,N_2033);
and U7730 (N_7730,N_1083,N_262);
nand U7731 (N_7731,N_4687,N_776);
nor U7732 (N_7732,N_4228,N_908);
or U7733 (N_7733,N_1364,N_335);
and U7734 (N_7734,N_1025,N_1885);
nand U7735 (N_7735,N_4261,N_1654);
nand U7736 (N_7736,N_2782,N_69);
nor U7737 (N_7737,N_4814,N_3007);
nand U7738 (N_7738,N_4803,N_540);
xnor U7739 (N_7739,N_1970,N_4786);
and U7740 (N_7740,N_1459,N_353);
nand U7741 (N_7741,N_488,N_4924);
and U7742 (N_7742,N_4390,N_4099);
nor U7743 (N_7743,N_3549,N_2376);
nor U7744 (N_7744,N_798,N_2921);
xnor U7745 (N_7745,N_4365,N_1157);
xnor U7746 (N_7746,N_1770,N_773);
and U7747 (N_7747,N_3776,N_4255);
xnor U7748 (N_7748,N_4701,N_4206);
nor U7749 (N_7749,N_2767,N_1235);
xor U7750 (N_7750,N_4034,N_2568);
nand U7751 (N_7751,N_1396,N_4893);
and U7752 (N_7752,N_368,N_814);
or U7753 (N_7753,N_3664,N_1708);
nor U7754 (N_7754,N_4146,N_3877);
or U7755 (N_7755,N_1408,N_495);
and U7756 (N_7756,N_2691,N_3567);
or U7757 (N_7757,N_1354,N_4140);
or U7758 (N_7758,N_3981,N_2372);
xor U7759 (N_7759,N_2956,N_2714);
xnor U7760 (N_7760,N_3128,N_4750);
nand U7761 (N_7761,N_764,N_2069);
and U7762 (N_7762,N_4968,N_1668);
nand U7763 (N_7763,N_2045,N_2794);
and U7764 (N_7764,N_4932,N_1165);
and U7765 (N_7765,N_3519,N_3107);
nand U7766 (N_7766,N_3269,N_1614);
or U7767 (N_7767,N_1078,N_3122);
nor U7768 (N_7768,N_3558,N_10);
xnor U7769 (N_7769,N_4560,N_1120);
xor U7770 (N_7770,N_4191,N_91);
or U7771 (N_7771,N_2826,N_130);
xnor U7772 (N_7772,N_3578,N_425);
and U7773 (N_7773,N_3711,N_4442);
nand U7774 (N_7774,N_3740,N_2812);
and U7775 (N_7775,N_111,N_4522);
nand U7776 (N_7776,N_975,N_4979);
or U7777 (N_7777,N_151,N_4891);
or U7778 (N_7778,N_3028,N_1217);
nor U7779 (N_7779,N_2031,N_1999);
nor U7780 (N_7780,N_2390,N_3359);
nand U7781 (N_7781,N_540,N_1719);
xor U7782 (N_7782,N_20,N_775);
nor U7783 (N_7783,N_63,N_3373);
and U7784 (N_7784,N_4105,N_1894);
nand U7785 (N_7785,N_3668,N_559);
and U7786 (N_7786,N_3947,N_4224);
nand U7787 (N_7787,N_4512,N_2055);
nor U7788 (N_7788,N_1891,N_3932);
xor U7789 (N_7789,N_2997,N_2259);
and U7790 (N_7790,N_514,N_3284);
and U7791 (N_7791,N_4561,N_1022);
nand U7792 (N_7792,N_1576,N_4829);
nor U7793 (N_7793,N_3801,N_4738);
nand U7794 (N_7794,N_1359,N_4866);
nand U7795 (N_7795,N_3116,N_1318);
and U7796 (N_7796,N_1677,N_2090);
or U7797 (N_7797,N_3419,N_3745);
xor U7798 (N_7798,N_4636,N_4006);
nor U7799 (N_7799,N_4201,N_980);
nand U7800 (N_7800,N_4137,N_2866);
nor U7801 (N_7801,N_2985,N_1342);
and U7802 (N_7802,N_3889,N_2813);
or U7803 (N_7803,N_140,N_2106);
nor U7804 (N_7804,N_931,N_4415);
or U7805 (N_7805,N_4464,N_3491);
xnor U7806 (N_7806,N_3759,N_301);
and U7807 (N_7807,N_668,N_4402);
xor U7808 (N_7808,N_3889,N_2539);
or U7809 (N_7809,N_3312,N_3798);
nor U7810 (N_7810,N_2758,N_3255);
nor U7811 (N_7811,N_640,N_2393);
xnor U7812 (N_7812,N_3882,N_3970);
xor U7813 (N_7813,N_4002,N_2187);
xor U7814 (N_7814,N_3634,N_1348);
nor U7815 (N_7815,N_3350,N_3695);
nor U7816 (N_7816,N_1615,N_361);
or U7817 (N_7817,N_744,N_3478);
nand U7818 (N_7818,N_4872,N_106);
nor U7819 (N_7819,N_4091,N_3539);
xor U7820 (N_7820,N_127,N_253);
nor U7821 (N_7821,N_3959,N_4714);
and U7822 (N_7822,N_229,N_223);
nand U7823 (N_7823,N_2575,N_3636);
or U7824 (N_7824,N_979,N_1742);
or U7825 (N_7825,N_1894,N_685);
or U7826 (N_7826,N_4305,N_3926);
and U7827 (N_7827,N_2922,N_222);
nand U7828 (N_7828,N_1941,N_2861);
xor U7829 (N_7829,N_369,N_4757);
or U7830 (N_7830,N_353,N_1387);
xor U7831 (N_7831,N_1240,N_2223);
and U7832 (N_7832,N_726,N_1653);
nor U7833 (N_7833,N_2177,N_4634);
nand U7834 (N_7834,N_3951,N_12);
and U7835 (N_7835,N_1805,N_1680);
nand U7836 (N_7836,N_153,N_4582);
and U7837 (N_7837,N_3950,N_4687);
nand U7838 (N_7838,N_1510,N_4719);
and U7839 (N_7839,N_4894,N_3683);
or U7840 (N_7840,N_3669,N_4764);
nor U7841 (N_7841,N_4657,N_498);
or U7842 (N_7842,N_1239,N_3952);
and U7843 (N_7843,N_3020,N_3778);
nor U7844 (N_7844,N_2980,N_1225);
nor U7845 (N_7845,N_1214,N_2791);
nor U7846 (N_7846,N_2403,N_205);
and U7847 (N_7847,N_93,N_1788);
and U7848 (N_7848,N_4235,N_2531);
or U7849 (N_7849,N_1164,N_3368);
and U7850 (N_7850,N_3591,N_3300);
xnor U7851 (N_7851,N_506,N_1789);
and U7852 (N_7852,N_4698,N_889);
nor U7853 (N_7853,N_3598,N_4299);
nor U7854 (N_7854,N_4087,N_3738);
and U7855 (N_7855,N_2385,N_1960);
nand U7856 (N_7856,N_3393,N_3122);
and U7857 (N_7857,N_3200,N_4069);
nor U7858 (N_7858,N_1440,N_3860);
or U7859 (N_7859,N_4243,N_109);
and U7860 (N_7860,N_4490,N_860);
xnor U7861 (N_7861,N_1367,N_518);
nand U7862 (N_7862,N_4379,N_1730);
or U7863 (N_7863,N_4859,N_2576);
or U7864 (N_7864,N_562,N_1231);
nor U7865 (N_7865,N_319,N_4113);
nand U7866 (N_7866,N_881,N_2980);
nand U7867 (N_7867,N_4307,N_1161);
and U7868 (N_7868,N_1966,N_3393);
nor U7869 (N_7869,N_148,N_732);
or U7870 (N_7870,N_4299,N_1179);
nor U7871 (N_7871,N_4805,N_2591);
or U7872 (N_7872,N_3510,N_4630);
and U7873 (N_7873,N_970,N_2120);
and U7874 (N_7874,N_2018,N_2227);
and U7875 (N_7875,N_1452,N_4060);
xnor U7876 (N_7876,N_1516,N_2438);
and U7877 (N_7877,N_156,N_1971);
nand U7878 (N_7878,N_1993,N_638);
and U7879 (N_7879,N_3378,N_2521);
xnor U7880 (N_7880,N_621,N_3436);
or U7881 (N_7881,N_3382,N_4567);
xnor U7882 (N_7882,N_1234,N_173);
nor U7883 (N_7883,N_4764,N_201);
or U7884 (N_7884,N_2595,N_3638);
or U7885 (N_7885,N_1924,N_4136);
nor U7886 (N_7886,N_3911,N_2380);
xnor U7887 (N_7887,N_2874,N_1895);
or U7888 (N_7888,N_3396,N_2915);
and U7889 (N_7889,N_3622,N_1947);
or U7890 (N_7890,N_1146,N_3693);
xnor U7891 (N_7891,N_840,N_2713);
nor U7892 (N_7892,N_2855,N_3742);
nand U7893 (N_7893,N_672,N_582);
nor U7894 (N_7894,N_4751,N_2761);
and U7895 (N_7895,N_3654,N_4442);
or U7896 (N_7896,N_4473,N_2890);
xnor U7897 (N_7897,N_3938,N_3102);
or U7898 (N_7898,N_4124,N_2808);
and U7899 (N_7899,N_55,N_1555);
or U7900 (N_7900,N_646,N_2130);
and U7901 (N_7901,N_4414,N_4711);
nand U7902 (N_7902,N_1589,N_2132);
nor U7903 (N_7903,N_4538,N_729);
and U7904 (N_7904,N_4791,N_1323);
nand U7905 (N_7905,N_1766,N_2763);
xor U7906 (N_7906,N_1365,N_1202);
xnor U7907 (N_7907,N_4663,N_563);
and U7908 (N_7908,N_4682,N_4533);
and U7909 (N_7909,N_1206,N_3838);
nor U7910 (N_7910,N_1292,N_3747);
nand U7911 (N_7911,N_4242,N_575);
xor U7912 (N_7912,N_1449,N_1729);
and U7913 (N_7913,N_845,N_2098);
nand U7914 (N_7914,N_3860,N_1527);
and U7915 (N_7915,N_1429,N_3218);
nor U7916 (N_7916,N_1920,N_2313);
and U7917 (N_7917,N_2866,N_2168);
xor U7918 (N_7918,N_1894,N_3060);
nor U7919 (N_7919,N_4065,N_1801);
or U7920 (N_7920,N_3869,N_1491);
or U7921 (N_7921,N_1470,N_1840);
and U7922 (N_7922,N_3595,N_3973);
xnor U7923 (N_7923,N_1521,N_4872);
or U7924 (N_7924,N_2099,N_372);
and U7925 (N_7925,N_3619,N_4887);
and U7926 (N_7926,N_2526,N_493);
and U7927 (N_7927,N_2438,N_1139);
nor U7928 (N_7928,N_222,N_898);
nor U7929 (N_7929,N_2294,N_1425);
nand U7930 (N_7930,N_925,N_4520);
and U7931 (N_7931,N_368,N_903);
or U7932 (N_7932,N_3756,N_3183);
and U7933 (N_7933,N_2940,N_1244);
and U7934 (N_7934,N_3334,N_2914);
nor U7935 (N_7935,N_1203,N_98);
and U7936 (N_7936,N_4854,N_3143);
nor U7937 (N_7937,N_1726,N_1913);
xor U7938 (N_7938,N_3636,N_3825);
or U7939 (N_7939,N_38,N_2665);
nand U7940 (N_7940,N_3978,N_3371);
and U7941 (N_7941,N_4975,N_2292);
and U7942 (N_7942,N_3870,N_1447);
and U7943 (N_7943,N_346,N_2474);
nor U7944 (N_7944,N_2236,N_3177);
and U7945 (N_7945,N_2837,N_3161);
xor U7946 (N_7946,N_3925,N_3016);
and U7947 (N_7947,N_4068,N_4122);
xor U7948 (N_7948,N_2938,N_2802);
or U7949 (N_7949,N_1159,N_1281);
or U7950 (N_7950,N_3406,N_2621);
or U7951 (N_7951,N_2556,N_3496);
nor U7952 (N_7952,N_263,N_2299);
xnor U7953 (N_7953,N_1787,N_76);
nand U7954 (N_7954,N_3529,N_2399);
nor U7955 (N_7955,N_4632,N_4837);
nor U7956 (N_7956,N_1344,N_1745);
and U7957 (N_7957,N_1952,N_1884);
and U7958 (N_7958,N_3758,N_4672);
and U7959 (N_7959,N_4935,N_3750);
nand U7960 (N_7960,N_2660,N_4386);
nor U7961 (N_7961,N_1500,N_4691);
xor U7962 (N_7962,N_2230,N_4126);
nor U7963 (N_7963,N_4747,N_4494);
xor U7964 (N_7964,N_2233,N_2577);
or U7965 (N_7965,N_1377,N_4220);
nor U7966 (N_7966,N_68,N_4232);
xor U7967 (N_7967,N_3644,N_3343);
nor U7968 (N_7968,N_1602,N_3261);
and U7969 (N_7969,N_240,N_759);
or U7970 (N_7970,N_3939,N_1424);
xnor U7971 (N_7971,N_1143,N_3399);
nand U7972 (N_7972,N_4422,N_2437);
and U7973 (N_7973,N_2969,N_3910);
nand U7974 (N_7974,N_3242,N_4618);
and U7975 (N_7975,N_2766,N_2711);
or U7976 (N_7976,N_3688,N_3485);
xnor U7977 (N_7977,N_469,N_1858);
nor U7978 (N_7978,N_719,N_1229);
and U7979 (N_7979,N_3335,N_3289);
or U7980 (N_7980,N_3736,N_1969);
nor U7981 (N_7981,N_3883,N_3220);
xor U7982 (N_7982,N_2500,N_2739);
nand U7983 (N_7983,N_4332,N_3741);
nand U7984 (N_7984,N_677,N_3743);
nand U7985 (N_7985,N_2058,N_1695);
nand U7986 (N_7986,N_3496,N_383);
xnor U7987 (N_7987,N_2916,N_4638);
nor U7988 (N_7988,N_3889,N_4980);
xor U7989 (N_7989,N_4726,N_1605);
or U7990 (N_7990,N_288,N_1743);
and U7991 (N_7991,N_1926,N_894);
or U7992 (N_7992,N_1534,N_4650);
or U7993 (N_7993,N_2464,N_4997);
nand U7994 (N_7994,N_117,N_1745);
xor U7995 (N_7995,N_523,N_3650);
and U7996 (N_7996,N_1220,N_2689);
or U7997 (N_7997,N_2291,N_4360);
nand U7998 (N_7998,N_524,N_2515);
or U7999 (N_7999,N_4412,N_3028);
or U8000 (N_8000,N_2384,N_1033);
xor U8001 (N_8001,N_2196,N_4768);
nor U8002 (N_8002,N_24,N_546);
xnor U8003 (N_8003,N_865,N_248);
and U8004 (N_8004,N_3637,N_4850);
nor U8005 (N_8005,N_2040,N_3728);
or U8006 (N_8006,N_2778,N_456);
and U8007 (N_8007,N_1537,N_246);
or U8008 (N_8008,N_951,N_212);
or U8009 (N_8009,N_3727,N_1990);
nand U8010 (N_8010,N_1388,N_835);
xor U8011 (N_8011,N_3902,N_4005);
nor U8012 (N_8012,N_3448,N_1484);
nor U8013 (N_8013,N_3855,N_1419);
xor U8014 (N_8014,N_3529,N_4548);
and U8015 (N_8015,N_2813,N_3096);
and U8016 (N_8016,N_1911,N_2740);
and U8017 (N_8017,N_1081,N_3033);
and U8018 (N_8018,N_1843,N_3725);
xnor U8019 (N_8019,N_44,N_771);
nand U8020 (N_8020,N_60,N_2497);
or U8021 (N_8021,N_529,N_1520);
nand U8022 (N_8022,N_3873,N_3782);
nand U8023 (N_8023,N_3671,N_2619);
nor U8024 (N_8024,N_1048,N_3323);
nand U8025 (N_8025,N_113,N_4677);
nor U8026 (N_8026,N_4822,N_1797);
nor U8027 (N_8027,N_1583,N_3208);
or U8028 (N_8028,N_2601,N_3368);
or U8029 (N_8029,N_3021,N_4862);
nand U8030 (N_8030,N_2803,N_3040);
nor U8031 (N_8031,N_2638,N_1637);
nor U8032 (N_8032,N_3882,N_1960);
xor U8033 (N_8033,N_3618,N_4937);
nand U8034 (N_8034,N_256,N_2440);
xor U8035 (N_8035,N_1789,N_4080);
or U8036 (N_8036,N_1013,N_2104);
and U8037 (N_8037,N_2381,N_1359);
or U8038 (N_8038,N_3587,N_1156);
xor U8039 (N_8039,N_26,N_549);
nand U8040 (N_8040,N_4098,N_2993);
nor U8041 (N_8041,N_1251,N_1377);
or U8042 (N_8042,N_1650,N_3454);
nor U8043 (N_8043,N_3637,N_307);
or U8044 (N_8044,N_1390,N_293);
nor U8045 (N_8045,N_3782,N_420);
nand U8046 (N_8046,N_2661,N_3947);
and U8047 (N_8047,N_2010,N_4999);
or U8048 (N_8048,N_488,N_1549);
nand U8049 (N_8049,N_654,N_2987);
xor U8050 (N_8050,N_3248,N_3492);
or U8051 (N_8051,N_1779,N_3070);
and U8052 (N_8052,N_4810,N_1553);
nand U8053 (N_8053,N_3999,N_1351);
and U8054 (N_8054,N_4529,N_2131);
xor U8055 (N_8055,N_4937,N_4236);
or U8056 (N_8056,N_2937,N_3494);
or U8057 (N_8057,N_1730,N_1308);
nor U8058 (N_8058,N_3361,N_206);
and U8059 (N_8059,N_2095,N_3497);
nor U8060 (N_8060,N_495,N_2792);
nand U8061 (N_8061,N_18,N_3788);
xnor U8062 (N_8062,N_2012,N_820);
nand U8063 (N_8063,N_4677,N_2279);
or U8064 (N_8064,N_408,N_667);
xor U8065 (N_8065,N_541,N_2424);
xnor U8066 (N_8066,N_4162,N_4173);
and U8067 (N_8067,N_4458,N_3917);
xnor U8068 (N_8068,N_4471,N_445);
nand U8069 (N_8069,N_4417,N_232);
and U8070 (N_8070,N_2487,N_153);
and U8071 (N_8071,N_293,N_1792);
nor U8072 (N_8072,N_3448,N_548);
nor U8073 (N_8073,N_3382,N_4776);
nand U8074 (N_8074,N_4934,N_3417);
nand U8075 (N_8075,N_432,N_1668);
and U8076 (N_8076,N_4495,N_3131);
xnor U8077 (N_8077,N_1332,N_3833);
nor U8078 (N_8078,N_171,N_285);
and U8079 (N_8079,N_3838,N_2062);
and U8080 (N_8080,N_4051,N_4784);
nor U8081 (N_8081,N_1198,N_516);
nor U8082 (N_8082,N_3358,N_3801);
nand U8083 (N_8083,N_4965,N_2092);
or U8084 (N_8084,N_928,N_3772);
nand U8085 (N_8085,N_2609,N_2141);
xor U8086 (N_8086,N_562,N_1099);
nor U8087 (N_8087,N_1251,N_1090);
nand U8088 (N_8088,N_2725,N_117);
xor U8089 (N_8089,N_4194,N_4216);
xnor U8090 (N_8090,N_1032,N_824);
and U8091 (N_8091,N_3543,N_1960);
nor U8092 (N_8092,N_3591,N_4161);
or U8093 (N_8093,N_516,N_48);
and U8094 (N_8094,N_647,N_3116);
nand U8095 (N_8095,N_1281,N_2921);
or U8096 (N_8096,N_2057,N_4340);
nand U8097 (N_8097,N_2655,N_1774);
and U8098 (N_8098,N_605,N_3896);
nand U8099 (N_8099,N_3603,N_4691);
or U8100 (N_8100,N_4089,N_1667);
nor U8101 (N_8101,N_2740,N_934);
nor U8102 (N_8102,N_4149,N_158);
and U8103 (N_8103,N_2854,N_1806);
nand U8104 (N_8104,N_1655,N_4977);
xnor U8105 (N_8105,N_1804,N_3147);
xor U8106 (N_8106,N_941,N_456);
xor U8107 (N_8107,N_2604,N_1614);
or U8108 (N_8108,N_3827,N_1781);
and U8109 (N_8109,N_1161,N_4421);
xnor U8110 (N_8110,N_926,N_3159);
or U8111 (N_8111,N_152,N_952);
or U8112 (N_8112,N_1109,N_1275);
xor U8113 (N_8113,N_51,N_3402);
or U8114 (N_8114,N_4400,N_4757);
and U8115 (N_8115,N_3047,N_2904);
and U8116 (N_8116,N_4075,N_1810);
xor U8117 (N_8117,N_4462,N_4712);
nor U8118 (N_8118,N_2265,N_589);
nor U8119 (N_8119,N_3639,N_3911);
or U8120 (N_8120,N_3481,N_3261);
nor U8121 (N_8121,N_4247,N_1507);
nand U8122 (N_8122,N_3312,N_2729);
xor U8123 (N_8123,N_2988,N_2434);
nor U8124 (N_8124,N_161,N_1661);
and U8125 (N_8125,N_586,N_2451);
nand U8126 (N_8126,N_599,N_3347);
nand U8127 (N_8127,N_4527,N_530);
nor U8128 (N_8128,N_332,N_449);
and U8129 (N_8129,N_4232,N_1308);
xor U8130 (N_8130,N_2537,N_281);
or U8131 (N_8131,N_4130,N_3848);
or U8132 (N_8132,N_2091,N_3614);
xor U8133 (N_8133,N_4369,N_2746);
or U8134 (N_8134,N_3980,N_4487);
xnor U8135 (N_8135,N_939,N_499);
and U8136 (N_8136,N_2477,N_1497);
or U8137 (N_8137,N_673,N_4238);
and U8138 (N_8138,N_3456,N_3143);
or U8139 (N_8139,N_1769,N_2823);
xnor U8140 (N_8140,N_643,N_2395);
nand U8141 (N_8141,N_2636,N_4751);
or U8142 (N_8142,N_3407,N_2745);
or U8143 (N_8143,N_4853,N_1540);
or U8144 (N_8144,N_4278,N_4318);
xnor U8145 (N_8145,N_4987,N_2052);
nand U8146 (N_8146,N_37,N_4246);
nand U8147 (N_8147,N_1017,N_453);
and U8148 (N_8148,N_1746,N_2959);
nor U8149 (N_8149,N_3652,N_4232);
nand U8150 (N_8150,N_224,N_2034);
and U8151 (N_8151,N_1041,N_1470);
and U8152 (N_8152,N_743,N_1907);
nand U8153 (N_8153,N_781,N_2938);
xor U8154 (N_8154,N_3885,N_2838);
nor U8155 (N_8155,N_3254,N_2713);
and U8156 (N_8156,N_3637,N_649);
and U8157 (N_8157,N_4098,N_1063);
nand U8158 (N_8158,N_3820,N_1226);
nand U8159 (N_8159,N_3662,N_2749);
nor U8160 (N_8160,N_4141,N_1812);
and U8161 (N_8161,N_2509,N_3882);
xnor U8162 (N_8162,N_1681,N_865);
or U8163 (N_8163,N_4437,N_4059);
xor U8164 (N_8164,N_2194,N_3161);
or U8165 (N_8165,N_4953,N_726);
and U8166 (N_8166,N_2462,N_1297);
nand U8167 (N_8167,N_4934,N_2235);
nand U8168 (N_8168,N_2783,N_2377);
xnor U8169 (N_8169,N_1749,N_4111);
nor U8170 (N_8170,N_4317,N_2564);
xnor U8171 (N_8171,N_1585,N_3885);
and U8172 (N_8172,N_3587,N_268);
or U8173 (N_8173,N_1423,N_1396);
nor U8174 (N_8174,N_14,N_4519);
xnor U8175 (N_8175,N_3778,N_121);
and U8176 (N_8176,N_2989,N_4574);
nor U8177 (N_8177,N_4737,N_4365);
nand U8178 (N_8178,N_2690,N_2579);
xor U8179 (N_8179,N_3138,N_1437);
nor U8180 (N_8180,N_2710,N_4574);
xnor U8181 (N_8181,N_2539,N_1518);
or U8182 (N_8182,N_46,N_15);
and U8183 (N_8183,N_4914,N_1509);
xor U8184 (N_8184,N_2546,N_2527);
nand U8185 (N_8185,N_1102,N_3729);
nor U8186 (N_8186,N_578,N_1481);
xnor U8187 (N_8187,N_4300,N_4696);
and U8188 (N_8188,N_1400,N_639);
nand U8189 (N_8189,N_4275,N_1839);
nor U8190 (N_8190,N_4731,N_770);
xnor U8191 (N_8191,N_4322,N_722);
xor U8192 (N_8192,N_3959,N_725);
nor U8193 (N_8193,N_4932,N_2156);
nor U8194 (N_8194,N_1429,N_2526);
or U8195 (N_8195,N_444,N_4028);
xnor U8196 (N_8196,N_1873,N_4896);
or U8197 (N_8197,N_1007,N_441);
nor U8198 (N_8198,N_3623,N_4081);
xnor U8199 (N_8199,N_1136,N_2871);
xor U8200 (N_8200,N_3677,N_649);
nor U8201 (N_8201,N_4582,N_3753);
nand U8202 (N_8202,N_3876,N_4731);
or U8203 (N_8203,N_3496,N_4774);
and U8204 (N_8204,N_16,N_3139);
or U8205 (N_8205,N_4201,N_1298);
nor U8206 (N_8206,N_3464,N_738);
nand U8207 (N_8207,N_4057,N_4491);
and U8208 (N_8208,N_4757,N_4810);
nor U8209 (N_8209,N_3755,N_3167);
or U8210 (N_8210,N_3644,N_574);
and U8211 (N_8211,N_4371,N_706);
xnor U8212 (N_8212,N_944,N_3789);
nand U8213 (N_8213,N_2243,N_2628);
xnor U8214 (N_8214,N_1819,N_2751);
and U8215 (N_8215,N_3800,N_936);
nor U8216 (N_8216,N_2778,N_3681);
xnor U8217 (N_8217,N_251,N_1040);
xor U8218 (N_8218,N_2262,N_4321);
nor U8219 (N_8219,N_297,N_1518);
and U8220 (N_8220,N_3964,N_4395);
or U8221 (N_8221,N_2682,N_1298);
xnor U8222 (N_8222,N_1504,N_4267);
xnor U8223 (N_8223,N_879,N_3823);
and U8224 (N_8224,N_890,N_2781);
or U8225 (N_8225,N_4185,N_578);
xor U8226 (N_8226,N_4662,N_2035);
xnor U8227 (N_8227,N_4112,N_4434);
nor U8228 (N_8228,N_4415,N_4837);
or U8229 (N_8229,N_304,N_2044);
xor U8230 (N_8230,N_2437,N_2565);
and U8231 (N_8231,N_4347,N_3784);
nor U8232 (N_8232,N_2492,N_1744);
xnor U8233 (N_8233,N_2208,N_4686);
xnor U8234 (N_8234,N_3935,N_3447);
nor U8235 (N_8235,N_4016,N_1982);
nand U8236 (N_8236,N_2741,N_1783);
nor U8237 (N_8237,N_1987,N_3543);
or U8238 (N_8238,N_686,N_1403);
and U8239 (N_8239,N_4682,N_1573);
and U8240 (N_8240,N_4212,N_756);
or U8241 (N_8241,N_1933,N_2347);
or U8242 (N_8242,N_731,N_4779);
nand U8243 (N_8243,N_4561,N_2814);
or U8244 (N_8244,N_4825,N_492);
or U8245 (N_8245,N_1228,N_4677);
or U8246 (N_8246,N_4790,N_82);
and U8247 (N_8247,N_3994,N_3757);
nor U8248 (N_8248,N_1423,N_4157);
and U8249 (N_8249,N_4720,N_771);
nor U8250 (N_8250,N_3145,N_3718);
nand U8251 (N_8251,N_1622,N_96);
nor U8252 (N_8252,N_2879,N_1497);
nor U8253 (N_8253,N_4154,N_709);
nand U8254 (N_8254,N_1800,N_3510);
or U8255 (N_8255,N_286,N_1075);
nand U8256 (N_8256,N_2678,N_3879);
nor U8257 (N_8257,N_4074,N_2265);
or U8258 (N_8258,N_2278,N_192);
nor U8259 (N_8259,N_4642,N_1696);
and U8260 (N_8260,N_4536,N_2399);
xor U8261 (N_8261,N_961,N_4117);
xor U8262 (N_8262,N_4535,N_284);
nand U8263 (N_8263,N_4255,N_606);
nand U8264 (N_8264,N_258,N_3914);
xnor U8265 (N_8265,N_3723,N_2505);
and U8266 (N_8266,N_1322,N_1204);
nor U8267 (N_8267,N_4992,N_1295);
or U8268 (N_8268,N_4231,N_3709);
and U8269 (N_8269,N_4162,N_1756);
nand U8270 (N_8270,N_1565,N_4493);
xor U8271 (N_8271,N_3299,N_987);
or U8272 (N_8272,N_3382,N_878);
or U8273 (N_8273,N_449,N_2680);
or U8274 (N_8274,N_4142,N_2237);
and U8275 (N_8275,N_3348,N_1794);
nand U8276 (N_8276,N_4754,N_1972);
and U8277 (N_8277,N_3434,N_4183);
nand U8278 (N_8278,N_1630,N_3836);
nand U8279 (N_8279,N_4920,N_943);
xnor U8280 (N_8280,N_4053,N_3839);
and U8281 (N_8281,N_3719,N_414);
and U8282 (N_8282,N_4885,N_1869);
and U8283 (N_8283,N_535,N_67);
or U8284 (N_8284,N_3633,N_853);
or U8285 (N_8285,N_2664,N_4942);
xnor U8286 (N_8286,N_2255,N_2102);
nand U8287 (N_8287,N_234,N_1756);
or U8288 (N_8288,N_3960,N_2078);
nor U8289 (N_8289,N_4435,N_3085);
nand U8290 (N_8290,N_169,N_774);
or U8291 (N_8291,N_216,N_2691);
nand U8292 (N_8292,N_2991,N_3786);
nand U8293 (N_8293,N_4594,N_4354);
xnor U8294 (N_8294,N_3065,N_3787);
xor U8295 (N_8295,N_219,N_2999);
and U8296 (N_8296,N_4404,N_4574);
xnor U8297 (N_8297,N_916,N_3165);
nand U8298 (N_8298,N_4405,N_774);
nand U8299 (N_8299,N_3021,N_4809);
xor U8300 (N_8300,N_2125,N_4228);
nor U8301 (N_8301,N_4926,N_1148);
nand U8302 (N_8302,N_3413,N_3610);
nor U8303 (N_8303,N_4824,N_3440);
and U8304 (N_8304,N_869,N_205);
nor U8305 (N_8305,N_3787,N_137);
nand U8306 (N_8306,N_2173,N_1932);
or U8307 (N_8307,N_1262,N_652);
nand U8308 (N_8308,N_4634,N_2083);
and U8309 (N_8309,N_4853,N_4673);
nor U8310 (N_8310,N_2333,N_1904);
or U8311 (N_8311,N_454,N_600);
nand U8312 (N_8312,N_497,N_1133);
and U8313 (N_8313,N_232,N_4749);
nor U8314 (N_8314,N_1895,N_1131);
and U8315 (N_8315,N_255,N_4432);
xor U8316 (N_8316,N_4604,N_576);
nor U8317 (N_8317,N_1878,N_2884);
or U8318 (N_8318,N_4558,N_1813);
or U8319 (N_8319,N_2091,N_2192);
nand U8320 (N_8320,N_4903,N_4116);
nor U8321 (N_8321,N_2277,N_3442);
nand U8322 (N_8322,N_4296,N_1135);
or U8323 (N_8323,N_1951,N_4563);
nand U8324 (N_8324,N_2294,N_642);
nand U8325 (N_8325,N_1570,N_2622);
and U8326 (N_8326,N_4155,N_3634);
nand U8327 (N_8327,N_494,N_3703);
or U8328 (N_8328,N_109,N_3279);
nand U8329 (N_8329,N_3218,N_2462);
or U8330 (N_8330,N_3118,N_146);
or U8331 (N_8331,N_796,N_1029);
xor U8332 (N_8332,N_1442,N_2350);
xnor U8333 (N_8333,N_4972,N_492);
or U8334 (N_8334,N_520,N_150);
nor U8335 (N_8335,N_4619,N_3526);
or U8336 (N_8336,N_3827,N_4759);
xnor U8337 (N_8337,N_2277,N_3372);
nand U8338 (N_8338,N_4166,N_2757);
nand U8339 (N_8339,N_3271,N_730);
nor U8340 (N_8340,N_3807,N_3117);
and U8341 (N_8341,N_1496,N_1926);
or U8342 (N_8342,N_133,N_829);
and U8343 (N_8343,N_1150,N_2812);
nand U8344 (N_8344,N_1803,N_1942);
xnor U8345 (N_8345,N_1796,N_4738);
nor U8346 (N_8346,N_4953,N_4765);
xnor U8347 (N_8347,N_968,N_1042);
or U8348 (N_8348,N_1812,N_3178);
nor U8349 (N_8349,N_1414,N_1228);
xor U8350 (N_8350,N_2707,N_2610);
nand U8351 (N_8351,N_3650,N_487);
nor U8352 (N_8352,N_4371,N_3356);
xnor U8353 (N_8353,N_3436,N_3218);
nand U8354 (N_8354,N_4274,N_3028);
xor U8355 (N_8355,N_2523,N_3251);
and U8356 (N_8356,N_984,N_1562);
xnor U8357 (N_8357,N_3426,N_432);
or U8358 (N_8358,N_4101,N_509);
nor U8359 (N_8359,N_4717,N_3445);
and U8360 (N_8360,N_112,N_2692);
and U8361 (N_8361,N_2132,N_1060);
or U8362 (N_8362,N_2719,N_776);
xnor U8363 (N_8363,N_4826,N_4638);
xnor U8364 (N_8364,N_1642,N_1356);
nor U8365 (N_8365,N_2197,N_1500);
xor U8366 (N_8366,N_3024,N_4418);
xnor U8367 (N_8367,N_2346,N_1819);
nand U8368 (N_8368,N_2526,N_3793);
nor U8369 (N_8369,N_331,N_4518);
xnor U8370 (N_8370,N_499,N_4468);
and U8371 (N_8371,N_130,N_147);
nor U8372 (N_8372,N_2520,N_3129);
or U8373 (N_8373,N_4003,N_3944);
xnor U8374 (N_8374,N_240,N_4265);
or U8375 (N_8375,N_2005,N_2699);
and U8376 (N_8376,N_272,N_2551);
and U8377 (N_8377,N_2524,N_1609);
nand U8378 (N_8378,N_3583,N_652);
or U8379 (N_8379,N_3194,N_844);
xor U8380 (N_8380,N_1166,N_4802);
or U8381 (N_8381,N_3442,N_1583);
and U8382 (N_8382,N_1327,N_1137);
or U8383 (N_8383,N_727,N_746);
or U8384 (N_8384,N_1874,N_929);
xor U8385 (N_8385,N_4798,N_490);
nor U8386 (N_8386,N_3672,N_1679);
nand U8387 (N_8387,N_4393,N_2855);
xor U8388 (N_8388,N_4058,N_3207);
nor U8389 (N_8389,N_482,N_57);
and U8390 (N_8390,N_2234,N_3380);
or U8391 (N_8391,N_4596,N_3249);
and U8392 (N_8392,N_362,N_1678);
nor U8393 (N_8393,N_4967,N_3196);
nor U8394 (N_8394,N_2889,N_601);
or U8395 (N_8395,N_2962,N_3466);
nand U8396 (N_8396,N_4131,N_2368);
nand U8397 (N_8397,N_317,N_1295);
xnor U8398 (N_8398,N_4479,N_3621);
nor U8399 (N_8399,N_3108,N_4812);
xnor U8400 (N_8400,N_4316,N_2754);
or U8401 (N_8401,N_298,N_2874);
nor U8402 (N_8402,N_647,N_4940);
nand U8403 (N_8403,N_4651,N_3609);
xor U8404 (N_8404,N_1417,N_531);
or U8405 (N_8405,N_83,N_4015);
nand U8406 (N_8406,N_3071,N_1744);
nand U8407 (N_8407,N_1213,N_1947);
xor U8408 (N_8408,N_1392,N_1973);
nor U8409 (N_8409,N_320,N_2656);
nor U8410 (N_8410,N_2544,N_4225);
nor U8411 (N_8411,N_1481,N_1732);
xnor U8412 (N_8412,N_3697,N_1618);
nand U8413 (N_8413,N_3352,N_288);
or U8414 (N_8414,N_354,N_2989);
or U8415 (N_8415,N_3464,N_4268);
nor U8416 (N_8416,N_4568,N_899);
or U8417 (N_8417,N_3594,N_3208);
and U8418 (N_8418,N_3866,N_877);
xor U8419 (N_8419,N_2077,N_855);
xor U8420 (N_8420,N_4028,N_2483);
xnor U8421 (N_8421,N_600,N_2101);
xor U8422 (N_8422,N_790,N_4034);
and U8423 (N_8423,N_2220,N_3075);
or U8424 (N_8424,N_2920,N_60);
nor U8425 (N_8425,N_1310,N_1564);
nand U8426 (N_8426,N_2104,N_3500);
or U8427 (N_8427,N_164,N_1159);
or U8428 (N_8428,N_2371,N_2904);
nor U8429 (N_8429,N_2461,N_454);
nand U8430 (N_8430,N_1413,N_1709);
xor U8431 (N_8431,N_2446,N_2743);
nor U8432 (N_8432,N_605,N_1120);
nand U8433 (N_8433,N_681,N_1964);
nor U8434 (N_8434,N_1553,N_1902);
or U8435 (N_8435,N_2930,N_521);
and U8436 (N_8436,N_3833,N_548);
and U8437 (N_8437,N_2150,N_254);
or U8438 (N_8438,N_1225,N_1319);
xor U8439 (N_8439,N_3794,N_1236);
nor U8440 (N_8440,N_487,N_2131);
nor U8441 (N_8441,N_3828,N_1128);
nor U8442 (N_8442,N_2350,N_3474);
or U8443 (N_8443,N_4845,N_3307);
nor U8444 (N_8444,N_4334,N_4014);
or U8445 (N_8445,N_4824,N_2537);
nor U8446 (N_8446,N_1801,N_2883);
and U8447 (N_8447,N_3957,N_3588);
nor U8448 (N_8448,N_4351,N_873);
xor U8449 (N_8449,N_2530,N_2954);
or U8450 (N_8450,N_282,N_2912);
nor U8451 (N_8451,N_1793,N_3732);
nor U8452 (N_8452,N_2007,N_3841);
nor U8453 (N_8453,N_1799,N_1540);
and U8454 (N_8454,N_4592,N_1991);
xnor U8455 (N_8455,N_2678,N_69);
or U8456 (N_8456,N_2195,N_216);
and U8457 (N_8457,N_4760,N_3932);
nand U8458 (N_8458,N_348,N_1253);
and U8459 (N_8459,N_3008,N_64);
and U8460 (N_8460,N_2870,N_3155);
and U8461 (N_8461,N_3630,N_3846);
xnor U8462 (N_8462,N_822,N_3533);
nor U8463 (N_8463,N_4984,N_4407);
nand U8464 (N_8464,N_2984,N_69);
xnor U8465 (N_8465,N_3201,N_4522);
nand U8466 (N_8466,N_2713,N_3310);
or U8467 (N_8467,N_3206,N_4575);
or U8468 (N_8468,N_3413,N_4821);
nor U8469 (N_8469,N_2694,N_3516);
nand U8470 (N_8470,N_4174,N_3717);
xnor U8471 (N_8471,N_2337,N_1282);
nor U8472 (N_8472,N_4862,N_3269);
nor U8473 (N_8473,N_4850,N_3066);
or U8474 (N_8474,N_3883,N_3493);
and U8475 (N_8475,N_2280,N_1340);
nor U8476 (N_8476,N_98,N_4477);
or U8477 (N_8477,N_1363,N_4997);
xor U8478 (N_8478,N_859,N_4887);
nor U8479 (N_8479,N_1631,N_2081);
or U8480 (N_8480,N_1936,N_808);
nor U8481 (N_8481,N_48,N_115);
and U8482 (N_8482,N_523,N_3805);
and U8483 (N_8483,N_1807,N_3364);
or U8484 (N_8484,N_4237,N_2920);
nor U8485 (N_8485,N_3548,N_1178);
xnor U8486 (N_8486,N_1853,N_3061);
nand U8487 (N_8487,N_2822,N_3907);
and U8488 (N_8488,N_3030,N_1861);
and U8489 (N_8489,N_3482,N_4470);
or U8490 (N_8490,N_1322,N_657);
nor U8491 (N_8491,N_3121,N_3473);
or U8492 (N_8492,N_1092,N_1225);
nand U8493 (N_8493,N_1108,N_4516);
or U8494 (N_8494,N_752,N_479);
nand U8495 (N_8495,N_4918,N_577);
nor U8496 (N_8496,N_1348,N_2421);
xnor U8497 (N_8497,N_695,N_2227);
and U8498 (N_8498,N_4962,N_943);
and U8499 (N_8499,N_2528,N_2233);
or U8500 (N_8500,N_596,N_150);
and U8501 (N_8501,N_3116,N_3723);
and U8502 (N_8502,N_3917,N_3929);
xnor U8503 (N_8503,N_3593,N_4748);
xnor U8504 (N_8504,N_4370,N_4932);
nor U8505 (N_8505,N_4526,N_95);
nor U8506 (N_8506,N_3246,N_1217);
xor U8507 (N_8507,N_4133,N_3955);
nor U8508 (N_8508,N_2119,N_1336);
and U8509 (N_8509,N_2813,N_1233);
nor U8510 (N_8510,N_1068,N_1917);
nand U8511 (N_8511,N_2299,N_266);
nor U8512 (N_8512,N_4533,N_2699);
and U8513 (N_8513,N_250,N_1832);
nand U8514 (N_8514,N_327,N_4374);
nor U8515 (N_8515,N_472,N_3130);
nand U8516 (N_8516,N_4801,N_3449);
xnor U8517 (N_8517,N_2724,N_40);
and U8518 (N_8518,N_4731,N_4952);
and U8519 (N_8519,N_1799,N_98);
nor U8520 (N_8520,N_2350,N_1164);
or U8521 (N_8521,N_1048,N_527);
xnor U8522 (N_8522,N_2381,N_4385);
and U8523 (N_8523,N_4834,N_2511);
nor U8524 (N_8524,N_1016,N_2161);
nor U8525 (N_8525,N_2038,N_3770);
and U8526 (N_8526,N_4319,N_2338);
nand U8527 (N_8527,N_4624,N_737);
xor U8528 (N_8528,N_3255,N_576);
nor U8529 (N_8529,N_1107,N_3651);
nand U8530 (N_8530,N_1063,N_1782);
nand U8531 (N_8531,N_4749,N_4030);
and U8532 (N_8532,N_668,N_4636);
and U8533 (N_8533,N_3221,N_3640);
nor U8534 (N_8534,N_2124,N_2660);
and U8535 (N_8535,N_1222,N_1550);
xor U8536 (N_8536,N_2699,N_3678);
xor U8537 (N_8537,N_3651,N_1974);
or U8538 (N_8538,N_926,N_3357);
and U8539 (N_8539,N_2057,N_1711);
and U8540 (N_8540,N_3159,N_1595);
nor U8541 (N_8541,N_4629,N_1467);
xnor U8542 (N_8542,N_3195,N_368);
and U8543 (N_8543,N_1613,N_3089);
nand U8544 (N_8544,N_4388,N_3671);
nor U8545 (N_8545,N_1049,N_3938);
or U8546 (N_8546,N_1821,N_1173);
nand U8547 (N_8547,N_2713,N_2575);
nand U8548 (N_8548,N_201,N_4283);
nand U8549 (N_8549,N_283,N_130);
or U8550 (N_8550,N_3577,N_3809);
xnor U8551 (N_8551,N_2661,N_2740);
and U8552 (N_8552,N_2588,N_346);
or U8553 (N_8553,N_2250,N_3006);
and U8554 (N_8554,N_904,N_2338);
nand U8555 (N_8555,N_19,N_3996);
nand U8556 (N_8556,N_2829,N_2066);
and U8557 (N_8557,N_4733,N_4525);
and U8558 (N_8558,N_2902,N_2201);
or U8559 (N_8559,N_4468,N_3980);
nand U8560 (N_8560,N_1385,N_3903);
or U8561 (N_8561,N_3652,N_2645);
or U8562 (N_8562,N_3827,N_4712);
and U8563 (N_8563,N_4409,N_573);
xor U8564 (N_8564,N_3347,N_2609);
or U8565 (N_8565,N_2439,N_2399);
xor U8566 (N_8566,N_410,N_2612);
xor U8567 (N_8567,N_1069,N_889);
nand U8568 (N_8568,N_2498,N_1025);
or U8569 (N_8569,N_3537,N_114);
xnor U8570 (N_8570,N_1734,N_3075);
and U8571 (N_8571,N_3548,N_2980);
or U8572 (N_8572,N_1594,N_2435);
and U8573 (N_8573,N_1533,N_3637);
nor U8574 (N_8574,N_1452,N_3071);
nor U8575 (N_8575,N_2030,N_1137);
nand U8576 (N_8576,N_451,N_104);
and U8577 (N_8577,N_2905,N_303);
nand U8578 (N_8578,N_3694,N_419);
nand U8579 (N_8579,N_1799,N_51);
nand U8580 (N_8580,N_3742,N_2138);
and U8581 (N_8581,N_3754,N_4637);
or U8582 (N_8582,N_2915,N_300);
nor U8583 (N_8583,N_526,N_762);
or U8584 (N_8584,N_2238,N_4264);
or U8585 (N_8585,N_972,N_337);
nand U8586 (N_8586,N_448,N_1896);
nor U8587 (N_8587,N_3153,N_1498);
xor U8588 (N_8588,N_3826,N_1945);
nand U8589 (N_8589,N_2887,N_262);
nor U8590 (N_8590,N_4328,N_3867);
or U8591 (N_8591,N_4421,N_3418);
nand U8592 (N_8592,N_165,N_3199);
and U8593 (N_8593,N_3315,N_4466);
xnor U8594 (N_8594,N_4432,N_806);
nor U8595 (N_8595,N_4572,N_2091);
xor U8596 (N_8596,N_1277,N_3443);
nand U8597 (N_8597,N_3976,N_4752);
and U8598 (N_8598,N_1477,N_261);
nand U8599 (N_8599,N_2197,N_133);
or U8600 (N_8600,N_2206,N_778);
or U8601 (N_8601,N_716,N_1960);
xor U8602 (N_8602,N_1104,N_4077);
or U8603 (N_8603,N_1050,N_1661);
xor U8604 (N_8604,N_2172,N_2564);
and U8605 (N_8605,N_138,N_1494);
or U8606 (N_8606,N_1866,N_2731);
nor U8607 (N_8607,N_3066,N_2569);
and U8608 (N_8608,N_2043,N_3606);
xnor U8609 (N_8609,N_4846,N_2800);
nand U8610 (N_8610,N_1342,N_1099);
or U8611 (N_8611,N_3076,N_4699);
nand U8612 (N_8612,N_4367,N_2387);
or U8613 (N_8613,N_1036,N_3070);
nand U8614 (N_8614,N_630,N_2817);
nand U8615 (N_8615,N_3630,N_4489);
nand U8616 (N_8616,N_2428,N_4038);
nor U8617 (N_8617,N_1612,N_3814);
xnor U8618 (N_8618,N_2825,N_2966);
and U8619 (N_8619,N_3839,N_3691);
or U8620 (N_8620,N_1253,N_3543);
nor U8621 (N_8621,N_1497,N_2722);
and U8622 (N_8622,N_3732,N_4786);
nor U8623 (N_8623,N_2749,N_1258);
or U8624 (N_8624,N_2078,N_678);
xor U8625 (N_8625,N_3866,N_872);
nand U8626 (N_8626,N_2774,N_4763);
and U8627 (N_8627,N_4175,N_1463);
xor U8628 (N_8628,N_3670,N_467);
nand U8629 (N_8629,N_2313,N_2549);
nor U8630 (N_8630,N_2269,N_4973);
or U8631 (N_8631,N_1929,N_2997);
or U8632 (N_8632,N_1907,N_1045);
or U8633 (N_8633,N_1208,N_3434);
or U8634 (N_8634,N_3661,N_1266);
or U8635 (N_8635,N_2895,N_3662);
or U8636 (N_8636,N_1977,N_1702);
or U8637 (N_8637,N_598,N_1875);
or U8638 (N_8638,N_3368,N_4092);
or U8639 (N_8639,N_33,N_1455);
or U8640 (N_8640,N_125,N_37);
nor U8641 (N_8641,N_3045,N_1605);
nor U8642 (N_8642,N_608,N_567);
nand U8643 (N_8643,N_1871,N_2808);
or U8644 (N_8644,N_1442,N_869);
nand U8645 (N_8645,N_3398,N_1622);
nor U8646 (N_8646,N_3480,N_1475);
or U8647 (N_8647,N_4831,N_136);
nand U8648 (N_8648,N_1421,N_2948);
and U8649 (N_8649,N_4904,N_4104);
or U8650 (N_8650,N_4677,N_3861);
xor U8651 (N_8651,N_4727,N_3432);
or U8652 (N_8652,N_4903,N_4933);
xor U8653 (N_8653,N_583,N_4660);
or U8654 (N_8654,N_3918,N_2334);
xor U8655 (N_8655,N_802,N_4883);
and U8656 (N_8656,N_71,N_1370);
nand U8657 (N_8657,N_1990,N_953);
nand U8658 (N_8658,N_3975,N_1825);
xor U8659 (N_8659,N_497,N_743);
or U8660 (N_8660,N_3030,N_4717);
nand U8661 (N_8661,N_1180,N_318);
and U8662 (N_8662,N_1318,N_4593);
nor U8663 (N_8663,N_3246,N_2079);
or U8664 (N_8664,N_3072,N_4815);
xnor U8665 (N_8665,N_1872,N_54);
nand U8666 (N_8666,N_1699,N_800);
xor U8667 (N_8667,N_4476,N_1142);
nor U8668 (N_8668,N_1143,N_4734);
or U8669 (N_8669,N_4718,N_1871);
or U8670 (N_8670,N_4095,N_1857);
nand U8671 (N_8671,N_1960,N_1957);
or U8672 (N_8672,N_181,N_3065);
and U8673 (N_8673,N_2729,N_1581);
and U8674 (N_8674,N_777,N_4745);
nor U8675 (N_8675,N_2570,N_1967);
nor U8676 (N_8676,N_3525,N_2836);
nor U8677 (N_8677,N_194,N_1797);
nor U8678 (N_8678,N_2355,N_4310);
xor U8679 (N_8679,N_2202,N_3956);
or U8680 (N_8680,N_4622,N_2666);
and U8681 (N_8681,N_3381,N_3573);
or U8682 (N_8682,N_828,N_3973);
nand U8683 (N_8683,N_1007,N_3102);
or U8684 (N_8684,N_3628,N_2782);
nand U8685 (N_8685,N_7,N_4754);
nand U8686 (N_8686,N_3454,N_3056);
nor U8687 (N_8687,N_187,N_4426);
xor U8688 (N_8688,N_4345,N_3113);
and U8689 (N_8689,N_2714,N_3371);
or U8690 (N_8690,N_3383,N_860);
nor U8691 (N_8691,N_4338,N_4439);
nor U8692 (N_8692,N_2933,N_1265);
or U8693 (N_8693,N_454,N_2521);
and U8694 (N_8694,N_4927,N_3191);
and U8695 (N_8695,N_2932,N_3860);
xnor U8696 (N_8696,N_1023,N_3381);
or U8697 (N_8697,N_1491,N_2126);
nor U8698 (N_8698,N_1137,N_995);
nor U8699 (N_8699,N_3102,N_3548);
and U8700 (N_8700,N_456,N_4969);
nor U8701 (N_8701,N_3014,N_2182);
nor U8702 (N_8702,N_1980,N_292);
and U8703 (N_8703,N_4241,N_2562);
or U8704 (N_8704,N_2076,N_2607);
and U8705 (N_8705,N_1491,N_466);
or U8706 (N_8706,N_52,N_3445);
and U8707 (N_8707,N_3080,N_3120);
nor U8708 (N_8708,N_718,N_2075);
and U8709 (N_8709,N_4815,N_1915);
xnor U8710 (N_8710,N_4470,N_4114);
nand U8711 (N_8711,N_1430,N_3861);
nand U8712 (N_8712,N_2985,N_1235);
nor U8713 (N_8713,N_353,N_2967);
or U8714 (N_8714,N_1173,N_2017);
xnor U8715 (N_8715,N_506,N_2946);
or U8716 (N_8716,N_762,N_3184);
nand U8717 (N_8717,N_1121,N_2387);
nor U8718 (N_8718,N_754,N_2109);
xor U8719 (N_8719,N_1058,N_4323);
and U8720 (N_8720,N_496,N_2987);
or U8721 (N_8721,N_2562,N_4818);
xor U8722 (N_8722,N_4534,N_1119);
and U8723 (N_8723,N_2628,N_3966);
nand U8724 (N_8724,N_3240,N_4460);
and U8725 (N_8725,N_2931,N_324);
nand U8726 (N_8726,N_2934,N_1894);
or U8727 (N_8727,N_405,N_3032);
xor U8728 (N_8728,N_3235,N_977);
nand U8729 (N_8729,N_3930,N_2327);
nand U8730 (N_8730,N_4729,N_1870);
xnor U8731 (N_8731,N_2211,N_125);
nor U8732 (N_8732,N_2565,N_198);
and U8733 (N_8733,N_2478,N_15);
xor U8734 (N_8734,N_3534,N_2609);
or U8735 (N_8735,N_958,N_1003);
and U8736 (N_8736,N_3165,N_3091);
and U8737 (N_8737,N_3773,N_4292);
nand U8738 (N_8738,N_2396,N_3684);
nor U8739 (N_8739,N_3228,N_3285);
and U8740 (N_8740,N_97,N_4194);
and U8741 (N_8741,N_4508,N_3763);
or U8742 (N_8742,N_1134,N_3868);
nand U8743 (N_8743,N_1367,N_629);
or U8744 (N_8744,N_3995,N_4293);
or U8745 (N_8745,N_3401,N_912);
or U8746 (N_8746,N_1968,N_1283);
or U8747 (N_8747,N_3671,N_1046);
nand U8748 (N_8748,N_4559,N_2461);
nor U8749 (N_8749,N_4863,N_3247);
or U8750 (N_8750,N_4920,N_1018);
nand U8751 (N_8751,N_336,N_1670);
nor U8752 (N_8752,N_773,N_99);
nand U8753 (N_8753,N_4746,N_3362);
nand U8754 (N_8754,N_4614,N_3184);
xor U8755 (N_8755,N_3625,N_857);
xnor U8756 (N_8756,N_4186,N_4524);
xnor U8757 (N_8757,N_3918,N_2409);
nand U8758 (N_8758,N_963,N_18);
nand U8759 (N_8759,N_827,N_3964);
nor U8760 (N_8760,N_559,N_2000);
xor U8761 (N_8761,N_60,N_2807);
xnor U8762 (N_8762,N_638,N_1684);
xnor U8763 (N_8763,N_2552,N_968);
nor U8764 (N_8764,N_4826,N_1599);
xor U8765 (N_8765,N_4687,N_4486);
nor U8766 (N_8766,N_4460,N_856);
or U8767 (N_8767,N_3440,N_1145);
nand U8768 (N_8768,N_3922,N_1489);
nand U8769 (N_8769,N_3725,N_1198);
xnor U8770 (N_8770,N_4896,N_3960);
and U8771 (N_8771,N_3493,N_3713);
nor U8772 (N_8772,N_3914,N_3837);
or U8773 (N_8773,N_1168,N_3457);
and U8774 (N_8774,N_4644,N_2847);
nor U8775 (N_8775,N_38,N_1186);
nand U8776 (N_8776,N_1687,N_2457);
xor U8777 (N_8777,N_818,N_1201);
xor U8778 (N_8778,N_1630,N_1216);
nor U8779 (N_8779,N_2560,N_3438);
nor U8780 (N_8780,N_2127,N_2024);
or U8781 (N_8781,N_2207,N_3503);
or U8782 (N_8782,N_4147,N_2952);
xor U8783 (N_8783,N_4616,N_1754);
or U8784 (N_8784,N_4881,N_2391);
xnor U8785 (N_8785,N_874,N_4381);
xor U8786 (N_8786,N_1562,N_768);
and U8787 (N_8787,N_1596,N_4792);
nor U8788 (N_8788,N_63,N_3433);
or U8789 (N_8789,N_1606,N_2922);
and U8790 (N_8790,N_843,N_3971);
or U8791 (N_8791,N_3040,N_1303);
nand U8792 (N_8792,N_1612,N_3276);
nand U8793 (N_8793,N_4494,N_1445);
nand U8794 (N_8794,N_1553,N_2161);
nor U8795 (N_8795,N_1377,N_2330);
and U8796 (N_8796,N_4982,N_1816);
nand U8797 (N_8797,N_1935,N_4959);
and U8798 (N_8798,N_4860,N_3021);
or U8799 (N_8799,N_1363,N_4378);
xor U8800 (N_8800,N_1848,N_2153);
or U8801 (N_8801,N_3585,N_3012);
nor U8802 (N_8802,N_1069,N_4533);
xnor U8803 (N_8803,N_3048,N_720);
or U8804 (N_8804,N_1599,N_4198);
or U8805 (N_8805,N_1603,N_2771);
or U8806 (N_8806,N_748,N_651);
or U8807 (N_8807,N_2143,N_782);
nor U8808 (N_8808,N_1369,N_3679);
xor U8809 (N_8809,N_4183,N_268);
or U8810 (N_8810,N_3704,N_1685);
nand U8811 (N_8811,N_4069,N_2455);
xor U8812 (N_8812,N_213,N_1626);
xor U8813 (N_8813,N_1440,N_2882);
nand U8814 (N_8814,N_3120,N_3773);
xnor U8815 (N_8815,N_3496,N_4303);
or U8816 (N_8816,N_4344,N_3890);
or U8817 (N_8817,N_922,N_2996);
and U8818 (N_8818,N_4078,N_37);
and U8819 (N_8819,N_1114,N_3513);
nor U8820 (N_8820,N_2496,N_4001);
xnor U8821 (N_8821,N_1302,N_4544);
and U8822 (N_8822,N_786,N_4534);
nand U8823 (N_8823,N_990,N_1485);
xnor U8824 (N_8824,N_1888,N_1643);
xnor U8825 (N_8825,N_1320,N_888);
nand U8826 (N_8826,N_888,N_1605);
or U8827 (N_8827,N_3010,N_1563);
nor U8828 (N_8828,N_1703,N_204);
nand U8829 (N_8829,N_4876,N_2122);
and U8830 (N_8830,N_3859,N_1319);
nor U8831 (N_8831,N_204,N_2049);
nand U8832 (N_8832,N_876,N_2020);
xor U8833 (N_8833,N_2290,N_3503);
and U8834 (N_8834,N_113,N_2118);
xor U8835 (N_8835,N_3299,N_1225);
nand U8836 (N_8836,N_2439,N_2007);
and U8837 (N_8837,N_895,N_277);
or U8838 (N_8838,N_3389,N_1998);
or U8839 (N_8839,N_3151,N_1175);
nand U8840 (N_8840,N_4476,N_4191);
and U8841 (N_8841,N_3329,N_129);
nand U8842 (N_8842,N_4054,N_4096);
nor U8843 (N_8843,N_1052,N_3870);
xor U8844 (N_8844,N_2177,N_2164);
xnor U8845 (N_8845,N_4447,N_440);
xnor U8846 (N_8846,N_1579,N_1965);
xnor U8847 (N_8847,N_1987,N_2750);
or U8848 (N_8848,N_1973,N_4361);
xor U8849 (N_8849,N_38,N_2243);
xor U8850 (N_8850,N_3639,N_4817);
and U8851 (N_8851,N_121,N_3648);
or U8852 (N_8852,N_4297,N_2589);
xnor U8853 (N_8853,N_3235,N_2778);
nand U8854 (N_8854,N_4048,N_1588);
nand U8855 (N_8855,N_1890,N_946);
or U8856 (N_8856,N_291,N_914);
and U8857 (N_8857,N_2536,N_420);
nand U8858 (N_8858,N_2290,N_1613);
xor U8859 (N_8859,N_4715,N_2341);
xor U8860 (N_8860,N_1460,N_4426);
xor U8861 (N_8861,N_2060,N_3373);
nor U8862 (N_8862,N_3105,N_1042);
xnor U8863 (N_8863,N_2920,N_455);
nor U8864 (N_8864,N_1615,N_1026);
nor U8865 (N_8865,N_3319,N_2704);
or U8866 (N_8866,N_3238,N_4799);
nor U8867 (N_8867,N_4941,N_266);
nand U8868 (N_8868,N_1984,N_4999);
xor U8869 (N_8869,N_3998,N_1517);
nor U8870 (N_8870,N_3599,N_3176);
nor U8871 (N_8871,N_4407,N_761);
nand U8872 (N_8872,N_4275,N_1920);
or U8873 (N_8873,N_1565,N_4132);
nor U8874 (N_8874,N_2396,N_4938);
and U8875 (N_8875,N_2201,N_979);
and U8876 (N_8876,N_881,N_1747);
nor U8877 (N_8877,N_785,N_4723);
xnor U8878 (N_8878,N_3845,N_998);
nand U8879 (N_8879,N_865,N_2624);
or U8880 (N_8880,N_4786,N_1381);
xnor U8881 (N_8881,N_3547,N_183);
nand U8882 (N_8882,N_336,N_1059);
and U8883 (N_8883,N_900,N_3164);
xnor U8884 (N_8884,N_2952,N_515);
or U8885 (N_8885,N_3063,N_2531);
nand U8886 (N_8886,N_3926,N_1085);
nor U8887 (N_8887,N_1219,N_4413);
xnor U8888 (N_8888,N_675,N_2282);
nand U8889 (N_8889,N_4324,N_2260);
nor U8890 (N_8890,N_744,N_168);
nor U8891 (N_8891,N_661,N_3438);
xor U8892 (N_8892,N_224,N_3745);
and U8893 (N_8893,N_3089,N_2021);
xnor U8894 (N_8894,N_911,N_4194);
xor U8895 (N_8895,N_1794,N_4392);
and U8896 (N_8896,N_1141,N_564);
nor U8897 (N_8897,N_1207,N_2352);
or U8898 (N_8898,N_3457,N_1862);
and U8899 (N_8899,N_259,N_2394);
xnor U8900 (N_8900,N_381,N_463);
nand U8901 (N_8901,N_2310,N_819);
xnor U8902 (N_8902,N_3702,N_1801);
and U8903 (N_8903,N_4751,N_4012);
nor U8904 (N_8904,N_3830,N_2976);
nor U8905 (N_8905,N_4354,N_560);
or U8906 (N_8906,N_4055,N_3214);
xnor U8907 (N_8907,N_1658,N_1878);
or U8908 (N_8908,N_838,N_2394);
or U8909 (N_8909,N_3834,N_3993);
or U8910 (N_8910,N_120,N_548);
nor U8911 (N_8911,N_4437,N_2106);
xor U8912 (N_8912,N_3585,N_4559);
nand U8913 (N_8913,N_712,N_4088);
or U8914 (N_8914,N_4343,N_3567);
xnor U8915 (N_8915,N_2738,N_1049);
nor U8916 (N_8916,N_937,N_4151);
or U8917 (N_8917,N_1489,N_605);
nor U8918 (N_8918,N_4336,N_4946);
xnor U8919 (N_8919,N_1836,N_4667);
or U8920 (N_8920,N_37,N_2770);
nand U8921 (N_8921,N_414,N_1642);
nand U8922 (N_8922,N_4116,N_1978);
and U8923 (N_8923,N_2820,N_1578);
xnor U8924 (N_8924,N_4551,N_4625);
nand U8925 (N_8925,N_1739,N_4952);
and U8926 (N_8926,N_1660,N_975);
or U8927 (N_8927,N_4595,N_201);
nand U8928 (N_8928,N_3719,N_439);
nor U8929 (N_8929,N_3019,N_3486);
nand U8930 (N_8930,N_3424,N_3620);
nand U8931 (N_8931,N_2508,N_3260);
xnor U8932 (N_8932,N_2956,N_386);
or U8933 (N_8933,N_1936,N_590);
xnor U8934 (N_8934,N_1898,N_4859);
nand U8935 (N_8935,N_4319,N_580);
and U8936 (N_8936,N_1215,N_722);
nor U8937 (N_8937,N_4117,N_208);
xnor U8938 (N_8938,N_41,N_23);
and U8939 (N_8939,N_1369,N_2926);
nor U8940 (N_8940,N_1059,N_1478);
nand U8941 (N_8941,N_825,N_88);
and U8942 (N_8942,N_1623,N_2660);
or U8943 (N_8943,N_4455,N_548);
xor U8944 (N_8944,N_129,N_3045);
nand U8945 (N_8945,N_3544,N_1791);
or U8946 (N_8946,N_3345,N_3179);
and U8947 (N_8947,N_3844,N_848);
xor U8948 (N_8948,N_645,N_1751);
or U8949 (N_8949,N_2623,N_4161);
and U8950 (N_8950,N_273,N_2479);
xor U8951 (N_8951,N_3770,N_2238);
xnor U8952 (N_8952,N_3191,N_316);
nand U8953 (N_8953,N_2426,N_3735);
nand U8954 (N_8954,N_3320,N_4045);
xor U8955 (N_8955,N_1518,N_4540);
or U8956 (N_8956,N_1648,N_764);
nand U8957 (N_8957,N_2160,N_1448);
nand U8958 (N_8958,N_354,N_3399);
and U8959 (N_8959,N_3380,N_646);
nor U8960 (N_8960,N_22,N_321);
nor U8961 (N_8961,N_3105,N_4161);
nor U8962 (N_8962,N_163,N_192);
nor U8963 (N_8963,N_4,N_1849);
xor U8964 (N_8964,N_1927,N_3321);
xor U8965 (N_8965,N_609,N_3530);
xnor U8966 (N_8966,N_260,N_1206);
nand U8967 (N_8967,N_1606,N_4582);
nor U8968 (N_8968,N_82,N_3354);
or U8969 (N_8969,N_3255,N_3958);
nand U8970 (N_8970,N_1957,N_4528);
nand U8971 (N_8971,N_778,N_1139);
xnor U8972 (N_8972,N_2005,N_1051);
or U8973 (N_8973,N_121,N_2398);
xor U8974 (N_8974,N_2287,N_4678);
and U8975 (N_8975,N_13,N_878);
nor U8976 (N_8976,N_3685,N_1129);
nor U8977 (N_8977,N_1616,N_706);
nor U8978 (N_8978,N_1153,N_2744);
nand U8979 (N_8979,N_2793,N_650);
nor U8980 (N_8980,N_1140,N_2052);
xor U8981 (N_8981,N_1800,N_2509);
xor U8982 (N_8982,N_4436,N_1126);
or U8983 (N_8983,N_315,N_3178);
or U8984 (N_8984,N_592,N_4938);
or U8985 (N_8985,N_543,N_3077);
xor U8986 (N_8986,N_1542,N_3290);
and U8987 (N_8987,N_733,N_3237);
xnor U8988 (N_8988,N_1043,N_768);
xnor U8989 (N_8989,N_2239,N_4919);
nor U8990 (N_8990,N_1892,N_1487);
xnor U8991 (N_8991,N_540,N_2073);
nor U8992 (N_8992,N_617,N_787);
nor U8993 (N_8993,N_2442,N_4800);
or U8994 (N_8994,N_1273,N_1403);
or U8995 (N_8995,N_4267,N_1512);
xnor U8996 (N_8996,N_2357,N_2901);
and U8997 (N_8997,N_683,N_4510);
nor U8998 (N_8998,N_4603,N_1282);
or U8999 (N_8999,N_3773,N_2313);
nand U9000 (N_9000,N_4662,N_2368);
xnor U9001 (N_9001,N_2684,N_2353);
or U9002 (N_9002,N_3538,N_31);
nand U9003 (N_9003,N_3663,N_3304);
nor U9004 (N_9004,N_3231,N_1534);
nor U9005 (N_9005,N_809,N_4548);
and U9006 (N_9006,N_3078,N_2538);
nor U9007 (N_9007,N_3003,N_2729);
xor U9008 (N_9008,N_3222,N_999);
nor U9009 (N_9009,N_2889,N_1085);
nor U9010 (N_9010,N_4529,N_883);
xor U9011 (N_9011,N_4810,N_2220);
nor U9012 (N_9012,N_2442,N_2631);
and U9013 (N_9013,N_608,N_2308);
and U9014 (N_9014,N_1629,N_1757);
xnor U9015 (N_9015,N_3060,N_1786);
nor U9016 (N_9016,N_4500,N_3024);
nor U9017 (N_9017,N_2389,N_476);
nor U9018 (N_9018,N_2447,N_1755);
or U9019 (N_9019,N_1882,N_548);
xor U9020 (N_9020,N_3840,N_537);
xor U9021 (N_9021,N_3506,N_3447);
and U9022 (N_9022,N_660,N_4393);
or U9023 (N_9023,N_3033,N_3831);
or U9024 (N_9024,N_944,N_781);
and U9025 (N_9025,N_238,N_3070);
xnor U9026 (N_9026,N_2655,N_2775);
or U9027 (N_9027,N_971,N_3976);
or U9028 (N_9028,N_4804,N_3940);
nor U9029 (N_9029,N_3642,N_1741);
nor U9030 (N_9030,N_1657,N_3530);
and U9031 (N_9031,N_3329,N_4149);
and U9032 (N_9032,N_2986,N_3999);
nand U9033 (N_9033,N_2009,N_2533);
nor U9034 (N_9034,N_4314,N_4689);
nor U9035 (N_9035,N_4058,N_1228);
nor U9036 (N_9036,N_3155,N_4741);
and U9037 (N_9037,N_4974,N_1135);
nor U9038 (N_9038,N_2413,N_3230);
and U9039 (N_9039,N_90,N_1792);
and U9040 (N_9040,N_1323,N_854);
nand U9041 (N_9041,N_3566,N_223);
and U9042 (N_9042,N_3518,N_1453);
and U9043 (N_9043,N_4043,N_3429);
nand U9044 (N_9044,N_3334,N_4651);
nand U9045 (N_9045,N_1182,N_3334);
nand U9046 (N_9046,N_595,N_4280);
nor U9047 (N_9047,N_2859,N_1880);
nor U9048 (N_9048,N_1425,N_4186);
and U9049 (N_9049,N_3491,N_3763);
nand U9050 (N_9050,N_4577,N_2836);
nor U9051 (N_9051,N_4787,N_1118);
and U9052 (N_9052,N_1398,N_1206);
nand U9053 (N_9053,N_547,N_1977);
and U9054 (N_9054,N_1255,N_746);
and U9055 (N_9055,N_1756,N_1492);
xor U9056 (N_9056,N_3266,N_3056);
nor U9057 (N_9057,N_2282,N_2498);
and U9058 (N_9058,N_2746,N_95);
or U9059 (N_9059,N_2533,N_1016);
or U9060 (N_9060,N_2984,N_4618);
xnor U9061 (N_9061,N_4219,N_971);
xor U9062 (N_9062,N_3502,N_2948);
and U9063 (N_9063,N_3526,N_710);
or U9064 (N_9064,N_3799,N_4731);
nor U9065 (N_9065,N_4443,N_839);
nor U9066 (N_9066,N_4406,N_108);
nor U9067 (N_9067,N_3399,N_3973);
nand U9068 (N_9068,N_3936,N_2550);
and U9069 (N_9069,N_3733,N_2542);
nand U9070 (N_9070,N_2321,N_1263);
or U9071 (N_9071,N_3488,N_622);
xor U9072 (N_9072,N_2902,N_4352);
nand U9073 (N_9073,N_3602,N_3268);
nor U9074 (N_9074,N_1235,N_3480);
nand U9075 (N_9075,N_616,N_51);
nor U9076 (N_9076,N_4143,N_1941);
or U9077 (N_9077,N_3467,N_573);
xor U9078 (N_9078,N_2620,N_3458);
nor U9079 (N_9079,N_3683,N_1568);
or U9080 (N_9080,N_1042,N_3963);
nor U9081 (N_9081,N_4276,N_4003);
nand U9082 (N_9082,N_2703,N_388);
and U9083 (N_9083,N_3276,N_3541);
nor U9084 (N_9084,N_1322,N_980);
and U9085 (N_9085,N_2265,N_348);
or U9086 (N_9086,N_1853,N_4356);
nor U9087 (N_9087,N_4428,N_4685);
xor U9088 (N_9088,N_1524,N_2224);
xor U9089 (N_9089,N_1645,N_1045);
and U9090 (N_9090,N_3369,N_3124);
xnor U9091 (N_9091,N_4233,N_3930);
nand U9092 (N_9092,N_3789,N_3140);
nor U9093 (N_9093,N_3293,N_3430);
and U9094 (N_9094,N_745,N_2121);
xnor U9095 (N_9095,N_1383,N_3839);
xor U9096 (N_9096,N_1722,N_3190);
nand U9097 (N_9097,N_1944,N_1594);
nand U9098 (N_9098,N_2810,N_3933);
nor U9099 (N_9099,N_1187,N_3577);
nor U9100 (N_9100,N_4879,N_2580);
nor U9101 (N_9101,N_1215,N_4457);
and U9102 (N_9102,N_4218,N_3521);
or U9103 (N_9103,N_1361,N_2608);
and U9104 (N_9104,N_2512,N_839);
and U9105 (N_9105,N_1017,N_2309);
nor U9106 (N_9106,N_2702,N_4452);
nor U9107 (N_9107,N_4240,N_2043);
or U9108 (N_9108,N_4655,N_4233);
xnor U9109 (N_9109,N_1434,N_993);
or U9110 (N_9110,N_878,N_1569);
and U9111 (N_9111,N_4672,N_3052);
and U9112 (N_9112,N_143,N_1583);
nor U9113 (N_9113,N_1950,N_3620);
xor U9114 (N_9114,N_3304,N_3226);
and U9115 (N_9115,N_2083,N_4087);
xnor U9116 (N_9116,N_3146,N_4840);
or U9117 (N_9117,N_1861,N_2411);
nand U9118 (N_9118,N_3933,N_2454);
nor U9119 (N_9119,N_3816,N_3380);
nor U9120 (N_9120,N_4390,N_810);
nand U9121 (N_9121,N_3933,N_413);
or U9122 (N_9122,N_2312,N_2836);
xor U9123 (N_9123,N_774,N_4858);
and U9124 (N_9124,N_3474,N_3447);
or U9125 (N_9125,N_4532,N_888);
nand U9126 (N_9126,N_3713,N_3484);
nor U9127 (N_9127,N_1710,N_3911);
nand U9128 (N_9128,N_2734,N_3642);
or U9129 (N_9129,N_3233,N_4740);
or U9130 (N_9130,N_3727,N_684);
xnor U9131 (N_9131,N_1389,N_4019);
or U9132 (N_9132,N_2614,N_4540);
or U9133 (N_9133,N_3812,N_109);
nand U9134 (N_9134,N_2898,N_3802);
or U9135 (N_9135,N_1725,N_4791);
nand U9136 (N_9136,N_1725,N_1546);
xnor U9137 (N_9137,N_3327,N_3986);
nor U9138 (N_9138,N_4430,N_4520);
and U9139 (N_9139,N_1490,N_966);
nand U9140 (N_9140,N_3144,N_4356);
nor U9141 (N_9141,N_3182,N_4182);
nor U9142 (N_9142,N_4285,N_1983);
nor U9143 (N_9143,N_3314,N_4101);
xor U9144 (N_9144,N_1099,N_1007);
or U9145 (N_9145,N_4599,N_4543);
or U9146 (N_9146,N_1427,N_4545);
nand U9147 (N_9147,N_1971,N_3639);
nor U9148 (N_9148,N_4803,N_2339);
xor U9149 (N_9149,N_4210,N_1905);
and U9150 (N_9150,N_2638,N_1692);
or U9151 (N_9151,N_2766,N_3200);
nor U9152 (N_9152,N_425,N_3519);
or U9153 (N_9153,N_1628,N_4596);
and U9154 (N_9154,N_2943,N_2445);
nand U9155 (N_9155,N_4458,N_571);
xnor U9156 (N_9156,N_2811,N_1785);
nor U9157 (N_9157,N_39,N_3319);
or U9158 (N_9158,N_4825,N_2014);
nand U9159 (N_9159,N_2670,N_145);
nand U9160 (N_9160,N_1591,N_2119);
nand U9161 (N_9161,N_1093,N_4129);
and U9162 (N_9162,N_1909,N_1205);
nor U9163 (N_9163,N_3238,N_361);
nor U9164 (N_9164,N_2984,N_2171);
nor U9165 (N_9165,N_2463,N_1252);
nand U9166 (N_9166,N_2626,N_3907);
or U9167 (N_9167,N_2607,N_2207);
and U9168 (N_9168,N_2066,N_1711);
nand U9169 (N_9169,N_2873,N_1942);
nand U9170 (N_9170,N_2126,N_4648);
and U9171 (N_9171,N_4813,N_3345);
nor U9172 (N_9172,N_4134,N_4040);
or U9173 (N_9173,N_1860,N_3691);
and U9174 (N_9174,N_1659,N_3016);
nor U9175 (N_9175,N_1056,N_470);
or U9176 (N_9176,N_561,N_4280);
or U9177 (N_9177,N_2943,N_2688);
and U9178 (N_9178,N_4328,N_4469);
and U9179 (N_9179,N_2509,N_690);
and U9180 (N_9180,N_1585,N_1784);
and U9181 (N_9181,N_792,N_3986);
nor U9182 (N_9182,N_4938,N_4085);
and U9183 (N_9183,N_2680,N_4808);
nor U9184 (N_9184,N_3645,N_2025);
and U9185 (N_9185,N_3514,N_2174);
nor U9186 (N_9186,N_3623,N_4537);
or U9187 (N_9187,N_1970,N_2942);
nor U9188 (N_9188,N_387,N_1718);
or U9189 (N_9189,N_1122,N_1616);
or U9190 (N_9190,N_864,N_899);
xor U9191 (N_9191,N_3702,N_3348);
or U9192 (N_9192,N_2034,N_1826);
xor U9193 (N_9193,N_4259,N_3370);
xor U9194 (N_9194,N_1759,N_4772);
and U9195 (N_9195,N_1044,N_2844);
nor U9196 (N_9196,N_2138,N_3741);
or U9197 (N_9197,N_2569,N_1741);
nor U9198 (N_9198,N_2663,N_1033);
nor U9199 (N_9199,N_3489,N_1365);
xnor U9200 (N_9200,N_1333,N_165);
nor U9201 (N_9201,N_526,N_2437);
or U9202 (N_9202,N_1988,N_2816);
nand U9203 (N_9203,N_4152,N_3129);
or U9204 (N_9204,N_2262,N_4097);
xor U9205 (N_9205,N_4597,N_4473);
or U9206 (N_9206,N_311,N_117);
nand U9207 (N_9207,N_2364,N_36);
nand U9208 (N_9208,N_400,N_2283);
nand U9209 (N_9209,N_4969,N_528);
and U9210 (N_9210,N_4772,N_4864);
or U9211 (N_9211,N_3901,N_4110);
nor U9212 (N_9212,N_2018,N_1255);
xor U9213 (N_9213,N_2846,N_740);
xnor U9214 (N_9214,N_311,N_2971);
nand U9215 (N_9215,N_4314,N_2326);
and U9216 (N_9216,N_1462,N_1308);
nand U9217 (N_9217,N_4372,N_4148);
and U9218 (N_9218,N_1518,N_923);
nand U9219 (N_9219,N_127,N_1705);
and U9220 (N_9220,N_4177,N_4539);
nand U9221 (N_9221,N_2964,N_1656);
xor U9222 (N_9222,N_4381,N_1335);
or U9223 (N_9223,N_3070,N_4453);
nand U9224 (N_9224,N_2939,N_628);
and U9225 (N_9225,N_3158,N_973);
nand U9226 (N_9226,N_1745,N_3197);
or U9227 (N_9227,N_1771,N_2183);
nand U9228 (N_9228,N_1268,N_3581);
nor U9229 (N_9229,N_1599,N_4696);
and U9230 (N_9230,N_4730,N_3256);
xnor U9231 (N_9231,N_4767,N_4986);
nor U9232 (N_9232,N_3490,N_755);
nor U9233 (N_9233,N_3060,N_4564);
nor U9234 (N_9234,N_2508,N_2582);
xnor U9235 (N_9235,N_3457,N_3418);
and U9236 (N_9236,N_3627,N_1784);
and U9237 (N_9237,N_882,N_4166);
xor U9238 (N_9238,N_4912,N_3328);
nand U9239 (N_9239,N_3485,N_4323);
nor U9240 (N_9240,N_2379,N_2866);
or U9241 (N_9241,N_3907,N_1157);
xnor U9242 (N_9242,N_3100,N_878);
and U9243 (N_9243,N_2581,N_1026);
and U9244 (N_9244,N_4990,N_921);
nand U9245 (N_9245,N_4245,N_2652);
and U9246 (N_9246,N_3187,N_3086);
nor U9247 (N_9247,N_3145,N_3994);
xor U9248 (N_9248,N_4625,N_4674);
xor U9249 (N_9249,N_2769,N_1326);
nor U9250 (N_9250,N_2845,N_4201);
or U9251 (N_9251,N_3486,N_1188);
nand U9252 (N_9252,N_866,N_933);
and U9253 (N_9253,N_2308,N_3951);
and U9254 (N_9254,N_1568,N_3875);
and U9255 (N_9255,N_2073,N_1982);
nand U9256 (N_9256,N_1355,N_4205);
nor U9257 (N_9257,N_4824,N_1948);
xor U9258 (N_9258,N_3865,N_4674);
nor U9259 (N_9259,N_4655,N_4566);
nor U9260 (N_9260,N_1186,N_1592);
xnor U9261 (N_9261,N_1577,N_4916);
nand U9262 (N_9262,N_2436,N_1768);
nor U9263 (N_9263,N_4527,N_2925);
xnor U9264 (N_9264,N_3845,N_4071);
nor U9265 (N_9265,N_1266,N_1790);
nor U9266 (N_9266,N_3459,N_522);
and U9267 (N_9267,N_1715,N_1584);
nor U9268 (N_9268,N_3192,N_1036);
or U9269 (N_9269,N_3010,N_3579);
nand U9270 (N_9270,N_4217,N_4071);
or U9271 (N_9271,N_2656,N_3907);
nor U9272 (N_9272,N_4400,N_1750);
nor U9273 (N_9273,N_1448,N_2652);
nor U9274 (N_9274,N_25,N_4710);
xnor U9275 (N_9275,N_3398,N_2901);
or U9276 (N_9276,N_690,N_12);
or U9277 (N_9277,N_3769,N_4833);
nor U9278 (N_9278,N_3764,N_3905);
and U9279 (N_9279,N_1122,N_4398);
nor U9280 (N_9280,N_242,N_1124);
and U9281 (N_9281,N_3116,N_4077);
xnor U9282 (N_9282,N_3029,N_1144);
or U9283 (N_9283,N_2064,N_1256);
and U9284 (N_9284,N_1671,N_78);
nand U9285 (N_9285,N_3824,N_4623);
nor U9286 (N_9286,N_1231,N_241);
nand U9287 (N_9287,N_3114,N_2435);
and U9288 (N_9288,N_1983,N_4515);
or U9289 (N_9289,N_1684,N_3007);
nor U9290 (N_9290,N_4477,N_1186);
nand U9291 (N_9291,N_1444,N_3756);
or U9292 (N_9292,N_575,N_2685);
nor U9293 (N_9293,N_3008,N_3186);
nand U9294 (N_9294,N_2836,N_1070);
nor U9295 (N_9295,N_1797,N_3971);
xor U9296 (N_9296,N_2988,N_4592);
xnor U9297 (N_9297,N_517,N_532);
and U9298 (N_9298,N_1318,N_11);
xnor U9299 (N_9299,N_3627,N_3744);
or U9300 (N_9300,N_1073,N_621);
and U9301 (N_9301,N_2533,N_4547);
and U9302 (N_9302,N_651,N_302);
xnor U9303 (N_9303,N_4678,N_141);
xnor U9304 (N_9304,N_2254,N_1898);
nor U9305 (N_9305,N_2346,N_227);
and U9306 (N_9306,N_746,N_853);
or U9307 (N_9307,N_1279,N_891);
nand U9308 (N_9308,N_2868,N_2811);
and U9309 (N_9309,N_1584,N_972);
xor U9310 (N_9310,N_1199,N_2940);
xor U9311 (N_9311,N_4325,N_66);
or U9312 (N_9312,N_2213,N_4284);
xor U9313 (N_9313,N_4001,N_3711);
xnor U9314 (N_9314,N_4046,N_1737);
nand U9315 (N_9315,N_258,N_2591);
and U9316 (N_9316,N_4297,N_2492);
nand U9317 (N_9317,N_1373,N_3256);
nand U9318 (N_9318,N_2796,N_3675);
nand U9319 (N_9319,N_1629,N_3764);
nor U9320 (N_9320,N_4198,N_34);
xor U9321 (N_9321,N_4804,N_2798);
xnor U9322 (N_9322,N_233,N_4534);
nor U9323 (N_9323,N_1815,N_4691);
nor U9324 (N_9324,N_4880,N_2015);
or U9325 (N_9325,N_4028,N_4873);
xnor U9326 (N_9326,N_1395,N_4885);
nand U9327 (N_9327,N_1980,N_2459);
nor U9328 (N_9328,N_1649,N_189);
nand U9329 (N_9329,N_2376,N_1029);
nor U9330 (N_9330,N_4034,N_1279);
xnor U9331 (N_9331,N_4552,N_3652);
or U9332 (N_9332,N_79,N_2891);
nor U9333 (N_9333,N_2122,N_4920);
xor U9334 (N_9334,N_3417,N_1392);
or U9335 (N_9335,N_2896,N_568);
or U9336 (N_9336,N_1281,N_4778);
nand U9337 (N_9337,N_1495,N_3545);
or U9338 (N_9338,N_476,N_4466);
nor U9339 (N_9339,N_1494,N_865);
or U9340 (N_9340,N_1925,N_3987);
or U9341 (N_9341,N_611,N_1525);
or U9342 (N_9342,N_2017,N_2087);
nand U9343 (N_9343,N_2233,N_1555);
xor U9344 (N_9344,N_3813,N_3290);
xor U9345 (N_9345,N_3895,N_4156);
and U9346 (N_9346,N_2887,N_3260);
and U9347 (N_9347,N_89,N_4198);
xor U9348 (N_9348,N_4013,N_4218);
or U9349 (N_9349,N_1333,N_191);
nor U9350 (N_9350,N_4248,N_4777);
xor U9351 (N_9351,N_915,N_3116);
xnor U9352 (N_9352,N_3462,N_1036);
or U9353 (N_9353,N_4245,N_740);
nor U9354 (N_9354,N_1541,N_3552);
and U9355 (N_9355,N_2040,N_1003);
nand U9356 (N_9356,N_2974,N_864);
xor U9357 (N_9357,N_1574,N_1371);
xnor U9358 (N_9358,N_3096,N_3236);
nor U9359 (N_9359,N_1845,N_1201);
or U9360 (N_9360,N_3997,N_2135);
nand U9361 (N_9361,N_540,N_2429);
nand U9362 (N_9362,N_526,N_1139);
or U9363 (N_9363,N_1651,N_373);
nor U9364 (N_9364,N_4931,N_1880);
or U9365 (N_9365,N_840,N_959);
or U9366 (N_9366,N_4841,N_1509);
nand U9367 (N_9367,N_564,N_1366);
nand U9368 (N_9368,N_1522,N_2978);
xor U9369 (N_9369,N_1537,N_4);
and U9370 (N_9370,N_4283,N_3213);
and U9371 (N_9371,N_3263,N_1280);
or U9372 (N_9372,N_1751,N_2906);
or U9373 (N_9373,N_118,N_3709);
or U9374 (N_9374,N_1627,N_3800);
or U9375 (N_9375,N_821,N_4762);
or U9376 (N_9376,N_519,N_1104);
nor U9377 (N_9377,N_201,N_2521);
xnor U9378 (N_9378,N_18,N_3445);
or U9379 (N_9379,N_4021,N_3598);
nand U9380 (N_9380,N_259,N_4779);
nand U9381 (N_9381,N_333,N_3201);
xor U9382 (N_9382,N_1097,N_630);
and U9383 (N_9383,N_139,N_3839);
or U9384 (N_9384,N_4058,N_647);
nand U9385 (N_9385,N_291,N_1606);
xor U9386 (N_9386,N_4188,N_2824);
nand U9387 (N_9387,N_1812,N_875);
nor U9388 (N_9388,N_2251,N_974);
and U9389 (N_9389,N_4516,N_3819);
nand U9390 (N_9390,N_1917,N_1854);
xor U9391 (N_9391,N_2307,N_4758);
or U9392 (N_9392,N_3040,N_1275);
and U9393 (N_9393,N_956,N_1639);
and U9394 (N_9394,N_2384,N_3331);
xnor U9395 (N_9395,N_410,N_903);
nor U9396 (N_9396,N_2989,N_3573);
nand U9397 (N_9397,N_2218,N_4356);
or U9398 (N_9398,N_1784,N_941);
xnor U9399 (N_9399,N_3698,N_1494);
nor U9400 (N_9400,N_3283,N_340);
or U9401 (N_9401,N_3687,N_1536);
nand U9402 (N_9402,N_1211,N_2696);
xnor U9403 (N_9403,N_508,N_1729);
and U9404 (N_9404,N_2411,N_2631);
and U9405 (N_9405,N_4446,N_4033);
nor U9406 (N_9406,N_916,N_2696);
and U9407 (N_9407,N_2637,N_1657);
or U9408 (N_9408,N_2985,N_4369);
or U9409 (N_9409,N_194,N_1647);
and U9410 (N_9410,N_3506,N_4957);
nor U9411 (N_9411,N_4770,N_4149);
and U9412 (N_9412,N_4735,N_654);
xnor U9413 (N_9413,N_323,N_3384);
nand U9414 (N_9414,N_2408,N_2153);
nor U9415 (N_9415,N_3161,N_48);
nand U9416 (N_9416,N_810,N_577);
nand U9417 (N_9417,N_3230,N_3692);
xor U9418 (N_9418,N_4239,N_4351);
nor U9419 (N_9419,N_2573,N_2617);
nand U9420 (N_9420,N_2268,N_3844);
xnor U9421 (N_9421,N_3243,N_1949);
xor U9422 (N_9422,N_2169,N_2);
xnor U9423 (N_9423,N_3036,N_629);
or U9424 (N_9424,N_849,N_2252);
and U9425 (N_9425,N_1715,N_1623);
nor U9426 (N_9426,N_1312,N_1191);
or U9427 (N_9427,N_1954,N_1465);
xor U9428 (N_9428,N_3679,N_4483);
and U9429 (N_9429,N_3225,N_2260);
nand U9430 (N_9430,N_3502,N_1095);
or U9431 (N_9431,N_2654,N_3859);
and U9432 (N_9432,N_388,N_4319);
nor U9433 (N_9433,N_4689,N_93);
or U9434 (N_9434,N_4180,N_3396);
nor U9435 (N_9435,N_1678,N_1156);
nand U9436 (N_9436,N_502,N_2519);
or U9437 (N_9437,N_276,N_813);
and U9438 (N_9438,N_1631,N_3277);
nand U9439 (N_9439,N_4792,N_3252);
xnor U9440 (N_9440,N_4431,N_2666);
nand U9441 (N_9441,N_258,N_4744);
or U9442 (N_9442,N_1535,N_1807);
or U9443 (N_9443,N_918,N_1497);
xnor U9444 (N_9444,N_3637,N_447);
xnor U9445 (N_9445,N_1904,N_3345);
or U9446 (N_9446,N_3189,N_781);
nor U9447 (N_9447,N_1503,N_4160);
or U9448 (N_9448,N_2491,N_3185);
and U9449 (N_9449,N_1894,N_1859);
xor U9450 (N_9450,N_4840,N_941);
and U9451 (N_9451,N_338,N_2330);
xnor U9452 (N_9452,N_4601,N_2265);
and U9453 (N_9453,N_1101,N_3997);
nand U9454 (N_9454,N_577,N_1665);
and U9455 (N_9455,N_1188,N_2392);
or U9456 (N_9456,N_2247,N_3934);
nand U9457 (N_9457,N_3749,N_4318);
nand U9458 (N_9458,N_4316,N_3292);
nor U9459 (N_9459,N_3378,N_3337);
or U9460 (N_9460,N_4423,N_2943);
xor U9461 (N_9461,N_1675,N_4952);
nor U9462 (N_9462,N_3195,N_4230);
xnor U9463 (N_9463,N_1668,N_4713);
nand U9464 (N_9464,N_4416,N_3663);
or U9465 (N_9465,N_3191,N_4741);
or U9466 (N_9466,N_1903,N_428);
xnor U9467 (N_9467,N_2468,N_1504);
and U9468 (N_9468,N_3397,N_2857);
or U9469 (N_9469,N_4636,N_1069);
nand U9470 (N_9470,N_4686,N_3413);
xor U9471 (N_9471,N_644,N_329);
xor U9472 (N_9472,N_2352,N_2254);
nand U9473 (N_9473,N_3081,N_3881);
nand U9474 (N_9474,N_139,N_585);
nor U9475 (N_9475,N_2442,N_296);
and U9476 (N_9476,N_2752,N_4552);
and U9477 (N_9477,N_3641,N_4065);
xnor U9478 (N_9478,N_1520,N_770);
nand U9479 (N_9479,N_1830,N_3406);
and U9480 (N_9480,N_46,N_4905);
xnor U9481 (N_9481,N_1503,N_109);
nand U9482 (N_9482,N_488,N_4388);
nor U9483 (N_9483,N_2747,N_55);
xnor U9484 (N_9484,N_4567,N_1223);
xnor U9485 (N_9485,N_1868,N_77);
or U9486 (N_9486,N_2045,N_2454);
nand U9487 (N_9487,N_4825,N_1207);
nand U9488 (N_9488,N_4560,N_1613);
nand U9489 (N_9489,N_3475,N_858);
and U9490 (N_9490,N_4524,N_4566);
xnor U9491 (N_9491,N_4255,N_2988);
nor U9492 (N_9492,N_2170,N_507);
nand U9493 (N_9493,N_2531,N_4028);
and U9494 (N_9494,N_2910,N_2927);
nand U9495 (N_9495,N_1039,N_1365);
nor U9496 (N_9496,N_3360,N_162);
and U9497 (N_9497,N_3250,N_4927);
xor U9498 (N_9498,N_3336,N_347);
nor U9499 (N_9499,N_3473,N_1211);
and U9500 (N_9500,N_1310,N_4733);
or U9501 (N_9501,N_1062,N_4626);
nor U9502 (N_9502,N_813,N_4606);
nor U9503 (N_9503,N_1134,N_1611);
and U9504 (N_9504,N_1067,N_2659);
or U9505 (N_9505,N_1736,N_60);
and U9506 (N_9506,N_2822,N_457);
nand U9507 (N_9507,N_292,N_4804);
xnor U9508 (N_9508,N_1966,N_2801);
and U9509 (N_9509,N_1830,N_2245);
xnor U9510 (N_9510,N_3078,N_3915);
xor U9511 (N_9511,N_4071,N_1229);
xnor U9512 (N_9512,N_2481,N_2729);
nand U9513 (N_9513,N_1326,N_1676);
xor U9514 (N_9514,N_1544,N_4794);
or U9515 (N_9515,N_2812,N_194);
xnor U9516 (N_9516,N_1240,N_4524);
nand U9517 (N_9517,N_712,N_1764);
xnor U9518 (N_9518,N_1596,N_2230);
nor U9519 (N_9519,N_1080,N_3001);
and U9520 (N_9520,N_451,N_2590);
and U9521 (N_9521,N_4927,N_603);
nor U9522 (N_9522,N_397,N_854);
xor U9523 (N_9523,N_460,N_2819);
nor U9524 (N_9524,N_2084,N_325);
nor U9525 (N_9525,N_597,N_1088);
and U9526 (N_9526,N_4463,N_1000);
and U9527 (N_9527,N_3875,N_3142);
xnor U9528 (N_9528,N_3652,N_766);
nor U9529 (N_9529,N_3108,N_2619);
nand U9530 (N_9530,N_3649,N_3535);
nand U9531 (N_9531,N_3877,N_582);
xor U9532 (N_9532,N_3979,N_2367);
nand U9533 (N_9533,N_3622,N_1731);
and U9534 (N_9534,N_4924,N_2726);
nand U9535 (N_9535,N_1324,N_3312);
and U9536 (N_9536,N_3327,N_3723);
xnor U9537 (N_9537,N_2336,N_4396);
and U9538 (N_9538,N_809,N_4122);
nand U9539 (N_9539,N_3258,N_301);
nor U9540 (N_9540,N_30,N_2004);
and U9541 (N_9541,N_1711,N_2122);
nor U9542 (N_9542,N_2427,N_1051);
nor U9543 (N_9543,N_342,N_2084);
nand U9544 (N_9544,N_548,N_1474);
or U9545 (N_9545,N_2317,N_3571);
or U9546 (N_9546,N_1209,N_4431);
nand U9547 (N_9547,N_443,N_1863);
and U9548 (N_9548,N_2791,N_1703);
nor U9549 (N_9549,N_3786,N_784);
nor U9550 (N_9550,N_3361,N_1764);
nand U9551 (N_9551,N_3122,N_4323);
and U9552 (N_9552,N_1374,N_4760);
and U9553 (N_9553,N_722,N_1976);
nor U9554 (N_9554,N_100,N_3797);
nand U9555 (N_9555,N_3367,N_3964);
nand U9556 (N_9556,N_2872,N_1201);
and U9557 (N_9557,N_4941,N_2137);
or U9558 (N_9558,N_2155,N_2034);
nor U9559 (N_9559,N_2493,N_1943);
nor U9560 (N_9560,N_464,N_4712);
and U9561 (N_9561,N_1967,N_870);
or U9562 (N_9562,N_4848,N_2189);
nand U9563 (N_9563,N_1780,N_2241);
xor U9564 (N_9564,N_2505,N_182);
xnor U9565 (N_9565,N_1050,N_4097);
and U9566 (N_9566,N_78,N_4276);
xnor U9567 (N_9567,N_1050,N_2121);
and U9568 (N_9568,N_754,N_4432);
nor U9569 (N_9569,N_723,N_2448);
or U9570 (N_9570,N_3711,N_3476);
or U9571 (N_9571,N_2776,N_1911);
xor U9572 (N_9572,N_3758,N_2651);
nand U9573 (N_9573,N_3736,N_3002);
nor U9574 (N_9574,N_3454,N_41);
nand U9575 (N_9575,N_3681,N_377);
nor U9576 (N_9576,N_1023,N_2369);
nand U9577 (N_9577,N_2511,N_1541);
nand U9578 (N_9578,N_814,N_1469);
xor U9579 (N_9579,N_3381,N_817);
nand U9580 (N_9580,N_2500,N_1421);
nor U9581 (N_9581,N_2556,N_2103);
and U9582 (N_9582,N_1285,N_4240);
xnor U9583 (N_9583,N_1587,N_2953);
nand U9584 (N_9584,N_4224,N_736);
or U9585 (N_9585,N_3286,N_2184);
xor U9586 (N_9586,N_2966,N_614);
nand U9587 (N_9587,N_3550,N_1343);
xor U9588 (N_9588,N_4500,N_978);
xnor U9589 (N_9589,N_3773,N_2199);
or U9590 (N_9590,N_4094,N_4036);
xnor U9591 (N_9591,N_2308,N_534);
and U9592 (N_9592,N_2874,N_4894);
or U9593 (N_9593,N_2356,N_4118);
and U9594 (N_9594,N_2913,N_4115);
xor U9595 (N_9595,N_4624,N_1538);
nand U9596 (N_9596,N_3263,N_2823);
nand U9597 (N_9597,N_2326,N_983);
nand U9598 (N_9598,N_1519,N_4361);
xor U9599 (N_9599,N_4960,N_2572);
nand U9600 (N_9600,N_2502,N_628);
and U9601 (N_9601,N_3540,N_3867);
nand U9602 (N_9602,N_3564,N_1152);
or U9603 (N_9603,N_216,N_3996);
and U9604 (N_9604,N_2464,N_2131);
nor U9605 (N_9605,N_3835,N_2081);
xor U9606 (N_9606,N_3384,N_3180);
xnor U9607 (N_9607,N_113,N_2928);
xnor U9608 (N_9608,N_3070,N_3580);
xnor U9609 (N_9609,N_735,N_4146);
xnor U9610 (N_9610,N_4871,N_3972);
xnor U9611 (N_9611,N_1474,N_3157);
nor U9612 (N_9612,N_3814,N_4520);
and U9613 (N_9613,N_4246,N_2384);
or U9614 (N_9614,N_381,N_1248);
nand U9615 (N_9615,N_643,N_2588);
or U9616 (N_9616,N_3411,N_8);
nand U9617 (N_9617,N_3004,N_6);
nor U9618 (N_9618,N_4027,N_107);
nand U9619 (N_9619,N_10,N_303);
nor U9620 (N_9620,N_2845,N_1053);
xor U9621 (N_9621,N_1084,N_864);
or U9622 (N_9622,N_1372,N_2452);
and U9623 (N_9623,N_2139,N_2468);
nor U9624 (N_9624,N_1869,N_3073);
or U9625 (N_9625,N_2560,N_1288);
xnor U9626 (N_9626,N_4300,N_194);
and U9627 (N_9627,N_1649,N_1080);
nor U9628 (N_9628,N_3459,N_2945);
nand U9629 (N_9629,N_714,N_2546);
xnor U9630 (N_9630,N_4851,N_2177);
nor U9631 (N_9631,N_154,N_3785);
nand U9632 (N_9632,N_121,N_2381);
or U9633 (N_9633,N_4197,N_1658);
nor U9634 (N_9634,N_1946,N_2612);
nand U9635 (N_9635,N_3634,N_3484);
nand U9636 (N_9636,N_195,N_290);
xnor U9637 (N_9637,N_1868,N_3966);
and U9638 (N_9638,N_223,N_4548);
nand U9639 (N_9639,N_2091,N_80);
xor U9640 (N_9640,N_939,N_544);
or U9641 (N_9641,N_1688,N_4358);
nand U9642 (N_9642,N_4350,N_4214);
nor U9643 (N_9643,N_4977,N_1170);
nor U9644 (N_9644,N_1124,N_3446);
and U9645 (N_9645,N_3947,N_3133);
nand U9646 (N_9646,N_3279,N_3142);
nor U9647 (N_9647,N_1819,N_4002);
nor U9648 (N_9648,N_2995,N_4140);
or U9649 (N_9649,N_4058,N_4352);
and U9650 (N_9650,N_190,N_4461);
nand U9651 (N_9651,N_4282,N_3687);
or U9652 (N_9652,N_2488,N_1182);
xnor U9653 (N_9653,N_2006,N_4210);
nor U9654 (N_9654,N_92,N_1548);
or U9655 (N_9655,N_4176,N_746);
nor U9656 (N_9656,N_3833,N_3735);
nand U9657 (N_9657,N_2060,N_4611);
and U9658 (N_9658,N_1613,N_308);
and U9659 (N_9659,N_4772,N_2349);
or U9660 (N_9660,N_4089,N_2853);
and U9661 (N_9661,N_646,N_1162);
xnor U9662 (N_9662,N_1224,N_1977);
xnor U9663 (N_9663,N_1989,N_3480);
xor U9664 (N_9664,N_3443,N_233);
xor U9665 (N_9665,N_3017,N_123);
xnor U9666 (N_9666,N_1190,N_95);
and U9667 (N_9667,N_1029,N_462);
and U9668 (N_9668,N_586,N_4830);
xnor U9669 (N_9669,N_3956,N_790);
and U9670 (N_9670,N_3653,N_4693);
or U9671 (N_9671,N_1638,N_1510);
xor U9672 (N_9672,N_4103,N_2936);
and U9673 (N_9673,N_4283,N_376);
and U9674 (N_9674,N_424,N_30);
xor U9675 (N_9675,N_2081,N_1508);
and U9676 (N_9676,N_208,N_4147);
xor U9677 (N_9677,N_1778,N_3747);
xor U9678 (N_9678,N_2452,N_4854);
nor U9679 (N_9679,N_2815,N_3368);
or U9680 (N_9680,N_916,N_1130);
xor U9681 (N_9681,N_4633,N_2770);
or U9682 (N_9682,N_2347,N_1087);
or U9683 (N_9683,N_2620,N_2919);
nor U9684 (N_9684,N_3011,N_816);
nor U9685 (N_9685,N_69,N_588);
nor U9686 (N_9686,N_1262,N_2179);
nor U9687 (N_9687,N_4095,N_3842);
or U9688 (N_9688,N_1970,N_3408);
nand U9689 (N_9689,N_3032,N_2770);
xor U9690 (N_9690,N_4363,N_1663);
xnor U9691 (N_9691,N_1156,N_2465);
nor U9692 (N_9692,N_3340,N_1565);
and U9693 (N_9693,N_1416,N_1543);
nand U9694 (N_9694,N_4091,N_4909);
nand U9695 (N_9695,N_3767,N_2622);
nand U9696 (N_9696,N_2270,N_2446);
nand U9697 (N_9697,N_2458,N_4149);
or U9698 (N_9698,N_4957,N_2636);
and U9699 (N_9699,N_4547,N_217);
and U9700 (N_9700,N_3217,N_333);
and U9701 (N_9701,N_3501,N_3667);
nor U9702 (N_9702,N_4594,N_1309);
and U9703 (N_9703,N_4547,N_4136);
xnor U9704 (N_9704,N_1388,N_1830);
and U9705 (N_9705,N_4481,N_626);
or U9706 (N_9706,N_1318,N_2333);
nor U9707 (N_9707,N_1197,N_945);
and U9708 (N_9708,N_1268,N_754);
xor U9709 (N_9709,N_3594,N_773);
or U9710 (N_9710,N_4252,N_2373);
nand U9711 (N_9711,N_3790,N_967);
nor U9712 (N_9712,N_3997,N_220);
nand U9713 (N_9713,N_3269,N_515);
or U9714 (N_9714,N_2228,N_280);
and U9715 (N_9715,N_37,N_2378);
and U9716 (N_9716,N_3463,N_1976);
and U9717 (N_9717,N_1535,N_3990);
nor U9718 (N_9718,N_4894,N_3469);
or U9719 (N_9719,N_3935,N_4004);
nand U9720 (N_9720,N_3289,N_2667);
xnor U9721 (N_9721,N_1417,N_274);
xor U9722 (N_9722,N_4545,N_3094);
or U9723 (N_9723,N_1646,N_2566);
nor U9724 (N_9724,N_2352,N_2606);
xor U9725 (N_9725,N_598,N_4585);
nor U9726 (N_9726,N_1897,N_276);
nand U9727 (N_9727,N_2525,N_1550);
or U9728 (N_9728,N_3588,N_248);
or U9729 (N_9729,N_4051,N_3131);
nor U9730 (N_9730,N_4673,N_2007);
xor U9731 (N_9731,N_2304,N_3378);
nor U9732 (N_9732,N_1078,N_663);
or U9733 (N_9733,N_2270,N_231);
nor U9734 (N_9734,N_4285,N_3824);
nand U9735 (N_9735,N_2940,N_268);
and U9736 (N_9736,N_1896,N_4776);
and U9737 (N_9737,N_3696,N_1628);
and U9738 (N_9738,N_1583,N_1820);
nor U9739 (N_9739,N_2178,N_2886);
and U9740 (N_9740,N_4882,N_1587);
xnor U9741 (N_9741,N_1723,N_2321);
nand U9742 (N_9742,N_993,N_2691);
and U9743 (N_9743,N_2109,N_306);
nor U9744 (N_9744,N_5,N_4270);
and U9745 (N_9745,N_3079,N_3013);
nand U9746 (N_9746,N_1873,N_4250);
nor U9747 (N_9747,N_4061,N_2903);
nor U9748 (N_9748,N_4263,N_3848);
nand U9749 (N_9749,N_382,N_2715);
xor U9750 (N_9750,N_4330,N_1381);
and U9751 (N_9751,N_4689,N_1828);
nand U9752 (N_9752,N_1758,N_4704);
or U9753 (N_9753,N_1398,N_4833);
nor U9754 (N_9754,N_4806,N_4537);
or U9755 (N_9755,N_4701,N_3878);
xor U9756 (N_9756,N_3833,N_1860);
nand U9757 (N_9757,N_4357,N_3628);
and U9758 (N_9758,N_1227,N_3623);
nor U9759 (N_9759,N_2433,N_4425);
and U9760 (N_9760,N_1581,N_395);
and U9761 (N_9761,N_4527,N_1675);
xor U9762 (N_9762,N_4089,N_3691);
nand U9763 (N_9763,N_1723,N_1549);
and U9764 (N_9764,N_4943,N_2870);
xor U9765 (N_9765,N_3044,N_3509);
nor U9766 (N_9766,N_3131,N_4407);
nand U9767 (N_9767,N_4331,N_3582);
and U9768 (N_9768,N_3827,N_4884);
and U9769 (N_9769,N_394,N_1117);
and U9770 (N_9770,N_4094,N_4966);
xor U9771 (N_9771,N_531,N_2797);
xor U9772 (N_9772,N_3290,N_865);
nor U9773 (N_9773,N_2755,N_2095);
and U9774 (N_9774,N_3834,N_1964);
xor U9775 (N_9775,N_2738,N_3536);
xor U9776 (N_9776,N_609,N_2273);
and U9777 (N_9777,N_2812,N_2474);
or U9778 (N_9778,N_234,N_1619);
nand U9779 (N_9779,N_2281,N_675);
or U9780 (N_9780,N_851,N_4824);
or U9781 (N_9781,N_1150,N_3642);
xnor U9782 (N_9782,N_2569,N_2142);
nand U9783 (N_9783,N_1081,N_3020);
nor U9784 (N_9784,N_1800,N_2734);
nand U9785 (N_9785,N_280,N_148);
nor U9786 (N_9786,N_3754,N_3056);
or U9787 (N_9787,N_4987,N_90);
and U9788 (N_9788,N_4642,N_1536);
or U9789 (N_9789,N_878,N_2381);
or U9790 (N_9790,N_3389,N_232);
nand U9791 (N_9791,N_2888,N_2290);
and U9792 (N_9792,N_2230,N_3159);
xnor U9793 (N_9793,N_2733,N_3710);
nand U9794 (N_9794,N_2633,N_2210);
or U9795 (N_9795,N_3719,N_3371);
nand U9796 (N_9796,N_4690,N_3087);
xnor U9797 (N_9797,N_1538,N_2652);
nand U9798 (N_9798,N_221,N_2595);
xnor U9799 (N_9799,N_4395,N_2535);
nand U9800 (N_9800,N_805,N_2542);
nor U9801 (N_9801,N_4609,N_308);
xnor U9802 (N_9802,N_4305,N_3426);
xor U9803 (N_9803,N_4184,N_759);
or U9804 (N_9804,N_2846,N_887);
nand U9805 (N_9805,N_2714,N_4456);
nor U9806 (N_9806,N_315,N_4032);
or U9807 (N_9807,N_2894,N_2621);
or U9808 (N_9808,N_1013,N_1618);
nand U9809 (N_9809,N_1233,N_4373);
xnor U9810 (N_9810,N_2119,N_4422);
nand U9811 (N_9811,N_541,N_1312);
and U9812 (N_9812,N_3111,N_2052);
nand U9813 (N_9813,N_1476,N_1847);
or U9814 (N_9814,N_1973,N_1340);
and U9815 (N_9815,N_645,N_2608);
or U9816 (N_9816,N_3617,N_713);
and U9817 (N_9817,N_2932,N_293);
or U9818 (N_9818,N_728,N_4032);
nand U9819 (N_9819,N_1466,N_4269);
and U9820 (N_9820,N_2724,N_1062);
or U9821 (N_9821,N_20,N_808);
and U9822 (N_9822,N_201,N_3239);
or U9823 (N_9823,N_597,N_833);
nand U9824 (N_9824,N_4843,N_4361);
and U9825 (N_9825,N_4756,N_2789);
xnor U9826 (N_9826,N_1902,N_4151);
nand U9827 (N_9827,N_118,N_4209);
and U9828 (N_9828,N_311,N_2349);
nand U9829 (N_9829,N_1313,N_3354);
or U9830 (N_9830,N_2646,N_62);
or U9831 (N_9831,N_4783,N_3582);
xor U9832 (N_9832,N_1803,N_1776);
nand U9833 (N_9833,N_3204,N_163);
and U9834 (N_9834,N_3812,N_2009);
and U9835 (N_9835,N_276,N_3621);
nand U9836 (N_9836,N_1824,N_4186);
or U9837 (N_9837,N_4122,N_2112);
nand U9838 (N_9838,N_1377,N_4701);
xor U9839 (N_9839,N_2440,N_3603);
nor U9840 (N_9840,N_964,N_1752);
nand U9841 (N_9841,N_4276,N_3068);
and U9842 (N_9842,N_1632,N_4096);
nor U9843 (N_9843,N_2570,N_4123);
xor U9844 (N_9844,N_4651,N_3312);
nand U9845 (N_9845,N_535,N_3622);
and U9846 (N_9846,N_1699,N_1489);
nor U9847 (N_9847,N_2593,N_590);
nand U9848 (N_9848,N_2308,N_2292);
xor U9849 (N_9849,N_4402,N_2886);
nand U9850 (N_9850,N_3530,N_1679);
nor U9851 (N_9851,N_825,N_4640);
and U9852 (N_9852,N_2228,N_3382);
nand U9853 (N_9853,N_2513,N_1404);
nand U9854 (N_9854,N_353,N_4721);
and U9855 (N_9855,N_1764,N_2736);
or U9856 (N_9856,N_4321,N_3150);
nand U9857 (N_9857,N_727,N_771);
nand U9858 (N_9858,N_1230,N_3273);
or U9859 (N_9859,N_2655,N_2926);
or U9860 (N_9860,N_2463,N_3480);
nor U9861 (N_9861,N_372,N_1959);
or U9862 (N_9862,N_4936,N_2686);
or U9863 (N_9863,N_4681,N_2450);
and U9864 (N_9864,N_4686,N_3432);
or U9865 (N_9865,N_2120,N_3190);
nand U9866 (N_9866,N_187,N_875);
xor U9867 (N_9867,N_4685,N_3089);
xor U9868 (N_9868,N_1305,N_4814);
and U9869 (N_9869,N_887,N_1315);
and U9870 (N_9870,N_1210,N_4528);
or U9871 (N_9871,N_2704,N_4693);
nor U9872 (N_9872,N_338,N_826);
nor U9873 (N_9873,N_3344,N_4746);
and U9874 (N_9874,N_1770,N_379);
xor U9875 (N_9875,N_1229,N_3294);
and U9876 (N_9876,N_953,N_4797);
nor U9877 (N_9877,N_4299,N_2791);
nor U9878 (N_9878,N_1349,N_3179);
nand U9879 (N_9879,N_4059,N_3746);
nand U9880 (N_9880,N_738,N_1626);
or U9881 (N_9881,N_4547,N_2418);
nand U9882 (N_9882,N_3890,N_698);
and U9883 (N_9883,N_3241,N_1606);
or U9884 (N_9884,N_3074,N_971);
and U9885 (N_9885,N_723,N_1721);
nand U9886 (N_9886,N_4529,N_1903);
or U9887 (N_9887,N_1069,N_3661);
nor U9888 (N_9888,N_2450,N_253);
nand U9889 (N_9889,N_4910,N_4539);
nand U9890 (N_9890,N_184,N_4509);
or U9891 (N_9891,N_3499,N_215);
and U9892 (N_9892,N_3333,N_1137);
xor U9893 (N_9893,N_1955,N_1939);
nand U9894 (N_9894,N_1641,N_3490);
nand U9895 (N_9895,N_3939,N_849);
nand U9896 (N_9896,N_1016,N_2890);
or U9897 (N_9897,N_3860,N_4751);
xnor U9898 (N_9898,N_833,N_729);
nor U9899 (N_9899,N_4534,N_3862);
or U9900 (N_9900,N_3238,N_2908);
and U9901 (N_9901,N_1730,N_3131);
nand U9902 (N_9902,N_1816,N_1739);
or U9903 (N_9903,N_2551,N_4215);
nor U9904 (N_9904,N_696,N_736);
and U9905 (N_9905,N_206,N_2082);
and U9906 (N_9906,N_2387,N_2618);
or U9907 (N_9907,N_3767,N_3501);
nand U9908 (N_9908,N_2312,N_3055);
and U9909 (N_9909,N_243,N_1086);
nand U9910 (N_9910,N_638,N_2157);
xor U9911 (N_9911,N_1777,N_4685);
and U9912 (N_9912,N_94,N_790);
and U9913 (N_9913,N_2077,N_975);
or U9914 (N_9914,N_1080,N_1112);
or U9915 (N_9915,N_2621,N_1948);
nor U9916 (N_9916,N_2954,N_617);
and U9917 (N_9917,N_2139,N_1);
and U9918 (N_9918,N_4564,N_3509);
nand U9919 (N_9919,N_1974,N_2246);
or U9920 (N_9920,N_1075,N_4751);
xnor U9921 (N_9921,N_1998,N_1765);
nor U9922 (N_9922,N_3606,N_3190);
xor U9923 (N_9923,N_4710,N_643);
or U9924 (N_9924,N_3948,N_2629);
nor U9925 (N_9925,N_3142,N_2786);
xnor U9926 (N_9926,N_1124,N_1908);
nor U9927 (N_9927,N_645,N_1376);
xnor U9928 (N_9928,N_3120,N_1843);
nand U9929 (N_9929,N_4920,N_3843);
and U9930 (N_9930,N_1685,N_3910);
and U9931 (N_9931,N_3231,N_2062);
nor U9932 (N_9932,N_3665,N_3734);
nand U9933 (N_9933,N_3657,N_283);
and U9934 (N_9934,N_4539,N_2014);
or U9935 (N_9935,N_1179,N_3735);
nand U9936 (N_9936,N_1522,N_4114);
nand U9937 (N_9937,N_2323,N_1576);
or U9938 (N_9938,N_2036,N_3925);
and U9939 (N_9939,N_1977,N_4553);
nor U9940 (N_9940,N_3871,N_3213);
and U9941 (N_9941,N_4121,N_3983);
xor U9942 (N_9942,N_639,N_3127);
nand U9943 (N_9943,N_4811,N_3044);
xor U9944 (N_9944,N_1062,N_2182);
nand U9945 (N_9945,N_12,N_1034);
or U9946 (N_9946,N_1693,N_2389);
xor U9947 (N_9947,N_4919,N_2296);
and U9948 (N_9948,N_1309,N_2648);
nor U9949 (N_9949,N_4041,N_3263);
nor U9950 (N_9950,N_1138,N_814);
nand U9951 (N_9951,N_4619,N_4442);
nor U9952 (N_9952,N_2228,N_4290);
nor U9953 (N_9953,N_1516,N_2118);
nand U9954 (N_9954,N_425,N_185);
and U9955 (N_9955,N_3037,N_4455);
and U9956 (N_9956,N_3739,N_2434);
nor U9957 (N_9957,N_703,N_4434);
nand U9958 (N_9958,N_2833,N_1101);
nand U9959 (N_9959,N_1678,N_4508);
nor U9960 (N_9960,N_1537,N_3636);
nor U9961 (N_9961,N_3351,N_33);
and U9962 (N_9962,N_3467,N_2935);
xor U9963 (N_9963,N_2478,N_3607);
or U9964 (N_9964,N_4733,N_1643);
or U9965 (N_9965,N_2561,N_1994);
nor U9966 (N_9966,N_1005,N_4376);
xor U9967 (N_9967,N_4501,N_2863);
nand U9968 (N_9968,N_1946,N_276);
nor U9969 (N_9969,N_2564,N_1548);
or U9970 (N_9970,N_3051,N_2370);
and U9971 (N_9971,N_2615,N_90);
nand U9972 (N_9972,N_418,N_3213);
xnor U9973 (N_9973,N_922,N_253);
nor U9974 (N_9974,N_2231,N_621);
xor U9975 (N_9975,N_1381,N_1286);
nor U9976 (N_9976,N_3662,N_1634);
nor U9977 (N_9977,N_40,N_4239);
nor U9978 (N_9978,N_4950,N_4082);
or U9979 (N_9979,N_2671,N_3235);
and U9980 (N_9980,N_2255,N_3258);
and U9981 (N_9981,N_3087,N_2072);
and U9982 (N_9982,N_1536,N_3496);
nor U9983 (N_9983,N_823,N_1894);
and U9984 (N_9984,N_1,N_1563);
xor U9985 (N_9985,N_3670,N_3673);
nand U9986 (N_9986,N_1596,N_3020);
nand U9987 (N_9987,N_2753,N_557);
xor U9988 (N_9988,N_857,N_4028);
nor U9989 (N_9989,N_227,N_3232);
nor U9990 (N_9990,N_2646,N_2388);
or U9991 (N_9991,N_267,N_1643);
or U9992 (N_9992,N_3261,N_4779);
nand U9993 (N_9993,N_2932,N_1689);
xnor U9994 (N_9994,N_3224,N_519);
or U9995 (N_9995,N_3488,N_2166);
or U9996 (N_9996,N_2692,N_4193);
or U9997 (N_9997,N_4460,N_544);
or U9998 (N_9998,N_1219,N_926);
or U9999 (N_9999,N_2968,N_993);
nand U10000 (N_10000,N_5241,N_6194);
nor U10001 (N_10001,N_5035,N_8667);
nand U10002 (N_10002,N_9807,N_9461);
nor U10003 (N_10003,N_9874,N_8665);
or U10004 (N_10004,N_6973,N_7794);
nor U10005 (N_10005,N_5583,N_6570);
xor U10006 (N_10006,N_6774,N_8773);
xor U10007 (N_10007,N_6036,N_8711);
or U10008 (N_10008,N_8053,N_5744);
nand U10009 (N_10009,N_8004,N_8298);
or U10010 (N_10010,N_6168,N_5254);
nor U10011 (N_10011,N_5234,N_6849);
or U10012 (N_10012,N_7319,N_7363);
nand U10013 (N_10013,N_9720,N_6881);
or U10014 (N_10014,N_6381,N_9855);
nand U10015 (N_10015,N_5835,N_8978);
nor U10016 (N_10016,N_7809,N_6580);
xor U10017 (N_10017,N_5888,N_5502);
and U10018 (N_10018,N_8821,N_6903);
nor U10019 (N_10019,N_7665,N_5595);
or U10020 (N_10020,N_6992,N_8726);
xor U10021 (N_10021,N_5388,N_9484);
nor U10022 (N_10022,N_5738,N_6968);
xor U10023 (N_10023,N_7923,N_5478);
xnor U10024 (N_10024,N_6200,N_9933);
xnor U10025 (N_10025,N_7943,N_9574);
or U10026 (N_10026,N_5173,N_7273);
xor U10027 (N_10027,N_8729,N_6598);
nor U10028 (N_10028,N_7237,N_8620);
xnor U10029 (N_10029,N_8939,N_9288);
nor U10030 (N_10030,N_5473,N_6606);
and U10031 (N_10031,N_8799,N_8803);
nand U10032 (N_10032,N_9932,N_7783);
xnor U10033 (N_10033,N_7953,N_5812);
and U10034 (N_10034,N_5218,N_7342);
xor U10035 (N_10035,N_8231,N_9451);
nor U10036 (N_10036,N_8548,N_9169);
xnor U10037 (N_10037,N_8842,N_8109);
xor U10038 (N_10038,N_7045,N_8964);
nand U10039 (N_10039,N_5316,N_7598);
and U10040 (N_10040,N_5811,N_5760);
or U10041 (N_10041,N_5135,N_6436);
or U10042 (N_10042,N_6408,N_9246);
and U10043 (N_10043,N_7121,N_9093);
xnor U10044 (N_10044,N_8673,N_7846);
or U10045 (N_10045,N_9852,N_7079);
or U10046 (N_10046,N_5436,N_5825);
nor U10047 (N_10047,N_8341,N_5906);
and U10048 (N_10048,N_6496,N_7546);
nand U10049 (N_10049,N_8283,N_7714);
and U10050 (N_10050,N_7967,N_7865);
nand U10051 (N_10051,N_5965,N_5985);
or U10052 (N_10052,N_9604,N_8865);
and U10053 (N_10053,N_9543,N_6063);
nor U10054 (N_10054,N_7299,N_7084);
or U10055 (N_10055,N_5975,N_7352);
or U10056 (N_10056,N_7455,N_9437);
or U10057 (N_10057,N_6893,N_8500);
or U10058 (N_10058,N_6607,N_9673);
and U10059 (N_10059,N_5109,N_9866);
or U10060 (N_10060,N_8443,N_6080);
xnor U10061 (N_10061,N_9469,N_5930);
nor U10062 (N_10062,N_8621,N_6747);
or U10063 (N_10063,N_9072,N_7025);
nor U10064 (N_10064,N_9555,N_6501);
or U10065 (N_10065,N_7011,N_9234);
nor U10066 (N_10066,N_5924,N_8728);
xnor U10067 (N_10067,N_7097,N_9167);
or U10068 (N_10068,N_7589,N_7344);
and U10069 (N_10069,N_5293,N_9754);
xnor U10070 (N_10070,N_9697,N_5966);
xnor U10071 (N_10071,N_6843,N_6572);
nand U10072 (N_10072,N_9609,N_9044);
nand U10073 (N_10073,N_9515,N_9032);
nor U10074 (N_10074,N_7381,N_5394);
nor U10075 (N_10075,N_6712,N_6478);
nand U10076 (N_10076,N_6970,N_8202);
nor U10077 (N_10077,N_6779,N_6584);
and U10078 (N_10078,N_9009,N_6518);
or U10079 (N_10079,N_7805,N_6096);
nor U10080 (N_10080,N_8382,N_5377);
nor U10081 (N_10081,N_6845,N_8346);
or U10082 (N_10082,N_5743,N_9858);
xor U10083 (N_10083,N_8181,N_8407);
or U10084 (N_10084,N_7904,N_8596);
nor U10085 (N_10085,N_9337,N_6961);
nand U10086 (N_10086,N_5069,N_9711);
or U10087 (N_10087,N_9019,N_7631);
and U10088 (N_10088,N_7807,N_5984);
or U10089 (N_10089,N_8076,N_6829);
xor U10090 (N_10090,N_6621,N_6998);
and U10091 (N_10091,N_7075,N_8313);
nand U10092 (N_10092,N_7855,N_9987);
and U10093 (N_10093,N_7551,N_8126);
xor U10094 (N_10094,N_8863,N_6180);
nand U10095 (N_10095,N_6497,N_5442);
xor U10096 (N_10096,N_7107,N_8826);
or U10097 (N_10097,N_8215,N_9064);
nor U10098 (N_10098,N_9343,N_9323);
nand U10099 (N_10099,N_5079,N_8314);
nand U10100 (N_10100,N_7530,N_8132);
nor U10101 (N_10101,N_8217,N_7788);
xnor U10102 (N_10102,N_7415,N_6474);
or U10103 (N_10103,N_7061,N_5193);
xnor U10104 (N_10104,N_5149,N_7478);
xor U10105 (N_10105,N_9204,N_7833);
nor U10106 (N_10106,N_6615,N_8575);
or U10107 (N_10107,N_7937,N_9724);
and U10108 (N_10108,N_6597,N_6406);
xnor U10109 (N_10109,N_8063,N_7161);
and U10110 (N_10110,N_9782,N_6816);
xnor U10111 (N_10111,N_5689,N_9519);
and U10112 (N_10112,N_5104,N_6334);
nand U10113 (N_10113,N_5127,N_5505);
nor U10114 (N_10114,N_7719,N_5251);
and U10115 (N_10115,N_5567,N_9809);
or U10116 (N_10116,N_6661,N_5164);
nand U10117 (N_10117,N_9528,N_9972);
xnor U10118 (N_10118,N_7938,N_6942);
or U10119 (N_10119,N_9974,N_6098);
nor U10120 (N_10120,N_6704,N_8157);
and U10121 (N_10121,N_9271,N_6311);
nor U10122 (N_10122,N_8660,N_7220);
nor U10123 (N_10123,N_9266,N_5384);
nor U10124 (N_10124,N_7502,N_5768);
nor U10125 (N_10125,N_9795,N_6703);
xor U10126 (N_10126,N_9481,N_5045);
nor U10127 (N_10127,N_7090,N_6950);
nand U10128 (N_10128,N_6795,N_7042);
nand U10129 (N_10129,N_8183,N_8151);
nor U10130 (N_10130,N_7667,N_6509);
xnor U10131 (N_10131,N_5031,N_7223);
and U10132 (N_10132,N_5716,N_9516);
nor U10133 (N_10133,N_7586,N_5510);
or U10134 (N_10134,N_7925,N_8748);
nor U10135 (N_10135,N_8207,N_7262);
nor U10136 (N_10136,N_6059,N_7158);
and U10137 (N_10137,N_9839,N_9835);
or U10138 (N_10138,N_6908,N_7173);
and U10139 (N_10139,N_8583,N_6548);
xnor U10140 (N_10140,N_6457,N_9701);
and U10141 (N_10141,N_9074,N_7741);
nand U10142 (N_10142,N_5654,N_7747);
and U10143 (N_10143,N_6367,N_9947);
xnor U10144 (N_10144,N_8384,N_8051);
and U10145 (N_10145,N_5209,N_5358);
nand U10146 (N_10146,N_7983,N_8211);
xor U10147 (N_10147,N_9853,N_7632);
nor U10148 (N_10148,N_9154,N_7677);
or U10149 (N_10149,N_6246,N_8391);
and U10150 (N_10150,N_6111,N_8242);
and U10151 (N_10151,N_5195,N_7847);
nor U10152 (N_10152,N_5183,N_6365);
nor U10153 (N_10153,N_9361,N_9401);
nor U10154 (N_10154,N_6789,N_7178);
xor U10155 (N_10155,N_8682,N_7543);
and U10156 (N_10156,N_9901,N_5468);
nor U10157 (N_10157,N_8533,N_8559);
xnor U10158 (N_10158,N_9063,N_6351);
nor U10159 (N_10159,N_7961,N_9182);
or U10160 (N_10160,N_7964,N_9746);
xor U10161 (N_10161,N_7170,N_8985);
and U10162 (N_10162,N_5685,N_9812);
nand U10163 (N_10163,N_5002,N_8037);
nor U10164 (N_10164,N_8235,N_9924);
and U10165 (N_10165,N_9836,N_9941);
nor U10166 (N_10166,N_7587,N_6181);
and U10167 (N_10167,N_8174,N_8072);
nor U10168 (N_10168,N_9233,N_8493);
xnor U10169 (N_10169,N_5423,N_6166);
nor U10170 (N_10170,N_6234,N_7601);
or U10171 (N_10171,N_7293,N_9070);
nand U10172 (N_10172,N_7375,N_6725);
xnor U10173 (N_10173,N_8928,N_7004);
nand U10174 (N_10174,N_9614,N_8038);
or U10175 (N_10175,N_6041,N_7447);
nor U10176 (N_10176,N_9375,N_8034);
xor U10177 (N_10177,N_7310,N_7804);
and U10178 (N_10178,N_7129,N_8988);
and U10179 (N_10179,N_6241,N_9573);
nand U10180 (N_10180,N_9774,N_6065);
or U10181 (N_10181,N_9315,N_6949);
nand U10182 (N_10182,N_9143,N_5203);
or U10183 (N_10183,N_5319,N_7898);
nand U10184 (N_10184,N_5256,N_6456);
nor U10185 (N_10185,N_9317,N_7909);
and U10186 (N_10186,N_7395,N_8400);
and U10187 (N_10187,N_8325,N_8497);
nand U10188 (N_10188,N_9970,N_5632);
or U10189 (N_10189,N_5162,N_8071);
nor U10190 (N_10190,N_6664,N_9050);
nor U10191 (N_10191,N_6730,N_5454);
or U10192 (N_10192,N_7990,N_6554);
nand U10193 (N_10193,N_5640,N_5585);
nor U10194 (N_10194,N_5681,N_6506);
xor U10195 (N_10195,N_7890,N_5868);
xnor U10196 (N_10196,N_5770,N_6197);
or U10197 (N_10197,N_5917,N_6448);
and U10198 (N_10198,N_5092,N_9714);
and U10199 (N_10199,N_5013,N_8653);
and U10200 (N_10200,N_6855,N_5165);
nand U10201 (N_10201,N_5114,N_9440);
and U10202 (N_10202,N_8809,N_8286);
or U10203 (N_10203,N_5662,N_7817);
nor U10204 (N_10204,N_6768,N_9973);
xor U10205 (N_10205,N_6438,N_8685);
xor U10206 (N_10206,N_6109,N_7740);
xor U10207 (N_10207,N_5573,N_7933);
or U10208 (N_10208,N_7142,N_5895);
or U10209 (N_10209,N_6411,N_5834);
nor U10210 (N_10210,N_8377,N_6485);
and U10211 (N_10211,N_5145,N_9572);
xnor U10212 (N_10212,N_9291,N_5056);
xnor U10213 (N_10213,N_5352,N_5605);
nor U10214 (N_10214,N_7032,N_6451);
or U10215 (N_10215,N_9173,N_6216);
nor U10216 (N_10216,N_6940,N_5467);
xnor U10217 (N_10217,N_9520,N_9388);
and U10218 (N_10218,N_6838,N_9163);
nand U10219 (N_10219,N_5444,N_9956);
or U10220 (N_10220,N_9518,N_7210);
nor U10221 (N_10221,N_5093,N_6978);
nor U10222 (N_10222,N_8791,N_8267);
and U10223 (N_10223,N_7263,N_6618);
or U10224 (N_10224,N_8851,N_9877);
xor U10225 (N_10225,N_8090,N_8700);
and U10226 (N_10226,N_5623,N_5350);
or U10227 (N_10227,N_5597,N_6188);
or U10228 (N_10228,N_9321,N_6716);
and U10229 (N_10229,N_8073,N_5022);
xor U10230 (N_10230,N_9022,N_6648);
xnor U10231 (N_10231,N_9152,N_9927);
nand U10232 (N_10232,N_5615,N_7491);
nor U10233 (N_10233,N_8044,N_7257);
nand U10234 (N_10234,N_5919,N_9067);
and U10235 (N_10235,N_8477,N_5530);
nand U10236 (N_10236,N_9674,N_8837);
nand U10237 (N_10237,N_8055,N_8420);
nand U10238 (N_10238,N_9301,N_7939);
xnor U10239 (N_10239,N_8833,N_7021);
or U10240 (N_10240,N_6426,N_5767);
nand U10241 (N_10241,N_9378,N_8259);
xor U10242 (N_10242,N_6171,N_6389);
nor U10243 (N_10243,N_7973,N_9483);
or U10244 (N_10244,N_5754,N_8425);
xor U10245 (N_10245,N_8776,N_7327);
nand U10246 (N_10246,N_8336,N_5869);
nand U10247 (N_10247,N_5469,N_8750);
xor U10248 (N_10248,N_6413,N_7056);
nor U10249 (N_10249,N_9625,N_9133);
or U10250 (N_10250,N_7572,N_7305);
or U10251 (N_10251,N_9558,N_7860);
nor U10252 (N_10252,N_6955,N_8937);
or U10253 (N_10253,N_5940,N_7020);
xnor U10254 (N_10254,N_8736,N_8710);
xor U10255 (N_10255,N_5484,N_8098);
or U10256 (N_10256,N_9448,N_8963);
xor U10257 (N_10257,N_7089,N_7311);
and U10258 (N_10258,N_5821,N_6594);
or U10259 (N_10259,N_7950,N_6515);
and U10260 (N_10260,N_7362,N_5515);
or U10261 (N_10261,N_7626,N_8180);
or U10262 (N_10262,N_8479,N_7073);
xor U10263 (N_10263,N_5958,N_9758);
nand U10264 (N_10264,N_6387,N_9996);
and U10265 (N_10265,N_5606,N_7348);
nor U10266 (N_10266,N_5243,N_9254);
nand U10267 (N_10267,N_6896,N_9938);
xnor U10268 (N_10268,N_9539,N_7493);
xnor U10269 (N_10269,N_6639,N_6672);
and U10270 (N_10270,N_9703,N_7731);
and U10271 (N_10271,N_9700,N_6342);
or U10272 (N_10272,N_6671,N_8948);
nor U10273 (N_10273,N_5983,N_9811);
nand U10274 (N_10274,N_5898,N_5936);
xor U10275 (N_10275,N_6354,N_5520);
xor U10276 (N_10276,N_7516,N_9220);
and U10277 (N_10277,N_7463,N_6294);
and U10278 (N_10278,N_8262,N_6419);
nor U10279 (N_10279,N_8698,N_8455);
nand U10280 (N_10280,N_9312,N_5758);
nand U10281 (N_10281,N_9100,N_5798);
nand U10282 (N_10282,N_8370,N_8800);
nand U10283 (N_10283,N_6860,N_9814);
nor U10284 (N_10284,N_8033,N_7600);
xor U10285 (N_10285,N_6244,N_9759);
nand U10286 (N_10286,N_6008,N_8714);
xor U10287 (N_10287,N_6839,N_7970);
nand U10288 (N_10288,N_9073,N_6283);
nor U10289 (N_10289,N_5498,N_7554);
and U10290 (N_10290,N_5020,N_7760);
and U10291 (N_10291,N_8946,N_7251);
nand U10292 (N_10292,N_8565,N_6376);
and U10293 (N_10293,N_9578,N_8993);
or U10294 (N_10294,N_9407,N_5196);
and U10295 (N_10295,N_5732,N_6072);
xor U10296 (N_10296,N_9715,N_5118);
nor U10297 (N_10297,N_8816,N_7825);
nand U10298 (N_10298,N_6803,N_6910);
nor U10299 (N_10299,N_5551,N_6382);
nor U10300 (N_10300,N_8793,N_9414);
and U10301 (N_10301,N_9706,N_7686);
xor U10302 (N_10302,N_7144,N_8647);
nand U10303 (N_10303,N_5494,N_7769);
xnor U10304 (N_10304,N_9688,N_8441);
nand U10305 (N_10305,N_5393,N_9250);
nand U10306 (N_10306,N_5348,N_6604);
and U10307 (N_10307,N_9303,N_7398);
nor U10308 (N_10308,N_6991,N_5616);
or U10309 (N_10309,N_5518,N_6946);
and U10310 (N_10310,N_5892,N_9242);
nor U10311 (N_10311,N_6744,N_5201);
nand U10312 (N_10312,N_6693,N_7037);
xnor U10313 (N_10313,N_6601,N_7364);
nor U10314 (N_10314,N_5911,N_8986);
xnor U10315 (N_10315,N_7414,N_5542);
xor U10316 (N_10316,N_8705,N_5126);
nor U10317 (N_10317,N_5920,N_8403);
nor U10318 (N_10318,N_8416,N_7213);
nor U10319 (N_10319,N_9522,N_6536);
xnor U10320 (N_10320,N_6928,N_6453);
or U10321 (N_10321,N_8942,N_6170);
or U10322 (N_10322,N_9579,N_6767);
nand U10323 (N_10323,N_7709,N_9966);
xor U10324 (N_10324,N_7561,N_7474);
and U10325 (N_10325,N_9957,N_7687);
nand U10326 (N_10326,N_8987,N_7372);
nand U10327 (N_10327,N_5432,N_9319);
nor U10328 (N_10328,N_9374,N_6617);
or U10329 (N_10329,N_6062,N_5641);
xnor U10330 (N_10330,N_5012,N_9731);
and U10331 (N_10331,N_9707,N_8068);
or U10332 (N_10332,N_9244,N_5894);
and U10333 (N_10333,N_5717,N_8465);
xor U10334 (N_10334,N_8999,N_6090);
and U10335 (N_10335,N_5095,N_8467);
or U10336 (N_10336,N_6434,N_7620);
or U10337 (N_10337,N_8553,N_5928);
nand U10338 (N_10338,N_5333,N_7854);
and U10339 (N_10339,N_8704,N_7347);
nand U10340 (N_10340,N_8149,N_7080);
nor U10341 (N_10341,N_9626,N_6460);
or U10342 (N_10342,N_7797,N_9637);
nor U10343 (N_10343,N_9824,N_7205);
nand U10344 (N_10344,N_6414,N_8900);
and U10345 (N_10345,N_5817,N_7457);
xor U10346 (N_10346,N_6801,N_7922);
nand U10347 (N_10347,N_7991,N_9257);
or U10348 (N_10348,N_8227,N_8878);
nor U10349 (N_10349,N_7418,N_5793);
and U10350 (N_10350,N_6455,N_5438);
nand U10351 (N_10351,N_6306,N_6251);
or U10352 (N_10352,N_7459,N_8846);
and U10353 (N_10353,N_5680,N_9241);
or U10354 (N_10354,N_7615,N_9536);
nor U10355 (N_10355,N_9619,N_8131);
xnor U10356 (N_10356,N_7942,N_9110);
nor U10357 (N_10357,N_7419,N_7317);
nor U10358 (N_10358,N_8175,N_8229);
or U10359 (N_10359,N_8220,N_7053);
nor U10360 (N_10360,N_6746,N_8507);
and U10361 (N_10361,N_6471,N_6179);
nor U10362 (N_10362,N_8200,N_9971);
nand U10363 (N_10363,N_6544,N_9583);
and U10364 (N_10364,N_7296,N_6060);
nand U10365 (N_10365,N_9175,N_6108);
and U10366 (N_10366,N_8790,N_6899);
or U10367 (N_10367,N_9949,N_8630);
and U10368 (N_10368,N_6900,N_7052);
nor U10369 (N_10369,N_5239,N_9931);
xor U10370 (N_10370,N_8196,N_8476);
or U10371 (N_10371,N_6235,N_7279);
xor U10372 (N_10372,N_8342,N_5722);
xnor U10373 (N_10373,N_9411,N_8095);
and U10374 (N_10374,N_8708,N_7893);
or U10375 (N_10375,N_6284,N_7320);
and U10376 (N_10376,N_6424,N_7533);
nand U10377 (N_10377,N_9545,N_7863);
nor U10378 (N_10378,N_8323,N_5021);
xor U10379 (N_10379,N_6809,N_5765);
nor U10380 (N_10380,N_5777,N_6163);
xor U10381 (N_10381,N_6960,N_9306);
xor U10382 (N_10382,N_8592,N_5005);
nand U10383 (N_10383,N_6433,N_6360);
and U10384 (N_10384,N_7048,N_6590);
or U10385 (N_10385,N_6252,N_7895);
nor U10386 (N_10386,N_8623,N_9320);
and U10387 (N_10387,N_7088,N_8780);
xnor U10388 (N_10388,N_7399,N_5369);
nor U10389 (N_10389,N_7108,N_7337);
xor U10390 (N_10390,N_8079,N_7444);
and U10391 (N_10391,N_8464,N_5736);
or U10392 (N_10392,N_8086,N_6954);
nand U10393 (N_10393,N_7204,N_6773);
xor U10394 (N_10394,N_8321,N_6752);
xor U10395 (N_10395,N_9251,N_5219);
or U10396 (N_10396,N_8664,N_9792);
or U10397 (N_10397,N_5877,N_9935);
nand U10398 (N_10398,N_7270,N_9681);
nor U10399 (N_10399,N_8114,N_7252);
nor U10400 (N_10400,N_6454,N_6611);
nor U10401 (N_10401,N_6461,N_7450);
xnor U10402 (N_10402,N_8699,N_7932);
xor U10403 (N_10403,N_9645,N_8074);
or U10404 (N_10404,N_7638,N_9851);
or U10405 (N_10405,N_8250,N_6393);
xor U10406 (N_10406,N_6821,N_7475);
and U10407 (N_10407,N_5688,N_7148);
or U10408 (N_10408,N_6858,N_8929);
xnor U10409 (N_10409,N_5084,N_7712);
nand U10410 (N_10410,N_9562,N_7800);
and U10411 (N_10411,N_7031,N_8922);
or U10412 (N_10412,N_8632,N_5426);
nand U10413 (N_10413,N_5840,N_8741);
and U10414 (N_10414,N_5405,N_7694);
nor U10415 (N_10415,N_9729,N_9381);
nand U10416 (N_10416,N_5627,N_5946);
nor U10417 (N_10417,N_6675,N_5582);
or U10418 (N_10418,N_6201,N_9622);
and U10419 (N_10419,N_6957,N_8348);
xor U10420 (N_10420,N_7189,N_6634);
nand U10421 (N_10421,N_6917,N_8895);
nand U10422 (N_10422,N_6793,N_5187);
or U10423 (N_10423,N_5143,N_6596);
xor U10424 (N_10424,N_7197,N_9921);
and U10425 (N_10425,N_5321,N_6965);
and U10426 (N_10426,N_9391,N_7226);
and U10427 (N_10427,N_5971,N_7231);
nand U10428 (N_10428,N_9294,N_7646);
nand U10429 (N_10429,N_6591,N_6350);
nand U10430 (N_10430,N_5283,N_5603);
or U10431 (N_10431,N_5452,N_8398);
or U10432 (N_10432,N_7141,N_9471);
nand U10433 (N_10433,N_9066,N_6759);
and U10434 (N_10434,N_7321,N_9902);
nor U10435 (N_10435,N_8337,N_7951);
and U10436 (N_10436,N_7831,N_5327);
nand U10437 (N_10437,N_8617,N_8587);
or U10438 (N_10438,N_9593,N_5806);
and U10439 (N_10439,N_8440,N_9549);
or U10440 (N_10440,N_9465,N_6233);
nand U10441 (N_10441,N_5098,N_7394);
nor U10442 (N_10442,N_7190,N_7663);
nand U10443 (N_10443,N_9171,N_7338);
nand U10444 (N_10444,N_9444,N_5867);
and U10445 (N_10445,N_9040,N_6718);
or U10446 (N_10446,N_7382,N_5310);
nor U10447 (N_10447,N_5063,N_5277);
nor U10448 (N_10448,N_9685,N_9088);
xnor U10449 (N_10449,N_9580,N_9496);
or U10450 (N_10450,N_9393,N_6243);
nor U10451 (N_10451,N_8022,N_5950);
xnor U10452 (N_10452,N_8767,N_5692);
or U10453 (N_10453,N_8007,N_8540);
and U10454 (N_10454,N_7013,N_9455);
and U10455 (N_10455,N_5332,N_6528);
nor U10456 (N_10456,N_9313,N_6932);
and U10457 (N_10457,N_8569,N_6359);
or U10458 (N_10458,N_8772,N_9410);
nand U10459 (N_10459,N_5536,N_8709);
xor U10460 (N_10460,N_9843,N_7968);
xor U10461 (N_10461,N_6545,N_6610);
nand U10462 (N_10462,N_9342,N_6245);
xnor U10463 (N_10463,N_9125,N_7096);
nand U10464 (N_10464,N_7094,N_6627);
nand U10465 (N_10465,N_7410,N_6280);
xor U10466 (N_10466,N_7801,N_5087);
nor U10467 (N_10467,N_5745,N_6131);
or U10468 (N_10468,N_9398,N_8734);
nor U10469 (N_10469,N_7218,N_8334);
or U10470 (N_10470,N_8691,N_9155);
or U10471 (N_10471,N_6093,N_5148);
nor U10472 (N_10472,N_6546,N_6740);
nor U10473 (N_10473,N_5794,N_6489);
nor U10474 (N_10474,N_9751,N_7793);
and U10475 (N_10475,N_5231,N_8934);
xnor U10476 (N_10476,N_7460,N_9506);
nor U10477 (N_10477,N_5751,N_6362);
or U10478 (N_10478,N_5434,N_8100);
xor U10479 (N_10479,N_9239,N_8120);
or U10480 (N_10480,N_7850,N_5235);
or U10481 (N_10481,N_8144,N_6620);
or U10482 (N_10482,N_5074,N_9888);
and U10483 (N_10483,N_8147,N_5461);
nand U10484 (N_10484,N_6764,N_5150);
nor U10485 (N_10485,N_5082,N_5058);
and U10486 (N_10486,N_9979,N_7169);
nand U10487 (N_10487,N_8359,N_5194);
xnor U10488 (N_10488,N_9463,N_9862);
nand U10489 (N_10489,N_7582,N_8775);
and U10490 (N_10490,N_6567,N_8077);
and U10491 (N_10491,N_8406,N_7255);
or U10492 (N_10492,N_6324,N_9503);
nor U10493 (N_10493,N_7216,N_5847);
and U10494 (N_10494,N_9236,N_5827);
or U10495 (N_10495,N_9621,N_7892);
or U10496 (N_10496,N_6889,N_9926);
or U10497 (N_10497,N_5335,N_8651);
or U10498 (N_10498,N_9763,N_5657);
and U10499 (N_10499,N_6997,N_7675);
and U10500 (N_10500,N_8672,N_6348);
nand U10501 (N_10501,N_5419,N_5933);
xor U10502 (N_10502,N_7024,N_5485);
xnor U10503 (N_10503,N_8042,N_8208);
and U10504 (N_10504,N_7329,N_9679);
or U10505 (N_10505,N_8466,N_5483);
xor U10506 (N_10506,N_5374,N_5737);
nor U10507 (N_10507,N_9341,N_8491);
xnor U10508 (N_10508,N_7766,N_9737);
and U10509 (N_10509,N_5506,N_6558);
xor U10510 (N_10510,N_6663,N_8158);
and U10511 (N_10511,N_8686,N_8538);
xor U10512 (N_10512,N_5280,N_7770);
nand U10513 (N_10513,N_7885,N_9948);
nor U10514 (N_10514,N_8331,N_7127);
or U10515 (N_10515,N_8103,N_9493);
xor U10516 (N_10516,N_8518,N_9467);
nand U10517 (N_10517,N_5392,N_7465);
or U10518 (N_10518,N_7350,N_6944);
and U10519 (N_10519,N_9350,N_5206);
or U10520 (N_10520,N_8444,N_5937);
xnor U10521 (N_10521,N_5647,N_5226);
xor U10522 (N_10522,N_8532,N_7609);
xnor U10523 (N_10523,N_8327,N_6047);
and U10524 (N_10524,N_9771,N_9308);
nand U10525 (N_10525,N_5010,N_6307);
nor U10526 (N_10526,N_7866,N_9511);
and U10527 (N_10527,N_9743,N_7359);
or U10528 (N_10528,N_7625,N_5996);
nand U10529 (N_10529,N_5968,N_9177);
and U10530 (N_10530,N_9423,N_9247);
and U10531 (N_10531,N_7652,N_6190);
and U10532 (N_10532,N_5250,N_9432);
xnor U10533 (N_10533,N_6887,N_6666);
and U10534 (N_10534,N_7544,N_9605);
and U10535 (N_10535,N_7274,N_5182);
nor U10536 (N_10536,N_8367,N_5404);
nor U10537 (N_10537,N_6120,N_5653);
and U10538 (N_10538,N_9161,N_5489);
nand U10539 (N_10539,N_9429,N_7492);
nand U10540 (N_10540,N_7683,N_7556);
or U10541 (N_10541,N_9300,N_6609);
and U10542 (N_10542,N_8683,N_7406);
and U10543 (N_10543,N_8864,N_6346);
or U10544 (N_10544,N_6304,N_8302);
nor U10545 (N_10545,N_8607,N_7277);
or U10546 (N_10546,N_7453,N_7490);
nor U10547 (N_10547,N_9793,N_6626);
xnor U10548 (N_10548,N_5430,N_5912);
nor U10549 (N_10549,N_9749,N_7157);
nand U10550 (N_10550,N_6670,N_5078);
and U10551 (N_10551,N_7260,N_6846);
and U10552 (N_10552,N_6237,N_9179);
or U10553 (N_10553,N_5555,N_8930);
nand U10554 (N_10554,N_6015,N_5204);
and U10555 (N_10555,N_5880,N_5790);
or U10556 (N_10556,N_7945,N_9781);
nor U10557 (N_10557,N_6340,N_6754);
and U10558 (N_10558,N_7367,N_9036);
or U10559 (N_10559,N_8473,N_7351);
nor U10560 (N_10560,N_6922,N_9667);
xor U10561 (N_10561,N_9529,N_9213);
or U10562 (N_10562,N_6749,N_7594);
nand U10563 (N_10563,N_8023,N_9620);
or U10564 (N_10564,N_8571,N_9546);
or U10565 (N_10565,N_6966,N_7143);
xor U10566 (N_10566,N_6371,N_5887);
xor U10567 (N_10567,N_6707,N_6739);
and U10568 (N_10568,N_7796,N_7393);
or U10569 (N_10569,N_9332,N_6732);
xnor U10570 (N_10570,N_6758,N_9669);
nor U10571 (N_10571,N_6573,N_9076);
xor U10572 (N_10572,N_8340,N_7795);
and U10573 (N_10573,N_6943,N_7118);
nor U10574 (N_10574,N_5370,N_6193);
nor U10575 (N_10575,N_7839,N_7834);
nor U10576 (N_10576,N_8967,N_9396);
nand U10577 (N_10577,N_9145,N_5117);
nor U10578 (N_10578,N_8275,N_8138);
or U10579 (N_10579,N_8358,N_6464);
or U10580 (N_10580,N_5217,N_5962);
nand U10581 (N_10581,N_6248,N_9544);
nor U10582 (N_10582,N_6911,N_6138);
nor U10583 (N_10583,N_8974,N_6886);
xnor U10584 (N_10584,N_9592,N_5026);
nand U10585 (N_10585,N_5838,N_6052);
and U10586 (N_10586,N_9565,N_6134);
nand U10587 (N_10587,N_6476,N_7000);
xor U10588 (N_10588,N_9240,N_5252);
xor U10589 (N_10589,N_9080,N_9172);
nand U10590 (N_10590,N_9512,N_5029);
nor U10591 (N_10591,N_7124,N_9662);
nor U10592 (N_10592,N_8462,N_6702);
nor U10593 (N_10593,N_7717,N_9863);
nand U10594 (N_10594,N_5208,N_9911);
and U10595 (N_10595,N_9750,N_7470);
nor U10596 (N_10596,N_8115,N_8724);
and U10597 (N_10597,N_5364,N_9212);
nor U10598 (N_10598,N_8738,N_6164);
nor U10599 (N_10599,N_6089,N_5124);
nand U10600 (N_10600,N_8648,N_9105);
nor U10601 (N_10601,N_5938,N_5481);
nand U10602 (N_10602,N_8868,N_8902);
and U10603 (N_10603,N_9687,N_5034);
xor U10604 (N_10604,N_6724,N_9369);
and U10605 (N_10605,N_9256,N_7730);
xor U10606 (N_10606,N_9086,N_7732);
or U10607 (N_10607,N_6510,N_5646);
and U10608 (N_10608,N_7249,N_7332);
nand U10609 (N_10609,N_5272,N_9485);
and U10610 (N_10610,N_5671,N_7010);
nand U10611 (N_10611,N_6172,N_9425);
and U10612 (N_10612,N_6400,N_8067);
and U10613 (N_10613,N_8117,N_6019);
nor U10614 (N_10614,N_8778,N_6207);
nor U10615 (N_10615,N_7816,N_8782);
and U10616 (N_10616,N_9823,N_9416);
xor U10617 (N_10617,N_7106,N_6320);
or U10618 (N_10618,N_9770,N_9140);
nor U10619 (N_10619,N_5931,N_7312);
xnor U10620 (N_10620,N_6600,N_8417);
and U10621 (N_10621,N_9224,N_9816);
xor U10622 (N_10622,N_7006,N_5696);
and U10623 (N_10623,N_6088,N_6286);
or U10624 (N_10624,N_5477,N_9216);
nand U10625 (N_10625,N_8219,N_5480);
xnor U10626 (N_10626,N_7564,N_7505);
and U10627 (N_10627,N_6953,N_7256);
and U10628 (N_10628,N_5826,N_9727);
and U10629 (N_10629,N_6678,N_7313);
nor U10630 (N_10630,N_8489,N_7672);
and U10631 (N_10631,N_7168,N_8525);
nor U10632 (N_10632,N_7880,N_5897);
nand U10633 (N_10633,N_8128,N_7966);
and U10634 (N_10634,N_9116,N_8107);
xor U10635 (N_10635,N_5527,N_6975);
or U10636 (N_10636,N_5375,N_9801);
nor U10637 (N_10637,N_7286,N_8612);
nand U10638 (N_10638,N_8136,N_6083);
nand U10639 (N_10639,N_5638,N_6177);
nor U10640 (N_10640,N_5445,N_8347);
nor U10641 (N_10641,N_9051,N_8234);
xnor U10642 (N_10642,N_8223,N_6258);
or U10643 (N_10643,N_5500,N_9584);
xor U10644 (N_10644,N_7242,N_8189);
or U10645 (N_10645,N_5373,N_6289);
and U10646 (N_10646,N_5497,N_8769);
or U10647 (N_10647,N_9599,N_5832);
xnor U10648 (N_10648,N_8983,N_7281);
nand U10649 (N_10649,N_6101,N_6814);
nor U10650 (N_10650,N_9111,N_7110);
nand U10651 (N_10651,N_5042,N_5463);
nor U10652 (N_10652,N_7420,N_8840);
xor U10653 (N_10653,N_6504,N_8645);
and U10654 (N_10654,N_7978,N_8696);
and U10655 (N_10655,N_9891,N_9203);
nor U10656 (N_10656,N_5772,N_8585);
nor U10657 (N_10657,N_7391,N_7041);
or U10658 (N_10658,N_8920,N_8770);
nor U10659 (N_10659,N_7999,N_5474);
nor U10660 (N_10660,N_6361,N_5025);
or U10661 (N_10661,N_6913,N_8222);
or U10662 (N_10662,N_8566,N_6798);
or U10663 (N_10663,N_8326,N_6927);
xor U10664 (N_10664,N_9790,N_5698);
nand U10665 (N_10665,N_5720,N_5759);
xor U10666 (N_10666,N_6025,N_6733);
xor U10667 (N_10667,N_6227,N_5929);
or U10668 (N_10668,N_5190,N_9062);
and U10669 (N_10669,N_8602,N_7604);
nand U10670 (N_10670,N_8789,N_9037);
xnor U10671 (N_10671,N_9383,N_7182);
nor U10672 (N_10672,N_7083,N_5267);
nor U10673 (N_10673,N_5949,N_6931);
nand U10674 (N_10674,N_8927,N_5449);
xnor U10675 (N_10675,N_8752,N_5257);
and U10676 (N_10676,N_5132,N_9296);
nor U10677 (N_10677,N_6430,N_6077);
and U10678 (N_10678,N_5824,N_7117);
or U10679 (N_10679,N_9984,N_6004);
or U10680 (N_10680,N_7195,N_8387);
nor U10681 (N_10681,N_9961,N_8508);
xor U10682 (N_10682,N_9449,N_6325);
nor U10683 (N_10683,N_6395,N_8373);
nor U10684 (N_10684,N_7877,N_8968);
nand U10685 (N_10685,N_6330,N_6299);
and U10686 (N_10686,N_7449,N_7150);
and U10687 (N_10687,N_7103,N_6832);
nand U10688 (N_10688,N_5200,N_8371);
nor U10689 (N_10689,N_5863,N_9680);
or U10690 (N_10690,N_7944,N_7315);
nand U10691 (N_10691,N_8815,N_9499);
and U10692 (N_10692,N_6270,N_6058);
nor U10693 (N_10693,N_5347,N_7120);
nand U10694 (N_10694,N_6266,N_9202);
and U10695 (N_10695,N_8894,N_9730);
xnor U10696 (N_10696,N_5368,N_9732);
or U10697 (N_10697,N_5161,N_9907);
or U10698 (N_10698,N_6815,N_8870);
nor U10699 (N_10699,N_6870,N_8276);
xnor U10700 (N_10700,N_7913,N_9428);
nand U10701 (N_10701,N_6837,N_5067);
xnor U10702 (N_10702,N_6605,N_7534);
and U10703 (N_10703,N_5336,N_7918);
or U10704 (N_10704,N_6553,N_7668);
nor U10705 (N_10705,N_7776,N_6756);
and U10706 (N_10706,N_6697,N_8839);
nand U10707 (N_10707,N_6480,N_6353);
xor U10708 (N_10708,N_5532,N_9328);
nor U10709 (N_10709,N_9489,N_8427);
xnor U10710 (N_10710,N_7365,N_6442);
nor U10711 (N_10711,N_8437,N_6006);
nand U10712 (N_10712,N_6578,N_5202);
and U10713 (N_10713,N_7291,N_8355);
nor U10714 (N_10714,N_7115,N_9084);
nor U10715 (N_10715,N_6994,N_5372);
nor U10716 (N_10716,N_7355,N_9912);
nand U10717 (N_10717,N_8389,N_5574);
xor U10718 (N_10718,N_8309,N_6631);
and U10719 (N_10719,N_7592,N_7729);
xnor U10720 (N_10720,N_8505,N_5378);
and U10721 (N_10721,N_5191,N_7540);
nand U10722 (N_10722,N_8555,N_6364);
nand U10723 (N_10723,N_8290,N_8624);
nor U10724 (N_10724,N_9442,N_6689);
and U10725 (N_10725,N_7757,N_5151);
nor U10726 (N_10726,N_8641,N_8031);
nor U10727 (N_10727,N_8718,N_6269);
nor U10728 (N_10728,N_8643,N_7340);
nand U10729 (N_10729,N_6698,N_7175);
nand U10730 (N_10730,N_7507,N_8560);
and U10731 (N_10731,N_5901,N_8271);
xor U10732 (N_10732,N_6380,N_6741);
xor U10733 (N_10733,N_5547,N_9507);
or U10734 (N_10734,N_8882,N_7699);
nand U10735 (N_10735,N_5170,N_9367);
xor U10736 (N_10736,N_5227,N_8781);
and U10737 (N_10737,N_9417,N_7618);
xor U10738 (N_10738,N_5433,N_9478);
xnor U10739 (N_10739,N_6655,N_9311);
xnor U10740 (N_10740,N_8595,N_6982);
nor U10741 (N_10741,N_6923,N_5492);
nor U10742 (N_10742,N_9676,N_7876);
xor U10743 (N_10743,N_6031,N_7008);
xor U10744 (N_10744,N_6972,N_6042);
xor U10745 (N_10745,N_7298,N_9636);
and U10746 (N_10746,N_9387,N_6141);
or U10747 (N_10747,N_9055,N_5690);
nand U10748 (N_10748,N_6804,N_8352);
or U10749 (N_10749,N_8303,N_6776);
nor U10750 (N_10750,N_7250,N_8652);
or U10751 (N_10751,N_9985,N_9890);
nand U10752 (N_10752,N_8594,N_5599);
and U10753 (N_10753,N_7518,N_5778);
xnor U10754 (N_10754,N_7979,N_9760);
and U10755 (N_10755,N_9092,N_7159);
nand U10756 (N_10756,N_7498,N_7803);
and U10757 (N_10757,N_5609,N_8418);
nand U10758 (N_10758,N_9627,N_6013);
xor U10759 (N_10759,N_5159,N_7821);
or U10760 (N_10760,N_5308,N_9185);
nand U10761 (N_10761,N_8707,N_6017);
xor U10762 (N_10762,N_5213,N_6394);
and U10763 (N_10763,N_7995,N_9265);
nor U10764 (N_10764,N_7720,N_8792);
or U10765 (N_10765,N_7401,N_5269);
and U10766 (N_10766,N_7357,N_9310);
or U10767 (N_10767,N_9753,N_9989);
nor U10768 (N_10768,N_8552,N_6519);
xnor U10769 (N_10769,N_6370,N_8094);
xnor U10770 (N_10770,N_9603,N_5686);
nor U10771 (N_10771,N_6212,N_8947);
and U10772 (N_10772,N_8461,N_7614);
and U10773 (N_10773,N_7012,N_8362);
nor U10774 (N_10774,N_5829,N_9473);
nand U10775 (N_10775,N_8430,N_6677);
xor U10776 (N_10776,N_8627,N_8872);
nand U10777 (N_10777,N_5312,N_7781);
or U10778 (N_10778,N_5221,N_8159);
or U10779 (N_10779,N_8526,N_6175);
nand U10780 (N_10780,N_7659,N_8404);
and U10781 (N_10781,N_8092,N_8258);
nor U10782 (N_10782,N_8381,N_5669);
nand U10783 (N_10783,N_9766,N_9613);
or U10784 (N_10784,N_6977,N_9096);
nor U10785 (N_10785,N_7887,N_7099);
nand U10786 (N_10786,N_7916,N_9011);
nand U10787 (N_10787,N_9717,N_7085);
and U10788 (N_10788,N_5803,N_9677);
and U10789 (N_10789,N_6305,N_8997);
and U10790 (N_10790,N_7133,N_9245);
nor U10791 (N_10791,N_6391,N_7727);
and U10792 (N_10792,N_6336,N_7753);
and U10793 (N_10793,N_5349,N_8396);
nor U10794 (N_10794,N_9523,N_9958);
and U10795 (N_10795,N_8060,N_6690);
xnor U10796 (N_10796,N_6161,N_8763);
nor U10797 (N_10797,N_7098,N_6647);
nand U10798 (N_10798,N_7179,N_6431);
xor U10799 (N_10799,N_5541,N_8556);
or U10800 (N_10800,N_6356,N_7992);
and U10801 (N_10801,N_8659,N_6969);
nand U10802 (N_10802,N_7081,N_9166);
nor U10803 (N_10803,N_9418,N_9196);
and U10804 (N_10804,N_6295,N_8442);
or U10805 (N_10805,N_5664,N_6228);
nand U10806 (N_10806,N_9453,N_6344);
or U10807 (N_10807,N_7580,N_6993);
and U10808 (N_10808,N_5486,N_8256);
and U10809 (N_10809,N_7087,N_9464);
or U10810 (N_10810,N_7771,N_5475);
nand U10811 (N_10811,N_5554,N_9945);
xor U10812 (N_10812,N_9993,N_8935);
xor U10813 (N_10813,N_7774,N_6737);
nor U10814 (N_10814,N_8195,N_6824);
xnor U10815 (N_10815,N_7761,N_5376);
or U10816 (N_10816,N_7427,N_7912);
xor U10817 (N_10817,N_9231,N_9885);
nand U10818 (N_10818,N_6397,N_8419);
or U10819 (N_10819,N_5266,N_8470);
and U10820 (N_10820,N_7005,N_9394);
nand U10821 (N_10821,N_8143,N_8433);
xor U10822 (N_10822,N_7234,N_7328);
nor U10823 (N_10823,N_8351,N_9441);
nor U10824 (N_10824,N_8529,N_5197);
xor U10825 (N_10825,N_7965,N_8254);
xor U10826 (N_10826,N_9656,N_5414);
and U10827 (N_10827,N_7433,N_9533);
and U10828 (N_10828,N_5024,N_9864);
nor U10829 (N_10829,N_6551,N_9882);
nor U10830 (N_10830,N_9624,N_8260);
or U10831 (N_10831,N_9340,N_9537);
and U10832 (N_10832,N_7092,N_8247);
xor U10833 (N_10833,N_9803,N_8424);
or U10834 (N_10834,N_8716,N_9960);
and U10835 (N_10835,N_9109,N_8307);
nor U10836 (N_10836,N_7558,N_6575);
xor U10837 (N_10837,N_5820,N_6936);
xnor U10838 (N_10838,N_6314,N_6024);
and U10839 (N_10839,N_6819,N_7706);
nand U10840 (N_10840,N_5508,N_6770);
or U10841 (N_10841,N_8657,N_5747);
xnor U10842 (N_10842,N_8239,N_7562);
nor U10843 (N_10843,N_8926,N_8875);
and U10844 (N_10844,N_6326,N_9225);
nor U10845 (N_10845,N_7324,N_6009);
xor U10846 (N_10846,N_8614,N_6076);
or U10847 (N_10847,N_7272,N_5588);
nor U10848 (N_10848,N_6140,N_6673);
xor U10849 (N_10849,N_5273,N_5755);
or U10850 (N_10850,N_9316,N_6040);
nor U10851 (N_10851,N_8858,N_7208);
nor U10852 (N_10852,N_7875,N_5819);
or U10853 (N_10853,N_9318,N_8413);
nand U10854 (N_10854,N_9886,N_8291);
nand U10855 (N_10855,N_6958,N_6589);
nor U10856 (N_10856,N_7984,N_5978);
and U10857 (N_10857,N_8225,N_8747);
or U10858 (N_10858,N_7900,N_8567);
xnor U10859 (N_10859,N_7897,N_9517);
nand U10860 (N_10860,N_7400,N_7055);
and U10861 (N_10861,N_5522,N_8439);
and U10862 (N_10862,N_7280,N_7438);
xor U10863 (N_10863,N_9232,N_5320);
nand U10864 (N_10864,N_8305,N_7924);
nor U10865 (N_10865,N_5845,N_8768);
nand U10866 (N_10866,N_5925,N_7002);
nand U10867 (N_10867,N_8043,N_6230);
and U10868 (N_10868,N_8783,N_6349);
xor U10869 (N_10869,N_9936,N_5386);
nand U10870 (N_10870,N_6165,N_7700);
xor U10871 (N_10871,N_9042,N_7749);
xor U10872 (N_10872,N_7884,N_7640);
or U10873 (N_10873,N_8662,N_5397);
nand U10874 (N_10874,N_9214,N_9872);
nand U10875 (N_10875,N_7033,N_7545);
and U10876 (N_10876,N_8853,N_7039);
xnor U10877 (N_10877,N_6771,N_8224);
and U10878 (N_10878,N_8483,N_8511);
xor U10879 (N_10879,N_5904,N_6614);
and U10880 (N_10880,N_7428,N_5106);
xnor U10881 (N_10881,N_6151,N_8820);
and U10882 (N_10882,N_6633,N_8860);
or U10883 (N_10883,N_6043,N_8740);
nand U10884 (N_10884,N_5589,N_8787);
nand U10885 (N_10885,N_7301,N_6477);
nor U10886 (N_10886,N_9368,N_8448);
and U10887 (N_10887,N_8153,N_7001);
xnor U10888 (N_10888,N_7542,N_7806);
or U10889 (N_10889,N_5230,N_5543);
nor U10890 (N_10890,N_5175,N_8570);
nand U10891 (N_10891,N_6595,N_7323);
and U10892 (N_10892,N_8912,N_7405);
nand U10893 (N_10893,N_8322,N_8972);
nand U10894 (N_10894,N_6490,N_7959);
and U10895 (N_10895,N_9597,N_6687);
nor U10896 (N_10896,N_7648,N_9628);
nor U10897 (N_10897,N_7018,N_5003);
nor U10898 (N_10898,N_8176,N_5954);
or U10899 (N_10899,N_6676,N_8855);
xnor U10900 (N_10900,N_7246,N_5837);
nor U10901 (N_10901,N_8654,N_8344);
and U10902 (N_10902,N_7606,N_7126);
and U10903 (N_10903,N_7377,N_6835);
nand U10904 (N_10904,N_7068,N_8788);
nand U10905 (N_10905,N_6127,N_8777);
nor U10906 (N_10906,N_6762,N_5017);
nand U10907 (N_10907,N_5714,N_8994);
xnor U10908 (N_10908,N_9253,N_8481);
xnor U10909 (N_10909,N_7070,N_8152);
nand U10910 (N_10910,N_5972,N_9883);
and U10911 (N_10911,N_9191,N_6191);
xnor U10912 (N_10912,N_7826,N_6665);
xnor U10913 (N_10913,N_6688,N_7633);
nand U10914 (N_10914,N_5533,N_6291);
nand U10915 (N_10915,N_5782,N_5730);
and U10916 (N_10916,N_9168,N_5166);
or U10917 (N_10917,N_5905,N_6037);
and U10918 (N_10918,N_9569,N_7153);
and U10919 (N_10919,N_8784,N_9136);
and U10920 (N_10920,N_8925,N_6500);
nor U10921 (N_10921,N_8265,N_7316);
nand U10922 (N_10922,N_8866,N_5297);
or U10923 (N_10923,N_5859,N_9292);
and U10924 (N_10924,N_9787,N_9498);
xor U10925 (N_10925,N_8221,N_7630);
xor U10926 (N_10926,N_6107,N_8137);
xnor U10927 (N_10927,N_7074,N_8599);
nor U10928 (N_10928,N_7903,N_6254);
and U10929 (N_10929,N_8233,N_8304);
or U10930 (N_10930,N_6576,N_5389);
xor U10931 (N_10931,N_9608,N_9634);
or U10932 (N_10932,N_8029,N_8057);
and U10933 (N_10933,N_8006,N_6668);
and U10934 (N_10934,N_5493,N_9721);
nor U10935 (N_10935,N_5537,N_5579);
nand U10936 (N_10936,N_8454,N_9029);
and U10937 (N_10937,N_9048,N_5805);
or U10938 (N_10938,N_5674,N_5134);
or U10939 (N_10939,N_8932,N_8292);
nand U10940 (N_10940,N_5586,N_9348);
nand U10941 (N_10941,N_6250,N_8850);
and U10942 (N_10942,N_7674,N_8545);
or U10943 (N_10943,N_9160,N_7814);
or U10944 (N_10944,N_5503,N_6907);
nand U10945 (N_10945,N_5309,N_9646);
xor U10946 (N_10946,N_5775,N_8886);
and U10947 (N_10947,N_5947,N_6085);
nor U10948 (N_10948,N_5870,N_5675);
or U10949 (N_10949,N_8822,N_6805);
nand U10950 (N_10950,N_6711,N_6806);
nand U10951 (N_10951,N_8905,N_7636);
xor U10952 (N_10952,N_8758,N_8118);
nor U10953 (N_10953,N_7187,N_7627);
and U10954 (N_10954,N_8854,N_5282);
xnor U10955 (N_10955,N_9922,N_7275);
nand U10956 (N_10956,N_8487,N_9726);
or U10957 (N_10957,N_6728,N_9371);
and U10958 (N_10958,N_5365,N_6256);
nand U10959 (N_10959,N_9689,N_5886);
or U10960 (N_10960,N_5476,N_6268);
nand U10961 (N_10961,N_8411,N_5833);
or U10962 (N_10962,N_7896,N_8121);
nand U10963 (N_10963,N_6018,N_7697);
xnor U10964 (N_10964,N_6482,N_8956);
xnor U10965 (N_10965,N_9283,N_5090);
or U10966 (N_10966,N_5723,N_9120);
nor U10967 (N_10967,N_7422,N_9438);
nand U10968 (N_10968,N_5948,N_5198);
nor U10969 (N_10969,N_7192,N_7199);
and U10970 (N_10970,N_6919,N_8268);
nor U10971 (N_10971,N_5346,N_7693);
nor U10972 (N_10972,N_6674,N_5927);
or U10973 (N_10973,N_5472,N_7705);
nand U10974 (N_10974,N_7212,N_9327);
nor U10975 (N_10975,N_7331,N_8013);
or U10976 (N_10976,N_7645,N_7211);
and U10977 (N_10977,N_8828,N_8745);
and U10978 (N_10978,N_8356,N_8412);
xor U10979 (N_10979,N_7634,N_5883);
nor U10980 (N_10980,N_6531,N_9226);
and U10981 (N_10981,N_8261,N_8408);
xor U10982 (N_10982,N_5951,N_9828);
nor U10983 (N_10983,N_7128,N_9262);
xor U10984 (N_10984,N_6505,N_5762);
or U10985 (N_10985,N_6851,N_9248);
nand U10986 (N_10986,N_6947,N_6449);
and U10987 (N_10987,N_5168,N_6750);
nor U10988 (N_10988,N_9830,N_9287);
or U10989 (N_10989,N_6780,N_8284);
or U10990 (N_10990,N_5763,N_7838);
nor U10991 (N_10991,N_9379,N_8056);
and U10992 (N_10992,N_8488,N_5160);
xnor U10993 (N_10993,N_5258,N_7509);
or U10994 (N_10994,N_8656,N_8634);
and U10995 (N_10995,N_6176,N_9046);
or U10996 (N_10996,N_5222,N_5028);
xor U10997 (N_10997,N_8913,N_7681);
xnor U10998 (N_10998,N_8838,N_9796);
or U10999 (N_10999,N_8578,N_7987);
nor U11000 (N_11000,N_6694,N_7258);
or U11001 (N_11001,N_9983,N_8032);
xor U11002 (N_11002,N_6195,N_6588);
nand U11003 (N_11003,N_8324,N_8834);
xnor U11004 (N_11004,N_7623,N_7845);
xnor U11005 (N_11005,N_9149,N_9094);
nand U11006 (N_11006,N_5107,N_5299);
nor U11007 (N_11007,N_6064,N_6945);
nand U11008 (N_11008,N_6532,N_6651);
or U11009 (N_11009,N_9447,N_8564);
nor U11010 (N_11010,N_7015,N_6848);
xor U11011 (N_11011,N_9964,N_8070);
xor U11012 (N_11012,N_8881,N_6002);
nor U11013 (N_11013,N_6092,N_6984);
nor U11014 (N_11014,N_6319,N_6290);
nor U11015 (N_11015,N_9899,N_9953);
and U11016 (N_11016,N_7735,N_7467);
and U11017 (N_11017,N_9629,N_5270);
nor U11018 (N_11018,N_5682,N_5529);
nand U11019 (N_11019,N_6847,N_7289);
and U11020 (N_11020,N_5014,N_5097);
and U11021 (N_11021,N_5007,N_5560);
xnor U11022 (N_11022,N_9660,N_9894);
and U11023 (N_11023,N_7767,N_6162);
and U11024 (N_11024,N_9745,N_8949);
and U11025 (N_11025,N_6114,N_7768);
nand U11026 (N_11026,N_5044,N_9122);
or U11027 (N_11027,N_8808,N_8961);
and U11028 (N_11028,N_9238,N_7266);
xnor U11029 (N_11029,N_9041,N_9376);
nor U11030 (N_11030,N_5157,N_8295);
nor U11031 (N_11031,N_5960,N_6123);
or U11032 (N_11032,N_5075,N_9405);
xor U11033 (N_11033,N_9475,N_5167);
and U11034 (N_11034,N_7322,N_7506);
and U11035 (N_11035,N_8658,N_5290);
or U11036 (N_11036,N_9725,N_8890);
xor U11037 (N_11037,N_6409,N_7193);
and U11038 (N_11038,N_9869,N_5487);
or U11039 (N_11039,N_8568,N_6495);
and U11040 (N_11040,N_6224,N_7701);
and U11041 (N_11041,N_5670,N_5071);
nand U11042 (N_11042,N_8779,N_8577);
nor U11043 (N_11043,N_7908,N_9082);
xnor U11044 (N_11044,N_8339,N_9831);
nand U11045 (N_11045,N_7670,N_6068);
xnor U11046 (N_11046,N_8965,N_8299);
xor U11047 (N_11047,N_8129,N_6238);
nor U11048 (N_11048,N_5660,N_7628);
nand U11049 (N_11049,N_8524,N_8919);
or U11050 (N_11050,N_5418,N_8112);
or U11051 (N_11051,N_5741,N_7579);
nor U11052 (N_11052,N_6962,N_9492);
nand U11053 (N_11053,N_6844,N_6278);
and U11054 (N_11054,N_9077,N_6223);
nor U11055 (N_11055,N_6368,N_5893);
nand U11056 (N_11056,N_7928,N_7882);
and U11057 (N_11057,N_8062,N_8139);
nor U11058 (N_11058,N_9618,N_6549);
xnor U11059 (N_11059,N_6339,N_9285);
nor U11060 (N_11060,N_6446,N_7931);
or U11061 (N_11061,N_7136,N_7949);
nor U11062 (N_11062,N_5172,N_9060);
nor U11063 (N_11063,N_6499,N_5249);
xor U11064 (N_11064,N_7439,N_6769);
nand U11065 (N_11065,N_7650,N_5424);
nand U11066 (N_11066,N_5103,N_6316);
and U11067 (N_11067,N_6527,N_6069);
or U11068 (N_11068,N_9761,N_8397);
nand U11069 (N_11069,N_7510,N_9001);
xnor U11070 (N_11070,N_7662,N_8021);
or U11071 (N_11071,N_9776,N_8164);
nand U11072 (N_11072,N_5810,N_6403);
nor U11073 (N_11073,N_8959,N_5453);
xor U11074 (N_11074,N_7014,N_9861);
and U11075 (N_11075,N_7139,N_7066);
or U11076 (N_11076,N_9757,N_8241);
and U11077 (N_11077,N_5395,N_6802);
and U11078 (N_11078,N_8586,N_9521);
nand U11079 (N_11079,N_6777,N_9273);
xnor U11080 (N_11080,N_5174,N_5188);
and U11081 (N_11081,N_8445,N_7790);
nand U11082 (N_11082,N_9353,N_9012);
nor U11083 (N_11083,N_5594,N_7109);
or U11084 (N_11084,N_8896,N_7651);
or U11085 (N_11085,N_7227,N_5259);
nand U11086 (N_11086,N_6322,N_7960);
and U11087 (N_11087,N_6967,N_5344);
xor U11088 (N_11088,N_8490,N_8506);
xnor U11089 (N_11089,N_6187,N_8104);
nand U11090 (N_11090,N_8695,N_5215);
or U11091 (N_11091,N_9419,N_5791);
nor U11092 (N_11092,N_9955,N_5116);
or U11093 (N_11093,N_9392,N_9639);
and U11094 (N_11094,N_8675,N_8914);
or U11095 (N_11095,N_9335,N_6653);
and U11096 (N_11096,N_9802,N_8845);
nor U11097 (N_11097,N_7034,N_9325);
nor U11098 (N_11098,N_9095,N_9794);
and U11099 (N_11099,N_5713,N_5088);
nor U11100 (N_11100,N_7149,N_7370);
xor U11101 (N_11101,N_8475,N_5363);
nor U11102 (N_11102,N_7384,N_8824);
nand U11103 (N_11103,N_7023,N_9752);
xor U11104 (N_11104,N_8690,N_9713);
or U11105 (N_11105,N_6988,N_5673);
nor U11106 (N_11106,N_5525,N_9825);
and U11107 (N_11107,N_6684,N_9577);
and U11108 (N_11108,N_7711,N_7325);
nand U11109 (N_11109,N_8677,N_5715);
xnor U11110 (N_11110,N_8008,N_7486);
and U11111 (N_11111,N_6030,N_8823);
nand U11112 (N_11112,N_6481,N_7748);
and U11113 (N_11113,N_9460,N_8639);
nor U11114 (N_11114,N_9208,N_8020);
nor U11115 (N_11115,N_7715,N_6386);
nand U11116 (N_11116,N_7899,N_5862);
nand U11117 (N_11117,N_8499,N_7152);
and U11118 (N_11118,N_8521,N_5340);
or U11119 (N_11119,N_8861,N_9690);
and U11120 (N_11120,N_7940,N_8399);
or U11121 (N_11121,N_5733,N_5342);
xnor U11122 (N_11122,N_6612,N_7941);
nand U11123 (N_11123,N_8628,N_9982);
xor U11124 (N_11124,N_9270,N_5939);
xnor U11125 (N_11125,N_6247,N_9786);
nor U11126 (N_11126,N_9207,N_9859);
nor U11127 (N_11127,N_8099,N_7692);
and U11128 (N_11128,N_8049,N_7385);
or U11129 (N_11129,N_8534,N_5417);
and U11130 (N_11130,N_8201,N_9364);
nor U11131 (N_11131,N_7007,N_9799);
xor U11132 (N_11132,N_5860,N_7934);
and U11133 (N_11133,N_9913,N_7840);
or U11134 (N_11134,N_6700,N_6811);
and U11135 (N_11135,N_6439,N_7710);
or U11136 (N_11136,N_7685,N_6273);
xnor U11137 (N_11137,N_8807,N_6914);
nor U11138 (N_11138,N_8960,N_8543);
nand U11139 (N_11139,N_5855,N_8282);
xnor U11140 (N_11140,N_8832,N_7733);
nand U11141 (N_11141,N_5639,N_6566);
and U11142 (N_11142,N_9881,N_6520);
xnor U11143 (N_11143,N_8980,N_7302);
nor U11144 (N_11144,N_9146,N_5298);
nand U11145 (N_11145,N_5631,N_5379);
xor U11146 (N_11146,N_8210,N_6941);
or U11147 (N_11147,N_8045,N_5666);
nor U11148 (N_11148,N_9780,N_6935);
xnor U11149 (N_11149,N_5356,N_6199);
or U11150 (N_11150,N_6556,N_6147);
xor U11151 (N_11151,N_6986,N_6731);
nand U11152 (N_11152,N_5233,N_9820);
and U11153 (N_11153,N_9954,N_5544);
and U11154 (N_11154,N_8102,N_7813);
or U11155 (N_11155,N_8563,N_5304);
or U11156 (N_11156,N_6075,N_7164);
xnor U11157 (N_11157,N_8830,N_7154);
xnor U11158 (N_11158,N_5661,N_9997);
nor U11159 (N_11159,N_7739,N_9330);
nand U11160 (N_11160,N_7408,N_7151);
nand U11161 (N_11161,N_9452,N_7758);
nand U11162 (N_11162,N_9900,N_9879);
and U11163 (N_11163,N_9695,N_6117);
xor U11164 (N_11164,N_7798,N_9906);
nand U11165 (N_11165,N_8954,N_8876);
or U11166 (N_11166,N_9959,N_6429);
xnor U11167 (N_11167,N_8984,N_5725);
or U11168 (N_11168,N_7244,N_8165);
and U11169 (N_11169,N_5740,N_5648);
nor U11170 (N_11170,N_8765,N_6182);
nor U11171 (N_11171,N_6522,N_8520);
or U11172 (N_11172,N_7575,N_5693);
nand U11173 (N_11173,N_5808,N_8810);
xor U11174 (N_11174,N_7792,N_5281);
or U11175 (N_11175,N_9157,N_6055);
and U11176 (N_11176,N_7203,N_5974);
xnor U11177 (N_11177,N_6867,N_7946);
nor U11178 (N_11178,N_8168,N_6049);
xor U11179 (N_11179,N_6281,N_5119);
or U11180 (N_11180,N_8402,N_8889);
nand U11181 (N_11181,N_6208,N_9352);
nand U11182 (N_11182,N_6204,N_9286);
xor U11183 (N_11183,N_8214,N_5181);
nand U11184 (N_11184,N_9290,N_5147);
nor U11185 (N_11185,N_9930,N_8410);
or U11186 (N_11186,N_9181,N_6154);
or U11187 (N_11187,N_6144,N_8608);
and U11188 (N_11188,N_6582,N_7818);
and U11189 (N_11189,N_8266,N_5464);
nor U11190 (N_11190,N_5138,N_6133);
or U11191 (N_11191,N_5015,N_8613);
nor U11192 (N_11192,N_7607,N_9554);
and U11193 (N_11193,N_5550,N_6772);
xnor U11194 (N_11194,N_8142,N_6508);
and U11195 (N_11195,N_8754,N_6823);
nor U11196 (N_11196,N_8320,N_7515);
nand U11197 (N_11197,N_6262,N_6511);
nor U11198 (N_11198,N_7318,N_5205);
or U11199 (N_11199,N_5471,N_7417);
or U11200 (N_11200,N_6792,N_8943);
or U11201 (N_11201,N_7642,N_5455);
nor U11202 (N_11202,N_5129,N_5504);
xor U11203 (N_11203,N_7479,N_9363);
nor U11204 (N_11204,N_8124,N_5955);
and U11205 (N_11205,N_6999,N_5121);
or U11206 (N_11206,N_5096,N_5921);
or U11207 (N_11207,N_9905,N_9377);
and U11208 (N_11208,N_6150,N_6866);
and U11209 (N_11209,N_7658,N_6050);
xnor U11210 (N_11210,N_8590,N_5800);
xnor U11211 (N_11211,N_9134,N_7236);
or U11212 (N_11212,N_5531,N_9209);
xor U11213 (N_11213,N_8449,N_7481);
nand U11214 (N_11214,N_9887,N_8827);
xor U11215 (N_11215,N_9832,N_6906);
or U11216 (N_11216,N_8725,N_9736);
or U11217 (N_11217,N_9691,N_6184);
nand U11218 (N_11218,N_8852,N_9769);
and U11219 (N_11219,N_7552,N_8527);
nand U11220 (N_11220,N_9436,N_7867);
and U11221 (N_11221,N_9596,N_8246);
xor U11222 (N_11222,N_6308,N_6094);
and U11223 (N_11223,N_7503,N_7207);
and U11224 (N_11224,N_6491,N_9132);
nand U11225 (N_11225,N_7038,N_5501);
and U11226 (N_11226,N_9000,N_7985);
or U11227 (N_11227,N_7812,N_6807);
or U11228 (N_11228,N_5961,N_7354);
xnor U11229 (N_11229,N_8172,N_6643);
and U11230 (N_11230,N_9326,N_7174);
nand U11231 (N_11231,N_9013,N_9571);
nor U11232 (N_11232,N_7009,N_7435);
and U11233 (N_11233,N_9445,N_6445);
nand U11234 (N_11234,N_6363,N_6135);
or U11235 (N_11235,N_8973,N_7851);
xnor U11236 (N_11236,N_6046,N_6221);
nand U11237 (N_11237,N_8760,N_7736);
nand U11238 (N_11238,N_8514,N_9390);
nor U11239 (N_11239,N_5568,N_7183);
or U11240 (N_11240,N_6820,N_8040);
xor U11241 (N_11241,N_9479,N_5294);
nand U11242 (N_11242,N_9490,N_8187);
nand U11243 (N_11243,N_8544,N_9838);
xor U11244 (N_11244,N_9331,N_8720);
and U11245 (N_11245,N_9389,N_6656);
xnor U11246 (N_11246,N_6507,N_7823);
or U11247 (N_11247,N_8897,N_6895);
and U11248 (N_11248,N_7541,N_5942);
xnor U11249 (N_11249,N_6443,N_7177);
xnor U11250 (N_11250,N_9005,N_7202);
nand U11251 (N_11251,N_9514,N_9652);
nand U11252 (N_11252,N_7050,N_9909);
and U11253 (N_11253,N_8345,N_9264);
nand U11254 (N_11254,N_9008,N_7963);
nand U11255 (N_11255,N_8108,N_6654);
xor U11256 (N_11256,N_9446,N_8802);
and U11257 (N_11257,N_9977,N_6552);
nor U11258 (N_11258,N_5752,N_9039);
and U11259 (N_11259,N_9028,N_6005);
nand U11260 (N_11260,N_5572,N_6122);
xor U11261 (N_11261,N_5381,N_5416);
xor U11262 (N_11262,N_6682,N_5403);
and U11263 (N_11263,N_5524,N_9083);
nor U11264 (N_11264,N_8447,N_5570);
xnor U11265 (N_11265,N_8576,N_5511);
nor U11266 (N_11266,N_8908,N_6996);
nand U11267 (N_11267,N_9805,N_6032);
nor U11268 (N_11268,N_5634,N_8197);
nor U11269 (N_11269,N_7680,N_6384);
and U11270 (N_11270,N_6067,N_7112);
and U11271 (N_11271,N_7330,N_7167);
xnor U11272 (N_11272,N_8636,N_8547);
nand U11273 (N_11273,N_6976,N_7416);
nor U11274 (N_11274,N_6989,N_7477);
xor U11275 (N_11275,N_8650,N_5652);
nand U11276 (N_11276,N_5749,N_9223);
nand U11277 (N_11277,N_9665,N_8582);
and U11278 (N_11278,N_5460,N_5130);
nand U11279 (N_11279,N_6293,N_6763);
nor U11280 (N_11280,N_7043,N_7147);
and U11281 (N_11281,N_6765,N_7808);
nor U11282 (N_11282,N_6412,N_6276);
nand U11283 (N_11283,N_6475,N_9267);
nand U11284 (N_11284,N_8693,N_5177);
or U11285 (N_11285,N_8308,N_7921);
or U11286 (N_11286,N_5694,N_6255);
nor U11287 (N_11287,N_7402,N_6203);
and U11288 (N_11288,N_7639,N_5923);
or U11289 (N_11289,N_5509,N_9568);
xor U11290 (N_11290,N_6602,N_7412);
and U11291 (N_11291,N_5428,N_9474);
nand U11292 (N_11292,N_8901,N_8958);
nand U11293 (N_11293,N_9298,N_6753);
and U11294 (N_11294,N_6142,N_5622);
xnor U11295 (N_11295,N_7036,N_8035);
and U11296 (N_11296,N_5192,N_9020);
or U11297 (N_11297,N_6517,N_8909);
xnor U11298 (N_11298,N_6452,N_7268);
or U11299 (N_11299,N_9128,N_5781);
xnor U11300 (N_11300,N_6232,N_7181);
or U11301 (N_11301,N_8088,N_9056);
nor U11302 (N_11302,N_9183,N_9892);
and U11303 (N_11303,N_6784,N_7780);
nand U11304 (N_11304,N_5406,N_8438);
nor U11305 (N_11305,N_9486,N_5969);
or U11306 (N_11306,N_7264,N_8723);
xor U11307 (N_11307,N_5956,N_9016);
and U11308 (N_11308,N_7440,N_5932);
xor U11309 (N_11309,N_8281,N_8026);
nand U11310 (N_11310,N_5649,N_6355);
nor U11311 (N_11311,N_5289,N_9783);
and U11312 (N_11312,N_6402,N_9898);
xor U11313 (N_11313,N_6148,N_7716);
nand U11314 (N_11314,N_6001,N_5678);
nand U11315 (N_11315,N_8141,N_5865);
nor U11316 (N_11316,N_8240,N_6377);
nand U11317 (N_11317,N_7430,N_6086);
xnor U11318 (N_11318,N_5569,N_8155);
nor U11319 (N_11319,N_7578,N_6959);
or U11320 (N_11320,N_8274,N_5773);
nor U11321 (N_11321,N_5809,N_8771);
nand U11322 (N_11322,N_7661,N_6155);
xnor U11323 (N_11323,N_8061,N_9047);
nand U11324 (N_11324,N_6645,N_7894);
xnor U11325 (N_11325,N_6971,N_9219);
or U11326 (N_11326,N_8041,N_8338);
or U11327 (N_11327,N_9426,N_6444);
and U11328 (N_11328,N_5879,N_6952);
or U11329 (N_11329,N_6112,N_6577);
xor U11330 (N_11330,N_7487,N_5571);
xnor U11331 (N_11331,N_8423,N_5796);
nor U11332 (N_11332,N_5706,N_6547);
and U11333 (N_11333,N_5288,N_7849);
or U11334 (N_11334,N_5291,N_8054);
nand U11335 (N_11335,N_6565,N_8369);
and U11336 (N_11336,N_6810,N_8859);
or U11337 (N_11337,N_8735,N_8805);
or U11338 (N_11338,N_8432,N_7027);
or U11339 (N_11339,N_7901,N_9057);
nor U11340 (N_11340,N_8515,N_8361);
nor U11341 (N_11341,N_8880,N_6450);
or U11342 (N_11342,N_9059,N_5169);
and U11343 (N_11343,N_6110,N_7755);
nand U11344 (N_11344,N_7489,N_6317);
xor U11345 (N_11345,N_7241,N_6901);
nand U11346 (N_11346,N_8588,N_5990);
xor U11347 (N_11347,N_8426,N_6735);
nor U11348 (N_11348,N_8542,N_8005);
and U11349 (N_11349,N_9784,N_8130);
nand U11350 (N_11350,N_7621,N_5651);
xnor U11351 (N_11351,N_9365,N_5528);
and U11352 (N_11352,N_7288,N_7707);
nor U11353 (N_11353,N_7155,N_5225);
nor U11354 (N_11354,N_7571,N_6742);
nand U11355 (N_11355,N_5830,N_8561);
nor U11356 (N_11356,N_8395,N_6873);
nand U11357 (N_11357,N_5584,N_6883);
and U11358 (N_11358,N_5676,N_6755);
nand U11359 (N_11359,N_7969,N_7754);
nor U11360 (N_11360,N_6275,N_9334);
nor U11361 (N_11361,N_8123,N_5784);
nand U11362 (N_11362,N_9675,N_8898);
or U11363 (N_11363,N_8177,N_6297);
nand U11364 (N_11364,N_9702,N_7390);
nand U11365 (N_11365,N_6215,N_5359);
or U11366 (N_11366,N_7295,N_8883);
nor U11367 (N_11367,N_7848,N_8991);
nand U11368 (N_11368,N_5366,N_7119);
nor U11369 (N_11369,N_6309,N_5620);
and U11370 (N_11370,N_6296,N_6623);
and U11371 (N_11371,N_8213,N_8873);
and U11372 (N_11372,N_5598,N_6559);
nand U11373 (N_11373,N_9153,N_9259);
and U11374 (N_11374,N_5667,N_9329);
nand U11375 (N_11375,N_6892,N_5009);
xnor U11376 (N_11376,N_7678,N_9221);
xnor U11377 (N_11377,N_9821,N_5776);
nor U11378 (N_11378,N_8990,N_9975);
nor U11379 (N_11379,N_5779,N_5146);
and U11380 (N_11380,N_9482,N_7881);
nor U11381 (N_11381,N_6834,N_5702);
and U11382 (N_11382,N_6432,N_6073);
and U11383 (N_11383,N_6405,N_8706);
xor U11384 (N_11384,N_6603,N_6056);
xnor U11385 (N_11385,N_8678,N_8460);
nand U11386 (N_11386,N_5663,N_6550);
or U11387 (N_11387,N_8306,N_9819);
nand U11388 (N_11388,N_9106,N_5854);
or U11389 (N_11389,N_7191,N_8484);
xnor U11390 (N_11390,N_6705,N_8885);
nor U11391 (N_11391,N_8193,N_8145);
or U11392 (N_11392,N_7230,N_6790);
and U11393 (N_11393,N_7265,N_9633);
nor U11394 (N_11394,N_8933,N_7971);
nand U11395 (N_11395,N_9768,N_6885);
nor U11396 (N_11396,N_7309,N_5122);
nor U11397 (N_11397,N_6538,N_9091);
or U11398 (N_11398,N_6029,N_9274);
nand U11399 (N_11399,N_9547,N_7059);
xnor U11400 (N_11400,N_7858,N_5981);
or U11401 (N_11401,N_5987,N_9917);
and U11402 (N_11402,N_8512,N_7853);
xnor U11403 (N_11403,N_9431,N_8977);
xnor U11404 (N_11404,N_9261,N_8253);
xor U11405 (N_11405,N_8976,N_7998);
nor U11406 (N_11406,N_8495,N_5382);
and U11407 (N_11407,N_7517,N_9089);
or U11408 (N_11408,N_8082,N_6341);
xor U11409 (N_11409,N_9151,N_8199);
or U11410 (N_11410,N_5110,N_9773);
xnor U11411 (N_11411,N_5039,N_8940);
xnor U11412 (N_11412,N_5391,N_8589);
nand U11413 (N_11413,N_6524,N_9395);
nor U11414 (N_11414,N_8536,N_6106);
or U11415 (N_11415,N_9215,N_6632);
or U11416 (N_11416,N_8610,N_7841);
and U11417 (N_11417,N_7993,N_7869);
and U11418 (N_11418,N_5038,N_7194);
nand U11419 (N_11419,N_7574,N_8907);
and U11420 (N_11420,N_6220,N_8376);
and U11421 (N_11421,N_9476,N_8541);
nand U11422 (N_11422,N_6587,N_6555);
xor U11423 (N_11423,N_5287,N_7878);
and U11424 (N_11424,N_7371,N_5705);
nand U11425 (N_11425,N_9397,N_6463);
or U11426 (N_11426,N_5561,N_6301);
nand U11427 (N_11427,N_6119,N_7307);
nor U11428 (N_11428,N_9370,N_7603);
or U11429 (N_11429,N_9148,N_6494);
nor U11430 (N_11430,N_8941,N_5247);
nand U11431 (N_11431,N_5977,N_8692);
or U11432 (N_11432,N_6035,N_9551);
and U11433 (N_11433,N_9532,N_6757);
nor U11434 (N_11434,N_8394,N_5552);
or U11435 (N_11435,N_6440,N_5526);
and U11436 (N_11436,N_9413,N_9908);
or U11437 (N_11437,N_5271,N_5576);
nor U11438 (N_11438,N_6425,N_8616);
xor U11439 (N_11439,N_6407,N_8817);
nor U11440 (N_11440,N_7051,N_5727);
and U11441 (N_11441,N_7955,N_8378);
and U11442 (N_11442,N_7238,N_8701);
and U11443 (N_11443,N_9277,N_5521);
xnor U11444 (N_11444,N_7619,N_5618);
nor U11445 (N_11445,N_9403,N_6399);
or U11446 (N_11446,N_7040,N_5353);
nand U11447 (N_11447,N_8717,N_9218);
and U11448 (N_11448,N_9141,N_7843);
and U11449 (N_11449,N_6267,N_9178);
or U11450 (N_11450,N_5158,N_8528);
or U11451 (N_11451,N_6000,N_6264);
nor U11452 (N_11452,N_5446,N_8572);
nand U11453 (N_11453,N_8018,N_6159);
nor U11454 (N_11454,N_5236,N_9849);
or U11455 (N_11455,N_5875,N_8995);
nand U11456 (N_11456,N_6585,N_6337);
and U11457 (N_11457,N_7222,N_5008);
nor U11458 (N_11458,N_5326,N_9205);
nand U11459 (N_11459,N_5491,N_5091);
and U11460 (N_11460,N_5055,N_5899);
xnor U11461 (N_11461,N_8047,N_6375);
nor U11462 (N_11462,N_5300,N_8379);
nand U11463 (N_11463,N_9130,N_8923);
and U11464 (N_11464,N_5998,N_8257);
nand U11465 (N_11465,N_7269,N_6635);
xnor U11466 (N_11466,N_9590,N_5607);
nor U11467 (N_11467,N_6876,N_9305);
nand U11468 (N_11468,N_9114,N_8539);
nand U11469 (N_11469,N_9090,N_5677);
nand U11470 (N_11470,N_7425,N_6332);
and U11471 (N_11471,N_8204,N_7743);
nor U11472 (N_11472,N_5385,N_7198);
or U11473 (N_11473,N_7862,N_5851);
nand U11474 (N_11474,N_5402,N_6833);
xnor U11475 (N_11475,N_9201,N_5052);
nor U11476 (N_11476,N_8795,N_6313);
xor U11477 (N_11477,N_6415,N_8550);
and U11478 (N_11478,N_7461,N_5457);
nor U11479 (N_11479,N_6271,N_6012);
and U11480 (N_11480,N_8294,N_7981);
xnor U11481 (N_11481,N_5330,N_5628);
or U11482 (N_11482,N_5600,N_6310);
nand U11483 (N_11483,N_6272,N_6218);
or U11484 (N_11484,N_7426,N_8471);
nand U11485 (N_11485,N_8915,N_6091);
or U11486 (N_11486,N_5611,N_8739);
and U11487 (N_11487,N_8762,N_5189);
or U11488 (N_11488,N_7972,N_6640);
and U11489 (N_11489,N_5360,N_6888);
or U11490 (N_11490,N_8167,N_7214);
and U11491 (N_11491,N_8287,N_9718);
or U11492 (N_11492,N_7671,N_6198);
and U11493 (N_11493,N_8680,N_7986);
and U11494 (N_11494,N_8093,N_5006);
nor U11495 (N_11495,N_7201,N_9623);
and U11496 (N_11496,N_6563,N_5441);
or U11497 (N_11497,N_9710,N_7413);
nand U11498 (N_11498,N_6608,N_5645);
xnor U11499 (N_11499,N_7060,N_6542);
nor U11500 (N_11500,N_9602,N_7029);
xnor U11501 (N_11501,N_5672,N_7889);
and U11502 (N_11502,N_8178,N_9967);
xnor U11503 (N_11503,N_5970,N_5683);
and U11504 (N_11504,N_9929,N_5367);
or U11505 (N_11505,N_8727,N_5841);
nand U11506 (N_11506,N_7819,N_6699);
or U11507 (N_11507,N_6345,N_9777);
or U11508 (N_11508,N_6861,N_9052);
and U11509 (N_11509,N_8494,N_9237);
or U11510 (N_11510,N_9309,N_5822);
nor U11511 (N_11511,N_8169,N_9895);
nor U11512 (N_11512,N_6104,N_7947);
nand U11513 (N_11513,N_9085,N_6710);
and U11514 (N_11514,N_5306,N_9293);
nor U11515 (N_11515,N_5120,N_6437);
xnor U11516 (N_11516,N_8230,N_9560);
xnor U11517 (N_11517,N_9845,N_5064);
nor U11518 (N_11518,N_6211,N_9648);
xor U11519 (N_11519,N_7185,N_7775);
nand U11520 (N_11520,N_9026,N_5635);
and U11521 (N_11521,N_9880,N_6722);
and U11522 (N_11522,N_7162,N_6185);
and U11523 (N_11523,N_6723,N_5889);
or U11524 (N_11524,N_6003,N_9229);
nor U11525 (N_11525,N_5559,N_8216);
or U11526 (N_11526,N_8957,N_5060);
or U11527 (N_11527,N_9600,N_7830);
xnor U11528 (N_11528,N_5108,N_6118);
or U11529 (N_11529,N_9470,N_9275);
nand U11530 (N_11530,N_5991,N_6398);
or U11531 (N_11531,N_9385,N_5581);
xor U11532 (N_11532,N_8474,N_6523);
or U11533 (N_11533,N_7689,N_7245);
or U11534 (N_11534,N_7361,N_6462);
xnor U11535 (N_11535,N_5465,N_8436);
nor U11536 (N_11536,N_7704,N_7065);
or U11537 (N_11537,N_5864,N_9500);
and U11538 (N_11538,N_6930,N_7647);
nand U11539 (N_11539,N_6302,N_6196);
or U11540 (N_11540,N_8848,N_9557);
xnor U11541 (N_11541,N_7547,N_5100);
xor U11542 (N_11542,N_6571,N_5112);
or U11543 (N_11543,N_6113,N_9848);
xor U11544 (N_11544,N_9504,N_9942);
nand U11545 (N_11545,N_6841,N_9249);
nand U11546 (N_11546,N_6951,N_9098);
xnor U11547 (N_11547,N_7494,N_9857);
xor U11548 (N_11548,N_7335,N_5766);
nor U11549 (N_11549,N_7044,N_9351);
and U11550 (N_11550,N_9045,N_6323);
and U11551 (N_11551,N_7030,N_5665);
or U11552 (N_11552,N_6288,N_8374);
and U11553 (N_11553,N_6533,N_7954);
xor U11554 (N_11554,N_9322,N_7930);
xnor U11555 (N_11555,N_9535,N_5852);
xor U11556 (N_11556,N_7871,N_5139);
nand U11557 (N_11557,N_5184,N_9211);
nand U11558 (N_11558,N_9526,N_6422);
or U11559 (N_11559,N_5989,N_7695);
nor U11560 (N_11560,N_9800,N_9655);
xor U11561 (N_11561,N_8644,N_5185);
or U11562 (N_11562,N_7336,N_8458);
nor U11563 (N_11563,N_7590,N_7974);
and U11564 (N_11564,N_5995,N_6516);
or U11565 (N_11565,N_5709,N_8010);
nand U11566 (N_11566,N_8688,N_5787);
or U11567 (N_11567,N_7527,N_5357);
or U11568 (N_11568,N_8064,N_8573);
nand U11569 (N_11569,N_7980,N_9054);
nand U11570 (N_11570,N_6372,N_6492);
nand U11571 (N_11571,N_9255,N_7333);
and U11572 (N_11572,N_6315,N_8631);
xnor U11573 (N_11573,N_7276,N_8422);
or U11574 (N_11574,N_7585,N_9344);
or U11575 (N_11575,N_8357,N_7721);
or U11576 (N_11576,N_6979,N_9995);
nand U11577 (N_11577,N_7915,N_5999);
nor U11578 (N_11578,N_5343,N_6875);
nand U11579 (N_11579,N_6160,N_7660);
nand U11580 (N_11580,N_8392,N_6061);
nand U11581 (N_11581,N_5401,N_9594);
nand U11582 (N_11582,N_9919,N_7452);
nor U11583 (N_11583,N_8633,N_9916);
nor U11584 (N_11584,N_5617,N_5399);
nand U11585 (N_11585,N_6948,N_5240);
nor U11586 (N_11586,N_6157,N_9548);
nor U11587 (N_11587,N_9531,N_9566);
nand U11588 (N_11588,N_7483,N_9360);
and U11589 (N_11589,N_9644,N_8084);
or U11590 (N_11590,N_6691,N_5047);
xnor U11591 (N_11591,N_7512,N_8264);
nand U11592 (N_11592,N_6852,N_6335);
or U11593 (N_11593,N_9873,N_8468);
or U11594 (N_11594,N_8385,N_6937);
or U11595 (N_11595,N_8272,N_5604);
and U11596 (N_11596,N_5818,N_9443);
nand U11597 (N_11597,N_9491,N_5059);
nand U11598 (N_11598,N_8415,N_6872);
nand U11599 (N_11599,N_5001,N_7929);
xor U11600 (N_11600,N_5590,N_9373);
or U11601 (N_11601,N_6503,N_8584);
nand U11602 (N_11602,N_9643,N_7132);
or U11603 (N_11603,N_7773,N_9260);
xnor U11604 (N_11604,N_5210,N_7283);
or U11605 (N_11605,N_7852,N_8689);
and U11606 (N_11606,N_8597,N_9357);
nand U11607 (N_11607,N_5371,N_7022);
xor U11608 (N_11608,N_7282,N_7664);
and U11609 (N_11609,N_9053,N_5102);
nor U11610 (N_11610,N_9439,N_7501);
xor U11611 (N_11611,N_7441,N_5341);
xor U11612 (N_11612,N_5276,N_9978);
or U11613 (N_11613,N_9454,N_8097);
and U11614 (N_11614,N_6963,N_5644);
or U11615 (N_11615,N_7488,N_8857);
nand U11616 (N_11616,N_9069,N_6743);
xnor U11617 (N_11617,N_5004,N_7445);
nor U11618 (N_11618,N_5325,N_8255);
and U11619 (N_11619,N_5994,N_9692);
nand U11620 (N_11620,N_8562,N_5440);
nand U11621 (N_11621,N_9117,N_8836);
nor U11622 (N_11622,N_5650,N_7113);
or U11623 (N_11623,N_7682,N_6257);
or U11624 (N_11624,N_7130,N_6066);
nor U11625 (N_11625,N_9433,N_6646);
nor U11626 (N_11626,N_5076,N_7617);
nand U11627 (N_11627,N_9668,N_6783);
or U11628 (N_11628,N_9611,N_9356);
nor U11629 (N_11629,N_8333,N_7076);
xnor U11630 (N_11630,N_6799,N_5305);
nor U11631 (N_11631,N_7504,N_6183);
or U11632 (N_11632,N_9723,N_7442);
xor U11633 (N_11633,N_6292,N_8806);
nor U11634 (N_11634,N_8236,N_9434);
or U11635 (N_11635,N_5771,N_5945);
xor U11636 (N_11636,N_5262,N_5534);
xnor U11637 (N_11637,N_7708,N_5136);
or U11638 (N_11638,N_8951,N_9156);
nor U11639 (N_11639,N_8434,N_6726);
and U11640 (N_11640,N_8606,N_7857);
and U11641 (N_11641,N_8844,N_9764);
xnor U11642 (N_11642,N_6662,N_9598);
xnor U11643 (N_11643,N_9112,N_5878);
and U11644 (N_11644,N_5470,N_5040);
or U11645 (N_11645,N_5853,N_9556);
xor U11646 (N_11646,N_7856,N_7872);
xnor U11647 (N_11647,N_6933,N_5398);
xnor U11648 (N_11648,N_8794,N_6265);
or U11649 (N_11649,N_7785,N_8962);
nand U11650 (N_11650,N_8715,N_9472);
xor U11651 (N_11651,N_8537,N_8203);
nand U11652 (N_11652,N_7267,N_7837);
nor U11653 (N_11653,N_6352,N_5619);
nand U11654 (N_11654,N_7906,N_8546);
and U11655 (N_11655,N_7576,N_9638);
xnor U11656 (N_11656,N_8350,N_6736);
xnor U11657 (N_11657,N_5621,N_6853);
nand U11658 (N_11658,N_6592,N_9817);
xnor U11659 (N_11659,N_9950,N_9951);
xor U11660 (N_11660,N_5876,N_6125);
nor U11661 (N_11661,N_6379,N_5519);
nand U11662 (N_11662,N_7644,N_7528);
or U11663 (N_11663,N_5575,N_7584);
and U11664 (N_11664,N_9235,N_7437);
xnor U11665 (N_11665,N_6225,N_9487);
xnor U11666 (N_11666,N_9696,N_6868);
or U11667 (N_11667,N_9808,N_7046);
xnor U11668 (N_11668,N_6561,N_7549);
xnor U11669 (N_11669,N_5437,N_5253);
nor U11670 (N_11670,N_9524,N_9601);
xnor U11671 (N_11671,N_6862,N_5223);
xor U11672 (N_11672,N_5592,N_9940);
or U11673 (N_11673,N_8383,N_7608);
xnor U11674 (N_11674,N_7868,N_7523);
nor U11675 (N_11675,N_7221,N_7789);
xnor U11676 (N_11676,N_5792,N_7828);
xor U11677 (N_11677,N_9944,N_9186);
nor U11678 (N_11678,N_9101,N_5564);
nor U11679 (N_11679,N_5224,N_6708);
or U11680 (N_11680,N_6734,N_7456);
or U11681 (N_11681,N_5831,N_7140);
and U11682 (N_11682,N_7698,N_8315);
or U11683 (N_11683,N_5051,N_6287);
nor U11684 (N_11684,N_7888,N_8879);
xnor U11685 (N_11685,N_7137,N_8911);
nor U11686 (N_11686,N_7497,N_8186);
and U11687 (N_11687,N_9755,N_7436);
nor U11688 (N_11688,N_6796,N_9170);
xnor U11689 (N_11689,N_7047,N_5425);
or U11690 (N_11690,N_6738,N_8831);
nand U11691 (N_11691,N_9779,N_9263);
nor U11692 (N_11692,N_5142,N_7072);
nor U11693 (N_11693,N_9268,N_9004);
nand U11694 (N_11694,N_5345,N_9778);
xnor U11695 (N_11695,N_8601,N_9412);
and U11696 (N_11696,N_9347,N_7026);
xor U11697 (N_11697,N_6136,N_5400);
nand U11698 (N_11698,N_6540,N_6007);
nand U11699 (N_11699,N_8310,N_7538);
and U11700 (N_11700,N_7746,N_5630);
or U11701 (N_11701,N_7690,N_8492);
or U11702 (N_11702,N_5992,N_5137);
and U11703 (N_11703,N_5548,N_5565);
and U11704 (N_11704,N_6709,N_8509);
xor U11705 (N_11705,N_8835,N_6143);
or U11706 (N_11706,N_9480,N_9789);
xor U11707 (N_11707,N_5539,N_6636);
nor U11708 (N_11708,N_5459,N_8593);
xor U11709 (N_11709,N_5407,N_5099);
xor U11710 (N_11710,N_8903,N_5264);
nand U11711 (N_11711,N_9666,N_6818);
nand U11712 (N_11712,N_8945,N_8386);
nand U11713 (N_11713,N_7772,N_9198);
nor U11714 (N_11714,N_9031,N_6680);
and U11715 (N_11715,N_7003,N_7285);
nor U11716 (N_11716,N_6189,N_6850);
nor U11717 (N_11717,N_6137,N_7926);
nand U11718 (N_11718,N_5323,N_8372);
nor U11719 (N_11719,N_5801,N_6167);
xnor U11720 (N_11720,N_7563,N_5354);
nor U11721 (N_11721,N_7728,N_9846);
or U11722 (N_11722,N_7146,N_6874);
nand U11723 (N_11723,N_9230,N_9847);
xnor U11724 (N_11724,N_5019,N_7835);
nand U11725 (N_11725,N_6128,N_7424);
nand U11726 (N_11726,N_8228,N_7742);
nor U11727 (N_11727,N_5797,N_5513);
xnor U11728 (N_11728,N_5396,N_6153);
and U11729 (N_11729,N_7870,N_7815);
and U11730 (N_11730,N_5284,N_5557);
or U11731 (N_11731,N_9075,N_7799);
xor U11732 (N_11732,N_8300,N_5216);
and U11733 (N_11733,N_9705,N_5361);
and U11734 (N_11734,N_9366,N_9607);
nand U11735 (N_11735,N_5857,N_8288);
xnor U11736 (N_11736,N_7160,N_6775);
or U11737 (N_11737,N_6483,N_5612);
or U11738 (N_11738,N_7611,N_5318);
nor U11739 (N_11739,N_5842,N_5220);
and U11740 (N_11740,N_9999,N_5613);
nand U11741 (N_11741,N_7171,N_9510);
nor U11742 (N_11742,N_5337,N_6990);
nor U11743 (N_11743,N_6240,N_7369);
nor U11744 (N_11744,N_8192,N_7666);
and U11745 (N_11745,N_6209,N_9509);
xor U11746 (N_11746,N_6586,N_8523);
nand U11747 (N_11747,N_7726,N_9952);
nand U11748 (N_11748,N_7637,N_5456);
and U11749 (N_11749,N_9307,N_5307);
nand U11750 (N_11750,N_5053,N_6149);
or U11751 (N_11751,N_6918,N_6692);
xnor U11752 (N_11752,N_9382,N_8116);
xnor U11753 (N_11753,N_5786,N_6891);
and U11754 (N_11754,N_9658,N_5980);
and U11755 (N_11755,N_9508,N_6964);
xor U11756 (N_11756,N_8557,N_7308);
nand U11757 (N_11757,N_5679,N_9678);
xnor U11758 (N_11758,N_5973,N_9164);
or U11759 (N_11759,N_5934,N_8841);
xnor U11760 (N_11760,N_8289,N_6174);
nor U11761 (N_11761,N_6836,N_5691);
xor U11762 (N_11762,N_5431,N_7874);
nand U11763 (N_11763,N_8393,N_8598);
nand U11764 (N_11764,N_9007,N_9282);
xnor U11765 (N_11765,N_7725,N_9422);
or U11766 (N_11766,N_5027,N_5362);
and U11767 (N_11767,N_7902,N_8759);
xor U11768 (N_11768,N_6369,N_7443);
nor U11769 (N_11769,N_9279,N_5083);
nand U11770 (N_11770,N_7643,N_9206);
and U11771 (N_11771,N_6057,N_8353);
xor U11772 (N_11772,N_9570,N_8944);
and U11773 (N_11773,N_9657,N_7100);
xor U11774 (N_11774,N_7387,N_5703);
or U11775 (N_11775,N_8666,N_9552);
and U11776 (N_11776,N_8472,N_5260);
nand U11777 (N_11777,N_9097,N_7485);
and U11778 (N_11778,N_5753,N_5815);
nand U11779 (N_11779,N_5115,N_9991);
nor U11780 (N_11780,N_6721,N_6530);
and U11781 (N_11781,N_5593,N_9630);
nand U11782 (N_11782,N_8028,N_8096);
nor U11783 (N_11783,N_8924,N_9435);
nand U11784 (N_11784,N_6641,N_7873);
or U11785 (N_11785,N_9810,N_8530);
nor U11786 (N_11786,N_5900,N_8730);
nor U11787 (N_11787,N_6428,N_8871);
nand U11788 (N_11788,N_8366,N_8194);
xor U11789 (N_11789,N_8744,N_8916);
and U11790 (N_11790,N_5048,N_7560);
nand U11791 (N_11791,N_8048,N_5697);
and U11792 (N_11792,N_8110,N_8156);
or U11793 (N_11793,N_6898,N_9904);
nor U11794 (N_11794,N_9650,N_7184);
or U11795 (N_11795,N_5447,N_6637);
nand U11796 (N_11796,N_5799,N_6822);
nor U11797 (N_11797,N_8721,N_8453);
nor U11798 (N_11798,N_5601,N_6667);
or U11799 (N_11799,N_9842,N_7345);
or U11800 (N_11800,N_7787,N_6259);
nor U11801 (N_11801,N_9684,N_6987);
xor U11802 (N_11802,N_9640,N_8364);
nand U11803 (N_11803,N_9567,N_7676);
or U11804 (N_11804,N_8554,N_5199);
or U11805 (N_11805,N_9458,N_8085);
xnor U11806 (N_11806,N_6132,N_6020);
nand U11807 (N_11807,N_6865,N_5073);
and U11808 (N_11808,N_7188,N_5922);
xnor U11809 (N_11809,N_5578,N_8000);
and U11810 (N_11810,N_6210,N_5077);
nand U11811 (N_11811,N_8622,N_7105);
nor U11812 (N_11812,N_8579,N_9990);
nor U11813 (N_11813,N_5780,N_7779);
or U11814 (N_11814,N_8349,N_9739);
and U11815 (N_11815,N_6328,N_9943);
nor U11816 (N_11816,N_8046,N_8884);
and U11817 (N_11817,N_5626,N_5881);
nand U11818 (N_11818,N_7777,N_8146);
and U11819 (N_11819,N_7217,N_7396);
nor U11820 (N_11820,N_8513,N_5329);
nand U11821 (N_11821,N_7379,N_7304);
nand U11822 (N_11822,N_6418,N_9709);
xnor U11823 (N_11823,N_5726,N_8317);
and U11824 (N_11824,N_5421,N_7529);
nor U11825 (N_11825,N_8629,N_8456);
and U11826 (N_11826,N_8981,N_5275);
nor U11827 (N_11827,N_9798,N_5988);
nor U11828 (N_11828,N_5080,N_6934);
or U11829 (N_11829,N_9595,N_7469);
nor U11830 (N_11830,N_7569,N_5959);
and U11831 (N_11831,N_6513,N_5113);
xor U11832 (N_11832,N_8191,N_9121);
nor U11833 (N_11833,N_6706,N_6685);
nand U11834 (N_11834,N_8979,N_7383);
and U11835 (N_11835,N_8649,N_9030);
nor U11836 (N_11836,N_6541,N_7054);
xnor U11837 (N_11837,N_7057,N_9252);
nand U11838 (N_11838,N_5708,N_5458);
nand U11839 (N_11839,N_5871,N_9358);
or U11840 (N_11840,N_6396,N_6390);
or U11841 (N_11841,N_5050,N_5566);
or U11842 (N_11842,N_6642,N_8906);
xor U11843 (N_11843,N_9427,N_6622);
xnor U11844 (N_11844,N_8328,N_9878);
xnor U11845 (N_11845,N_9867,N_6427);
and U11846 (N_11846,N_5914,N_7935);
or U11847 (N_11847,N_7206,N_6441);
nor U11848 (N_11848,N_7473,N_7062);
nand U11849 (N_11849,N_6139,N_5957);
and U11850 (N_11850,N_7017,N_5952);
nor U11851 (N_11851,N_7524,N_9704);
xnor U11852 (N_11852,N_7975,N_9420);
and U11853 (N_11853,N_5633,N_5383);
nand U11854 (N_11854,N_8811,N_6785);
xor U11855 (N_11855,N_9841,N_8737);
or U11856 (N_11856,N_6385,N_5331);
or U11857 (N_11857,N_9174,N_8252);
nor U11858 (N_11858,N_8921,N_6920);
or U11859 (N_11859,N_8661,N_8891);
nor U11860 (N_11860,N_9027,N_9642);
xor U11861 (N_11861,N_7476,N_8679);
xnor U11862 (N_11862,N_9079,N_6479);
nor U11863 (N_11863,N_6095,N_7165);
nand U11864 (N_11864,N_9372,N_9870);
and U11865 (N_11865,N_7287,N_9561);
nand U11866 (N_11866,N_9017,N_5724);
nor U11867 (N_11867,N_5523,N_8119);
nor U11868 (N_11868,N_8135,N_5176);
and U11869 (N_11869,N_7593,N_8089);
and U11870 (N_11870,N_7300,N_9963);
or U11871 (N_11871,N_9672,N_9962);
or U11872 (N_11872,N_8269,N_5783);
xnor U11873 (N_11873,N_8273,N_9610);
nor U11874 (N_11874,N_9006,N_8615);
nor U11875 (N_11875,N_9497,N_7125);
and U11876 (N_11876,N_7429,N_5380);
and U11877 (N_11877,N_9649,N_7353);
xor U11878 (N_11878,N_9409,N_8232);
nor U11879 (N_11879,N_7239,N_7597);
and U11880 (N_11880,N_5614,N_6629);
and U11881 (N_11881,N_9742,N_5964);
nor U11882 (N_11882,N_7859,N_9025);
or U11883 (N_11883,N_9785,N_8756);
and U11884 (N_11884,N_6488,N_7292);
and U11885 (N_11885,N_6178,N_9939);
and U11886 (N_11886,N_5285,N_7482);
or U11887 (N_11887,N_8319,N_8050);
or U11888 (N_11888,N_7356,N_5292);
nand U11889 (N_11889,N_8435,N_6051);
xor U11890 (N_11890,N_7669,N_7111);
nor U11891 (N_11891,N_9065,N_7649);
nor U11892 (N_11892,N_5804,N_9135);
xnor U11893 (N_11893,N_5415,N_6044);
or U11894 (N_11894,N_6016,N_6831);
nor U11895 (N_11895,N_8150,N_7247);
nand U11896 (N_11896,N_8813,N_8893);
nor U11897 (N_11897,N_6854,N_6902);
xnor U11898 (N_11898,N_9324,N_6099);
nand U11899 (N_11899,N_7228,N_6715);
nor U11900 (N_11900,N_9302,N_7595);
or U11901 (N_11901,N_9284,N_8459);
nor U11902 (N_11902,N_9813,N_7172);
or U11903 (N_11903,N_5836,N_5742);
xnor U11904 (N_11904,N_7977,N_5030);
nor U11905 (N_11905,N_9456,N_6021);
nand U11906 (N_11906,N_6856,N_8753);
nand U11907 (N_11907,N_8580,N_6593);
xnor U11908 (N_11908,N_5499,N_6926);
and U11909 (N_11909,N_6921,N_6038);
or U11910 (N_11910,N_7910,N_9137);
xor U11911 (N_11911,N_8684,N_9826);
xor U11912 (N_11912,N_6048,N_6781);
nor U11913 (N_11913,N_9399,N_8009);
nand U11914 (N_11914,N_8522,N_5057);
nand U11915 (N_11915,N_8874,N_6423);
nor U11916 (N_11916,N_9038,N_8125);
xor U11917 (N_11917,N_6884,N_5844);
nor U11918 (N_11918,N_9834,N_8755);
or U11919 (N_11919,N_5643,N_9818);
nor U11920 (N_11920,N_7200,N_9147);
nor U11921 (N_11921,N_7346,N_5066);
or U11922 (N_11922,N_8611,N_7820);
or U11923 (N_11923,N_6242,N_7568);
xnor U11924 (N_11924,N_9969,N_7696);
xor U11925 (N_11925,N_6938,N_6879);
or U11926 (N_11926,N_5546,N_9920);
xnor U11927 (N_11927,N_6465,N_8519);
and U11928 (N_11928,N_5081,N_5413);
and U11929 (N_11929,N_8428,N_9683);
xnor U11930 (N_11930,N_6840,N_7616);
or U11931 (N_11931,N_5278,N_8245);
nand U11932 (N_11932,N_5943,N_6071);
nand U11933 (N_11933,N_6714,N_9457);
and U11934 (N_11934,N_7864,N_8002);
nor U11935 (N_11935,N_5885,N_6543);
nor U11936 (N_11936,N_5089,N_5488);
nor U11937 (N_11937,N_9190,N_7243);
or U11938 (N_11938,N_6679,N_9854);
xor U11939 (N_11939,N_5054,N_9897);
and U11940 (N_11940,N_5750,N_6078);
nand U11941 (N_11941,N_7224,N_8019);
nor U11942 (N_11942,N_9430,N_7134);
nand U11943 (N_11943,N_8819,N_6312);
nor U11944 (N_11944,N_8642,N_6074);
xnor U11945 (N_11945,N_5711,N_7526);
xor U11946 (N_11946,N_8749,N_6748);
and U11947 (N_11947,N_7071,N_8036);
nor U11948 (N_11948,N_7688,N_9534);
or U11949 (N_11949,N_8992,N_7407);
xor U11950 (N_11950,N_8148,N_9587);
or U11951 (N_11951,N_5046,N_9735);
nor U11952 (N_11952,N_7451,N_7271);
or U11953 (N_11953,N_5695,N_9192);
nor U11954 (N_11954,N_5788,N_7891);
nor U11955 (N_11955,N_7842,N_8899);
nand U11956 (N_11956,N_5896,N_6303);
xnor U11957 (N_11957,N_8368,N_9408);
and U11958 (N_11958,N_9553,N_9653);
or U11959 (N_11959,N_5658,N_7235);
nand U11960 (N_11960,N_5390,N_9165);
nand U11961 (N_11961,N_6033,N_8388);
nor U11962 (N_11962,N_5495,N_8184);
nor U11963 (N_11963,N_8113,N_6486);
nor U11964 (N_11964,N_8637,N_6658);
and U11965 (N_11965,N_9258,N_8401);
nand U11966 (N_11966,N_8003,N_9582);
nor U11967 (N_11967,N_6537,N_5496);
or U11968 (N_11968,N_5976,N_9061);
nand U11969 (N_11969,N_7778,N_5212);
nor U11970 (N_11970,N_6925,N_6980);
nand U11971 (N_11971,N_9314,N_6285);
and U11972 (N_11972,N_5756,N_9276);
nor U11973 (N_11973,N_9144,N_5913);
nand U11974 (N_11974,N_7176,N_6321);
xor U11975 (N_11975,N_9659,N_8558);
or U11976 (N_11976,N_6766,N_5926);
xnor U11977 (N_11977,N_9797,N_6701);
nor U11978 (N_11978,N_5000,N_6081);
or U11979 (N_11979,N_9043,N_7691);
nand U11980 (N_11980,N_5866,N_6791);
nand U11981 (N_11981,N_8971,N_6034);
nand U11982 (N_11982,N_6416,N_5229);
and U11983 (N_11983,N_7624,N_9217);
and U11984 (N_11984,N_6939,N_8016);
nand U11985 (N_11985,N_6717,N_5246);
xor U11986 (N_11986,N_6347,N_6084);
or U11987 (N_11987,N_9210,N_5062);
or U11988 (N_11988,N_7163,N_8179);
xor U11989 (N_11989,N_8173,N_9289);
and U11990 (N_11990,N_6329,N_7392);
nor U11991 (N_11991,N_9581,N_7988);
nor U11992 (N_11992,N_6827,N_9158);
and U11993 (N_11993,N_7522,N_5211);
and U11994 (N_11994,N_5846,N_8039);
and U11995 (N_11995,N_8966,N_7349);
nand U11996 (N_11996,N_7886,N_7791);
nor U11997 (N_11997,N_6458,N_9540);
and U11998 (N_11998,N_6373,N_6219);
nor U11999 (N_11999,N_6657,N_5085);
nor U12000 (N_12000,N_5577,N_6410);
nand U12001 (N_12001,N_7763,N_8796);
or U12002 (N_12002,N_5011,N_9384);
xor U12003 (N_12003,N_7653,N_5935);
xnor U12004 (N_12004,N_6213,N_7577);
nor U12005 (N_12005,N_8182,N_9336);
nor U12006 (N_12006,N_8027,N_9131);
nor U12007 (N_12007,N_7673,N_7762);
nand U12008 (N_12008,N_6863,N_5512);
and U12009 (N_12009,N_7905,N_8917);
xor U12010 (N_12010,N_7602,N_6526);
nand U12011 (N_12011,N_7752,N_7297);
nand U12012 (N_12012,N_7566,N_6686);
nor U12013 (N_12013,N_8170,N_7656);
xnor U12014 (N_12014,N_8829,N_8798);
nand U12015 (N_12015,N_6788,N_6124);
nor U12016 (N_12016,N_9606,N_6156);
nor U12017 (N_12017,N_6581,N_9734);
nand U12018 (N_12018,N_9349,N_5036);
nand U12019 (N_12019,N_9998,N_8888);
nand U12020 (N_12020,N_5141,N_9494);
nand U12021 (N_12021,N_8732,N_6842);
nand U12022 (N_12022,N_7920,N_8081);
nor U12023 (N_12023,N_6534,N_7233);
and U12024 (N_12024,N_5580,N_9415);
or U12025 (N_12025,N_6696,N_5105);
nand U12026 (N_12026,N_6417,N_8936);
nand U12027 (N_12027,N_8280,N_9188);
nand U12028 (N_12028,N_9049,N_5997);
xnor U12029 (N_12029,N_7948,N_9928);
nand U12030 (N_12030,N_7180,N_7539);
xnor U12031 (N_12031,N_8091,N_8869);
xor U12032 (N_12032,N_8162,N_8480);
nand U12033 (N_12033,N_6695,N_9527);
nand U12034 (N_12034,N_7466,N_5861);
or U12035 (N_12035,N_9767,N_9355);
nand U12036 (N_12036,N_6130,N_6298);
or U12037 (N_12037,N_7936,N_8931);
xnor U12038 (N_12038,N_5993,N_7019);
nor U12039 (N_12039,N_5757,N_6924);
xnor U12040 (N_12040,N_6249,N_9272);
nor U12041 (N_12041,N_9876,N_7016);
nand U12042 (N_12042,N_5295,N_8105);
or U12043 (N_12043,N_5687,N_5761);
nand U12044 (N_12044,N_8106,N_5152);
nor U12045 (N_12045,N_7104,N_6116);
and U12046 (N_12046,N_9126,N_5874);
xor U12047 (N_12047,N_7738,N_5507);
xnor U12048 (N_12048,N_6318,N_9359);
or U12049 (N_12049,N_9654,N_8482);
nand U12050 (N_12050,N_5903,N_7306);
nand U12051 (N_12051,N_9278,N_6560);
and U12052 (N_12052,N_6882,N_6229);
nor U12053 (N_12053,N_6484,N_8655);
nand U12054 (N_12054,N_7145,N_8160);
and U12055 (N_12055,N_9693,N_8703);
nor U12056 (N_12056,N_6562,N_6239);
or U12057 (N_12057,N_8083,N_8251);
xnor U12058 (N_12058,N_7832,N_7588);
and U12059 (N_12059,N_8496,N_7548);
nor U12060 (N_12060,N_6628,N_9513);
xnor U12061 (N_12061,N_9559,N_9976);
xnor U12062 (N_12062,N_8278,N_8625);
nor U12063 (N_12063,N_5301,N_5813);
or U12064 (N_12064,N_9304,N_8431);
nor U12065 (N_12065,N_5701,N_7622);
and U12066 (N_12066,N_9829,N_7339);
xor U12067 (N_12067,N_7248,N_9647);
nand U12068 (N_12068,N_6574,N_8669);
nand U12069 (N_12069,N_6274,N_6498);
nand U12070 (N_12070,N_5916,N_6333);
xor U12071 (N_12071,N_5443,N_8635);
xor U12072 (N_12072,N_9994,N_8646);
nand U12073 (N_12073,N_6760,N_8774);
nand U12074 (N_12074,N_6564,N_5721);
xor U12075 (N_12075,N_8414,N_6169);
and U12076 (N_12076,N_5915,N_9837);
and U12077 (N_12077,N_5558,N_9462);
nand U12078 (N_12078,N_7745,N_7513);
nor U12079 (N_12079,N_9421,N_5237);
or U12080 (N_12080,N_9980,N_7976);
xor U12081 (N_12081,N_9868,N_7583);
and U12082 (N_12082,N_8277,N_6808);
or U12083 (N_12083,N_9651,N_8297);
nor U12084 (N_12084,N_9946,N_7657);
nand U12085 (N_12085,N_9380,N_9127);
and U12086 (N_12086,N_9856,N_5731);
xor U12087 (N_12087,N_7919,N_8982);
or U12088 (N_12088,N_6787,N_6830);
nor U12089 (N_12089,N_8955,N_7077);
xnor U12090 (N_12090,N_9115,N_6644);
nor U12091 (N_12091,N_6909,N_7684);
xnor U12092 (N_12092,N_7500,N_9850);
nor U12093 (N_12093,N_6028,N_7641);
xor U12094 (N_12094,N_8989,N_8676);
nor U12095 (N_12095,N_6358,N_5538);
nand U12096 (N_12096,N_9400,N_5155);
or U12097 (N_12097,N_7389,N_7836);
nand U12098 (N_12098,N_7764,N_6624);
and U12099 (N_12099,N_9664,N_8757);
xor U12100 (N_12100,N_8785,N_8311);
nand U12101 (N_12101,N_5735,N_8166);
or U12102 (N_12102,N_8722,N_5562);
nand U12103 (N_12103,N_9631,N_7956);
nand U12104 (N_12104,N_7724,N_5700);
or U12105 (N_12105,N_7086,N_7432);
nand U12106 (N_12106,N_5587,N_9686);
nor U12107 (N_12107,N_9345,N_7811);
or U12108 (N_12108,N_8316,N_9589);
nand U12109 (N_12109,N_6103,N_7612);
or U12110 (N_12110,N_5764,N_6719);
nor U12111 (N_12111,N_9860,N_7550);
xnor U12112 (N_12112,N_5016,N_6472);
xor U12113 (N_12113,N_9195,N_8354);
xor U12114 (N_12114,N_7514,N_7829);
xnor U12115 (N_12115,N_7314,N_6022);
nor U12116 (N_12116,N_7565,N_5659);
or U12117 (N_12117,N_9199,N_9021);
nand U12118 (N_12118,N_9564,N_9612);
nand U12119 (N_12119,N_6327,N_9563);
or U12120 (N_12120,N_5979,N_5314);
xor U12121 (N_12121,N_7028,N_9840);
or U12122 (N_12122,N_7599,N_8365);
or U12123 (N_12123,N_6864,N_7559);
xor U12124 (N_12124,N_9362,N_6467);
nand U12125 (N_12125,N_6039,N_9339);
xor U12126 (N_12126,N_7844,N_6338);
nand U12127 (N_12127,N_9015,N_5910);
xnor U12128 (N_12128,N_7596,N_8249);
xnor U12129 (N_12129,N_6152,N_6625);
or U12130 (N_12130,N_5420,N_8671);
or U12131 (N_12131,N_8185,N_5131);
and U12132 (N_12132,N_8025,N_8618);
nor U12133 (N_12133,N_5033,N_9495);
nor U12134 (N_12134,N_7718,N_6388);
or U12135 (N_12135,N_9716,N_9903);
nand U12136 (N_12136,N_9107,N_9150);
nand U12137 (N_12137,N_5268,N_6470);
nand U12138 (N_12138,N_5858,N_6214);
nor U12139 (N_12139,N_7434,N_5409);
nor U12140 (N_12140,N_5637,N_7917);
or U12141 (N_12141,N_5439,N_5111);
and U12142 (N_12142,N_5704,N_8746);
and U12143 (N_12143,N_8619,N_6121);
xor U12144 (N_12144,N_5902,N_6974);
xor U12145 (N_12145,N_8733,N_7431);
xnor U12146 (N_12146,N_5242,N_9788);
xnor U12147 (N_12147,N_7782,N_9748);
xor U12148 (N_12148,N_9915,N_8953);
nor U12149 (N_12149,N_8127,N_7049);
and U12150 (N_12150,N_8702,N_9333);
and U12151 (N_12151,N_6192,N_9002);
xor U12152 (N_12152,N_5072,N_8581);
nand U12153 (N_12153,N_5816,N_6146);
nor U12154 (N_12154,N_8263,N_7386);
nand U12155 (N_12155,N_8161,N_9728);
nor U12156 (N_12156,N_8421,N_6638);
and U12157 (N_12157,N_8640,N_5037);
xor U12158 (N_12158,N_6813,N_5807);
or U12159 (N_12159,N_5315,N_8600);
or U12160 (N_12160,N_6374,N_9893);
nor U12161 (N_12161,N_6277,N_8450);
nand U12162 (N_12162,N_6929,N_8591);
or U12163 (N_12163,N_7994,N_8209);
nor U12164 (N_12164,N_9663,N_6599);
nor U12165 (N_12165,N_6011,N_8069);
nand U12166 (N_12166,N_8486,N_6079);
xor U12167 (N_12167,N_7480,N_8052);
or U12168 (N_12168,N_9694,N_5624);
xor U12169 (N_12169,N_9722,N_8786);
and U12170 (N_12170,N_6260,N_5101);
xnor U12171 (N_12171,N_9386,N_8867);
or U12172 (N_12172,N_8111,N_5610);
xor U12173 (N_12173,N_7861,N_6812);
nand U12174 (N_12174,N_9193,N_9058);
xor U12175 (N_12175,N_9118,N_8375);
nor U12176 (N_12176,N_7982,N_8014);
or U12177 (N_12177,N_9747,N_9586);
nor U12178 (N_12178,N_6459,N_7091);
or U12179 (N_12179,N_5140,N_8205);
nand U12180 (N_12180,N_9875,N_6466);
nor U12181 (N_12181,N_5123,N_6023);
or U12182 (N_12182,N_9138,N_6797);
xnor U12183 (N_12183,N_5549,N_9937);
nand U12184 (N_12184,N_6331,N_8011);
and U12185 (N_12185,N_8188,N_6145);
or U12186 (N_12186,N_7454,N_5718);
xor U12187 (N_12187,N_6826,N_6097);
and U12188 (N_12188,N_5699,N_6857);
or U12189 (N_12189,N_7536,N_5207);
xnor U12190 (N_12190,N_9023,N_8731);
nand U12191 (N_12191,N_9124,N_5049);
and U12192 (N_12192,N_7360,N_5065);
or U12193 (N_12193,N_7734,N_9123);
nand U12194 (N_12194,N_8604,N_5411);
nor U12195 (N_12195,N_6912,N_7411);
or U12196 (N_12196,N_8452,N_7471);
nand U12197 (N_12197,N_7723,N_8335);
nand U12198 (N_12198,N_6539,N_7750);
and U12199 (N_12199,N_9884,N_7958);
nand U12200 (N_12200,N_5274,N_5154);
nor U12201 (N_12201,N_9184,N_8638);
and U12202 (N_12202,N_9159,N_6027);
xor U12203 (N_12203,N_6226,N_8293);
xnor U12204 (N_12204,N_8478,N_5516);
xnor U12205 (N_12205,N_7069,N_9910);
and U12206 (N_12206,N_9189,N_8761);
and U12207 (N_12207,N_7765,N_8910);
or U12208 (N_12208,N_8551,N_9988);
nor U12209 (N_12209,N_7555,N_6514);
nand U12210 (N_12210,N_6468,N_9477);
xor U12211 (N_12211,N_6102,N_8764);
or U12212 (N_12212,N_7879,N_9087);
nand U12213 (N_12213,N_9762,N_6649);
and U12214 (N_12214,N_8198,N_6915);
and U12215 (N_12215,N_8078,N_7102);
and U12216 (N_12216,N_7519,N_8498);
xnor U12217 (N_12217,N_6300,N_5178);
nor U12218 (N_12218,N_8237,N_7114);
xor U12219 (N_12219,N_8066,N_5684);
nor U12220 (N_12220,N_7290,N_8998);
or U12221 (N_12221,N_5591,N_9459);
or U12222 (N_12222,N_6878,N_5180);
nand U12223 (N_12223,N_9661,N_8030);
and U12224 (N_12224,N_8510,N_8743);
or U12225 (N_12225,N_9918,N_5163);
xor U12226 (N_12226,N_8892,N_5338);
and U12227 (N_12227,N_5296,N_6383);
and U12228 (N_12228,N_5982,N_8059);
nor U12229 (N_12229,N_9699,N_8343);
nor U12230 (N_12230,N_9772,N_5517);
nor U12231 (N_12231,N_7802,N_6619);
nor U12232 (N_12232,N_5710,N_6173);
and U12233 (N_12233,N_8856,N_8457);
nor U12234 (N_12234,N_8301,N_9981);
nor U12235 (N_12235,N_5302,N_6366);
xnor U12236 (N_12236,N_8122,N_7521);
nand U12237 (N_12237,N_5068,N_9889);
or U12238 (N_12238,N_5769,N_7138);
nand U12239 (N_12239,N_5739,N_6282);
or U12240 (N_12240,N_5839,N_8380);
and U12241 (N_12241,N_6253,N_5918);
xor U12242 (N_12242,N_9142,N_9670);
nor U12243 (N_12243,N_7135,N_5856);
xnor U12244 (N_12244,N_7570,N_9187);
or U12245 (N_12245,N_5128,N_6205);
nor U12246 (N_12246,N_7737,N_6681);
or U12247 (N_12247,N_6652,N_9243);
nor U12248 (N_12248,N_6435,N_7095);
and U12249 (N_12249,N_5545,N_7520);
nand U12250 (N_12250,N_5795,N_8687);
nand U12251 (N_12251,N_8847,N_7229);
or U12252 (N_12252,N_5355,N_8015);
xnor U12253 (N_12253,N_7573,N_6727);
and U12254 (N_12254,N_5023,N_5553);
or U12255 (N_12255,N_6579,N_7464);
and U12256 (N_12256,N_8058,N_5625);
or U12257 (N_12257,N_6087,N_7278);
or U12258 (N_12258,N_9865,N_5263);
xor U12259 (N_12259,N_9197,N_7225);
and U12260 (N_12260,N_9585,N_6616);
or U12261 (N_12261,N_8501,N_8024);
xnor U12262 (N_12262,N_7341,N_5823);
nor U12263 (N_12263,N_9108,N_8238);
nand U12264 (N_12264,N_7629,N_6568);
xor U12265 (N_12265,N_6669,N_9139);
nor U12266 (N_12266,N_8605,N_5563);
xor U12267 (N_12267,N_9406,N_8849);
xnor U12268 (N_12268,N_7254,N_7591);
xnor U12269 (N_12269,N_8243,N_5719);
and U12270 (N_12270,N_6401,N_6070);
nor U12271 (N_12271,N_8751,N_6956);
xnor U12272 (N_12272,N_7421,N_8719);
or U12273 (N_12273,N_7116,N_9632);
and U12274 (N_12274,N_9740,N_6343);
xor U12275 (N_12275,N_6487,N_6782);
xor U12276 (N_12276,N_6761,N_7810);
nand U12277 (N_12277,N_6535,N_7403);
nor U12278 (N_12278,N_9099,N_7824);
and U12279 (N_12279,N_8075,N_6981);
nor U12280 (N_12280,N_8463,N_5279);
or U12281 (N_12281,N_5490,N_5729);
nand U12282 (N_12282,N_9162,N_5041);
nand U12283 (N_12283,N_7215,N_8996);
and U12284 (N_12284,N_9354,N_9671);
nor U12285 (N_12285,N_8975,N_5556);
nor U12286 (N_12286,N_5629,N_8134);
nor U12287 (N_12287,N_6404,N_8531);
and U12288 (N_12288,N_6502,N_9450);
and U12289 (N_12289,N_5466,N_6105);
and U12290 (N_12290,N_5802,N_5953);
and U12291 (N_12291,N_9018,N_8950);
xnor U12292 (N_12292,N_9299,N_6521);
nand U12293 (N_12293,N_7303,N_5540);
xnor U12294 (N_12294,N_9775,N_7989);
xnor U12295 (N_12295,N_7196,N_9180);
nor U12296 (N_12296,N_8218,N_9822);
and U12297 (N_12297,N_5882,N_5435);
nand U12298 (N_12298,N_6745,N_9804);
and U12299 (N_12299,N_5642,N_9119);
xor U12300 (N_12300,N_8818,N_7927);
nor U12301 (N_12301,N_5479,N_8312);
nand U12302 (N_12302,N_9081,N_6794);
nor U12303 (N_12303,N_6817,N_9200);
or U12304 (N_12304,N_8504,N_5907);
nor U12305 (N_12305,N_6613,N_6010);
nand U12306 (N_12306,N_6751,N_6569);
or U12307 (N_12307,N_5086,N_7186);
or U12308 (N_12308,N_8952,N_8363);
or U12309 (N_12309,N_5094,N_7064);
nor U12310 (N_12310,N_7343,N_5944);
nand U12311 (N_12311,N_7366,N_9033);
or U12312 (N_12312,N_9550,N_7499);
and U12313 (N_12313,N_6222,N_9014);
and U12314 (N_12314,N_6877,N_9024);
xnor U12315 (N_12315,N_9010,N_9765);
nand U12316 (N_12316,N_5873,N_7537);
nor U12317 (N_12317,N_5265,N_8285);
xnor U12318 (N_12318,N_7610,N_9071);
and U12319 (N_12319,N_7827,N_7553);
and U12320 (N_12320,N_5387,N_5018);
and U12321 (N_12321,N_6261,N_6473);
xnor U12322 (N_12322,N_5133,N_9501);
xnor U12323 (N_12323,N_6126,N_9295);
nand U12324 (N_12324,N_6447,N_7240);
nand U12325 (N_12325,N_7911,N_5963);
and U12326 (N_12326,N_5238,N_9003);
nand U12327 (N_12327,N_9923,N_5608);
nand U12328 (N_12328,N_5313,N_6683);
or U12329 (N_12329,N_7679,N_8801);
nand U12330 (N_12330,N_6129,N_8516);
and U12331 (N_12331,N_9698,N_6026);
or U12332 (N_12332,N_8087,N_9806);
and U12333 (N_12333,N_7374,N_7078);
xnor U12334 (N_12334,N_9269,N_9505);
nand U12335 (N_12335,N_9525,N_5043);
nand U12336 (N_12336,N_5967,N_8409);
and U12337 (N_12337,N_6529,N_7209);
nand U12338 (N_12338,N_7655,N_8390);
nor U12339 (N_12339,N_6828,N_7082);
and U12340 (N_12340,N_9925,N_5890);
nor U12341 (N_12341,N_7822,N_9402);
nor U12342 (N_12342,N_9194,N_5785);
and U12343 (N_12343,N_7093,N_5908);
and U12344 (N_12344,N_9035,N_9934);
nand U12345 (N_12345,N_6236,N_5849);
nand U12346 (N_12346,N_9682,N_5351);
nand U12347 (N_12347,N_9542,N_7446);
nor U12348 (N_12348,N_5843,N_9129);
and U12349 (N_12349,N_7581,N_6995);
or U12350 (N_12350,N_8332,N_6778);
nor U12351 (N_12351,N_7404,N_8663);
and U12352 (N_12352,N_7409,N_7468);
xnor U12353 (N_12353,N_7531,N_9756);
and U12354 (N_12354,N_5322,N_7358);
and U12355 (N_12355,N_5214,N_6053);
nand U12356 (N_12356,N_5328,N_8626);
or U12357 (N_12357,N_6525,N_5451);
or U12358 (N_12358,N_9338,N_5228);
nand U12359 (N_12359,N_9641,N_6082);
nand U12360 (N_12360,N_6583,N_8101);
or U12361 (N_12361,N_8970,N_5032);
xnor U12362 (N_12362,N_9833,N_6469);
or U12363 (N_12363,N_9466,N_6392);
nand U12364 (N_12364,N_8609,N_9738);
or U12365 (N_12365,N_5707,N_7703);
and U12366 (N_12366,N_5186,N_6650);
nand U12367 (N_12367,N_5244,N_8485);
xnor U12368 (N_12368,N_6115,N_6859);
nand U12369 (N_12369,N_5668,N_5303);
nand U12370 (N_12370,N_7123,N_5636);
nand U12371 (N_12371,N_7458,N_8429);
nand U12372 (N_12372,N_5656,N_6786);
or U12373 (N_12373,N_8938,N_8330);
nor U12374 (N_12374,N_7996,N_5462);
and U12375 (N_12375,N_6880,N_6630);
nor U12376 (N_12376,N_6916,N_6660);
or U12377 (N_12377,N_8502,N_9102);
nand U12378 (N_12378,N_8694,N_5429);
xnor U12379 (N_12379,N_9280,N_9346);
and U12380 (N_12380,N_7759,N_5872);
nor U12381 (N_12381,N_5448,N_7784);
nand U12382 (N_12382,N_7326,N_9733);
nand U12383 (N_12383,N_9615,N_8080);
and U12384 (N_12384,N_7294,N_7156);
nor U12385 (N_12385,N_8877,N_9530);
nand U12386 (N_12386,N_9078,N_5125);
and U12387 (N_12387,N_7368,N_9635);
nand U12388 (N_12388,N_7035,N_8154);
or U12389 (N_12389,N_5410,N_9103);
or U12390 (N_12390,N_6378,N_5602);
nand U12391 (N_12391,N_9986,N_8171);
nand U12392 (N_12392,N_9815,N_9844);
xnor U12393 (N_12393,N_5144,N_5286);
nand U12394 (N_12394,N_8405,N_6890);
and U12395 (N_12395,N_5828,N_7423);
xnor U12396 (N_12396,N_6983,N_7997);
or U12397 (N_12397,N_7751,N_7508);
or U12398 (N_12398,N_9228,N_8140);
xor U12399 (N_12399,N_9968,N_5789);
nor U12400 (N_12400,N_5311,N_8446);
and U12401 (N_12401,N_9719,N_5339);
or U12402 (N_12402,N_8206,N_7122);
xnor U12403 (N_12403,N_5450,N_8843);
or U12404 (N_12404,N_7380,N_5255);
or U12405 (N_12405,N_8133,N_6100);
nand U12406 (N_12406,N_6158,N_5748);
and U12407 (N_12407,N_8797,N_7219);
xor U12408 (N_12408,N_5734,N_9227);
nor U12409 (N_12409,N_8244,N_7744);
nor U12410 (N_12410,N_9591,N_6202);
xnor U12411 (N_12411,N_7535,N_6825);
and U12412 (N_12412,N_9068,N_9744);
xnor U12413 (N_12413,N_5412,N_5232);
nand U12414 (N_12414,N_5156,N_8670);
nand U12415 (N_12415,N_6421,N_5850);
or U12416 (N_12416,N_6512,N_8887);
or U12417 (N_12417,N_7883,N_6905);
or U12418 (N_12418,N_9281,N_7058);
xnor U12419 (N_12419,N_7702,N_7261);
nor U12420 (N_12420,N_5324,N_9404);
xnor U12421 (N_12421,N_7567,N_9576);
and U12422 (N_12422,N_7496,N_6014);
and U12423 (N_12423,N_8742,N_7484);
nor U12424 (N_12424,N_6493,N_5848);
nor U12425 (N_12425,N_6871,N_8603);
nor U12426 (N_12426,N_6420,N_7166);
or U12427 (N_12427,N_8329,N_8674);
nand U12428 (N_12428,N_8226,N_9896);
xnor U12429 (N_12429,N_7388,N_8503);
xnor U12430 (N_12430,N_6186,N_9488);
or U12431 (N_12431,N_7907,N_9914);
nand U12432 (N_12432,N_8668,N_7376);
and U12433 (N_12433,N_5986,N_5245);
or U12434 (N_12434,N_5334,N_9222);
nand U12435 (N_12435,N_7654,N_8012);
or U12436 (N_12436,N_5317,N_5941);
nand U12437 (N_12437,N_7635,N_5153);
nand U12438 (N_12438,N_9741,N_5179);
or U12439 (N_12439,N_6357,N_7373);
nor U12440 (N_12440,N_5746,N_5884);
xor U12441 (N_12441,N_8574,N_5728);
and U12442 (N_12442,N_6217,N_6869);
nor U12443 (N_12443,N_7232,N_9708);
xnor U12444 (N_12444,N_6659,N_6897);
nor U12445 (N_12445,N_6894,N_8001);
nand U12446 (N_12446,N_7378,N_8904);
xnor U12447 (N_12447,N_5655,N_9871);
or U12448 (N_12448,N_6054,N_7786);
xor U12449 (N_12449,N_9176,N_8712);
and U12450 (N_12450,N_5070,N_8360);
xnor U12451 (N_12451,N_7952,N_7284);
nor U12452 (N_12452,N_8279,N_5171);
nor U12453 (N_12453,N_5774,N_9827);
nand U12454 (N_12454,N_7613,N_7448);
nor U12455 (N_12455,N_9575,N_9588);
nor U12456 (N_12456,N_8017,N_5514);
nand U12457 (N_12457,N_7532,N_7259);
xnor U12458 (N_12458,N_5422,N_8163);
xnor U12459 (N_12459,N_5408,N_7472);
nor U12460 (N_12460,N_6206,N_7962);
nand U12461 (N_12461,N_5909,N_5482);
and U12462 (N_12462,N_8469,N_6263);
xor U12463 (N_12463,N_7525,N_6800);
nand U12464 (N_12464,N_8190,N_7605);
xor U12465 (N_12465,N_9616,N_9712);
xor U12466 (N_12466,N_7397,N_6279);
or U12467 (N_12467,N_9617,N_6045);
and U12468 (N_12468,N_8804,N_6557);
and U12469 (N_12469,N_8296,N_9113);
nor U12470 (N_12470,N_5535,N_8969);
nor U12471 (N_12471,N_8697,N_8812);
and U12472 (N_12472,N_8248,N_7713);
or U12473 (N_12473,N_8814,N_7063);
and U12474 (N_12474,N_8862,N_5814);
xor U12475 (N_12475,N_5248,N_9468);
nor U12476 (N_12476,N_7131,N_7334);
nor U12477 (N_12477,N_8065,N_6231);
xor U12478 (N_12478,N_7253,N_5712);
and U12479 (N_12479,N_8825,N_8766);
nand U12480 (N_12480,N_9297,N_7722);
nand U12481 (N_12481,N_8318,N_9541);
or U12482 (N_12482,N_7101,N_6904);
nor U12483 (N_12483,N_7067,N_5427);
or U12484 (N_12484,N_8270,N_8451);
nand U12485 (N_12485,N_7957,N_8535);
nand U12486 (N_12486,N_7462,N_9034);
xor U12487 (N_12487,N_7756,N_6720);
or U12488 (N_12488,N_9424,N_8713);
nor U12489 (N_12489,N_5596,N_6985);
xor U12490 (N_12490,N_5261,N_6713);
and U12491 (N_12491,N_9538,N_8918);
and U12492 (N_12492,N_6729,N_9965);
and U12493 (N_12493,N_7557,N_8517);
nor U12494 (N_12494,N_8212,N_9791);
nand U12495 (N_12495,N_5891,N_7495);
or U12496 (N_12496,N_5061,N_8681);
and U12497 (N_12497,N_7511,N_9992);
or U12498 (N_12498,N_9104,N_8549);
or U12499 (N_12499,N_7914,N_9502);
nor U12500 (N_12500,N_8718,N_9096);
and U12501 (N_12501,N_7030,N_8571);
and U12502 (N_12502,N_7238,N_5586);
nor U12503 (N_12503,N_8701,N_8730);
or U12504 (N_12504,N_8641,N_9075);
nand U12505 (N_12505,N_9413,N_6691);
xnor U12506 (N_12506,N_7624,N_5006);
xnor U12507 (N_12507,N_9445,N_5837);
and U12508 (N_12508,N_9622,N_7938);
nor U12509 (N_12509,N_8942,N_5653);
xor U12510 (N_12510,N_8826,N_7955);
or U12511 (N_12511,N_5282,N_8848);
or U12512 (N_12512,N_6613,N_9535);
nand U12513 (N_12513,N_6277,N_6287);
xnor U12514 (N_12514,N_5173,N_8758);
nor U12515 (N_12515,N_8469,N_9690);
and U12516 (N_12516,N_7213,N_7515);
nor U12517 (N_12517,N_5919,N_6266);
and U12518 (N_12518,N_9019,N_7174);
and U12519 (N_12519,N_6182,N_6885);
xor U12520 (N_12520,N_5252,N_7354);
and U12521 (N_12521,N_5274,N_9598);
or U12522 (N_12522,N_6272,N_6837);
nor U12523 (N_12523,N_5890,N_7529);
or U12524 (N_12524,N_9211,N_7910);
xor U12525 (N_12525,N_9831,N_7523);
nand U12526 (N_12526,N_5598,N_9303);
and U12527 (N_12527,N_7649,N_8124);
nand U12528 (N_12528,N_9133,N_7993);
and U12529 (N_12529,N_7843,N_5094);
and U12530 (N_12530,N_7894,N_8499);
xor U12531 (N_12531,N_5765,N_9831);
nand U12532 (N_12532,N_5785,N_5654);
xnor U12533 (N_12533,N_5364,N_7251);
xnor U12534 (N_12534,N_5668,N_9906);
and U12535 (N_12535,N_8437,N_9024);
and U12536 (N_12536,N_7171,N_8157);
nor U12537 (N_12537,N_6440,N_5885);
xnor U12538 (N_12538,N_5534,N_8772);
or U12539 (N_12539,N_6200,N_6346);
xnor U12540 (N_12540,N_9421,N_7994);
xnor U12541 (N_12541,N_6817,N_9042);
or U12542 (N_12542,N_7707,N_8429);
and U12543 (N_12543,N_7032,N_5879);
and U12544 (N_12544,N_5144,N_7531);
nor U12545 (N_12545,N_8296,N_8974);
nor U12546 (N_12546,N_8047,N_6178);
and U12547 (N_12547,N_7266,N_7347);
xor U12548 (N_12548,N_7906,N_5995);
xnor U12549 (N_12549,N_9553,N_9395);
and U12550 (N_12550,N_7129,N_6367);
xnor U12551 (N_12551,N_5657,N_9873);
nand U12552 (N_12552,N_6783,N_9085);
or U12553 (N_12553,N_8300,N_6637);
or U12554 (N_12554,N_5531,N_5931);
or U12555 (N_12555,N_5443,N_9790);
xnor U12556 (N_12556,N_7189,N_7662);
xor U12557 (N_12557,N_7480,N_6585);
and U12558 (N_12558,N_7656,N_9707);
or U12559 (N_12559,N_6649,N_9813);
xnor U12560 (N_12560,N_5295,N_9469);
nand U12561 (N_12561,N_7786,N_8894);
xnor U12562 (N_12562,N_5005,N_5475);
and U12563 (N_12563,N_7947,N_7462);
xor U12564 (N_12564,N_5271,N_8633);
nor U12565 (N_12565,N_7125,N_6537);
nand U12566 (N_12566,N_8312,N_8469);
or U12567 (N_12567,N_6746,N_8293);
xor U12568 (N_12568,N_5650,N_7469);
xnor U12569 (N_12569,N_5662,N_8510);
xnor U12570 (N_12570,N_5924,N_8271);
and U12571 (N_12571,N_9174,N_7425);
or U12572 (N_12572,N_7653,N_5909);
nor U12573 (N_12573,N_7213,N_5944);
and U12574 (N_12574,N_6632,N_7599);
and U12575 (N_12575,N_6416,N_7090);
nor U12576 (N_12576,N_9598,N_8548);
and U12577 (N_12577,N_5498,N_8376);
nor U12578 (N_12578,N_6933,N_6035);
xor U12579 (N_12579,N_7717,N_8609);
or U12580 (N_12580,N_6251,N_6271);
or U12581 (N_12581,N_8542,N_9725);
nor U12582 (N_12582,N_9407,N_5277);
nand U12583 (N_12583,N_9973,N_7895);
or U12584 (N_12584,N_6147,N_9656);
nor U12585 (N_12585,N_6722,N_6798);
xor U12586 (N_12586,N_6764,N_7296);
nand U12587 (N_12587,N_8262,N_6336);
and U12588 (N_12588,N_9640,N_5452);
xnor U12589 (N_12589,N_7968,N_6813);
nand U12590 (N_12590,N_6125,N_8964);
nand U12591 (N_12591,N_5629,N_9355);
and U12592 (N_12592,N_6223,N_9772);
xnor U12593 (N_12593,N_6720,N_5734);
xor U12594 (N_12594,N_6686,N_7042);
nand U12595 (N_12595,N_7951,N_7170);
or U12596 (N_12596,N_7450,N_9108);
and U12597 (N_12597,N_9063,N_6666);
and U12598 (N_12598,N_6588,N_6429);
and U12599 (N_12599,N_6311,N_7071);
nand U12600 (N_12600,N_6100,N_8343);
or U12601 (N_12601,N_5701,N_7925);
or U12602 (N_12602,N_5347,N_9617);
xnor U12603 (N_12603,N_8957,N_9303);
or U12604 (N_12604,N_5563,N_9034);
and U12605 (N_12605,N_8153,N_5322);
xnor U12606 (N_12606,N_6796,N_7928);
nor U12607 (N_12607,N_6940,N_6777);
nand U12608 (N_12608,N_7182,N_5684);
and U12609 (N_12609,N_6285,N_5591);
nor U12610 (N_12610,N_5694,N_6930);
nand U12611 (N_12611,N_5566,N_7602);
and U12612 (N_12612,N_8457,N_9138);
xor U12613 (N_12613,N_6500,N_7608);
nand U12614 (N_12614,N_9527,N_7707);
or U12615 (N_12615,N_6987,N_5856);
nor U12616 (N_12616,N_6717,N_5143);
nor U12617 (N_12617,N_6674,N_8136);
and U12618 (N_12618,N_5049,N_6694);
xnor U12619 (N_12619,N_7232,N_5365);
xor U12620 (N_12620,N_5576,N_5820);
and U12621 (N_12621,N_6067,N_7368);
nand U12622 (N_12622,N_7142,N_9020);
xnor U12623 (N_12623,N_6415,N_7571);
xor U12624 (N_12624,N_7343,N_9939);
or U12625 (N_12625,N_7438,N_5064);
or U12626 (N_12626,N_8657,N_8822);
nor U12627 (N_12627,N_6337,N_7906);
xor U12628 (N_12628,N_7490,N_9193);
or U12629 (N_12629,N_6117,N_7374);
nand U12630 (N_12630,N_5485,N_9632);
nor U12631 (N_12631,N_9021,N_5643);
or U12632 (N_12632,N_9124,N_5235);
nor U12633 (N_12633,N_5612,N_8414);
and U12634 (N_12634,N_7346,N_5805);
nor U12635 (N_12635,N_9390,N_9468);
nand U12636 (N_12636,N_7160,N_7968);
nor U12637 (N_12637,N_6483,N_9389);
nand U12638 (N_12638,N_5847,N_5157);
and U12639 (N_12639,N_8419,N_6277);
nor U12640 (N_12640,N_5731,N_5899);
and U12641 (N_12641,N_8870,N_5003);
xnor U12642 (N_12642,N_5593,N_6686);
nand U12643 (N_12643,N_5710,N_9346);
and U12644 (N_12644,N_8099,N_7981);
xor U12645 (N_12645,N_9805,N_5182);
or U12646 (N_12646,N_5522,N_6024);
xnor U12647 (N_12647,N_9823,N_6807);
and U12648 (N_12648,N_7467,N_6653);
or U12649 (N_12649,N_8821,N_7503);
nand U12650 (N_12650,N_9339,N_9528);
nor U12651 (N_12651,N_5370,N_6183);
nand U12652 (N_12652,N_8452,N_5142);
xnor U12653 (N_12653,N_5601,N_9872);
nand U12654 (N_12654,N_5805,N_5766);
or U12655 (N_12655,N_6810,N_9555);
xnor U12656 (N_12656,N_7797,N_6497);
nor U12657 (N_12657,N_8574,N_9861);
or U12658 (N_12658,N_9414,N_7372);
xor U12659 (N_12659,N_6761,N_9991);
xnor U12660 (N_12660,N_6847,N_9718);
xnor U12661 (N_12661,N_7751,N_9166);
or U12662 (N_12662,N_7800,N_9096);
or U12663 (N_12663,N_8442,N_7638);
or U12664 (N_12664,N_9860,N_9347);
and U12665 (N_12665,N_7484,N_9662);
nand U12666 (N_12666,N_6222,N_9102);
or U12667 (N_12667,N_6101,N_6058);
and U12668 (N_12668,N_5375,N_9918);
and U12669 (N_12669,N_9419,N_8308);
xor U12670 (N_12670,N_9551,N_7949);
and U12671 (N_12671,N_7841,N_9671);
nor U12672 (N_12672,N_6620,N_6058);
xor U12673 (N_12673,N_7523,N_6257);
xor U12674 (N_12674,N_7141,N_5293);
and U12675 (N_12675,N_8549,N_6948);
or U12676 (N_12676,N_7839,N_5245);
nand U12677 (N_12677,N_6859,N_8101);
nand U12678 (N_12678,N_8644,N_6613);
or U12679 (N_12679,N_5651,N_7569);
xor U12680 (N_12680,N_7493,N_8450);
or U12681 (N_12681,N_7739,N_9076);
nor U12682 (N_12682,N_8266,N_7874);
or U12683 (N_12683,N_7800,N_7170);
and U12684 (N_12684,N_9947,N_6328);
nand U12685 (N_12685,N_5635,N_6334);
xor U12686 (N_12686,N_8402,N_9874);
nand U12687 (N_12687,N_9496,N_7358);
nor U12688 (N_12688,N_6488,N_8769);
xnor U12689 (N_12689,N_5272,N_9740);
or U12690 (N_12690,N_7036,N_8140);
xnor U12691 (N_12691,N_9082,N_9600);
and U12692 (N_12692,N_8036,N_6720);
xor U12693 (N_12693,N_9102,N_9762);
xor U12694 (N_12694,N_5739,N_7615);
nor U12695 (N_12695,N_7391,N_5339);
or U12696 (N_12696,N_7936,N_9863);
nor U12697 (N_12697,N_5592,N_9619);
xnor U12698 (N_12698,N_8148,N_7493);
or U12699 (N_12699,N_6074,N_6133);
nor U12700 (N_12700,N_5961,N_8441);
or U12701 (N_12701,N_7476,N_5077);
nand U12702 (N_12702,N_6296,N_8674);
xnor U12703 (N_12703,N_9573,N_5529);
or U12704 (N_12704,N_6564,N_9663);
or U12705 (N_12705,N_7405,N_7211);
nor U12706 (N_12706,N_7377,N_5891);
or U12707 (N_12707,N_8465,N_5611);
nand U12708 (N_12708,N_6838,N_5503);
xnor U12709 (N_12709,N_7087,N_9027);
nand U12710 (N_12710,N_9075,N_8283);
or U12711 (N_12711,N_6560,N_6923);
nand U12712 (N_12712,N_5163,N_9277);
nand U12713 (N_12713,N_9687,N_5314);
or U12714 (N_12714,N_9406,N_6549);
nor U12715 (N_12715,N_9257,N_8844);
nor U12716 (N_12716,N_8199,N_9122);
or U12717 (N_12717,N_7676,N_6897);
and U12718 (N_12718,N_8182,N_5773);
and U12719 (N_12719,N_5304,N_9081);
nor U12720 (N_12720,N_7144,N_7521);
nor U12721 (N_12721,N_6396,N_9496);
xnor U12722 (N_12722,N_5723,N_9484);
and U12723 (N_12723,N_5599,N_5172);
nand U12724 (N_12724,N_8277,N_8088);
xor U12725 (N_12725,N_5647,N_5939);
or U12726 (N_12726,N_7113,N_7620);
or U12727 (N_12727,N_6032,N_9482);
xor U12728 (N_12728,N_5600,N_8981);
nor U12729 (N_12729,N_8404,N_8785);
and U12730 (N_12730,N_9513,N_9478);
and U12731 (N_12731,N_7672,N_7128);
nor U12732 (N_12732,N_6216,N_6078);
xor U12733 (N_12733,N_8790,N_5336);
nor U12734 (N_12734,N_9422,N_5748);
and U12735 (N_12735,N_7546,N_8367);
or U12736 (N_12736,N_6944,N_6866);
or U12737 (N_12737,N_8435,N_7367);
xor U12738 (N_12738,N_5423,N_5120);
and U12739 (N_12739,N_9820,N_8853);
nand U12740 (N_12740,N_7448,N_6887);
nand U12741 (N_12741,N_5817,N_6134);
and U12742 (N_12742,N_9294,N_8428);
xor U12743 (N_12743,N_8414,N_7940);
xnor U12744 (N_12744,N_8334,N_8052);
or U12745 (N_12745,N_6605,N_9895);
xnor U12746 (N_12746,N_9195,N_7098);
and U12747 (N_12747,N_8036,N_6936);
xor U12748 (N_12748,N_6891,N_8062);
or U12749 (N_12749,N_8034,N_5506);
xor U12750 (N_12750,N_9116,N_7055);
xor U12751 (N_12751,N_8622,N_5368);
xor U12752 (N_12752,N_6011,N_7004);
nand U12753 (N_12753,N_9991,N_5461);
and U12754 (N_12754,N_6938,N_6330);
nand U12755 (N_12755,N_6048,N_5438);
nand U12756 (N_12756,N_6063,N_7211);
and U12757 (N_12757,N_6614,N_5104);
or U12758 (N_12758,N_9040,N_9278);
and U12759 (N_12759,N_8663,N_9274);
or U12760 (N_12760,N_5236,N_6322);
nand U12761 (N_12761,N_9324,N_7685);
and U12762 (N_12762,N_6586,N_6283);
nand U12763 (N_12763,N_8160,N_8177);
xor U12764 (N_12764,N_8599,N_7657);
nor U12765 (N_12765,N_9560,N_8938);
or U12766 (N_12766,N_7323,N_5771);
or U12767 (N_12767,N_6666,N_8839);
and U12768 (N_12768,N_8265,N_8704);
and U12769 (N_12769,N_6931,N_9913);
or U12770 (N_12770,N_7067,N_8938);
and U12771 (N_12771,N_5050,N_8059);
nor U12772 (N_12772,N_6303,N_9556);
nand U12773 (N_12773,N_5215,N_8187);
nand U12774 (N_12774,N_8620,N_5392);
or U12775 (N_12775,N_5342,N_7656);
and U12776 (N_12776,N_7248,N_7542);
nand U12777 (N_12777,N_7179,N_7196);
xnor U12778 (N_12778,N_5633,N_7714);
and U12779 (N_12779,N_8862,N_6575);
and U12780 (N_12780,N_5641,N_8541);
nand U12781 (N_12781,N_9754,N_9952);
and U12782 (N_12782,N_9137,N_5586);
and U12783 (N_12783,N_7727,N_5427);
nor U12784 (N_12784,N_5492,N_6415);
nand U12785 (N_12785,N_8235,N_7904);
and U12786 (N_12786,N_9836,N_7181);
nor U12787 (N_12787,N_6482,N_7629);
and U12788 (N_12788,N_9631,N_8995);
xnor U12789 (N_12789,N_8365,N_6292);
xnor U12790 (N_12790,N_7459,N_6539);
and U12791 (N_12791,N_7208,N_7754);
nor U12792 (N_12792,N_6672,N_5139);
nor U12793 (N_12793,N_6756,N_5700);
or U12794 (N_12794,N_8929,N_9815);
or U12795 (N_12795,N_9230,N_5155);
xnor U12796 (N_12796,N_6659,N_7301);
and U12797 (N_12797,N_8318,N_9523);
and U12798 (N_12798,N_7179,N_9872);
nor U12799 (N_12799,N_7704,N_6466);
or U12800 (N_12800,N_8567,N_8424);
or U12801 (N_12801,N_5164,N_9657);
xnor U12802 (N_12802,N_9091,N_6418);
and U12803 (N_12803,N_7027,N_9620);
xor U12804 (N_12804,N_5994,N_7699);
nand U12805 (N_12805,N_5173,N_6185);
and U12806 (N_12806,N_8103,N_8044);
and U12807 (N_12807,N_7464,N_5102);
and U12808 (N_12808,N_5306,N_9932);
xor U12809 (N_12809,N_7585,N_9537);
xnor U12810 (N_12810,N_5301,N_9920);
xor U12811 (N_12811,N_9851,N_9504);
or U12812 (N_12812,N_6988,N_5092);
nand U12813 (N_12813,N_8094,N_7902);
nand U12814 (N_12814,N_9147,N_7167);
nand U12815 (N_12815,N_6820,N_8689);
nor U12816 (N_12816,N_9376,N_7248);
or U12817 (N_12817,N_6427,N_7478);
and U12818 (N_12818,N_7848,N_9795);
and U12819 (N_12819,N_8320,N_9694);
and U12820 (N_12820,N_9558,N_7455);
or U12821 (N_12821,N_8265,N_7571);
or U12822 (N_12822,N_8313,N_8310);
xnor U12823 (N_12823,N_6878,N_7403);
nor U12824 (N_12824,N_5939,N_6073);
and U12825 (N_12825,N_7618,N_7273);
nand U12826 (N_12826,N_7014,N_7691);
nand U12827 (N_12827,N_8309,N_9392);
nor U12828 (N_12828,N_9857,N_6889);
xnor U12829 (N_12829,N_7916,N_7666);
or U12830 (N_12830,N_7135,N_7167);
xnor U12831 (N_12831,N_6659,N_6859);
nor U12832 (N_12832,N_5120,N_6333);
and U12833 (N_12833,N_7595,N_8423);
nor U12834 (N_12834,N_6555,N_6241);
xnor U12835 (N_12835,N_8881,N_9784);
xor U12836 (N_12836,N_6711,N_6996);
nand U12837 (N_12837,N_7758,N_6000);
xnor U12838 (N_12838,N_6926,N_6626);
nor U12839 (N_12839,N_6266,N_8070);
and U12840 (N_12840,N_5747,N_9357);
or U12841 (N_12841,N_5019,N_9389);
nand U12842 (N_12842,N_6414,N_5127);
xor U12843 (N_12843,N_9309,N_6668);
nand U12844 (N_12844,N_5455,N_5694);
and U12845 (N_12845,N_9784,N_8361);
nor U12846 (N_12846,N_9005,N_7649);
and U12847 (N_12847,N_9556,N_7719);
nand U12848 (N_12848,N_7103,N_6845);
or U12849 (N_12849,N_5550,N_7797);
or U12850 (N_12850,N_6151,N_6510);
or U12851 (N_12851,N_6549,N_8560);
xor U12852 (N_12852,N_8226,N_9867);
xor U12853 (N_12853,N_6808,N_5333);
and U12854 (N_12854,N_9758,N_6148);
or U12855 (N_12855,N_8515,N_6317);
nand U12856 (N_12856,N_9781,N_9447);
nor U12857 (N_12857,N_6916,N_5190);
nor U12858 (N_12858,N_5602,N_5078);
xnor U12859 (N_12859,N_8952,N_6700);
nand U12860 (N_12860,N_8607,N_6693);
nor U12861 (N_12861,N_5112,N_8410);
nor U12862 (N_12862,N_7958,N_7914);
and U12863 (N_12863,N_7525,N_7930);
xnor U12864 (N_12864,N_5198,N_8561);
nor U12865 (N_12865,N_6331,N_6774);
nand U12866 (N_12866,N_5289,N_8647);
and U12867 (N_12867,N_7786,N_5307);
nor U12868 (N_12868,N_6951,N_7176);
nor U12869 (N_12869,N_5183,N_7372);
xnor U12870 (N_12870,N_8962,N_6420);
nand U12871 (N_12871,N_7372,N_8198);
nor U12872 (N_12872,N_9296,N_8671);
xor U12873 (N_12873,N_6129,N_8046);
xor U12874 (N_12874,N_5380,N_6935);
nor U12875 (N_12875,N_6810,N_7145);
or U12876 (N_12876,N_5987,N_6735);
xor U12877 (N_12877,N_5833,N_5543);
and U12878 (N_12878,N_9841,N_5972);
and U12879 (N_12879,N_5723,N_8426);
or U12880 (N_12880,N_9129,N_6725);
and U12881 (N_12881,N_7490,N_7770);
or U12882 (N_12882,N_9968,N_6014);
nand U12883 (N_12883,N_8146,N_8612);
xor U12884 (N_12884,N_6803,N_6668);
xnor U12885 (N_12885,N_6488,N_9034);
nand U12886 (N_12886,N_5845,N_8170);
nor U12887 (N_12887,N_6507,N_5378);
nor U12888 (N_12888,N_8615,N_8642);
and U12889 (N_12889,N_8680,N_5967);
and U12890 (N_12890,N_5719,N_7893);
and U12891 (N_12891,N_5066,N_8696);
or U12892 (N_12892,N_5937,N_5335);
nand U12893 (N_12893,N_6777,N_6525);
nor U12894 (N_12894,N_6786,N_9722);
nand U12895 (N_12895,N_8479,N_5110);
and U12896 (N_12896,N_7642,N_9033);
xnor U12897 (N_12897,N_7281,N_8952);
and U12898 (N_12898,N_6403,N_5915);
nand U12899 (N_12899,N_8153,N_5331);
nor U12900 (N_12900,N_5090,N_6154);
or U12901 (N_12901,N_8526,N_8230);
and U12902 (N_12902,N_9863,N_5242);
nor U12903 (N_12903,N_7489,N_5448);
or U12904 (N_12904,N_7747,N_5017);
nand U12905 (N_12905,N_7967,N_5052);
and U12906 (N_12906,N_7136,N_8225);
nor U12907 (N_12907,N_7848,N_9408);
or U12908 (N_12908,N_9268,N_6210);
nor U12909 (N_12909,N_9171,N_9338);
nand U12910 (N_12910,N_5414,N_9828);
nor U12911 (N_12911,N_9091,N_8662);
and U12912 (N_12912,N_5639,N_7887);
nor U12913 (N_12913,N_6174,N_7677);
nor U12914 (N_12914,N_5557,N_6308);
or U12915 (N_12915,N_5120,N_6969);
or U12916 (N_12916,N_9983,N_8645);
nand U12917 (N_12917,N_6370,N_5945);
nand U12918 (N_12918,N_8818,N_8694);
nor U12919 (N_12919,N_8970,N_7101);
or U12920 (N_12920,N_6466,N_5384);
and U12921 (N_12921,N_7048,N_7097);
and U12922 (N_12922,N_8642,N_7370);
xnor U12923 (N_12923,N_7333,N_9856);
nor U12924 (N_12924,N_8293,N_7943);
nor U12925 (N_12925,N_9676,N_7561);
or U12926 (N_12926,N_6935,N_7333);
or U12927 (N_12927,N_7257,N_8165);
and U12928 (N_12928,N_8558,N_7573);
and U12929 (N_12929,N_7290,N_9091);
nand U12930 (N_12930,N_5514,N_9976);
nor U12931 (N_12931,N_8304,N_5850);
and U12932 (N_12932,N_8480,N_6111);
xnor U12933 (N_12933,N_8620,N_5555);
and U12934 (N_12934,N_8814,N_5992);
xor U12935 (N_12935,N_7581,N_8041);
nor U12936 (N_12936,N_6702,N_8813);
nand U12937 (N_12937,N_6321,N_6732);
or U12938 (N_12938,N_9386,N_8881);
and U12939 (N_12939,N_9836,N_9741);
xnor U12940 (N_12940,N_5665,N_6063);
nor U12941 (N_12941,N_7139,N_8503);
nand U12942 (N_12942,N_7012,N_5067);
or U12943 (N_12943,N_8894,N_7230);
xor U12944 (N_12944,N_6336,N_8144);
xnor U12945 (N_12945,N_7671,N_8451);
xnor U12946 (N_12946,N_8738,N_7129);
xnor U12947 (N_12947,N_9160,N_6303);
nand U12948 (N_12948,N_7663,N_8263);
nand U12949 (N_12949,N_9979,N_9981);
nand U12950 (N_12950,N_5399,N_9740);
and U12951 (N_12951,N_9263,N_9007);
nand U12952 (N_12952,N_7412,N_8071);
xor U12953 (N_12953,N_7532,N_8150);
or U12954 (N_12954,N_7896,N_7448);
nand U12955 (N_12955,N_7139,N_9398);
nand U12956 (N_12956,N_8605,N_6234);
or U12957 (N_12957,N_5069,N_8637);
xor U12958 (N_12958,N_6649,N_9127);
and U12959 (N_12959,N_7445,N_5164);
nor U12960 (N_12960,N_7222,N_9861);
xor U12961 (N_12961,N_9635,N_5175);
and U12962 (N_12962,N_7163,N_7017);
or U12963 (N_12963,N_8166,N_7788);
nand U12964 (N_12964,N_7789,N_8001);
nor U12965 (N_12965,N_7151,N_5069);
and U12966 (N_12966,N_8548,N_8295);
nand U12967 (N_12967,N_8811,N_7049);
and U12968 (N_12968,N_9666,N_7952);
xnor U12969 (N_12969,N_9620,N_8577);
nand U12970 (N_12970,N_6191,N_6234);
and U12971 (N_12971,N_5038,N_8889);
xor U12972 (N_12972,N_5998,N_6253);
nor U12973 (N_12973,N_8115,N_9071);
nor U12974 (N_12974,N_5281,N_8383);
or U12975 (N_12975,N_5206,N_5290);
or U12976 (N_12976,N_5338,N_6885);
and U12977 (N_12977,N_6007,N_6291);
nor U12978 (N_12978,N_9007,N_5909);
or U12979 (N_12979,N_8556,N_7366);
nor U12980 (N_12980,N_9096,N_9900);
or U12981 (N_12981,N_5815,N_8328);
xnor U12982 (N_12982,N_7094,N_7343);
nand U12983 (N_12983,N_5722,N_6559);
nand U12984 (N_12984,N_5101,N_6207);
nand U12985 (N_12985,N_6990,N_6504);
xnor U12986 (N_12986,N_7385,N_6133);
xnor U12987 (N_12987,N_5402,N_6203);
or U12988 (N_12988,N_8846,N_5035);
xnor U12989 (N_12989,N_8390,N_7885);
xor U12990 (N_12990,N_9165,N_8269);
or U12991 (N_12991,N_6539,N_7633);
nand U12992 (N_12992,N_7349,N_8092);
xor U12993 (N_12993,N_7470,N_5650);
nor U12994 (N_12994,N_5895,N_7026);
nor U12995 (N_12995,N_7248,N_8041);
xor U12996 (N_12996,N_6875,N_5369);
xnor U12997 (N_12997,N_5470,N_6920);
xor U12998 (N_12998,N_9336,N_5613);
xor U12999 (N_12999,N_8215,N_9260);
nand U13000 (N_13000,N_6310,N_7986);
and U13001 (N_13001,N_6089,N_7540);
nor U13002 (N_13002,N_9152,N_9365);
and U13003 (N_13003,N_5479,N_8829);
xor U13004 (N_13004,N_8351,N_6338);
and U13005 (N_13005,N_7846,N_5845);
nand U13006 (N_13006,N_7363,N_9437);
nor U13007 (N_13007,N_6827,N_6880);
or U13008 (N_13008,N_6142,N_7895);
xor U13009 (N_13009,N_8795,N_9270);
nand U13010 (N_13010,N_8923,N_7130);
or U13011 (N_13011,N_8958,N_6265);
xor U13012 (N_13012,N_5213,N_5873);
or U13013 (N_13013,N_7897,N_6728);
nor U13014 (N_13014,N_8634,N_9022);
nand U13015 (N_13015,N_5991,N_9902);
xnor U13016 (N_13016,N_5376,N_5193);
and U13017 (N_13017,N_7694,N_9077);
nor U13018 (N_13018,N_7909,N_5328);
nand U13019 (N_13019,N_5424,N_7736);
or U13020 (N_13020,N_9243,N_6515);
or U13021 (N_13021,N_8470,N_6002);
and U13022 (N_13022,N_5881,N_5227);
and U13023 (N_13023,N_5485,N_7732);
nor U13024 (N_13024,N_8123,N_6358);
and U13025 (N_13025,N_8304,N_7600);
nand U13026 (N_13026,N_7018,N_7762);
or U13027 (N_13027,N_7500,N_9102);
xnor U13028 (N_13028,N_9838,N_7268);
nand U13029 (N_13029,N_9158,N_9526);
nor U13030 (N_13030,N_7510,N_5652);
xor U13031 (N_13031,N_8588,N_5252);
nor U13032 (N_13032,N_7493,N_8426);
and U13033 (N_13033,N_5191,N_5271);
nor U13034 (N_13034,N_6620,N_6361);
and U13035 (N_13035,N_8540,N_5316);
nand U13036 (N_13036,N_5228,N_6127);
xor U13037 (N_13037,N_8137,N_9532);
nand U13038 (N_13038,N_8810,N_6264);
and U13039 (N_13039,N_8594,N_6573);
xnor U13040 (N_13040,N_6622,N_7910);
or U13041 (N_13041,N_9521,N_7826);
nand U13042 (N_13042,N_8832,N_6717);
nor U13043 (N_13043,N_9296,N_6814);
nor U13044 (N_13044,N_8290,N_7919);
nor U13045 (N_13045,N_6762,N_8138);
and U13046 (N_13046,N_6977,N_9059);
xor U13047 (N_13047,N_6475,N_6223);
xor U13048 (N_13048,N_9185,N_8018);
nand U13049 (N_13049,N_9764,N_6544);
or U13050 (N_13050,N_9405,N_9838);
and U13051 (N_13051,N_7300,N_5662);
and U13052 (N_13052,N_8922,N_7569);
xor U13053 (N_13053,N_8328,N_6814);
or U13054 (N_13054,N_9216,N_9439);
or U13055 (N_13055,N_9393,N_9174);
nand U13056 (N_13056,N_7908,N_8097);
and U13057 (N_13057,N_8909,N_6544);
nand U13058 (N_13058,N_5289,N_7698);
and U13059 (N_13059,N_6880,N_8557);
xor U13060 (N_13060,N_5113,N_5103);
nor U13061 (N_13061,N_7153,N_7019);
and U13062 (N_13062,N_8895,N_6378);
or U13063 (N_13063,N_9553,N_9443);
and U13064 (N_13064,N_9059,N_9889);
xor U13065 (N_13065,N_5690,N_5928);
nor U13066 (N_13066,N_8832,N_5670);
nand U13067 (N_13067,N_8666,N_9120);
nor U13068 (N_13068,N_7223,N_7271);
or U13069 (N_13069,N_6473,N_9259);
nand U13070 (N_13070,N_9517,N_9708);
xnor U13071 (N_13071,N_9545,N_5283);
xnor U13072 (N_13072,N_5339,N_7278);
xnor U13073 (N_13073,N_6303,N_8222);
nand U13074 (N_13074,N_9825,N_7923);
or U13075 (N_13075,N_6996,N_7325);
and U13076 (N_13076,N_9456,N_5115);
nor U13077 (N_13077,N_9698,N_7228);
xnor U13078 (N_13078,N_5525,N_9949);
nor U13079 (N_13079,N_9068,N_9185);
or U13080 (N_13080,N_7831,N_7991);
or U13081 (N_13081,N_9233,N_5013);
xor U13082 (N_13082,N_5777,N_5187);
and U13083 (N_13083,N_5142,N_7500);
or U13084 (N_13084,N_9744,N_5222);
nor U13085 (N_13085,N_7846,N_9350);
nand U13086 (N_13086,N_5300,N_6378);
nand U13087 (N_13087,N_9934,N_9495);
or U13088 (N_13088,N_8770,N_5626);
and U13089 (N_13089,N_8859,N_9143);
nor U13090 (N_13090,N_9214,N_6054);
nor U13091 (N_13091,N_7389,N_5723);
nor U13092 (N_13092,N_8880,N_8427);
or U13093 (N_13093,N_7610,N_7498);
nand U13094 (N_13094,N_5710,N_5331);
and U13095 (N_13095,N_6074,N_7798);
nand U13096 (N_13096,N_8209,N_6614);
nand U13097 (N_13097,N_5932,N_5003);
nand U13098 (N_13098,N_7545,N_5590);
xor U13099 (N_13099,N_5888,N_7146);
and U13100 (N_13100,N_6460,N_8022);
nor U13101 (N_13101,N_9002,N_9867);
nor U13102 (N_13102,N_6870,N_7946);
xor U13103 (N_13103,N_6994,N_9763);
or U13104 (N_13104,N_7775,N_7452);
or U13105 (N_13105,N_6688,N_9073);
or U13106 (N_13106,N_8846,N_5472);
nor U13107 (N_13107,N_9725,N_9470);
nor U13108 (N_13108,N_9316,N_7893);
nor U13109 (N_13109,N_6558,N_6137);
nand U13110 (N_13110,N_7590,N_7585);
or U13111 (N_13111,N_7951,N_5452);
and U13112 (N_13112,N_9087,N_7641);
nand U13113 (N_13113,N_5413,N_7291);
nand U13114 (N_13114,N_7296,N_6696);
nor U13115 (N_13115,N_7726,N_7535);
nand U13116 (N_13116,N_5027,N_5188);
xor U13117 (N_13117,N_6764,N_8215);
nor U13118 (N_13118,N_7017,N_5416);
nand U13119 (N_13119,N_7936,N_9511);
xnor U13120 (N_13120,N_9552,N_7733);
nor U13121 (N_13121,N_5431,N_8364);
or U13122 (N_13122,N_7327,N_6450);
xnor U13123 (N_13123,N_6153,N_6685);
nand U13124 (N_13124,N_8592,N_5143);
and U13125 (N_13125,N_6663,N_6535);
xnor U13126 (N_13126,N_5077,N_5766);
or U13127 (N_13127,N_9991,N_9229);
nor U13128 (N_13128,N_5242,N_7883);
xnor U13129 (N_13129,N_5722,N_7264);
xor U13130 (N_13130,N_7430,N_9127);
nor U13131 (N_13131,N_9728,N_9824);
or U13132 (N_13132,N_5302,N_6779);
nor U13133 (N_13133,N_8076,N_9496);
nand U13134 (N_13134,N_9696,N_9682);
nor U13135 (N_13135,N_8086,N_5359);
xor U13136 (N_13136,N_7093,N_9257);
nand U13137 (N_13137,N_6122,N_6961);
and U13138 (N_13138,N_8340,N_7042);
or U13139 (N_13139,N_7315,N_8855);
nand U13140 (N_13140,N_6412,N_9399);
or U13141 (N_13141,N_9389,N_7432);
and U13142 (N_13142,N_5746,N_6350);
nand U13143 (N_13143,N_6247,N_9662);
nand U13144 (N_13144,N_5660,N_9170);
nor U13145 (N_13145,N_8641,N_7128);
nand U13146 (N_13146,N_9655,N_9132);
or U13147 (N_13147,N_5706,N_8974);
nor U13148 (N_13148,N_6209,N_7791);
or U13149 (N_13149,N_9545,N_7955);
and U13150 (N_13150,N_5160,N_7558);
nand U13151 (N_13151,N_9429,N_5149);
xor U13152 (N_13152,N_8960,N_9433);
or U13153 (N_13153,N_6299,N_9578);
and U13154 (N_13154,N_8725,N_6209);
nor U13155 (N_13155,N_7206,N_8003);
and U13156 (N_13156,N_5465,N_9998);
or U13157 (N_13157,N_8787,N_9045);
nor U13158 (N_13158,N_7201,N_7019);
nor U13159 (N_13159,N_5504,N_8684);
nor U13160 (N_13160,N_5403,N_5620);
xnor U13161 (N_13161,N_7565,N_5251);
nand U13162 (N_13162,N_7272,N_8747);
xnor U13163 (N_13163,N_5466,N_9974);
nor U13164 (N_13164,N_5975,N_5243);
nand U13165 (N_13165,N_5986,N_7351);
nor U13166 (N_13166,N_9347,N_6834);
nor U13167 (N_13167,N_6441,N_5768);
xnor U13168 (N_13168,N_5293,N_8694);
xor U13169 (N_13169,N_8470,N_5046);
nor U13170 (N_13170,N_6407,N_8379);
nor U13171 (N_13171,N_6872,N_8707);
nand U13172 (N_13172,N_7191,N_7661);
nand U13173 (N_13173,N_9004,N_5555);
or U13174 (N_13174,N_5014,N_8191);
xnor U13175 (N_13175,N_6892,N_7402);
and U13176 (N_13176,N_8915,N_7783);
nor U13177 (N_13177,N_5299,N_9057);
or U13178 (N_13178,N_7976,N_6727);
xor U13179 (N_13179,N_7009,N_8417);
nor U13180 (N_13180,N_9460,N_5888);
nor U13181 (N_13181,N_5957,N_8765);
and U13182 (N_13182,N_5377,N_9325);
nand U13183 (N_13183,N_8977,N_6244);
xor U13184 (N_13184,N_8334,N_6717);
or U13185 (N_13185,N_9067,N_6661);
nor U13186 (N_13186,N_9368,N_9345);
or U13187 (N_13187,N_5068,N_9131);
and U13188 (N_13188,N_5981,N_5820);
nor U13189 (N_13189,N_9977,N_7311);
xor U13190 (N_13190,N_8791,N_7563);
xor U13191 (N_13191,N_5993,N_8175);
and U13192 (N_13192,N_5426,N_9173);
xor U13193 (N_13193,N_9151,N_7150);
and U13194 (N_13194,N_9505,N_7323);
xor U13195 (N_13195,N_5751,N_6299);
and U13196 (N_13196,N_6929,N_6360);
xor U13197 (N_13197,N_5509,N_6467);
nand U13198 (N_13198,N_5802,N_5011);
or U13199 (N_13199,N_7315,N_8911);
and U13200 (N_13200,N_5327,N_6556);
nand U13201 (N_13201,N_8560,N_7963);
or U13202 (N_13202,N_5079,N_7575);
nor U13203 (N_13203,N_8476,N_8273);
or U13204 (N_13204,N_8294,N_8543);
xnor U13205 (N_13205,N_7752,N_8811);
and U13206 (N_13206,N_6688,N_5540);
nor U13207 (N_13207,N_8067,N_9081);
and U13208 (N_13208,N_7309,N_6289);
or U13209 (N_13209,N_6969,N_5951);
or U13210 (N_13210,N_6899,N_7868);
nand U13211 (N_13211,N_8968,N_9868);
nand U13212 (N_13212,N_5419,N_7479);
nand U13213 (N_13213,N_6983,N_7878);
or U13214 (N_13214,N_6486,N_7086);
or U13215 (N_13215,N_5285,N_7880);
nand U13216 (N_13216,N_8283,N_8310);
nand U13217 (N_13217,N_7192,N_6204);
nand U13218 (N_13218,N_6005,N_8274);
nand U13219 (N_13219,N_5654,N_8182);
or U13220 (N_13220,N_9060,N_9108);
xnor U13221 (N_13221,N_8930,N_7892);
and U13222 (N_13222,N_9188,N_9638);
or U13223 (N_13223,N_5466,N_8361);
nand U13224 (N_13224,N_6570,N_9410);
or U13225 (N_13225,N_9814,N_9395);
or U13226 (N_13226,N_6771,N_6468);
nand U13227 (N_13227,N_6700,N_9853);
xnor U13228 (N_13228,N_8053,N_5617);
or U13229 (N_13229,N_9285,N_8346);
and U13230 (N_13230,N_5815,N_9808);
xor U13231 (N_13231,N_6870,N_8324);
nor U13232 (N_13232,N_9008,N_9520);
nor U13233 (N_13233,N_5565,N_5887);
or U13234 (N_13234,N_8530,N_9195);
nor U13235 (N_13235,N_6937,N_6862);
nand U13236 (N_13236,N_5177,N_9859);
nor U13237 (N_13237,N_5143,N_7131);
nor U13238 (N_13238,N_5224,N_5350);
and U13239 (N_13239,N_6157,N_7876);
or U13240 (N_13240,N_5112,N_9402);
and U13241 (N_13241,N_6753,N_6312);
nand U13242 (N_13242,N_7943,N_5025);
or U13243 (N_13243,N_8539,N_5997);
or U13244 (N_13244,N_8000,N_5575);
nor U13245 (N_13245,N_5635,N_7723);
xor U13246 (N_13246,N_6322,N_5631);
nor U13247 (N_13247,N_8139,N_7875);
xor U13248 (N_13248,N_7217,N_6416);
and U13249 (N_13249,N_8200,N_7466);
nand U13250 (N_13250,N_7983,N_7280);
xor U13251 (N_13251,N_6506,N_7292);
xor U13252 (N_13252,N_6496,N_6107);
and U13253 (N_13253,N_8896,N_9019);
and U13254 (N_13254,N_9370,N_6743);
or U13255 (N_13255,N_9112,N_6746);
nor U13256 (N_13256,N_7047,N_8622);
and U13257 (N_13257,N_8933,N_5208);
xnor U13258 (N_13258,N_9036,N_7614);
and U13259 (N_13259,N_7196,N_5492);
xor U13260 (N_13260,N_7384,N_7308);
xnor U13261 (N_13261,N_6016,N_6391);
xnor U13262 (N_13262,N_5447,N_5405);
nor U13263 (N_13263,N_7233,N_6433);
xnor U13264 (N_13264,N_6716,N_8412);
or U13265 (N_13265,N_9915,N_9231);
nor U13266 (N_13266,N_9374,N_8263);
xnor U13267 (N_13267,N_9579,N_9219);
nand U13268 (N_13268,N_8715,N_6836);
nor U13269 (N_13269,N_7568,N_9044);
and U13270 (N_13270,N_6164,N_5112);
or U13271 (N_13271,N_5866,N_5754);
nand U13272 (N_13272,N_9006,N_8566);
or U13273 (N_13273,N_8328,N_5939);
nand U13274 (N_13274,N_9444,N_6943);
xor U13275 (N_13275,N_9601,N_7084);
xor U13276 (N_13276,N_6848,N_7160);
xor U13277 (N_13277,N_6153,N_9142);
or U13278 (N_13278,N_5360,N_8932);
nand U13279 (N_13279,N_7927,N_5493);
or U13280 (N_13280,N_7964,N_6850);
nor U13281 (N_13281,N_5366,N_7258);
nor U13282 (N_13282,N_5664,N_6116);
nor U13283 (N_13283,N_5623,N_6499);
xnor U13284 (N_13284,N_7146,N_9545);
nand U13285 (N_13285,N_6718,N_6374);
nor U13286 (N_13286,N_5697,N_7004);
nand U13287 (N_13287,N_9673,N_5178);
or U13288 (N_13288,N_5239,N_5844);
and U13289 (N_13289,N_9214,N_8307);
or U13290 (N_13290,N_6735,N_8581);
or U13291 (N_13291,N_9718,N_8391);
nand U13292 (N_13292,N_9763,N_8505);
and U13293 (N_13293,N_6576,N_8428);
and U13294 (N_13294,N_7253,N_8010);
nor U13295 (N_13295,N_7914,N_8905);
xor U13296 (N_13296,N_5456,N_5971);
nand U13297 (N_13297,N_7750,N_5525);
nor U13298 (N_13298,N_5888,N_5990);
and U13299 (N_13299,N_7766,N_7319);
or U13300 (N_13300,N_6763,N_6060);
xnor U13301 (N_13301,N_6769,N_7708);
nor U13302 (N_13302,N_9172,N_7118);
nand U13303 (N_13303,N_5278,N_5929);
nand U13304 (N_13304,N_5100,N_6639);
xor U13305 (N_13305,N_6749,N_6264);
or U13306 (N_13306,N_9557,N_5930);
and U13307 (N_13307,N_5429,N_7248);
nand U13308 (N_13308,N_9349,N_8519);
nor U13309 (N_13309,N_7044,N_8368);
nor U13310 (N_13310,N_7052,N_5810);
nor U13311 (N_13311,N_5123,N_9775);
nand U13312 (N_13312,N_7361,N_5237);
or U13313 (N_13313,N_8192,N_6382);
nand U13314 (N_13314,N_7290,N_8574);
nor U13315 (N_13315,N_9383,N_7057);
nor U13316 (N_13316,N_6233,N_8984);
xor U13317 (N_13317,N_5858,N_8417);
or U13318 (N_13318,N_7536,N_8924);
nor U13319 (N_13319,N_8060,N_8314);
nor U13320 (N_13320,N_7969,N_9868);
and U13321 (N_13321,N_8943,N_7880);
nand U13322 (N_13322,N_7097,N_9346);
nand U13323 (N_13323,N_5983,N_6713);
and U13324 (N_13324,N_8525,N_7044);
and U13325 (N_13325,N_6957,N_6373);
nand U13326 (N_13326,N_5280,N_6393);
nor U13327 (N_13327,N_9236,N_7619);
or U13328 (N_13328,N_5454,N_5563);
or U13329 (N_13329,N_8364,N_9769);
and U13330 (N_13330,N_7056,N_5521);
xnor U13331 (N_13331,N_8294,N_9294);
nand U13332 (N_13332,N_8900,N_8253);
or U13333 (N_13333,N_8607,N_6370);
or U13334 (N_13334,N_8616,N_7256);
or U13335 (N_13335,N_8442,N_5995);
nor U13336 (N_13336,N_7933,N_8753);
nand U13337 (N_13337,N_7898,N_8067);
xnor U13338 (N_13338,N_6507,N_7460);
nand U13339 (N_13339,N_8882,N_5102);
nand U13340 (N_13340,N_5965,N_8450);
xor U13341 (N_13341,N_7635,N_9997);
or U13342 (N_13342,N_5348,N_7115);
and U13343 (N_13343,N_8746,N_8532);
nand U13344 (N_13344,N_5928,N_6560);
nor U13345 (N_13345,N_7667,N_6648);
or U13346 (N_13346,N_7022,N_5218);
or U13347 (N_13347,N_9752,N_7159);
or U13348 (N_13348,N_9168,N_7134);
or U13349 (N_13349,N_6026,N_6242);
xnor U13350 (N_13350,N_7449,N_6987);
nor U13351 (N_13351,N_6413,N_9338);
nor U13352 (N_13352,N_8988,N_8381);
nand U13353 (N_13353,N_6098,N_8010);
nor U13354 (N_13354,N_6452,N_7112);
nor U13355 (N_13355,N_6431,N_5461);
and U13356 (N_13356,N_6814,N_6772);
or U13357 (N_13357,N_5359,N_7102);
and U13358 (N_13358,N_9446,N_9239);
xnor U13359 (N_13359,N_5799,N_5927);
or U13360 (N_13360,N_7567,N_9278);
nand U13361 (N_13361,N_5003,N_9692);
nand U13362 (N_13362,N_9126,N_6053);
nand U13363 (N_13363,N_5716,N_5155);
nand U13364 (N_13364,N_5586,N_7489);
nand U13365 (N_13365,N_8160,N_6019);
xnor U13366 (N_13366,N_5523,N_8799);
nand U13367 (N_13367,N_8038,N_8452);
xnor U13368 (N_13368,N_6980,N_6809);
xnor U13369 (N_13369,N_5897,N_5318);
and U13370 (N_13370,N_8282,N_5437);
nor U13371 (N_13371,N_8041,N_6679);
xnor U13372 (N_13372,N_9463,N_6771);
xnor U13373 (N_13373,N_8316,N_8319);
or U13374 (N_13374,N_8842,N_5987);
or U13375 (N_13375,N_7114,N_5025);
nand U13376 (N_13376,N_6226,N_8993);
and U13377 (N_13377,N_7987,N_7334);
or U13378 (N_13378,N_9134,N_5357);
nand U13379 (N_13379,N_7840,N_5058);
nand U13380 (N_13380,N_6377,N_8898);
or U13381 (N_13381,N_9806,N_5048);
xor U13382 (N_13382,N_6883,N_9200);
and U13383 (N_13383,N_9267,N_5293);
and U13384 (N_13384,N_9776,N_9771);
xnor U13385 (N_13385,N_6406,N_9344);
and U13386 (N_13386,N_5771,N_5647);
xnor U13387 (N_13387,N_9129,N_7458);
nor U13388 (N_13388,N_6796,N_7335);
nand U13389 (N_13389,N_6050,N_9304);
nor U13390 (N_13390,N_8613,N_8257);
nand U13391 (N_13391,N_7546,N_9243);
nand U13392 (N_13392,N_5284,N_9099);
and U13393 (N_13393,N_6124,N_7342);
nor U13394 (N_13394,N_8338,N_8058);
or U13395 (N_13395,N_7010,N_5297);
nor U13396 (N_13396,N_8396,N_6214);
and U13397 (N_13397,N_6674,N_9366);
xor U13398 (N_13398,N_5605,N_9116);
or U13399 (N_13399,N_7007,N_6235);
or U13400 (N_13400,N_6657,N_7793);
or U13401 (N_13401,N_5505,N_8461);
xor U13402 (N_13402,N_7642,N_6484);
or U13403 (N_13403,N_9398,N_8279);
nand U13404 (N_13404,N_6739,N_7800);
nor U13405 (N_13405,N_9411,N_8691);
nand U13406 (N_13406,N_9959,N_5487);
xor U13407 (N_13407,N_7449,N_7374);
nor U13408 (N_13408,N_7318,N_5964);
nand U13409 (N_13409,N_7441,N_9218);
nor U13410 (N_13410,N_5454,N_5380);
and U13411 (N_13411,N_8877,N_7360);
or U13412 (N_13412,N_6637,N_6583);
nor U13413 (N_13413,N_6714,N_6298);
xnor U13414 (N_13414,N_8752,N_6979);
and U13415 (N_13415,N_6783,N_9155);
and U13416 (N_13416,N_9019,N_5301);
and U13417 (N_13417,N_9626,N_5066);
xor U13418 (N_13418,N_8478,N_6228);
and U13419 (N_13419,N_6903,N_5876);
xor U13420 (N_13420,N_8597,N_8954);
nor U13421 (N_13421,N_9151,N_5638);
xor U13422 (N_13422,N_8251,N_8856);
or U13423 (N_13423,N_5408,N_7994);
nand U13424 (N_13424,N_8608,N_7338);
and U13425 (N_13425,N_8017,N_5749);
nand U13426 (N_13426,N_7194,N_9014);
or U13427 (N_13427,N_5007,N_6563);
nor U13428 (N_13428,N_5724,N_6655);
nor U13429 (N_13429,N_6489,N_6573);
xnor U13430 (N_13430,N_9711,N_5330);
and U13431 (N_13431,N_8413,N_5839);
nand U13432 (N_13432,N_6035,N_9358);
nor U13433 (N_13433,N_6443,N_5562);
or U13434 (N_13434,N_6251,N_8637);
and U13435 (N_13435,N_6927,N_8587);
or U13436 (N_13436,N_6462,N_5593);
and U13437 (N_13437,N_5961,N_9717);
and U13438 (N_13438,N_5206,N_8339);
or U13439 (N_13439,N_9175,N_6112);
and U13440 (N_13440,N_7914,N_9426);
nand U13441 (N_13441,N_9689,N_7459);
xor U13442 (N_13442,N_9077,N_8872);
nor U13443 (N_13443,N_8589,N_7747);
and U13444 (N_13444,N_5098,N_7613);
xnor U13445 (N_13445,N_7325,N_8740);
or U13446 (N_13446,N_5666,N_8896);
nand U13447 (N_13447,N_7113,N_8052);
nand U13448 (N_13448,N_8085,N_8306);
and U13449 (N_13449,N_9628,N_6766);
and U13450 (N_13450,N_7321,N_9765);
and U13451 (N_13451,N_7378,N_9080);
and U13452 (N_13452,N_5493,N_5973);
nor U13453 (N_13453,N_6709,N_7140);
xnor U13454 (N_13454,N_5356,N_8956);
nor U13455 (N_13455,N_9384,N_5119);
nor U13456 (N_13456,N_8026,N_8616);
nand U13457 (N_13457,N_9785,N_7954);
nand U13458 (N_13458,N_7475,N_8822);
or U13459 (N_13459,N_6992,N_9937);
or U13460 (N_13460,N_5825,N_9325);
nand U13461 (N_13461,N_9127,N_8350);
and U13462 (N_13462,N_8175,N_6818);
or U13463 (N_13463,N_9092,N_5658);
xor U13464 (N_13464,N_7617,N_6850);
and U13465 (N_13465,N_8317,N_9916);
nand U13466 (N_13466,N_8536,N_8911);
nand U13467 (N_13467,N_5428,N_9722);
xnor U13468 (N_13468,N_9972,N_9539);
xnor U13469 (N_13469,N_7266,N_9000);
or U13470 (N_13470,N_6900,N_8654);
nand U13471 (N_13471,N_7866,N_6943);
or U13472 (N_13472,N_8570,N_8178);
xor U13473 (N_13473,N_5498,N_9440);
nor U13474 (N_13474,N_6983,N_9078);
xnor U13475 (N_13475,N_6498,N_7788);
and U13476 (N_13476,N_8859,N_5942);
xnor U13477 (N_13477,N_8305,N_9693);
or U13478 (N_13478,N_5381,N_8914);
nor U13479 (N_13479,N_9160,N_6814);
or U13480 (N_13480,N_7262,N_8072);
nand U13481 (N_13481,N_9424,N_8041);
nand U13482 (N_13482,N_9704,N_6395);
and U13483 (N_13483,N_6127,N_6172);
nor U13484 (N_13484,N_5986,N_7687);
and U13485 (N_13485,N_8924,N_6031);
nor U13486 (N_13486,N_8852,N_7658);
nand U13487 (N_13487,N_8488,N_6668);
and U13488 (N_13488,N_7826,N_5535);
nand U13489 (N_13489,N_5602,N_6034);
nand U13490 (N_13490,N_9298,N_5501);
nand U13491 (N_13491,N_9590,N_9377);
and U13492 (N_13492,N_5927,N_8845);
nand U13493 (N_13493,N_5680,N_6645);
or U13494 (N_13494,N_5415,N_8369);
or U13495 (N_13495,N_6640,N_6876);
or U13496 (N_13496,N_8626,N_6548);
nor U13497 (N_13497,N_7953,N_7404);
nand U13498 (N_13498,N_7787,N_6797);
nor U13499 (N_13499,N_8992,N_8270);
or U13500 (N_13500,N_8465,N_5314);
and U13501 (N_13501,N_5575,N_9538);
nand U13502 (N_13502,N_6984,N_9031);
nand U13503 (N_13503,N_5543,N_9304);
nor U13504 (N_13504,N_5940,N_5301);
xor U13505 (N_13505,N_5393,N_7237);
nor U13506 (N_13506,N_5169,N_7854);
xor U13507 (N_13507,N_9624,N_8905);
nor U13508 (N_13508,N_9552,N_7302);
nand U13509 (N_13509,N_8382,N_6728);
xor U13510 (N_13510,N_5087,N_6711);
xnor U13511 (N_13511,N_9186,N_7923);
and U13512 (N_13512,N_9233,N_7408);
xor U13513 (N_13513,N_8689,N_8981);
nand U13514 (N_13514,N_7763,N_5363);
xor U13515 (N_13515,N_5134,N_9769);
and U13516 (N_13516,N_7837,N_8018);
and U13517 (N_13517,N_7574,N_8036);
xor U13518 (N_13518,N_9745,N_7505);
nor U13519 (N_13519,N_8444,N_8586);
and U13520 (N_13520,N_7169,N_7170);
xnor U13521 (N_13521,N_6017,N_7585);
nor U13522 (N_13522,N_9308,N_7008);
nand U13523 (N_13523,N_5582,N_6798);
nand U13524 (N_13524,N_7190,N_5288);
xor U13525 (N_13525,N_7716,N_8619);
nor U13526 (N_13526,N_7032,N_5909);
xnor U13527 (N_13527,N_8330,N_6693);
or U13528 (N_13528,N_5384,N_5702);
nor U13529 (N_13529,N_5580,N_8424);
and U13530 (N_13530,N_8004,N_6965);
and U13531 (N_13531,N_9021,N_6782);
or U13532 (N_13532,N_5818,N_6051);
or U13533 (N_13533,N_7782,N_9625);
xor U13534 (N_13534,N_6301,N_9175);
nand U13535 (N_13535,N_7950,N_7398);
nor U13536 (N_13536,N_9190,N_7232);
nand U13537 (N_13537,N_6865,N_7395);
and U13538 (N_13538,N_6640,N_6853);
nor U13539 (N_13539,N_5794,N_7497);
or U13540 (N_13540,N_7971,N_9712);
nor U13541 (N_13541,N_8255,N_6889);
nand U13542 (N_13542,N_7947,N_7132);
or U13543 (N_13543,N_9846,N_5837);
or U13544 (N_13544,N_6251,N_6848);
nand U13545 (N_13545,N_9031,N_6197);
nand U13546 (N_13546,N_5905,N_7696);
nor U13547 (N_13547,N_8597,N_7158);
xnor U13548 (N_13548,N_7514,N_7480);
and U13549 (N_13549,N_9167,N_7302);
or U13550 (N_13550,N_6576,N_6652);
or U13551 (N_13551,N_7106,N_9668);
and U13552 (N_13552,N_5428,N_8951);
nand U13553 (N_13553,N_6573,N_8783);
xnor U13554 (N_13554,N_8415,N_9911);
or U13555 (N_13555,N_7740,N_7241);
and U13556 (N_13556,N_6613,N_7495);
nand U13557 (N_13557,N_7131,N_7164);
or U13558 (N_13558,N_9647,N_7216);
nand U13559 (N_13559,N_6947,N_6743);
xor U13560 (N_13560,N_6457,N_6780);
nand U13561 (N_13561,N_8963,N_9478);
and U13562 (N_13562,N_7121,N_5725);
or U13563 (N_13563,N_7594,N_9394);
xnor U13564 (N_13564,N_5622,N_6447);
xor U13565 (N_13565,N_7431,N_6850);
nor U13566 (N_13566,N_6846,N_6316);
and U13567 (N_13567,N_6015,N_7431);
xnor U13568 (N_13568,N_9658,N_5821);
xor U13569 (N_13569,N_8749,N_9482);
nand U13570 (N_13570,N_7004,N_5481);
nor U13571 (N_13571,N_9402,N_7927);
nor U13572 (N_13572,N_5322,N_8134);
and U13573 (N_13573,N_6809,N_5499);
xor U13574 (N_13574,N_6706,N_9535);
or U13575 (N_13575,N_5387,N_9993);
nand U13576 (N_13576,N_8261,N_9561);
xor U13577 (N_13577,N_6787,N_8281);
xor U13578 (N_13578,N_9218,N_7908);
nor U13579 (N_13579,N_7000,N_5937);
nand U13580 (N_13580,N_9452,N_8868);
and U13581 (N_13581,N_5226,N_7359);
nor U13582 (N_13582,N_7352,N_5357);
or U13583 (N_13583,N_7831,N_7334);
and U13584 (N_13584,N_9060,N_6773);
xor U13585 (N_13585,N_6428,N_5951);
nor U13586 (N_13586,N_5020,N_8167);
nand U13587 (N_13587,N_7456,N_9083);
nand U13588 (N_13588,N_6714,N_7404);
or U13589 (N_13589,N_7410,N_8062);
nor U13590 (N_13590,N_6113,N_6544);
xor U13591 (N_13591,N_5156,N_5846);
or U13592 (N_13592,N_9969,N_6820);
and U13593 (N_13593,N_8552,N_6756);
xor U13594 (N_13594,N_7846,N_6146);
nand U13595 (N_13595,N_8312,N_5772);
nand U13596 (N_13596,N_7878,N_7903);
and U13597 (N_13597,N_6748,N_6593);
nand U13598 (N_13598,N_8263,N_7332);
nand U13599 (N_13599,N_6244,N_5650);
nand U13600 (N_13600,N_7986,N_9302);
nand U13601 (N_13601,N_9845,N_9958);
and U13602 (N_13602,N_8947,N_8090);
xnor U13603 (N_13603,N_6089,N_7311);
nand U13604 (N_13604,N_5355,N_6842);
and U13605 (N_13605,N_6111,N_5509);
nor U13606 (N_13606,N_6939,N_6571);
nand U13607 (N_13607,N_7694,N_5583);
xnor U13608 (N_13608,N_7047,N_9177);
and U13609 (N_13609,N_6879,N_8686);
and U13610 (N_13610,N_8083,N_7715);
or U13611 (N_13611,N_9135,N_6020);
and U13612 (N_13612,N_7652,N_6321);
nand U13613 (N_13613,N_7467,N_6175);
xnor U13614 (N_13614,N_7806,N_9136);
and U13615 (N_13615,N_5966,N_9961);
xnor U13616 (N_13616,N_5806,N_6794);
or U13617 (N_13617,N_7442,N_7326);
and U13618 (N_13618,N_6309,N_9834);
and U13619 (N_13619,N_5263,N_9224);
nand U13620 (N_13620,N_8943,N_8508);
and U13621 (N_13621,N_5335,N_6533);
nor U13622 (N_13622,N_8099,N_7154);
and U13623 (N_13623,N_8524,N_7295);
xor U13624 (N_13624,N_9022,N_7341);
and U13625 (N_13625,N_5381,N_6606);
nor U13626 (N_13626,N_9020,N_6222);
xnor U13627 (N_13627,N_5985,N_6975);
nand U13628 (N_13628,N_8425,N_9937);
xor U13629 (N_13629,N_8719,N_8915);
or U13630 (N_13630,N_5267,N_6287);
nor U13631 (N_13631,N_8888,N_8790);
nand U13632 (N_13632,N_8234,N_7058);
or U13633 (N_13633,N_5093,N_9961);
nor U13634 (N_13634,N_7474,N_7799);
nor U13635 (N_13635,N_5878,N_9920);
or U13636 (N_13636,N_9006,N_7480);
and U13637 (N_13637,N_5494,N_5856);
nand U13638 (N_13638,N_8780,N_9497);
and U13639 (N_13639,N_9191,N_9151);
and U13640 (N_13640,N_6590,N_6060);
or U13641 (N_13641,N_7839,N_5183);
xnor U13642 (N_13642,N_9799,N_9420);
or U13643 (N_13643,N_8295,N_7766);
and U13644 (N_13644,N_6066,N_9532);
xnor U13645 (N_13645,N_5600,N_9830);
and U13646 (N_13646,N_8013,N_9893);
xnor U13647 (N_13647,N_9690,N_8105);
nand U13648 (N_13648,N_9397,N_7244);
nor U13649 (N_13649,N_8352,N_5578);
xor U13650 (N_13650,N_5149,N_7357);
nand U13651 (N_13651,N_8288,N_7581);
or U13652 (N_13652,N_6684,N_8549);
nor U13653 (N_13653,N_6643,N_9517);
and U13654 (N_13654,N_7960,N_7040);
nor U13655 (N_13655,N_6849,N_6124);
and U13656 (N_13656,N_8630,N_9724);
xor U13657 (N_13657,N_5944,N_7111);
and U13658 (N_13658,N_5835,N_8085);
xnor U13659 (N_13659,N_5272,N_6140);
nor U13660 (N_13660,N_7298,N_5190);
xor U13661 (N_13661,N_5477,N_7999);
xnor U13662 (N_13662,N_6203,N_7178);
nand U13663 (N_13663,N_9691,N_6496);
nand U13664 (N_13664,N_8529,N_7208);
nor U13665 (N_13665,N_8401,N_5106);
or U13666 (N_13666,N_7151,N_7033);
and U13667 (N_13667,N_8508,N_9446);
nor U13668 (N_13668,N_6136,N_9489);
or U13669 (N_13669,N_5980,N_8308);
xnor U13670 (N_13670,N_6581,N_8643);
nor U13671 (N_13671,N_9964,N_7229);
nor U13672 (N_13672,N_6443,N_7784);
nand U13673 (N_13673,N_9552,N_5396);
or U13674 (N_13674,N_9550,N_6984);
xor U13675 (N_13675,N_9424,N_6634);
nand U13676 (N_13676,N_9905,N_5734);
nand U13677 (N_13677,N_8442,N_6079);
or U13678 (N_13678,N_9774,N_7379);
and U13679 (N_13679,N_8612,N_7524);
and U13680 (N_13680,N_8077,N_8664);
nor U13681 (N_13681,N_7247,N_5196);
and U13682 (N_13682,N_7328,N_7619);
and U13683 (N_13683,N_6126,N_8061);
nor U13684 (N_13684,N_7808,N_6760);
and U13685 (N_13685,N_8869,N_9894);
nand U13686 (N_13686,N_5366,N_5114);
and U13687 (N_13687,N_7710,N_8103);
nor U13688 (N_13688,N_6980,N_9470);
nand U13689 (N_13689,N_8413,N_6315);
and U13690 (N_13690,N_9983,N_9636);
nand U13691 (N_13691,N_8812,N_8499);
nand U13692 (N_13692,N_5957,N_8428);
nor U13693 (N_13693,N_5984,N_5599);
xor U13694 (N_13694,N_5443,N_5735);
nor U13695 (N_13695,N_9142,N_8397);
and U13696 (N_13696,N_7045,N_9253);
xnor U13697 (N_13697,N_5875,N_5614);
or U13698 (N_13698,N_5285,N_7262);
and U13699 (N_13699,N_5941,N_6591);
or U13700 (N_13700,N_5634,N_9542);
and U13701 (N_13701,N_8706,N_9844);
and U13702 (N_13702,N_5122,N_7846);
xnor U13703 (N_13703,N_9171,N_9113);
nand U13704 (N_13704,N_9907,N_9290);
or U13705 (N_13705,N_8810,N_7504);
or U13706 (N_13706,N_7949,N_5423);
and U13707 (N_13707,N_5681,N_9198);
xor U13708 (N_13708,N_7795,N_8533);
nor U13709 (N_13709,N_8234,N_6973);
or U13710 (N_13710,N_7751,N_9320);
nand U13711 (N_13711,N_5972,N_8059);
or U13712 (N_13712,N_9791,N_8302);
and U13713 (N_13713,N_6112,N_5646);
or U13714 (N_13714,N_5815,N_6984);
xnor U13715 (N_13715,N_9820,N_5929);
nor U13716 (N_13716,N_9991,N_5988);
nand U13717 (N_13717,N_5234,N_9833);
or U13718 (N_13718,N_9838,N_6644);
nand U13719 (N_13719,N_5041,N_7223);
nor U13720 (N_13720,N_8489,N_6446);
or U13721 (N_13721,N_8532,N_5897);
nand U13722 (N_13722,N_9790,N_7213);
and U13723 (N_13723,N_7381,N_8368);
nor U13724 (N_13724,N_6027,N_5537);
nor U13725 (N_13725,N_9438,N_8658);
and U13726 (N_13726,N_8900,N_9543);
nand U13727 (N_13727,N_7023,N_6415);
nand U13728 (N_13728,N_8570,N_8843);
xor U13729 (N_13729,N_8660,N_8321);
and U13730 (N_13730,N_7851,N_5543);
and U13731 (N_13731,N_9028,N_8411);
or U13732 (N_13732,N_9035,N_5051);
nor U13733 (N_13733,N_6857,N_8037);
nand U13734 (N_13734,N_5080,N_8959);
and U13735 (N_13735,N_9322,N_7389);
nand U13736 (N_13736,N_9495,N_9181);
xor U13737 (N_13737,N_8381,N_9154);
nor U13738 (N_13738,N_9500,N_5495);
xor U13739 (N_13739,N_7700,N_9925);
nand U13740 (N_13740,N_8161,N_8081);
or U13741 (N_13741,N_5795,N_5300);
or U13742 (N_13742,N_8512,N_5412);
nor U13743 (N_13743,N_7429,N_9201);
and U13744 (N_13744,N_8346,N_7189);
nor U13745 (N_13745,N_7998,N_5719);
nor U13746 (N_13746,N_8436,N_7390);
and U13747 (N_13747,N_7317,N_6452);
xnor U13748 (N_13748,N_9979,N_8630);
or U13749 (N_13749,N_7520,N_6038);
nor U13750 (N_13750,N_5167,N_9967);
nand U13751 (N_13751,N_6598,N_6146);
or U13752 (N_13752,N_7414,N_8001);
and U13753 (N_13753,N_6926,N_9156);
nor U13754 (N_13754,N_9535,N_6135);
xnor U13755 (N_13755,N_7879,N_7836);
and U13756 (N_13756,N_7333,N_5240);
nand U13757 (N_13757,N_7918,N_6976);
and U13758 (N_13758,N_6554,N_9945);
and U13759 (N_13759,N_7374,N_6446);
and U13760 (N_13760,N_8983,N_9098);
or U13761 (N_13761,N_6150,N_7626);
nor U13762 (N_13762,N_8997,N_9901);
or U13763 (N_13763,N_9217,N_5752);
xor U13764 (N_13764,N_8824,N_5399);
or U13765 (N_13765,N_9275,N_5571);
or U13766 (N_13766,N_8638,N_9730);
or U13767 (N_13767,N_6889,N_5817);
and U13768 (N_13768,N_9838,N_5703);
nand U13769 (N_13769,N_5003,N_7634);
and U13770 (N_13770,N_8276,N_6423);
nand U13771 (N_13771,N_6460,N_6342);
nor U13772 (N_13772,N_7045,N_6779);
nand U13773 (N_13773,N_8341,N_8077);
nor U13774 (N_13774,N_5185,N_6614);
nand U13775 (N_13775,N_5705,N_9388);
nor U13776 (N_13776,N_7368,N_9613);
nand U13777 (N_13777,N_9705,N_6202);
xnor U13778 (N_13778,N_5981,N_8239);
xor U13779 (N_13779,N_7062,N_8371);
xor U13780 (N_13780,N_6063,N_7375);
nand U13781 (N_13781,N_8206,N_5488);
and U13782 (N_13782,N_7698,N_8391);
nor U13783 (N_13783,N_7327,N_7554);
nand U13784 (N_13784,N_5629,N_7068);
nor U13785 (N_13785,N_7066,N_7822);
nor U13786 (N_13786,N_7912,N_8257);
xor U13787 (N_13787,N_6783,N_8274);
nor U13788 (N_13788,N_8257,N_5186);
nand U13789 (N_13789,N_6530,N_9647);
or U13790 (N_13790,N_9333,N_6689);
and U13791 (N_13791,N_9355,N_5826);
nand U13792 (N_13792,N_5856,N_9917);
or U13793 (N_13793,N_6611,N_6271);
and U13794 (N_13794,N_6406,N_9964);
xor U13795 (N_13795,N_7444,N_9251);
and U13796 (N_13796,N_9294,N_6832);
nor U13797 (N_13797,N_6802,N_7806);
nand U13798 (N_13798,N_7253,N_7992);
and U13799 (N_13799,N_6453,N_7911);
xnor U13800 (N_13800,N_9645,N_8267);
nand U13801 (N_13801,N_7807,N_6299);
nand U13802 (N_13802,N_5799,N_8638);
and U13803 (N_13803,N_9387,N_7701);
nand U13804 (N_13804,N_6342,N_6584);
or U13805 (N_13805,N_5375,N_8528);
xor U13806 (N_13806,N_7416,N_6757);
and U13807 (N_13807,N_7148,N_6139);
nand U13808 (N_13808,N_9604,N_7090);
or U13809 (N_13809,N_5555,N_8622);
or U13810 (N_13810,N_7562,N_5600);
nor U13811 (N_13811,N_9755,N_8837);
or U13812 (N_13812,N_9503,N_9853);
or U13813 (N_13813,N_8253,N_8344);
xnor U13814 (N_13814,N_7379,N_9654);
nor U13815 (N_13815,N_7034,N_9678);
or U13816 (N_13816,N_9905,N_6118);
nor U13817 (N_13817,N_9029,N_7395);
or U13818 (N_13818,N_5250,N_5275);
nor U13819 (N_13819,N_9818,N_6906);
nor U13820 (N_13820,N_7212,N_5847);
xor U13821 (N_13821,N_9292,N_7521);
xnor U13822 (N_13822,N_5187,N_9837);
nand U13823 (N_13823,N_9136,N_5639);
nor U13824 (N_13824,N_7483,N_6664);
and U13825 (N_13825,N_5714,N_9812);
and U13826 (N_13826,N_5703,N_7595);
and U13827 (N_13827,N_5418,N_5319);
xor U13828 (N_13828,N_6879,N_9526);
nor U13829 (N_13829,N_9642,N_6050);
nor U13830 (N_13830,N_7927,N_8055);
or U13831 (N_13831,N_8971,N_6604);
nor U13832 (N_13832,N_6659,N_5327);
or U13833 (N_13833,N_6763,N_9812);
nor U13834 (N_13834,N_6537,N_6878);
nor U13835 (N_13835,N_5292,N_8924);
nand U13836 (N_13836,N_5147,N_6204);
or U13837 (N_13837,N_6514,N_9490);
xnor U13838 (N_13838,N_8695,N_5181);
nor U13839 (N_13839,N_6503,N_7001);
and U13840 (N_13840,N_9553,N_5586);
and U13841 (N_13841,N_7754,N_6740);
or U13842 (N_13842,N_5255,N_7643);
xor U13843 (N_13843,N_5089,N_8230);
nor U13844 (N_13844,N_5886,N_7273);
xnor U13845 (N_13845,N_9928,N_9884);
or U13846 (N_13846,N_7866,N_6481);
nand U13847 (N_13847,N_6302,N_8453);
or U13848 (N_13848,N_9282,N_8382);
nand U13849 (N_13849,N_7451,N_9230);
nand U13850 (N_13850,N_9912,N_8422);
and U13851 (N_13851,N_9082,N_6459);
or U13852 (N_13852,N_6160,N_6806);
nand U13853 (N_13853,N_6818,N_8607);
xor U13854 (N_13854,N_7657,N_5959);
and U13855 (N_13855,N_7707,N_8480);
and U13856 (N_13856,N_7776,N_8367);
nor U13857 (N_13857,N_5104,N_8745);
xnor U13858 (N_13858,N_7948,N_5587);
nor U13859 (N_13859,N_6137,N_6183);
and U13860 (N_13860,N_6164,N_7929);
or U13861 (N_13861,N_8989,N_7330);
xor U13862 (N_13862,N_5732,N_7979);
nand U13863 (N_13863,N_8803,N_8412);
nand U13864 (N_13864,N_8465,N_7028);
and U13865 (N_13865,N_6106,N_6006);
and U13866 (N_13866,N_9854,N_6576);
nand U13867 (N_13867,N_9560,N_8262);
nor U13868 (N_13868,N_7438,N_9800);
or U13869 (N_13869,N_5066,N_7947);
nand U13870 (N_13870,N_9670,N_5201);
nor U13871 (N_13871,N_8341,N_6958);
xnor U13872 (N_13872,N_7772,N_7406);
and U13873 (N_13873,N_9617,N_7899);
nor U13874 (N_13874,N_8033,N_6128);
nand U13875 (N_13875,N_7474,N_8630);
xor U13876 (N_13876,N_6849,N_6822);
xnor U13877 (N_13877,N_6761,N_8860);
or U13878 (N_13878,N_5522,N_6828);
xnor U13879 (N_13879,N_9168,N_8325);
xor U13880 (N_13880,N_6676,N_6124);
and U13881 (N_13881,N_9151,N_8203);
xor U13882 (N_13882,N_7719,N_6095);
and U13883 (N_13883,N_8407,N_5528);
nand U13884 (N_13884,N_8366,N_9710);
xnor U13885 (N_13885,N_5169,N_7824);
xor U13886 (N_13886,N_8929,N_5168);
xor U13887 (N_13887,N_8537,N_8341);
nor U13888 (N_13888,N_9430,N_8515);
nand U13889 (N_13889,N_7874,N_7887);
nand U13890 (N_13890,N_9827,N_6855);
or U13891 (N_13891,N_6373,N_6710);
nand U13892 (N_13892,N_6691,N_5683);
or U13893 (N_13893,N_5373,N_8746);
or U13894 (N_13894,N_5206,N_7182);
nor U13895 (N_13895,N_7842,N_6266);
nand U13896 (N_13896,N_9583,N_7888);
xor U13897 (N_13897,N_9051,N_6844);
or U13898 (N_13898,N_6476,N_6143);
or U13899 (N_13899,N_7381,N_9949);
xnor U13900 (N_13900,N_6243,N_9443);
nand U13901 (N_13901,N_6156,N_7921);
nor U13902 (N_13902,N_5828,N_8144);
xor U13903 (N_13903,N_7832,N_8072);
or U13904 (N_13904,N_7148,N_7916);
nand U13905 (N_13905,N_8784,N_7612);
and U13906 (N_13906,N_6404,N_7819);
or U13907 (N_13907,N_5337,N_8347);
nor U13908 (N_13908,N_5880,N_6971);
and U13909 (N_13909,N_7658,N_5461);
xnor U13910 (N_13910,N_5310,N_5890);
nand U13911 (N_13911,N_5273,N_7798);
and U13912 (N_13912,N_9815,N_7407);
or U13913 (N_13913,N_7344,N_9340);
or U13914 (N_13914,N_8146,N_6021);
and U13915 (N_13915,N_8980,N_7663);
and U13916 (N_13916,N_5649,N_8982);
and U13917 (N_13917,N_7797,N_8409);
nand U13918 (N_13918,N_7028,N_8851);
or U13919 (N_13919,N_9511,N_6169);
xnor U13920 (N_13920,N_6011,N_8477);
nand U13921 (N_13921,N_9946,N_8190);
nand U13922 (N_13922,N_5789,N_8696);
and U13923 (N_13923,N_7109,N_8108);
nor U13924 (N_13924,N_5688,N_5914);
nand U13925 (N_13925,N_7265,N_8381);
and U13926 (N_13926,N_8307,N_5027);
and U13927 (N_13927,N_8564,N_9343);
nor U13928 (N_13928,N_5303,N_9599);
xor U13929 (N_13929,N_9197,N_5845);
nor U13930 (N_13930,N_8433,N_8307);
nand U13931 (N_13931,N_9321,N_7069);
or U13932 (N_13932,N_6518,N_6635);
xor U13933 (N_13933,N_5338,N_9997);
and U13934 (N_13934,N_7597,N_9045);
nand U13935 (N_13935,N_7285,N_6613);
nand U13936 (N_13936,N_8066,N_6939);
and U13937 (N_13937,N_8802,N_8576);
nand U13938 (N_13938,N_5113,N_7118);
xnor U13939 (N_13939,N_6819,N_7095);
nand U13940 (N_13940,N_7927,N_8003);
nand U13941 (N_13941,N_5493,N_5174);
or U13942 (N_13942,N_7772,N_7719);
or U13943 (N_13943,N_5241,N_8605);
nand U13944 (N_13944,N_7391,N_7076);
and U13945 (N_13945,N_9386,N_9199);
and U13946 (N_13946,N_5747,N_8540);
nand U13947 (N_13947,N_9270,N_7128);
nand U13948 (N_13948,N_7279,N_5233);
xnor U13949 (N_13949,N_5217,N_9012);
nor U13950 (N_13950,N_7569,N_5473);
or U13951 (N_13951,N_5596,N_7818);
or U13952 (N_13952,N_9092,N_6550);
nor U13953 (N_13953,N_5227,N_9185);
nor U13954 (N_13954,N_6524,N_7389);
nand U13955 (N_13955,N_5805,N_7135);
nor U13956 (N_13956,N_5890,N_8358);
nor U13957 (N_13957,N_7968,N_6651);
nand U13958 (N_13958,N_5980,N_7664);
and U13959 (N_13959,N_5398,N_7983);
nor U13960 (N_13960,N_5422,N_5123);
and U13961 (N_13961,N_9790,N_6708);
nor U13962 (N_13962,N_8917,N_8182);
or U13963 (N_13963,N_5010,N_5758);
nand U13964 (N_13964,N_5489,N_5735);
nor U13965 (N_13965,N_5656,N_7669);
xor U13966 (N_13966,N_7819,N_5769);
nand U13967 (N_13967,N_9644,N_7412);
nand U13968 (N_13968,N_5718,N_9552);
and U13969 (N_13969,N_9037,N_9492);
or U13970 (N_13970,N_7458,N_8623);
nand U13971 (N_13971,N_7412,N_6640);
xor U13972 (N_13972,N_6635,N_9371);
nor U13973 (N_13973,N_5274,N_8879);
nand U13974 (N_13974,N_5874,N_5945);
or U13975 (N_13975,N_5567,N_6701);
or U13976 (N_13976,N_9802,N_8718);
nand U13977 (N_13977,N_9669,N_9009);
nand U13978 (N_13978,N_8636,N_7138);
nor U13979 (N_13979,N_7729,N_9640);
xor U13980 (N_13980,N_5757,N_7251);
xnor U13981 (N_13981,N_6460,N_7367);
xnor U13982 (N_13982,N_9193,N_7105);
and U13983 (N_13983,N_8631,N_5309);
nor U13984 (N_13984,N_5292,N_6090);
or U13985 (N_13985,N_5022,N_6044);
or U13986 (N_13986,N_5262,N_8044);
xor U13987 (N_13987,N_5515,N_5092);
or U13988 (N_13988,N_8636,N_6578);
nand U13989 (N_13989,N_6727,N_5610);
nor U13990 (N_13990,N_7192,N_7756);
nand U13991 (N_13991,N_5703,N_9631);
nand U13992 (N_13992,N_7508,N_6033);
or U13993 (N_13993,N_6041,N_6438);
or U13994 (N_13994,N_8718,N_9289);
nand U13995 (N_13995,N_6098,N_5646);
xnor U13996 (N_13996,N_7738,N_7536);
xnor U13997 (N_13997,N_9167,N_9360);
xor U13998 (N_13998,N_8763,N_6033);
or U13999 (N_13999,N_7723,N_9199);
or U14000 (N_14000,N_8226,N_8896);
or U14001 (N_14001,N_5984,N_6485);
and U14002 (N_14002,N_9419,N_6453);
xnor U14003 (N_14003,N_7920,N_6386);
or U14004 (N_14004,N_6351,N_8457);
nand U14005 (N_14005,N_9556,N_9348);
nand U14006 (N_14006,N_6771,N_9110);
and U14007 (N_14007,N_5941,N_8216);
xnor U14008 (N_14008,N_9872,N_6192);
nor U14009 (N_14009,N_6710,N_5241);
nand U14010 (N_14010,N_7233,N_9200);
and U14011 (N_14011,N_9238,N_7325);
or U14012 (N_14012,N_9568,N_8448);
xnor U14013 (N_14013,N_5282,N_6283);
nor U14014 (N_14014,N_6412,N_8647);
nor U14015 (N_14015,N_5276,N_8976);
nor U14016 (N_14016,N_9485,N_6188);
or U14017 (N_14017,N_7778,N_7929);
xor U14018 (N_14018,N_6301,N_6253);
and U14019 (N_14019,N_8566,N_8816);
or U14020 (N_14020,N_7576,N_5782);
or U14021 (N_14021,N_8097,N_9303);
and U14022 (N_14022,N_9348,N_6773);
or U14023 (N_14023,N_9219,N_7179);
xor U14024 (N_14024,N_7725,N_7861);
nor U14025 (N_14025,N_7641,N_6986);
or U14026 (N_14026,N_7398,N_6166);
nor U14027 (N_14027,N_9063,N_7600);
and U14028 (N_14028,N_9126,N_5544);
nor U14029 (N_14029,N_9271,N_7878);
and U14030 (N_14030,N_8062,N_8293);
and U14031 (N_14031,N_9733,N_9871);
xnor U14032 (N_14032,N_9685,N_7690);
or U14033 (N_14033,N_5403,N_9457);
xor U14034 (N_14034,N_8458,N_5323);
xor U14035 (N_14035,N_6870,N_6435);
or U14036 (N_14036,N_7572,N_8732);
nor U14037 (N_14037,N_7949,N_9589);
xor U14038 (N_14038,N_8273,N_6101);
and U14039 (N_14039,N_7440,N_7139);
nand U14040 (N_14040,N_6208,N_6723);
nor U14041 (N_14041,N_6503,N_5699);
xnor U14042 (N_14042,N_6419,N_5635);
or U14043 (N_14043,N_8796,N_8400);
nand U14044 (N_14044,N_9170,N_8228);
and U14045 (N_14045,N_6351,N_6865);
nor U14046 (N_14046,N_5559,N_8071);
nor U14047 (N_14047,N_6738,N_9661);
or U14048 (N_14048,N_7169,N_6509);
nand U14049 (N_14049,N_6727,N_5745);
and U14050 (N_14050,N_9731,N_6989);
xnor U14051 (N_14051,N_6951,N_7270);
xor U14052 (N_14052,N_6609,N_8140);
nor U14053 (N_14053,N_6868,N_8673);
or U14054 (N_14054,N_8549,N_7845);
nand U14055 (N_14055,N_8853,N_8963);
nand U14056 (N_14056,N_6849,N_6651);
nor U14057 (N_14057,N_9583,N_6976);
xnor U14058 (N_14058,N_8320,N_5991);
nor U14059 (N_14059,N_8685,N_6744);
xnor U14060 (N_14060,N_9927,N_5501);
and U14061 (N_14061,N_5560,N_6059);
nor U14062 (N_14062,N_7713,N_6524);
nand U14063 (N_14063,N_9429,N_5975);
or U14064 (N_14064,N_9978,N_9283);
or U14065 (N_14065,N_9782,N_9575);
nand U14066 (N_14066,N_5552,N_7272);
or U14067 (N_14067,N_7592,N_7521);
xnor U14068 (N_14068,N_7906,N_7421);
or U14069 (N_14069,N_9334,N_9567);
nand U14070 (N_14070,N_6409,N_5851);
xnor U14071 (N_14071,N_6482,N_5949);
xor U14072 (N_14072,N_9174,N_6719);
nor U14073 (N_14073,N_8158,N_8956);
xnor U14074 (N_14074,N_9033,N_6537);
nor U14075 (N_14075,N_5624,N_5912);
xnor U14076 (N_14076,N_7179,N_9560);
or U14077 (N_14077,N_8256,N_8300);
nor U14078 (N_14078,N_6450,N_6881);
nor U14079 (N_14079,N_7903,N_7219);
nand U14080 (N_14080,N_7914,N_8728);
nor U14081 (N_14081,N_6588,N_6896);
or U14082 (N_14082,N_7329,N_8137);
xor U14083 (N_14083,N_7573,N_9790);
nor U14084 (N_14084,N_6780,N_8604);
nor U14085 (N_14085,N_9620,N_5423);
xor U14086 (N_14086,N_8727,N_7560);
or U14087 (N_14087,N_8503,N_7738);
or U14088 (N_14088,N_8108,N_7727);
xor U14089 (N_14089,N_7543,N_8275);
or U14090 (N_14090,N_6940,N_9946);
nand U14091 (N_14091,N_7603,N_8507);
and U14092 (N_14092,N_8185,N_5336);
or U14093 (N_14093,N_8843,N_9475);
or U14094 (N_14094,N_9283,N_7888);
xor U14095 (N_14095,N_6890,N_8812);
and U14096 (N_14096,N_8799,N_7795);
or U14097 (N_14097,N_6992,N_5839);
or U14098 (N_14098,N_6022,N_5407);
xnor U14099 (N_14099,N_7815,N_6389);
nor U14100 (N_14100,N_8947,N_7353);
xnor U14101 (N_14101,N_6304,N_9521);
and U14102 (N_14102,N_6923,N_9697);
and U14103 (N_14103,N_6364,N_8859);
nor U14104 (N_14104,N_7961,N_6272);
or U14105 (N_14105,N_6324,N_7875);
or U14106 (N_14106,N_6843,N_8597);
or U14107 (N_14107,N_6662,N_6954);
or U14108 (N_14108,N_8970,N_8842);
or U14109 (N_14109,N_8671,N_6873);
and U14110 (N_14110,N_9458,N_8434);
nand U14111 (N_14111,N_8179,N_6837);
and U14112 (N_14112,N_9809,N_7675);
xnor U14113 (N_14113,N_7782,N_8479);
nand U14114 (N_14114,N_5140,N_7056);
xnor U14115 (N_14115,N_9712,N_9468);
nand U14116 (N_14116,N_7085,N_6082);
or U14117 (N_14117,N_7382,N_7395);
or U14118 (N_14118,N_6399,N_5363);
nor U14119 (N_14119,N_9340,N_6127);
nand U14120 (N_14120,N_9722,N_9791);
or U14121 (N_14121,N_5614,N_7723);
or U14122 (N_14122,N_8798,N_5252);
or U14123 (N_14123,N_6204,N_8438);
xor U14124 (N_14124,N_8401,N_5836);
or U14125 (N_14125,N_5209,N_8630);
and U14126 (N_14126,N_8983,N_9583);
and U14127 (N_14127,N_5088,N_7050);
nor U14128 (N_14128,N_7700,N_9173);
and U14129 (N_14129,N_5242,N_8150);
and U14130 (N_14130,N_8191,N_8403);
nor U14131 (N_14131,N_9175,N_8975);
and U14132 (N_14132,N_7302,N_7054);
or U14133 (N_14133,N_8055,N_6796);
nor U14134 (N_14134,N_8920,N_5706);
nor U14135 (N_14135,N_9091,N_5645);
nor U14136 (N_14136,N_5374,N_7987);
nand U14137 (N_14137,N_5525,N_8019);
nor U14138 (N_14138,N_8909,N_8952);
xor U14139 (N_14139,N_8281,N_5830);
nand U14140 (N_14140,N_5778,N_5250);
nand U14141 (N_14141,N_7098,N_5459);
and U14142 (N_14142,N_9944,N_9760);
or U14143 (N_14143,N_6883,N_8277);
nand U14144 (N_14144,N_6884,N_8098);
xor U14145 (N_14145,N_9482,N_7182);
nor U14146 (N_14146,N_5855,N_7136);
or U14147 (N_14147,N_9437,N_7591);
nor U14148 (N_14148,N_7585,N_8527);
xor U14149 (N_14149,N_8524,N_9084);
xnor U14150 (N_14150,N_6085,N_8651);
nand U14151 (N_14151,N_7136,N_9739);
nand U14152 (N_14152,N_6903,N_8183);
or U14153 (N_14153,N_8453,N_6037);
xnor U14154 (N_14154,N_5080,N_7823);
and U14155 (N_14155,N_7093,N_5419);
nor U14156 (N_14156,N_5896,N_9081);
or U14157 (N_14157,N_7003,N_9136);
or U14158 (N_14158,N_9218,N_5640);
xnor U14159 (N_14159,N_9118,N_8599);
nand U14160 (N_14160,N_5767,N_7785);
and U14161 (N_14161,N_5075,N_9624);
nand U14162 (N_14162,N_5425,N_5256);
or U14163 (N_14163,N_5013,N_8911);
nor U14164 (N_14164,N_7639,N_8065);
and U14165 (N_14165,N_5657,N_9057);
nand U14166 (N_14166,N_9563,N_9147);
and U14167 (N_14167,N_8764,N_7097);
nor U14168 (N_14168,N_7562,N_5351);
or U14169 (N_14169,N_5856,N_9012);
or U14170 (N_14170,N_5912,N_5817);
xnor U14171 (N_14171,N_6725,N_8414);
nand U14172 (N_14172,N_6954,N_5754);
and U14173 (N_14173,N_6589,N_5776);
or U14174 (N_14174,N_6400,N_6770);
nor U14175 (N_14175,N_5582,N_6001);
xnor U14176 (N_14176,N_6101,N_9221);
or U14177 (N_14177,N_6843,N_5000);
nand U14178 (N_14178,N_9137,N_9401);
and U14179 (N_14179,N_8614,N_6272);
and U14180 (N_14180,N_5083,N_8863);
xnor U14181 (N_14181,N_7683,N_7124);
nor U14182 (N_14182,N_7928,N_7275);
and U14183 (N_14183,N_5198,N_6167);
or U14184 (N_14184,N_8239,N_5527);
nand U14185 (N_14185,N_5495,N_7725);
or U14186 (N_14186,N_5792,N_6272);
or U14187 (N_14187,N_9305,N_6550);
xor U14188 (N_14188,N_8564,N_8213);
xnor U14189 (N_14189,N_6324,N_7644);
xor U14190 (N_14190,N_7962,N_5639);
and U14191 (N_14191,N_5077,N_8704);
nand U14192 (N_14192,N_8155,N_7263);
nand U14193 (N_14193,N_6402,N_7948);
and U14194 (N_14194,N_7862,N_5415);
or U14195 (N_14195,N_5714,N_6870);
xnor U14196 (N_14196,N_6083,N_7297);
xnor U14197 (N_14197,N_5112,N_7471);
xor U14198 (N_14198,N_9897,N_8866);
and U14199 (N_14199,N_9292,N_5479);
and U14200 (N_14200,N_6092,N_7867);
nor U14201 (N_14201,N_7907,N_6127);
nor U14202 (N_14202,N_8776,N_6971);
nor U14203 (N_14203,N_8987,N_6182);
or U14204 (N_14204,N_8114,N_8729);
or U14205 (N_14205,N_6707,N_8519);
or U14206 (N_14206,N_6713,N_5347);
or U14207 (N_14207,N_8848,N_6289);
nor U14208 (N_14208,N_5507,N_7273);
xor U14209 (N_14209,N_6928,N_7612);
nor U14210 (N_14210,N_6451,N_5678);
or U14211 (N_14211,N_6086,N_8317);
nor U14212 (N_14212,N_5188,N_8052);
nor U14213 (N_14213,N_9019,N_5883);
nor U14214 (N_14214,N_8974,N_5531);
and U14215 (N_14215,N_8818,N_6769);
or U14216 (N_14216,N_8967,N_6728);
xor U14217 (N_14217,N_8155,N_9756);
nand U14218 (N_14218,N_7992,N_5835);
xor U14219 (N_14219,N_5841,N_5994);
nor U14220 (N_14220,N_8169,N_5973);
xnor U14221 (N_14221,N_6059,N_8929);
or U14222 (N_14222,N_9842,N_6016);
nand U14223 (N_14223,N_8199,N_5623);
nor U14224 (N_14224,N_9226,N_6582);
nor U14225 (N_14225,N_6842,N_6427);
xor U14226 (N_14226,N_8086,N_6396);
nand U14227 (N_14227,N_9163,N_9197);
nor U14228 (N_14228,N_8871,N_7672);
nand U14229 (N_14229,N_9511,N_8632);
and U14230 (N_14230,N_5722,N_6710);
nor U14231 (N_14231,N_7120,N_5360);
or U14232 (N_14232,N_5544,N_7296);
nor U14233 (N_14233,N_9208,N_6741);
or U14234 (N_14234,N_8920,N_5780);
nor U14235 (N_14235,N_7765,N_7150);
and U14236 (N_14236,N_7710,N_8105);
and U14237 (N_14237,N_9570,N_5464);
or U14238 (N_14238,N_7029,N_5478);
and U14239 (N_14239,N_8937,N_6628);
nand U14240 (N_14240,N_9594,N_9982);
nor U14241 (N_14241,N_5168,N_9928);
xor U14242 (N_14242,N_5177,N_5621);
nand U14243 (N_14243,N_8022,N_6462);
xor U14244 (N_14244,N_9822,N_5974);
nor U14245 (N_14245,N_5261,N_6869);
xnor U14246 (N_14246,N_9923,N_9641);
nor U14247 (N_14247,N_7007,N_9119);
or U14248 (N_14248,N_6041,N_8330);
nand U14249 (N_14249,N_8906,N_8405);
nand U14250 (N_14250,N_9459,N_7693);
nor U14251 (N_14251,N_7729,N_8621);
nand U14252 (N_14252,N_5600,N_9115);
nor U14253 (N_14253,N_7606,N_9530);
or U14254 (N_14254,N_7682,N_5486);
xnor U14255 (N_14255,N_6266,N_8772);
nand U14256 (N_14256,N_6286,N_8883);
or U14257 (N_14257,N_9194,N_8672);
xor U14258 (N_14258,N_9522,N_7961);
nand U14259 (N_14259,N_9902,N_8132);
nand U14260 (N_14260,N_9126,N_7060);
nor U14261 (N_14261,N_6317,N_7816);
nor U14262 (N_14262,N_9808,N_9767);
nand U14263 (N_14263,N_9128,N_7977);
xor U14264 (N_14264,N_8373,N_7328);
xor U14265 (N_14265,N_8642,N_8711);
and U14266 (N_14266,N_6535,N_8082);
xor U14267 (N_14267,N_9009,N_8706);
nand U14268 (N_14268,N_5148,N_8542);
nor U14269 (N_14269,N_9806,N_6951);
xnor U14270 (N_14270,N_7611,N_5693);
xnor U14271 (N_14271,N_8848,N_5797);
or U14272 (N_14272,N_5170,N_6999);
and U14273 (N_14273,N_6018,N_9466);
xor U14274 (N_14274,N_6954,N_7104);
xnor U14275 (N_14275,N_8056,N_6312);
nand U14276 (N_14276,N_9221,N_6882);
xnor U14277 (N_14277,N_5865,N_8117);
and U14278 (N_14278,N_9575,N_7504);
xnor U14279 (N_14279,N_7948,N_6404);
and U14280 (N_14280,N_8276,N_6916);
nor U14281 (N_14281,N_7849,N_8780);
and U14282 (N_14282,N_8816,N_9403);
or U14283 (N_14283,N_8541,N_5945);
and U14284 (N_14284,N_6407,N_5861);
nor U14285 (N_14285,N_6410,N_9533);
or U14286 (N_14286,N_9180,N_7370);
xnor U14287 (N_14287,N_9320,N_8440);
or U14288 (N_14288,N_7817,N_7708);
nand U14289 (N_14289,N_7590,N_7169);
nor U14290 (N_14290,N_7561,N_6260);
nor U14291 (N_14291,N_5148,N_5097);
or U14292 (N_14292,N_5666,N_6432);
nor U14293 (N_14293,N_6551,N_9286);
or U14294 (N_14294,N_5554,N_9260);
or U14295 (N_14295,N_7114,N_7028);
nor U14296 (N_14296,N_6928,N_7946);
or U14297 (N_14297,N_9727,N_5869);
nand U14298 (N_14298,N_8334,N_6928);
and U14299 (N_14299,N_5247,N_5476);
nor U14300 (N_14300,N_9827,N_6149);
and U14301 (N_14301,N_6226,N_6806);
or U14302 (N_14302,N_7845,N_6155);
and U14303 (N_14303,N_7381,N_6885);
or U14304 (N_14304,N_9463,N_7115);
xnor U14305 (N_14305,N_7016,N_6171);
or U14306 (N_14306,N_5727,N_9223);
xnor U14307 (N_14307,N_6249,N_7207);
and U14308 (N_14308,N_9801,N_9590);
and U14309 (N_14309,N_9156,N_8018);
xor U14310 (N_14310,N_5009,N_7474);
nand U14311 (N_14311,N_9826,N_7365);
or U14312 (N_14312,N_8585,N_7207);
xor U14313 (N_14313,N_9363,N_6583);
or U14314 (N_14314,N_6515,N_5637);
or U14315 (N_14315,N_9015,N_5395);
and U14316 (N_14316,N_6207,N_5902);
or U14317 (N_14317,N_7102,N_8431);
and U14318 (N_14318,N_5860,N_6489);
nand U14319 (N_14319,N_8804,N_6346);
nor U14320 (N_14320,N_8606,N_8774);
nand U14321 (N_14321,N_5019,N_5186);
nand U14322 (N_14322,N_7111,N_9403);
and U14323 (N_14323,N_5906,N_6798);
nand U14324 (N_14324,N_8378,N_9356);
or U14325 (N_14325,N_5258,N_7353);
or U14326 (N_14326,N_7703,N_8144);
or U14327 (N_14327,N_5469,N_8808);
and U14328 (N_14328,N_5951,N_5616);
nor U14329 (N_14329,N_8651,N_8009);
or U14330 (N_14330,N_8598,N_6592);
nand U14331 (N_14331,N_7042,N_9003);
nor U14332 (N_14332,N_7849,N_7180);
nand U14333 (N_14333,N_8920,N_9285);
xnor U14334 (N_14334,N_5685,N_6909);
and U14335 (N_14335,N_5695,N_7657);
nor U14336 (N_14336,N_9283,N_5153);
nor U14337 (N_14337,N_6589,N_5645);
and U14338 (N_14338,N_7693,N_8026);
xnor U14339 (N_14339,N_9350,N_7856);
xor U14340 (N_14340,N_7864,N_9584);
or U14341 (N_14341,N_6399,N_7838);
or U14342 (N_14342,N_8001,N_5067);
and U14343 (N_14343,N_9609,N_8549);
nand U14344 (N_14344,N_7986,N_5633);
or U14345 (N_14345,N_6803,N_9356);
xnor U14346 (N_14346,N_5424,N_9048);
and U14347 (N_14347,N_7836,N_9112);
and U14348 (N_14348,N_9829,N_8705);
nor U14349 (N_14349,N_9983,N_7930);
nor U14350 (N_14350,N_6371,N_6050);
xnor U14351 (N_14351,N_7575,N_9093);
or U14352 (N_14352,N_7679,N_6604);
nor U14353 (N_14353,N_5985,N_8194);
xnor U14354 (N_14354,N_5232,N_8620);
xnor U14355 (N_14355,N_8551,N_7942);
nor U14356 (N_14356,N_6728,N_5682);
xnor U14357 (N_14357,N_7381,N_6074);
xor U14358 (N_14358,N_7182,N_5520);
and U14359 (N_14359,N_7410,N_5784);
nand U14360 (N_14360,N_6507,N_6774);
xor U14361 (N_14361,N_6174,N_7246);
xnor U14362 (N_14362,N_9967,N_9146);
nor U14363 (N_14363,N_8021,N_9079);
or U14364 (N_14364,N_6678,N_5433);
nor U14365 (N_14365,N_9874,N_9641);
or U14366 (N_14366,N_7196,N_7008);
nor U14367 (N_14367,N_5786,N_5461);
nand U14368 (N_14368,N_7215,N_9443);
nand U14369 (N_14369,N_8003,N_5179);
nor U14370 (N_14370,N_9618,N_9798);
and U14371 (N_14371,N_5217,N_5589);
or U14372 (N_14372,N_6103,N_5444);
or U14373 (N_14373,N_9665,N_8193);
xnor U14374 (N_14374,N_9833,N_8865);
and U14375 (N_14375,N_9477,N_6147);
nor U14376 (N_14376,N_6913,N_5316);
and U14377 (N_14377,N_9548,N_7428);
or U14378 (N_14378,N_8237,N_7886);
nor U14379 (N_14379,N_5242,N_7398);
nand U14380 (N_14380,N_9983,N_6712);
xnor U14381 (N_14381,N_6692,N_8984);
nor U14382 (N_14382,N_7344,N_7545);
and U14383 (N_14383,N_9765,N_7737);
nand U14384 (N_14384,N_8977,N_9464);
xor U14385 (N_14385,N_9665,N_5708);
nor U14386 (N_14386,N_8251,N_5724);
or U14387 (N_14387,N_6908,N_9237);
xnor U14388 (N_14388,N_8925,N_9530);
nor U14389 (N_14389,N_5796,N_8028);
nor U14390 (N_14390,N_8586,N_5704);
nand U14391 (N_14391,N_8551,N_9285);
nor U14392 (N_14392,N_7157,N_7493);
nor U14393 (N_14393,N_8018,N_8803);
and U14394 (N_14394,N_6182,N_7236);
xnor U14395 (N_14395,N_7137,N_5713);
or U14396 (N_14396,N_8071,N_7827);
nor U14397 (N_14397,N_8927,N_5961);
and U14398 (N_14398,N_8349,N_8200);
and U14399 (N_14399,N_9946,N_6226);
and U14400 (N_14400,N_9822,N_5565);
and U14401 (N_14401,N_5195,N_6123);
nor U14402 (N_14402,N_8568,N_7154);
or U14403 (N_14403,N_7890,N_7059);
and U14404 (N_14404,N_5152,N_9373);
xor U14405 (N_14405,N_7991,N_7731);
nand U14406 (N_14406,N_7532,N_9712);
nand U14407 (N_14407,N_8434,N_6497);
nor U14408 (N_14408,N_5130,N_5444);
or U14409 (N_14409,N_5634,N_9340);
nor U14410 (N_14410,N_6109,N_5762);
or U14411 (N_14411,N_8519,N_8398);
or U14412 (N_14412,N_8595,N_9163);
nor U14413 (N_14413,N_5876,N_9268);
nand U14414 (N_14414,N_6085,N_7178);
and U14415 (N_14415,N_9022,N_6346);
nor U14416 (N_14416,N_9851,N_7533);
nor U14417 (N_14417,N_7118,N_5211);
xor U14418 (N_14418,N_7998,N_5446);
nor U14419 (N_14419,N_6863,N_7674);
xor U14420 (N_14420,N_5904,N_7756);
and U14421 (N_14421,N_7155,N_8171);
or U14422 (N_14422,N_5057,N_5907);
nor U14423 (N_14423,N_8909,N_6372);
or U14424 (N_14424,N_7108,N_7233);
or U14425 (N_14425,N_7023,N_5469);
or U14426 (N_14426,N_5501,N_7583);
nand U14427 (N_14427,N_7980,N_5770);
nand U14428 (N_14428,N_8790,N_8239);
nor U14429 (N_14429,N_9996,N_5659);
nand U14430 (N_14430,N_7937,N_8793);
xnor U14431 (N_14431,N_9101,N_7596);
and U14432 (N_14432,N_7598,N_7549);
nor U14433 (N_14433,N_9819,N_5050);
and U14434 (N_14434,N_7187,N_5545);
nor U14435 (N_14435,N_6624,N_8623);
or U14436 (N_14436,N_5643,N_8460);
nand U14437 (N_14437,N_5758,N_6221);
or U14438 (N_14438,N_8576,N_8929);
xor U14439 (N_14439,N_8565,N_9901);
xor U14440 (N_14440,N_7524,N_8694);
xor U14441 (N_14441,N_6476,N_7363);
nand U14442 (N_14442,N_8566,N_5960);
and U14443 (N_14443,N_9979,N_5949);
or U14444 (N_14444,N_6213,N_5993);
and U14445 (N_14445,N_6722,N_8698);
nand U14446 (N_14446,N_7337,N_6220);
xnor U14447 (N_14447,N_9134,N_5401);
nor U14448 (N_14448,N_5969,N_8739);
and U14449 (N_14449,N_5254,N_6169);
or U14450 (N_14450,N_8224,N_5484);
or U14451 (N_14451,N_9912,N_6995);
and U14452 (N_14452,N_6141,N_5291);
nor U14453 (N_14453,N_7333,N_6879);
nand U14454 (N_14454,N_5980,N_9767);
nor U14455 (N_14455,N_7064,N_6355);
and U14456 (N_14456,N_8642,N_8569);
nand U14457 (N_14457,N_6173,N_9424);
or U14458 (N_14458,N_7676,N_8578);
xnor U14459 (N_14459,N_7870,N_9976);
nand U14460 (N_14460,N_5337,N_8381);
and U14461 (N_14461,N_9608,N_9406);
or U14462 (N_14462,N_6527,N_8128);
xor U14463 (N_14463,N_7395,N_6481);
and U14464 (N_14464,N_9942,N_9616);
nor U14465 (N_14465,N_8028,N_7693);
xnor U14466 (N_14466,N_5049,N_6622);
xor U14467 (N_14467,N_8607,N_9025);
xnor U14468 (N_14468,N_7971,N_8922);
nand U14469 (N_14469,N_5898,N_9695);
or U14470 (N_14470,N_6882,N_5936);
or U14471 (N_14471,N_5906,N_9918);
and U14472 (N_14472,N_8524,N_6546);
or U14473 (N_14473,N_5945,N_7833);
or U14474 (N_14474,N_8811,N_6003);
nor U14475 (N_14475,N_5883,N_7106);
xnor U14476 (N_14476,N_7578,N_8647);
nor U14477 (N_14477,N_8323,N_7848);
and U14478 (N_14478,N_7168,N_6723);
nand U14479 (N_14479,N_7809,N_9418);
nand U14480 (N_14480,N_9978,N_7010);
nand U14481 (N_14481,N_7234,N_8434);
or U14482 (N_14482,N_6168,N_6962);
nor U14483 (N_14483,N_9168,N_7233);
and U14484 (N_14484,N_7231,N_9426);
nand U14485 (N_14485,N_9519,N_8947);
nor U14486 (N_14486,N_6132,N_9625);
or U14487 (N_14487,N_8628,N_5051);
xor U14488 (N_14488,N_6011,N_6604);
xnor U14489 (N_14489,N_6601,N_6957);
nand U14490 (N_14490,N_6776,N_7091);
nor U14491 (N_14491,N_7735,N_6109);
xor U14492 (N_14492,N_6018,N_8245);
xor U14493 (N_14493,N_9307,N_5963);
nor U14494 (N_14494,N_8661,N_8858);
xor U14495 (N_14495,N_9417,N_9233);
nand U14496 (N_14496,N_7152,N_8067);
nand U14497 (N_14497,N_9018,N_8493);
xor U14498 (N_14498,N_5645,N_8277);
xnor U14499 (N_14499,N_9366,N_9938);
and U14500 (N_14500,N_5967,N_5908);
nor U14501 (N_14501,N_8786,N_5386);
nand U14502 (N_14502,N_6209,N_6130);
or U14503 (N_14503,N_9512,N_9069);
xor U14504 (N_14504,N_7721,N_6362);
nor U14505 (N_14505,N_7325,N_5940);
nand U14506 (N_14506,N_6678,N_6237);
and U14507 (N_14507,N_7397,N_6051);
and U14508 (N_14508,N_8076,N_5001);
or U14509 (N_14509,N_5843,N_9172);
nor U14510 (N_14510,N_8879,N_7627);
nand U14511 (N_14511,N_7866,N_8583);
nand U14512 (N_14512,N_6918,N_6462);
nand U14513 (N_14513,N_9459,N_7753);
or U14514 (N_14514,N_6767,N_9368);
nor U14515 (N_14515,N_8735,N_9524);
xnor U14516 (N_14516,N_5973,N_7451);
nand U14517 (N_14517,N_5619,N_9637);
nor U14518 (N_14518,N_7653,N_8581);
or U14519 (N_14519,N_6522,N_7649);
and U14520 (N_14520,N_8340,N_5157);
nand U14521 (N_14521,N_9509,N_6631);
or U14522 (N_14522,N_8232,N_8707);
or U14523 (N_14523,N_8903,N_9334);
or U14524 (N_14524,N_9375,N_9275);
nor U14525 (N_14525,N_7277,N_7950);
or U14526 (N_14526,N_5028,N_6427);
nor U14527 (N_14527,N_5780,N_5503);
and U14528 (N_14528,N_8580,N_6993);
nand U14529 (N_14529,N_5256,N_6947);
and U14530 (N_14530,N_6579,N_6138);
and U14531 (N_14531,N_7288,N_9342);
and U14532 (N_14532,N_6547,N_8772);
or U14533 (N_14533,N_9189,N_9517);
nand U14534 (N_14534,N_6926,N_5051);
xnor U14535 (N_14535,N_6059,N_9992);
nand U14536 (N_14536,N_8794,N_9137);
or U14537 (N_14537,N_5296,N_6192);
and U14538 (N_14538,N_6870,N_5316);
or U14539 (N_14539,N_8227,N_6402);
and U14540 (N_14540,N_9171,N_8903);
or U14541 (N_14541,N_5167,N_9360);
nand U14542 (N_14542,N_6661,N_9171);
or U14543 (N_14543,N_6476,N_9800);
and U14544 (N_14544,N_9552,N_5176);
xnor U14545 (N_14545,N_7139,N_6095);
nand U14546 (N_14546,N_9978,N_6524);
nor U14547 (N_14547,N_6289,N_8875);
xor U14548 (N_14548,N_8674,N_6191);
or U14549 (N_14549,N_9829,N_9899);
nand U14550 (N_14550,N_8217,N_6455);
xor U14551 (N_14551,N_7215,N_5171);
or U14552 (N_14552,N_9689,N_5398);
xor U14553 (N_14553,N_7847,N_9793);
or U14554 (N_14554,N_7488,N_9123);
and U14555 (N_14555,N_5737,N_5982);
and U14556 (N_14556,N_7119,N_5873);
xor U14557 (N_14557,N_6230,N_9340);
and U14558 (N_14558,N_5034,N_8928);
and U14559 (N_14559,N_5206,N_5052);
nand U14560 (N_14560,N_5382,N_7451);
xnor U14561 (N_14561,N_8259,N_5068);
and U14562 (N_14562,N_8123,N_7834);
nand U14563 (N_14563,N_8375,N_9648);
or U14564 (N_14564,N_5431,N_7679);
nand U14565 (N_14565,N_6981,N_6643);
and U14566 (N_14566,N_7728,N_5944);
and U14567 (N_14567,N_8903,N_9469);
nor U14568 (N_14568,N_5229,N_9672);
or U14569 (N_14569,N_6407,N_7196);
xor U14570 (N_14570,N_6071,N_5094);
nor U14571 (N_14571,N_5773,N_9616);
nor U14572 (N_14572,N_7357,N_6991);
xor U14573 (N_14573,N_7146,N_5648);
nor U14574 (N_14574,N_6868,N_6026);
nand U14575 (N_14575,N_7025,N_8436);
or U14576 (N_14576,N_9531,N_6028);
nand U14577 (N_14577,N_8217,N_7003);
xor U14578 (N_14578,N_6941,N_8700);
nand U14579 (N_14579,N_8218,N_7937);
xor U14580 (N_14580,N_5845,N_5079);
xor U14581 (N_14581,N_9551,N_5732);
xnor U14582 (N_14582,N_9558,N_5300);
or U14583 (N_14583,N_7565,N_6328);
nand U14584 (N_14584,N_9864,N_9239);
xnor U14585 (N_14585,N_8572,N_5130);
and U14586 (N_14586,N_7293,N_8785);
xor U14587 (N_14587,N_7125,N_5253);
nor U14588 (N_14588,N_5403,N_5068);
nand U14589 (N_14589,N_5647,N_6039);
nor U14590 (N_14590,N_6374,N_5084);
nand U14591 (N_14591,N_8612,N_9131);
xnor U14592 (N_14592,N_9274,N_5885);
or U14593 (N_14593,N_8554,N_6494);
xor U14594 (N_14594,N_9085,N_6678);
or U14595 (N_14595,N_6359,N_7175);
or U14596 (N_14596,N_9369,N_9164);
nor U14597 (N_14597,N_9334,N_6792);
nor U14598 (N_14598,N_6253,N_9765);
nor U14599 (N_14599,N_9031,N_7101);
nand U14600 (N_14600,N_6883,N_7368);
or U14601 (N_14601,N_6955,N_5967);
and U14602 (N_14602,N_8540,N_7302);
nand U14603 (N_14603,N_6470,N_9356);
xor U14604 (N_14604,N_5308,N_8213);
nor U14605 (N_14605,N_8944,N_6456);
nor U14606 (N_14606,N_6613,N_6847);
nand U14607 (N_14607,N_8261,N_8849);
xor U14608 (N_14608,N_5597,N_6211);
nand U14609 (N_14609,N_8325,N_7357);
nand U14610 (N_14610,N_8959,N_6777);
xor U14611 (N_14611,N_5273,N_8312);
xor U14612 (N_14612,N_9776,N_9428);
xor U14613 (N_14613,N_7324,N_9604);
xor U14614 (N_14614,N_7557,N_9890);
and U14615 (N_14615,N_7720,N_7018);
nand U14616 (N_14616,N_7951,N_8286);
and U14617 (N_14617,N_5714,N_5887);
nor U14618 (N_14618,N_6496,N_8818);
and U14619 (N_14619,N_6300,N_6614);
nand U14620 (N_14620,N_9372,N_9333);
xor U14621 (N_14621,N_6819,N_7132);
or U14622 (N_14622,N_8341,N_6084);
nand U14623 (N_14623,N_5902,N_6440);
nor U14624 (N_14624,N_5196,N_6022);
xor U14625 (N_14625,N_5264,N_9481);
nor U14626 (N_14626,N_5374,N_6163);
or U14627 (N_14627,N_9678,N_8949);
nor U14628 (N_14628,N_7590,N_9978);
or U14629 (N_14629,N_9103,N_7741);
or U14630 (N_14630,N_8623,N_8762);
or U14631 (N_14631,N_8031,N_7505);
nor U14632 (N_14632,N_8222,N_5035);
nand U14633 (N_14633,N_9642,N_7915);
xor U14634 (N_14634,N_8865,N_7549);
or U14635 (N_14635,N_5982,N_6249);
and U14636 (N_14636,N_6569,N_6632);
xor U14637 (N_14637,N_9739,N_6570);
nor U14638 (N_14638,N_9163,N_5062);
and U14639 (N_14639,N_9712,N_6757);
nand U14640 (N_14640,N_7866,N_7701);
xnor U14641 (N_14641,N_9699,N_9674);
and U14642 (N_14642,N_9865,N_5637);
and U14643 (N_14643,N_8710,N_8755);
or U14644 (N_14644,N_8973,N_5431);
xor U14645 (N_14645,N_5696,N_7697);
xnor U14646 (N_14646,N_9671,N_5394);
and U14647 (N_14647,N_6672,N_7891);
or U14648 (N_14648,N_8674,N_9233);
nand U14649 (N_14649,N_5958,N_5991);
and U14650 (N_14650,N_5181,N_7795);
xor U14651 (N_14651,N_8654,N_9969);
nand U14652 (N_14652,N_6124,N_9983);
nor U14653 (N_14653,N_8593,N_5587);
nor U14654 (N_14654,N_5933,N_6475);
nand U14655 (N_14655,N_5123,N_9959);
nand U14656 (N_14656,N_7603,N_7101);
nor U14657 (N_14657,N_5170,N_5619);
nor U14658 (N_14658,N_5375,N_8030);
nor U14659 (N_14659,N_5304,N_5150);
xnor U14660 (N_14660,N_7532,N_5474);
nand U14661 (N_14661,N_5169,N_5911);
nor U14662 (N_14662,N_5783,N_7656);
and U14663 (N_14663,N_9894,N_5011);
and U14664 (N_14664,N_9048,N_6196);
nor U14665 (N_14665,N_9672,N_8103);
nand U14666 (N_14666,N_5756,N_6363);
xor U14667 (N_14667,N_5000,N_7781);
nand U14668 (N_14668,N_8650,N_5965);
nand U14669 (N_14669,N_6800,N_6340);
or U14670 (N_14670,N_5499,N_8543);
xor U14671 (N_14671,N_8001,N_5532);
nand U14672 (N_14672,N_7638,N_6196);
and U14673 (N_14673,N_9553,N_6375);
or U14674 (N_14674,N_6780,N_6948);
nor U14675 (N_14675,N_6858,N_8553);
and U14676 (N_14676,N_5028,N_8653);
and U14677 (N_14677,N_6086,N_7837);
nor U14678 (N_14678,N_7276,N_6565);
xnor U14679 (N_14679,N_5410,N_8196);
nor U14680 (N_14680,N_7026,N_6046);
or U14681 (N_14681,N_8006,N_8046);
xnor U14682 (N_14682,N_5043,N_7594);
nand U14683 (N_14683,N_7553,N_9953);
nor U14684 (N_14684,N_5215,N_8639);
nor U14685 (N_14685,N_8092,N_5060);
nand U14686 (N_14686,N_5661,N_9955);
or U14687 (N_14687,N_5135,N_5420);
nand U14688 (N_14688,N_5706,N_5851);
nor U14689 (N_14689,N_6686,N_6102);
and U14690 (N_14690,N_9510,N_7240);
nand U14691 (N_14691,N_8978,N_5131);
nor U14692 (N_14692,N_8181,N_9400);
nand U14693 (N_14693,N_7101,N_9500);
nand U14694 (N_14694,N_5358,N_8577);
and U14695 (N_14695,N_5983,N_9058);
nor U14696 (N_14696,N_6012,N_8712);
or U14697 (N_14697,N_8665,N_5088);
or U14698 (N_14698,N_9046,N_6652);
nand U14699 (N_14699,N_5032,N_5766);
and U14700 (N_14700,N_5491,N_6978);
or U14701 (N_14701,N_5076,N_8421);
and U14702 (N_14702,N_7890,N_9637);
or U14703 (N_14703,N_9100,N_8901);
or U14704 (N_14704,N_9375,N_8591);
nand U14705 (N_14705,N_8511,N_7177);
xnor U14706 (N_14706,N_7629,N_6813);
xor U14707 (N_14707,N_5924,N_7764);
nand U14708 (N_14708,N_8408,N_6337);
nand U14709 (N_14709,N_9129,N_5966);
or U14710 (N_14710,N_6491,N_8154);
xnor U14711 (N_14711,N_8963,N_6913);
nand U14712 (N_14712,N_5919,N_5358);
nor U14713 (N_14713,N_5055,N_6943);
xor U14714 (N_14714,N_7199,N_6896);
or U14715 (N_14715,N_7051,N_6656);
and U14716 (N_14716,N_5044,N_8265);
and U14717 (N_14717,N_9716,N_7007);
nand U14718 (N_14718,N_7681,N_7271);
or U14719 (N_14719,N_8639,N_8180);
and U14720 (N_14720,N_8250,N_9661);
xor U14721 (N_14721,N_8126,N_5033);
or U14722 (N_14722,N_5248,N_7467);
or U14723 (N_14723,N_7314,N_7260);
nand U14724 (N_14724,N_8278,N_9469);
nor U14725 (N_14725,N_8055,N_5643);
or U14726 (N_14726,N_7420,N_5640);
and U14727 (N_14727,N_8382,N_6098);
nand U14728 (N_14728,N_9767,N_5650);
xnor U14729 (N_14729,N_5615,N_8482);
xor U14730 (N_14730,N_8958,N_5601);
nand U14731 (N_14731,N_9356,N_6997);
xor U14732 (N_14732,N_6401,N_6852);
nor U14733 (N_14733,N_5796,N_6411);
nor U14734 (N_14734,N_7376,N_9029);
xor U14735 (N_14735,N_7981,N_9573);
and U14736 (N_14736,N_9987,N_9607);
nand U14737 (N_14737,N_7454,N_7546);
nor U14738 (N_14738,N_9577,N_7793);
nand U14739 (N_14739,N_9778,N_9410);
xnor U14740 (N_14740,N_5854,N_7368);
nor U14741 (N_14741,N_6814,N_9407);
nand U14742 (N_14742,N_9915,N_9919);
or U14743 (N_14743,N_5512,N_8261);
and U14744 (N_14744,N_9106,N_7860);
or U14745 (N_14745,N_7193,N_8879);
xnor U14746 (N_14746,N_7300,N_7970);
nand U14747 (N_14747,N_8392,N_7319);
or U14748 (N_14748,N_5405,N_7769);
and U14749 (N_14749,N_9171,N_5338);
and U14750 (N_14750,N_9467,N_7385);
or U14751 (N_14751,N_7618,N_7325);
nand U14752 (N_14752,N_7741,N_8880);
nor U14753 (N_14753,N_6971,N_5069);
and U14754 (N_14754,N_8505,N_9705);
xor U14755 (N_14755,N_5508,N_9387);
and U14756 (N_14756,N_5510,N_9233);
nand U14757 (N_14757,N_6654,N_5434);
and U14758 (N_14758,N_6435,N_7370);
and U14759 (N_14759,N_5208,N_9759);
xnor U14760 (N_14760,N_6348,N_9327);
and U14761 (N_14761,N_8911,N_8763);
and U14762 (N_14762,N_9016,N_6570);
or U14763 (N_14763,N_7099,N_5061);
and U14764 (N_14764,N_5631,N_7356);
xnor U14765 (N_14765,N_6644,N_9417);
nor U14766 (N_14766,N_8314,N_8341);
or U14767 (N_14767,N_7614,N_8447);
xnor U14768 (N_14768,N_6806,N_9489);
and U14769 (N_14769,N_5853,N_5892);
nor U14770 (N_14770,N_9245,N_9296);
nand U14771 (N_14771,N_8317,N_5188);
or U14772 (N_14772,N_5657,N_6068);
nand U14773 (N_14773,N_9137,N_7877);
and U14774 (N_14774,N_6956,N_5111);
xor U14775 (N_14775,N_9971,N_8335);
and U14776 (N_14776,N_7947,N_8553);
xor U14777 (N_14777,N_6223,N_6848);
and U14778 (N_14778,N_6861,N_7430);
nor U14779 (N_14779,N_6303,N_6007);
nand U14780 (N_14780,N_7920,N_7791);
xor U14781 (N_14781,N_8133,N_5979);
nand U14782 (N_14782,N_8599,N_9761);
and U14783 (N_14783,N_8286,N_9084);
nand U14784 (N_14784,N_6871,N_6175);
and U14785 (N_14785,N_8158,N_5627);
nor U14786 (N_14786,N_7285,N_9204);
and U14787 (N_14787,N_5186,N_9806);
and U14788 (N_14788,N_8726,N_6331);
and U14789 (N_14789,N_5322,N_5202);
or U14790 (N_14790,N_9104,N_7733);
nor U14791 (N_14791,N_8573,N_5736);
and U14792 (N_14792,N_8151,N_7710);
or U14793 (N_14793,N_6336,N_9425);
nor U14794 (N_14794,N_5107,N_6303);
nor U14795 (N_14795,N_8754,N_5441);
nor U14796 (N_14796,N_8839,N_6747);
xnor U14797 (N_14797,N_6691,N_5241);
and U14798 (N_14798,N_9229,N_6152);
and U14799 (N_14799,N_5395,N_9075);
and U14800 (N_14800,N_5154,N_8065);
and U14801 (N_14801,N_5324,N_5504);
nand U14802 (N_14802,N_9127,N_7255);
nand U14803 (N_14803,N_9226,N_8497);
nand U14804 (N_14804,N_6818,N_9364);
or U14805 (N_14805,N_7527,N_8466);
and U14806 (N_14806,N_8591,N_5293);
or U14807 (N_14807,N_5735,N_9183);
nor U14808 (N_14808,N_5682,N_5568);
nor U14809 (N_14809,N_5461,N_9489);
nor U14810 (N_14810,N_7962,N_8647);
nor U14811 (N_14811,N_5891,N_6866);
xor U14812 (N_14812,N_7558,N_8850);
xor U14813 (N_14813,N_5659,N_8430);
xnor U14814 (N_14814,N_7048,N_7894);
and U14815 (N_14815,N_7989,N_6495);
nand U14816 (N_14816,N_5915,N_6575);
xor U14817 (N_14817,N_5549,N_7809);
nand U14818 (N_14818,N_9691,N_8401);
nand U14819 (N_14819,N_7739,N_5202);
nand U14820 (N_14820,N_7339,N_6502);
or U14821 (N_14821,N_8229,N_5683);
or U14822 (N_14822,N_7877,N_5364);
xnor U14823 (N_14823,N_8097,N_8941);
nand U14824 (N_14824,N_6290,N_6913);
or U14825 (N_14825,N_6106,N_5262);
or U14826 (N_14826,N_5227,N_6522);
nor U14827 (N_14827,N_6699,N_7476);
or U14828 (N_14828,N_8636,N_5695);
and U14829 (N_14829,N_8158,N_6360);
nand U14830 (N_14830,N_9072,N_5707);
or U14831 (N_14831,N_5997,N_9938);
xnor U14832 (N_14832,N_8168,N_5473);
and U14833 (N_14833,N_9350,N_7740);
and U14834 (N_14834,N_7352,N_5225);
nor U14835 (N_14835,N_6998,N_6533);
nor U14836 (N_14836,N_5313,N_5948);
or U14837 (N_14837,N_6753,N_7764);
or U14838 (N_14838,N_6106,N_9740);
nand U14839 (N_14839,N_9176,N_9875);
nand U14840 (N_14840,N_7338,N_7494);
xnor U14841 (N_14841,N_8715,N_7431);
nand U14842 (N_14842,N_8824,N_6045);
or U14843 (N_14843,N_9059,N_5550);
and U14844 (N_14844,N_7417,N_9541);
xnor U14845 (N_14845,N_9038,N_5576);
nand U14846 (N_14846,N_8654,N_8760);
xnor U14847 (N_14847,N_8119,N_8765);
xnor U14848 (N_14848,N_6157,N_8236);
nand U14849 (N_14849,N_8150,N_5130);
nand U14850 (N_14850,N_7286,N_8654);
nor U14851 (N_14851,N_8875,N_9122);
nor U14852 (N_14852,N_7560,N_6026);
nor U14853 (N_14853,N_6535,N_5823);
and U14854 (N_14854,N_5987,N_8120);
and U14855 (N_14855,N_6184,N_9286);
and U14856 (N_14856,N_8374,N_5821);
nand U14857 (N_14857,N_8387,N_9494);
or U14858 (N_14858,N_8027,N_7895);
nand U14859 (N_14859,N_5144,N_7083);
or U14860 (N_14860,N_5244,N_7692);
or U14861 (N_14861,N_5241,N_9633);
nor U14862 (N_14862,N_6676,N_8988);
nor U14863 (N_14863,N_9191,N_9969);
or U14864 (N_14864,N_5239,N_6701);
or U14865 (N_14865,N_9809,N_7758);
or U14866 (N_14866,N_7748,N_7992);
nor U14867 (N_14867,N_6616,N_6970);
and U14868 (N_14868,N_6776,N_6585);
nand U14869 (N_14869,N_9404,N_7262);
or U14870 (N_14870,N_5908,N_6315);
or U14871 (N_14871,N_9738,N_6665);
and U14872 (N_14872,N_5717,N_9072);
nand U14873 (N_14873,N_7605,N_9345);
xor U14874 (N_14874,N_6571,N_9854);
and U14875 (N_14875,N_9246,N_6049);
nor U14876 (N_14876,N_6572,N_5570);
xor U14877 (N_14877,N_6294,N_7809);
or U14878 (N_14878,N_5822,N_6554);
nand U14879 (N_14879,N_8787,N_6449);
xnor U14880 (N_14880,N_6836,N_9242);
xnor U14881 (N_14881,N_8136,N_9518);
or U14882 (N_14882,N_6806,N_8336);
nor U14883 (N_14883,N_8731,N_6079);
nor U14884 (N_14884,N_5508,N_5718);
and U14885 (N_14885,N_8196,N_9394);
and U14886 (N_14886,N_7372,N_9611);
and U14887 (N_14887,N_6977,N_7415);
and U14888 (N_14888,N_8629,N_9743);
xor U14889 (N_14889,N_5836,N_7840);
and U14890 (N_14890,N_6899,N_6014);
xor U14891 (N_14891,N_7724,N_7991);
or U14892 (N_14892,N_9942,N_7973);
and U14893 (N_14893,N_9136,N_5451);
nand U14894 (N_14894,N_8725,N_5955);
nor U14895 (N_14895,N_9206,N_9665);
nand U14896 (N_14896,N_8995,N_5475);
xor U14897 (N_14897,N_9420,N_7988);
nand U14898 (N_14898,N_5367,N_5802);
xnor U14899 (N_14899,N_8830,N_8712);
or U14900 (N_14900,N_9912,N_6919);
nor U14901 (N_14901,N_6909,N_9334);
nor U14902 (N_14902,N_6513,N_7555);
nor U14903 (N_14903,N_9480,N_8481);
xor U14904 (N_14904,N_5055,N_7002);
and U14905 (N_14905,N_7349,N_8565);
nor U14906 (N_14906,N_8278,N_7589);
nor U14907 (N_14907,N_6743,N_6297);
and U14908 (N_14908,N_7486,N_7306);
xor U14909 (N_14909,N_7929,N_8087);
nor U14910 (N_14910,N_5773,N_5440);
nor U14911 (N_14911,N_5822,N_9630);
xnor U14912 (N_14912,N_5020,N_5686);
nor U14913 (N_14913,N_8018,N_5951);
xnor U14914 (N_14914,N_8389,N_5068);
or U14915 (N_14915,N_9387,N_7061);
xor U14916 (N_14916,N_9749,N_6094);
and U14917 (N_14917,N_9034,N_7777);
nor U14918 (N_14918,N_9072,N_9129);
or U14919 (N_14919,N_7249,N_6859);
xor U14920 (N_14920,N_7946,N_8916);
xor U14921 (N_14921,N_6833,N_7928);
nand U14922 (N_14922,N_9576,N_5357);
xnor U14923 (N_14923,N_9341,N_7249);
xnor U14924 (N_14924,N_9677,N_7645);
or U14925 (N_14925,N_6344,N_8194);
nor U14926 (N_14926,N_9764,N_7167);
nand U14927 (N_14927,N_5391,N_5011);
and U14928 (N_14928,N_6604,N_6701);
nand U14929 (N_14929,N_7698,N_5451);
and U14930 (N_14930,N_8508,N_6794);
xor U14931 (N_14931,N_9050,N_6844);
nand U14932 (N_14932,N_6061,N_5178);
and U14933 (N_14933,N_5357,N_7950);
and U14934 (N_14934,N_9596,N_6033);
xnor U14935 (N_14935,N_8616,N_9132);
xor U14936 (N_14936,N_9227,N_5051);
or U14937 (N_14937,N_9805,N_6521);
or U14938 (N_14938,N_7171,N_5411);
nor U14939 (N_14939,N_6037,N_9696);
xnor U14940 (N_14940,N_9007,N_6973);
or U14941 (N_14941,N_9312,N_7427);
and U14942 (N_14942,N_7850,N_6357);
nand U14943 (N_14943,N_9306,N_8672);
or U14944 (N_14944,N_5911,N_5141);
and U14945 (N_14945,N_8244,N_9394);
or U14946 (N_14946,N_6589,N_6609);
xor U14947 (N_14947,N_6840,N_8368);
xnor U14948 (N_14948,N_8101,N_7027);
and U14949 (N_14949,N_8723,N_7118);
or U14950 (N_14950,N_8257,N_8787);
or U14951 (N_14951,N_7756,N_9627);
or U14952 (N_14952,N_5724,N_7728);
nand U14953 (N_14953,N_8285,N_9110);
and U14954 (N_14954,N_7222,N_9718);
nand U14955 (N_14955,N_8362,N_6233);
and U14956 (N_14956,N_9920,N_6490);
and U14957 (N_14957,N_7073,N_8717);
nand U14958 (N_14958,N_8849,N_9110);
and U14959 (N_14959,N_7991,N_7562);
nand U14960 (N_14960,N_5524,N_5111);
and U14961 (N_14961,N_6418,N_6967);
nand U14962 (N_14962,N_8219,N_5153);
xor U14963 (N_14963,N_8089,N_6575);
nand U14964 (N_14964,N_8171,N_9868);
or U14965 (N_14965,N_6814,N_8518);
nand U14966 (N_14966,N_7247,N_6246);
and U14967 (N_14967,N_9817,N_9632);
nor U14968 (N_14968,N_9502,N_6521);
or U14969 (N_14969,N_6023,N_9198);
nand U14970 (N_14970,N_6660,N_5015);
nor U14971 (N_14971,N_5845,N_7676);
or U14972 (N_14972,N_7677,N_9399);
xor U14973 (N_14973,N_7217,N_8840);
and U14974 (N_14974,N_9906,N_6945);
and U14975 (N_14975,N_6130,N_8394);
and U14976 (N_14976,N_7405,N_6237);
nand U14977 (N_14977,N_5401,N_6783);
nor U14978 (N_14978,N_8504,N_5835);
xnor U14979 (N_14979,N_8598,N_6589);
nand U14980 (N_14980,N_8694,N_9719);
and U14981 (N_14981,N_5376,N_8449);
or U14982 (N_14982,N_5569,N_6461);
and U14983 (N_14983,N_8667,N_6504);
and U14984 (N_14984,N_7281,N_9232);
and U14985 (N_14985,N_5526,N_7702);
or U14986 (N_14986,N_8296,N_8159);
nor U14987 (N_14987,N_9762,N_6202);
and U14988 (N_14988,N_7354,N_9100);
or U14989 (N_14989,N_8601,N_5460);
or U14990 (N_14990,N_6820,N_9746);
xor U14991 (N_14991,N_7137,N_7568);
nand U14992 (N_14992,N_7816,N_9136);
or U14993 (N_14993,N_9736,N_6903);
xor U14994 (N_14994,N_6912,N_7523);
nand U14995 (N_14995,N_9283,N_5224);
nand U14996 (N_14996,N_9354,N_9880);
or U14997 (N_14997,N_6220,N_9272);
and U14998 (N_14998,N_5062,N_8159);
xor U14999 (N_14999,N_6311,N_7488);
nor U15000 (N_15000,N_14760,N_13365);
nand U15001 (N_15001,N_10417,N_13347);
nand U15002 (N_15002,N_10313,N_11144);
and U15003 (N_15003,N_13684,N_12348);
nor U15004 (N_15004,N_13657,N_14818);
or U15005 (N_15005,N_10769,N_12825);
nand U15006 (N_15006,N_14362,N_10082);
nor U15007 (N_15007,N_13976,N_10038);
nor U15008 (N_15008,N_14605,N_11868);
nand U15009 (N_15009,N_14799,N_14715);
and U15010 (N_15010,N_12788,N_14003);
xnor U15011 (N_15011,N_12777,N_14025);
nor U15012 (N_15012,N_12417,N_14625);
nand U15013 (N_15013,N_10708,N_10399);
or U15014 (N_15014,N_14459,N_12643);
nand U15015 (N_15015,N_12418,N_10718);
or U15016 (N_15016,N_13852,N_12450);
and U15017 (N_15017,N_12970,N_11403);
xor U15018 (N_15018,N_12554,N_14915);
or U15019 (N_15019,N_13156,N_14132);
or U15020 (N_15020,N_12130,N_12475);
xnor U15021 (N_15021,N_12884,N_11156);
and U15022 (N_15022,N_14038,N_13120);
nand U15023 (N_15023,N_12594,N_12822);
nand U15024 (N_15024,N_13421,N_11973);
nand U15025 (N_15025,N_14214,N_12419);
and U15026 (N_15026,N_14897,N_10505);
and U15027 (N_15027,N_11240,N_14379);
nand U15028 (N_15028,N_13488,N_14883);
nor U15029 (N_15029,N_14954,N_12717);
nand U15030 (N_15030,N_12133,N_12156);
xnor U15031 (N_15031,N_12444,N_14851);
xnor U15032 (N_15032,N_11546,N_10960);
xor U15033 (N_15033,N_10688,N_13535);
nor U15034 (N_15034,N_12420,N_14040);
and U15035 (N_15035,N_13945,N_12945);
nor U15036 (N_15036,N_14706,N_14553);
nor U15037 (N_15037,N_11782,N_11257);
or U15038 (N_15038,N_13280,N_11463);
nor U15039 (N_15039,N_13300,N_14381);
nor U15040 (N_15040,N_10492,N_12654);
nor U15041 (N_15041,N_10012,N_13273);
and U15042 (N_15042,N_12863,N_10063);
nand U15043 (N_15043,N_12678,N_12966);
or U15044 (N_15044,N_11325,N_14039);
and U15045 (N_15045,N_13730,N_12843);
nand U15046 (N_15046,N_10620,N_11140);
nor U15047 (N_15047,N_12645,N_11623);
nor U15048 (N_15048,N_12281,N_12566);
xor U15049 (N_15049,N_14812,N_11956);
nand U15050 (N_15050,N_12710,N_14322);
or U15051 (N_15051,N_11547,N_11972);
nor U15052 (N_15052,N_10702,N_12109);
nand U15053 (N_15053,N_13638,N_10150);
or U15054 (N_15054,N_10430,N_13065);
nand U15055 (N_15055,N_11051,N_10065);
or U15056 (N_15056,N_13266,N_14659);
nor U15057 (N_15057,N_11747,N_12771);
nor U15058 (N_15058,N_14341,N_10717);
nand U15059 (N_15059,N_11872,N_10163);
xnor U15060 (N_15060,N_13599,N_10114);
and U15061 (N_15061,N_14218,N_12561);
xnor U15062 (N_15062,N_11723,N_13370);
nand U15063 (N_15063,N_11505,N_14245);
nand U15064 (N_15064,N_14704,N_13737);
nand U15065 (N_15065,N_11160,N_11298);
nand U15066 (N_15066,N_12347,N_10509);
or U15067 (N_15067,N_12448,N_12326);
nand U15068 (N_15068,N_10432,N_11545);
nor U15069 (N_15069,N_13743,N_14923);
and U15070 (N_15070,N_12657,N_13747);
or U15071 (N_15071,N_11145,N_13158);
or U15072 (N_15072,N_13765,N_10543);
nor U15073 (N_15073,N_13040,N_12699);
nor U15074 (N_15074,N_11243,N_12177);
nor U15075 (N_15075,N_14757,N_12545);
xnor U15076 (N_15076,N_12578,N_12687);
and U15077 (N_15077,N_13756,N_14085);
or U15078 (N_15078,N_10537,N_11447);
xnor U15079 (N_15079,N_14495,N_13694);
or U15080 (N_15080,N_10506,N_10843);
nand U15081 (N_15081,N_14853,N_10014);
and U15082 (N_15082,N_10085,N_11624);
nand U15083 (N_15083,N_13030,N_11724);
nand U15084 (N_15084,N_12662,N_10281);
nand U15085 (N_15085,N_14138,N_11955);
and U15086 (N_15086,N_12181,N_14167);
nor U15087 (N_15087,N_14781,N_12824);
and U15088 (N_15088,N_13003,N_10555);
xor U15089 (N_15089,N_10893,N_11016);
and U15090 (N_15090,N_13930,N_12129);
nand U15091 (N_15091,N_12095,N_13226);
and U15092 (N_15092,N_14217,N_10919);
and U15093 (N_15093,N_11562,N_14251);
and U15094 (N_15094,N_12559,N_13016);
nand U15095 (N_15095,N_12575,N_12622);
nor U15096 (N_15096,N_14616,N_14430);
xor U15097 (N_15097,N_11139,N_13782);
nor U15098 (N_15098,N_14096,N_11296);
xnor U15099 (N_15099,N_13736,N_13998);
or U15100 (N_15100,N_12006,N_14718);
xor U15101 (N_15101,N_10148,N_13850);
nor U15102 (N_15102,N_14857,N_11914);
xnor U15103 (N_15103,N_10673,N_10405);
nor U15104 (N_15104,N_12893,N_10308);
xnor U15105 (N_15105,N_13268,N_14325);
and U15106 (N_15106,N_13640,N_12873);
xnor U15107 (N_15107,N_12366,N_12954);
and U15108 (N_15108,N_14825,N_14403);
xnor U15109 (N_15109,N_14801,N_12530);
nor U15110 (N_15110,N_11580,N_14030);
and U15111 (N_15111,N_10050,N_13048);
nor U15112 (N_15112,N_13680,N_13794);
xor U15113 (N_15113,N_13742,N_10459);
nor U15114 (N_15114,N_11647,N_12330);
or U15115 (N_15115,N_13260,N_12915);
nor U15116 (N_15116,N_11945,N_10247);
nand U15117 (N_15117,N_12567,N_12431);
xnor U15118 (N_15118,N_13452,N_12106);
or U15119 (N_15119,N_14656,N_14670);
and U15120 (N_15120,N_12779,N_10475);
or U15121 (N_15121,N_14174,N_13231);
or U15122 (N_15122,N_13574,N_12042);
or U15123 (N_15123,N_13610,N_13228);
or U15124 (N_15124,N_13067,N_11382);
and U15125 (N_15125,N_11800,N_14017);
or U15126 (N_15126,N_11259,N_10263);
or U15127 (N_15127,N_11472,N_13405);
xor U15128 (N_15128,N_13677,N_10729);
or U15129 (N_15129,N_14224,N_14640);
and U15130 (N_15130,N_13066,N_11048);
nor U15131 (N_15131,N_13202,N_12105);
and U15132 (N_15132,N_13176,N_10116);
nor U15133 (N_15133,N_13670,N_14509);
nor U15134 (N_15134,N_12520,N_11757);
nand U15135 (N_15135,N_12034,N_10796);
and U15136 (N_15136,N_10149,N_14513);
xor U15137 (N_15137,N_12199,N_12671);
nand U15138 (N_15138,N_11763,N_10317);
nor U15139 (N_15139,N_10494,N_13554);
nand U15140 (N_15140,N_11556,N_11917);
nand U15141 (N_15141,N_11488,N_12638);
xor U15142 (N_15142,N_10978,N_13648);
nand U15143 (N_15143,N_13407,N_11925);
xor U15144 (N_15144,N_10278,N_12150);
xnor U15145 (N_15145,N_13965,N_13943);
nand U15146 (N_15146,N_11024,N_10618);
and U15147 (N_15147,N_11253,N_11086);
nand U15148 (N_15148,N_13198,N_12839);
xor U15149 (N_15149,N_11060,N_11558);
nand U15150 (N_15150,N_11702,N_11727);
or U15151 (N_15151,N_10300,N_11131);
nor U15152 (N_15152,N_14391,N_11158);
and U15153 (N_15153,N_12857,N_11531);
nand U15154 (N_15154,N_11828,N_11761);
xnor U15155 (N_15155,N_14772,N_11661);
nand U15156 (N_15156,N_11197,N_13536);
xnor U15157 (N_15157,N_10540,N_11813);
and U15158 (N_15158,N_13305,N_13614);
nor U15159 (N_15159,N_11745,N_12144);
xnor U15160 (N_15160,N_13064,N_11913);
and U15161 (N_15161,N_13315,N_10955);
and U15162 (N_15162,N_14621,N_13732);
and U15163 (N_15163,N_14433,N_10541);
xnor U15164 (N_15164,N_11184,N_10794);
nor U15165 (N_15165,N_11008,N_10023);
xor U15166 (N_15166,N_14061,N_13979);
nand U15167 (N_15167,N_14265,N_12886);
nor U15168 (N_15168,N_13051,N_12665);
and U15169 (N_15169,N_10306,N_12068);
or U15170 (N_15170,N_10360,N_14094);
xnor U15171 (N_15171,N_10061,N_10269);
nand U15172 (N_15172,N_11471,N_14454);
xnor U15173 (N_15173,N_10238,N_14767);
xor U15174 (N_15174,N_14962,N_10950);
nor U15175 (N_15175,N_13603,N_13106);
and U15176 (N_15176,N_14068,N_14112);
and U15177 (N_15177,N_10407,N_14216);
nand U15178 (N_15178,N_14371,N_13829);
nand U15179 (N_15179,N_12328,N_13672);
and U15180 (N_15180,N_14572,N_11818);
xnor U15181 (N_15181,N_12012,N_13279);
nor U15182 (N_15182,N_12772,N_14558);
nand U15183 (N_15183,N_12350,N_13096);
and U15184 (N_15184,N_11934,N_12850);
and U15185 (N_15185,N_14891,N_13556);
or U15186 (N_15186,N_14047,N_11045);
nor U15187 (N_15187,N_10707,N_10005);
xor U15188 (N_15188,N_10120,N_12607);
xor U15189 (N_15189,N_14782,N_12730);
or U15190 (N_15190,N_14761,N_10699);
xor U15191 (N_15191,N_10368,N_10725);
or U15192 (N_15192,N_13731,N_14678);
nor U15193 (N_15193,N_14508,N_13272);
xnor U15194 (N_15194,N_10513,N_14215);
or U15195 (N_15195,N_13702,N_14449);
xnor U15196 (N_15196,N_12615,N_13224);
nor U15197 (N_15197,N_14770,N_13163);
xnor U15198 (N_15198,N_13642,N_13100);
xor U15199 (N_15199,N_10554,N_14305);
xor U15200 (N_15200,N_14404,N_14351);
nor U15201 (N_15201,N_11438,N_11576);
and U15202 (N_15202,N_10333,N_11117);
nor U15203 (N_15203,N_14993,N_12739);
nand U15204 (N_15204,N_11735,N_12132);
or U15205 (N_15205,N_14398,N_10384);
and U15206 (N_15206,N_14827,N_14065);
nand U15207 (N_15207,N_10041,N_11338);
and U15208 (N_15208,N_12553,N_11864);
or U15209 (N_15209,N_11857,N_13439);
nand U15210 (N_15210,N_12927,N_13544);
nor U15211 (N_15211,N_12878,N_11808);
or U15212 (N_15212,N_13038,N_13446);
and U15213 (N_15213,N_12452,N_12291);
and U15214 (N_15214,N_14150,N_11555);
xnor U15215 (N_15215,N_11109,N_13581);
nand U15216 (N_15216,N_12190,N_10639);
or U15217 (N_15217,N_13502,N_10053);
nor U15218 (N_15218,N_10265,N_10452);
or U15219 (N_15219,N_12337,N_14453);
or U15220 (N_15220,N_10827,N_14570);
xor U15221 (N_15221,N_10434,N_12735);
nor U15222 (N_15222,N_12176,N_13873);
xor U15223 (N_15223,N_11173,N_14298);
nand U15224 (N_15224,N_11612,N_10856);
xnor U15225 (N_15225,N_14646,N_13057);
xnor U15226 (N_15226,N_12690,N_11900);
and U15227 (N_15227,N_14575,N_12149);
xnor U15228 (N_15228,N_10244,N_14498);
nor U15229 (N_15229,N_12406,N_10233);
xor U15230 (N_15230,N_12482,N_12941);
xnor U15231 (N_15231,N_14890,N_14144);
or U15232 (N_15232,N_12152,N_12365);
or U15233 (N_15233,N_14585,N_11931);
and U15234 (N_15234,N_12810,N_14483);
nor U15235 (N_15235,N_13652,N_11871);
or U15236 (N_15236,N_13424,N_11074);
and U15237 (N_15237,N_14233,N_10840);
nor U15238 (N_15238,N_13802,N_12702);
xor U15239 (N_15239,N_13585,N_14566);
and U15240 (N_15240,N_11742,N_12938);
or U15241 (N_15241,N_10568,N_13422);
xnor U15242 (N_15242,N_11346,N_12339);
or U15243 (N_15243,N_12200,N_10465);
and U15244 (N_15244,N_10448,N_10880);
nand U15245 (N_15245,N_13751,N_11066);
nor U15246 (N_15246,N_11908,N_13338);
nor U15247 (N_15247,N_14713,N_14653);
nor U15248 (N_15248,N_14166,N_14295);
xor U15249 (N_15249,N_10389,N_10208);
or U15250 (N_15250,N_13840,N_13104);
xnor U15251 (N_15251,N_13074,N_12496);
nor U15252 (N_15252,N_13810,N_11494);
nor U15253 (N_15253,N_11422,N_14568);
nor U15254 (N_15254,N_12243,N_10987);
xor U15255 (N_15255,N_12731,N_11714);
xnor U15256 (N_15256,N_10176,N_10654);
nor U15257 (N_15257,N_10370,N_10064);
or U15258 (N_15258,N_10635,N_10656);
and U15259 (N_15259,N_10387,N_11377);
and U15260 (N_15260,N_14945,N_10890);
or U15261 (N_15261,N_10571,N_12639);
or U15262 (N_15262,N_13068,N_12600);
or U15263 (N_15263,N_13575,N_11744);
and U15264 (N_15264,N_13649,N_10552);
nor U15265 (N_15265,N_13078,N_12841);
nor U15266 (N_15266,N_13658,N_12518);
nand U15267 (N_15267,N_12957,N_10188);
nor U15268 (N_15268,N_11272,N_11464);
or U15269 (N_15269,N_12844,N_14866);
xnor U15270 (N_15270,N_14474,N_13616);
nor U15271 (N_15271,N_12249,N_10312);
and U15272 (N_15272,N_11314,N_12959);
and U15273 (N_15273,N_14059,N_10478);
and U15274 (N_15274,N_11357,N_13253);
xnor U15275 (N_15275,N_12466,N_14643);
nand U15276 (N_15276,N_14358,N_12631);
nand U15277 (N_15277,N_10361,N_13663);
and U15278 (N_15278,N_10922,N_12276);
and U15279 (N_15279,N_12598,N_10304);
or U15280 (N_15280,N_10001,N_12103);
or U15281 (N_15281,N_10777,N_14856);
or U15282 (N_15282,N_13821,N_14824);
or U15283 (N_15283,N_14199,N_12216);
nor U15284 (N_15284,N_14735,N_11476);
xnor U15285 (N_15285,N_10069,N_13703);
xor U15286 (N_15286,N_14252,N_11376);
nor U15287 (N_15287,N_11087,N_11099);
and U15288 (N_15288,N_13590,N_12629);
xor U15289 (N_15289,N_14971,N_14301);
nand U15290 (N_15290,N_13270,N_11027);
xor U15291 (N_15291,N_12907,N_10415);
nand U15292 (N_15292,N_13897,N_11170);
nand U15293 (N_15293,N_11187,N_10756);
nor U15294 (N_15294,N_11866,N_13083);
nand U15295 (N_15295,N_12897,N_10489);
xnor U15296 (N_15296,N_12302,N_10825);
and U15297 (N_15297,N_13991,N_12627);
nor U15298 (N_15298,N_11462,N_10604);
and U15299 (N_15299,N_11411,N_11044);
nor U15300 (N_15300,N_13384,N_12499);
nor U15301 (N_15301,N_12207,N_14155);
nand U15302 (N_15302,N_13056,N_14516);
or U15303 (N_15303,N_11206,N_13942);
and U15304 (N_15304,N_10395,N_13167);
or U15305 (N_15305,N_12940,N_13902);
xor U15306 (N_15306,N_10047,N_12193);
and U15307 (N_15307,N_14342,N_11174);
nand U15308 (N_15308,N_12613,N_13341);
nor U15309 (N_15309,N_12107,N_13872);
nor U15310 (N_15310,N_14792,N_12061);
nand U15311 (N_15311,N_11572,N_14244);
and U15312 (N_15312,N_14839,N_12385);
and U15313 (N_15313,N_11273,N_10549);
xnor U15314 (N_15314,N_14023,N_14893);
and U15315 (N_15315,N_11846,N_14826);
nor U15316 (N_15316,N_10603,N_12037);
nand U15317 (N_15317,N_13608,N_11652);
and U15318 (N_15318,N_11706,N_13157);
nor U15319 (N_15319,N_11939,N_11870);
xnor U15320 (N_15320,N_11121,N_14170);
nand U15321 (N_15321,N_12165,N_11754);
or U15322 (N_15322,N_12770,N_14121);
xor U15323 (N_15323,N_14161,N_11736);
or U15324 (N_15324,N_14090,N_11903);
and U15325 (N_15325,N_11823,N_11313);
nor U15326 (N_15326,N_12025,N_11617);
xnor U15327 (N_15327,N_11785,N_11811);
nand U15328 (N_15328,N_13572,N_12506);
xnor U15329 (N_15329,N_13368,N_14935);
or U15330 (N_15330,N_10750,N_12972);
nor U15331 (N_15331,N_13843,N_10535);
and U15332 (N_15332,N_12397,N_11485);
nor U15333 (N_15333,N_12602,N_12202);
nand U15334 (N_15334,N_10301,N_10516);
xnor U15335 (N_15335,N_12542,N_13512);
or U15336 (N_15336,N_13801,N_10010);
nor U15337 (N_15337,N_13546,N_14504);
and U15338 (N_15338,N_10181,N_10159);
and U15339 (N_15339,N_14577,N_11593);
or U15340 (N_15340,N_14791,N_11538);
nor U15341 (N_15341,N_10598,N_14308);
xor U15342 (N_15342,N_12624,N_12231);
or U15343 (N_15343,N_12395,N_13822);
xnor U15344 (N_15344,N_14898,N_11839);
nand U15345 (N_15345,N_11461,N_10558);
nand U15346 (N_15346,N_10470,N_13006);
nand U15347 (N_15347,N_11695,N_11953);
nand U15348 (N_15348,N_14268,N_12059);
and U15349 (N_15349,N_11344,N_10206);
xnor U15350 (N_15350,N_13237,N_11862);
nor U15351 (N_15351,N_12313,N_12709);
or U15352 (N_15352,N_12087,N_11549);
xnor U15353 (N_15353,N_14376,N_10689);
or U15354 (N_15354,N_14887,N_14154);
nor U15355 (N_15355,N_13707,N_12977);
or U15356 (N_15356,N_11317,N_11178);
nand U15357 (N_15357,N_10590,N_14111);
nand U15358 (N_15358,N_12352,N_13673);
xnor U15359 (N_15359,N_13085,N_11067);
nor U15360 (N_15360,N_10884,N_12626);
nor U15361 (N_15361,N_10239,N_13857);
nor U15362 (N_15362,N_10381,N_14961);
nor U15363 (N_15363,N_14324,N_11428);
nand U15364 (N_15364,N_10497,N_10225);
xnor U15365 (N_15365,N_11798,N_14936);
and U15366 (N_15366,N_10040,N_11890);
and U15367 (N_15367,N_13238,N_11384);
xor U15368 (N_15368,N_14194,N_11295);
nand U15369 (N_15369,N_12075,N_14164);
nor U15370 (N_15370,N_12257,N_11380);
nand U15371 (N_15371,N_14406,N_14906);
nand U15372 (N_15372,N_11247,N_12445);
nor U15373 (N_15373,N_14554,N_10421);
xnor U15374 (N_15374,N_11921,N_10153);
or U15375 (N_15375,N_14844,N_14388);
nor U15376 (N_15376,N_13285,N_11473);
xnor U15377 (N_15377,N_12260,N_13613);
and U15378 (N_15378,N_11102,N_14714);
nor U15379 (N_15379,N_10406,N_13717);
and U15380 (N_15380,N_13968,N_13073);
nand U15381 (N_15381,N_13451,N_12074);
nor U15382 (N_15382,N_11017,N_14537);
and U15383 (N_15383,N_14581,N_10488);
nand U15384 (N_15384,N_14707,N_12015);
nor U15385 (N_15385,N_11129,N_13740);
xnor U15386 (N_15386,N_14445,N_10573);
and U15387 (N_15387,N_11692,N_11982);
nand U15388 (N_15388,N_10690,N_14650);
and U15389 (N_15389,N_12247,N_14796);
or U15390 (N_15390,N_13706,N_12002);
xor U15391 (N_15391,N_12171,N_14636);
xnor U15392 (N_15392,N_13570,N_11250);
nor U15393 (N_15393,N_12756,N_11269);
or U15394 (N_15394,N_13212,N_12534);
nand U15395 (N_15395,N_13054,N_14808);
xor U15396 (N_15396,N_12169,N_14266);
nor U15397 (N_15397,N_10696,N_12135);
nand U15398 (N_15398,N_12218,N_13661);
nand U15399 (N_15399,N_13007,N_10990);
nor U15400 (N_15400,N_10075,N_12659);
xnor U15401 (N_15401,N_14255,N_12924);
and U15402 (N_15402,N_10863,N_11437);
xnor U15403 (N_15403,N_14262,N_13859);
xor U15404 (N_15404,N_12707,N_11963);
xnor U15405 (N_15405,N_11025,N_13580);
nor U15406 (N_15406,N_13682,N_10439);
and U15407 (N_15407,N_14469,N_12222);
nand U15408 (N_15408,N_12642,N_14436);
xnor U15409 (N_15409,N_13256,N_13997);
xnor U15410 (N_15410,N_10902,N_13115);
nor U15411 (N_15411,N_12459,N_12405);
and U15412 (N_15412,N_11201,N_13427);
or U15413 (N_15413,N_10924,N_10227);
and U15414 (N_15414,N_12052,N_11423);
nor U15415 (N_15415,N_13077,N_10155);
nand U15416 (N_15416,N_14596,N_13209);
nand U15417 (N_15417,N_14004,N_10976);
nor U15418 (N_15418,N_13199,N_12043);
nor U15419 (N_15419,N_12791,N_13653);
xor U15420 (N_15420,N_14423,N_11780);
and U15421 (N_15421,N_14119,N_12947);
xnor U15422 (N_15422,N_14567,N_11588);
nor U15423 (N_15423,N_12693,N_13970);
or U15424 (N_15424,N_10039,N_10973);
xor U15425 (N_15425,N_12111,N_13362);
nor U15426 (N_15426,N_14285,N_11478);
nand U15427 (N_15427,N_14304,N_13444);
nand U15428 (N_15428,N_14086,N_14479);
nor U15429 (N_15429,N_13475,N_14192);
and U15430 (N_15430,N_10821,N_12262);
and U15431 (N_15431,N_10134,N_12384);
nor U15432 (N_15432,N_13388,N_11323);
and U15433 (N_15433,N_10511,N_13501);
nor U15434 (N_15434,N_14667,N_13147);
and U15435 (N_15435,N_14927,N_14947);
and U15436 (N_15436,N_13321,N_11978);
nand U15437 (N_15437,N_11354,N_12118);
or U15438 (N_15438,N_13931,N_13705);
xor U15439 (N_15439,N_12086,N_10298);
xor U15440 (N_15440,N_10129,N_14242);
nor U15441 (N_15441,N_11185,N_10780);
nand U15442 (N_15442,N_11957,N_11608);
nand U15443 (N_15443,N_13458,N_10425);
nand U15444 (N_15444,N_13937,N_12354);
nand U15445 (N_15445,N_12618,N_11777);
and U15446 (N_15446,N_13161,N_13477);
xor U15447 (N_15447,N_10316,N_10775);
and U15448 (N_15448,N_11372,N_11516);
or U15449 (N_15449,N_12592,N_12535);
xnor U15450 (N_15450,N_12625,N_14178);
and U15451 (N_15451,N_12568,N_12433);
nor U15452 (N_15452,N_12314,N_12827);
and U15453 (N_15453,N_12953,N_11451);
nor U15454 (N_15454,N_13103,N_14429);
or U15455 (N_15455,N_10779,N_14139);
xnor U15456 (N_15456,N_11509,N_11611);
xor U15457 (N_15457,N_11984,N_12484);
or U15458 (N_15458,N_13357,N_14908);
nor U15459 (N_15459,N_10904,N_11468);
nand U15460 (N_15460,N_14130,N_14066);
xnor U15461 (N_15461,N_14984,N_12532);
nor U15462 (N_15462,N_12019,N_11748);
nand U15463 (N_15463,N_12404,N_10123);
and U15464 (N_15464,N_13335,N_13623);
xor U15465 (N_15465,N_10240,N_13303);
and U15466 (N_15466,N_11071,N_10414);
or U15467 (N_15467,N_14559,N_10232);
nand U15468 (N_15468,N_10350,N_13646);
nand U15469 (N_15469,N_14968,N_12093);
and U15470 (N_15470,N_13042,N_14514);
xor U15471 (N_15471,N_10701,N_11856);
or U15472 (N_15472,N_11030,N_10192);
nor U15473 (N_15473,N_11579,N_13947);
or U15474 (N_15474,N_10789,N_11132);
xor U15475 (N_15475,N_13524,N_14867);
nand U15476 (N_15476,N_12266,N_11776);
xnor U15477 (N_15477,N_10803,N_11297);
xnor U15478 (N_15478,N_14146,N_11548);
and U15479 (N_15479,N_13060,N_10137);
nand U15480 (N_15480,N_11552,N_12370);
and U15481 (N_15481,N_14953,N_13785);
xnor U15482 (N_15482,N_13111,N_10234);
nor U15483 (N_15483,N_11924,N_13485);
nand U15484 (N_15484,N_13686,N_12428);
and U15485 (N_15485,N_13059,N_10520);
nor U15486 (N_15486,N_10800,N_14415);
nand U15487 (N_15487,N_10502,N_10963);
or U15488 (N_15488,N_14288,N_10022);
or U15489 (N_15489,N_12442,N_13645);
xnor U15490 (N_15490,N_10647,N_12585);
and U15491 (N_15491,N_13387,N_13254);
or U15492 (N_15492,N_14289,N_14614);
xnor U15493 (N_15493,N_14922,N_13641);
nand U15494 (N_15494,N_11733,N_11151);
or U15495 (N_15495,N_10091,N_11435);
and U15496 (N_15496,N_11838,N_12910);
nor U15497 (N_15497,N_14858,N_10746);
and U15498 (N_15498,N_13777,N_13814);
xor U15499 (N_15499,N_14565,N_14521);
and U15500 (N_15500,N_10899,N_11791);
nand U15501 (N_15501,N_12577,N_13329);
nand U15502 (N_15502,N_10180,N_14695);
nand U15503 (N_15503,N_11676,N_11070);
or U15504 (N_15504,N_12454,N_10382);
or U15505 (N_15505,N_10228,N_10168);
nor U15506 (N_15506,N_12390,N_14082);
nand U15507 (N_15507,N_14582,N_11557);
and U15508 (N_15508,N_14374,N_13183);
and U15509 (N_15509,N_11664,N_11679);
and U15510 (N_15510,N_14687,N_10527);
nor U15511 (N_15511,N_14197,N_11609);
nor U15512 (N_15512,N_10171,N_14569);
xor U15513 (N_15513,N_13708,N_12936);
nor U15514 (N_15514,N_14044,N_14422);
nand U15515 (N_15515,N_10575,N_12014);
xor U15516 (N_15516,N_11339,N_10663);
and U15517 (N_15517,N_10755,N_12005);
nand U15518 (N_15518,N_12774,N_14260);
or U15519 (N_15519,N_11162,N_10697);
and U15520 (N_15520,N_13709,N_10989);
and U15521 (N_15521,N_13214,N_10512);
nor U15522 (N_15522,N_12091,N_10706);
and U15523 (N_15523,N_14490,N_13200);
xor U15524 (N_15524,N_13724,N_14762);
xor U15525 (N_15525,N_11211,N_14529);
nand U15526 (N_15526,N_11453,N_10215);
xnor U15527 (N_15527,N_13168,N_13624);
and U15528 (N_15528,N_11831,N_12652);
nor U15529 (N_15529,N_13403,N_12661);
nor U15530 (N_15530,N_12733,N_10811);
nand U15531 (N_15531,N_11614,N_13276);
and U15532 (N_15532,N_10289,N_12300);
xnor U15533 (N_15533,N_13679,N_10337);
or U15534 (N_15534,N_11658,N_12937);
or U15535 (N_15535,N_13215,N_13851);
and U15536 (N_15536,N_11636,N_11210);
and U15537 (N_15537,N_11920,N_14123);
and U15538 (N_15538,N_10563,N_14624);
xor U15539 (N_15539,N_11672,N_11032);
nor U15540 (N_15540,N_14950,N_14136);
xnor U15541 (N_15541,N_14795,N_11493);
or U15542 (N_15542,N_12815,N_12838);
and U15543 (N_15543,N_13013,N_14912);
and U15544 (N_15544,N_13769,N_13109);
or U15545 (N_15545,N_11902,N_10714);
nor U15546 (N_15546,N_13671,N_11414);
xnor U15547 (N_15547,N_14287,N_14043);
nand U15548 (N_15548,N_12802,N_10641);
and U15549 (N_15549,N_14396,N_10562);
or U15550 (N_15550,N_10732,N_12254);
xor U15551 (N_15551,N_11628,N_13734);
xor U15552 (N_15552,N_12686,N_14250);
nand U15553 (N_15553,N_12425,N_10931);
or U15554 (N_15554,N_11741,N_14815);
or U15555 (N_15555,N_14871,N_11565);
or U15556 (N_15556,N_10889,N_13963);
nand U15557 (N_15557,N_12173,N_12446);
xnor U15558 (N_15558,N_13600,N_11039);
and U15559 (N_15559,N_12139,N_12901);
or U15560 (N_15560,N_12324,N_14160);
and U15561 (N_15561,N_12780,N_14691);
and U15562 (N_15562,N_14032,N_14332);
and U15563 (N_15563,N_12944,N_10837);
or U15564 (N_15564,N_13015,N_11564);
or U15565 (N_15565,N_13172,N_10348);
nand U15566 (N_15566,N_14008,N_10449);
nand U15567 (N_15567,N_11009,N_14081);
or U15568 (N_15568,N_12599,N_13337);
and U15569 (N_15569,N_14363,N_11918);
nor U15570 (N_15570,N_12641,N_12570);
nand U15571 (N_15571,N_12789,N_14705);
and U15572 (N_15572,N_10966,N_12698);
nand U15573 (N_15573,N_13223,N_14273);
nor U15574 (N_15574,N_14805,N_10757);
nor U15575 (N_15575,N_11993,N_10771);
and U15576 (N_15576,N_14875,N_14424);
and U15577 (N_15577,N_13956,N_10920);
nor U15578 (N_15578,N_12505,N_12519);
and U15579 (N_15579,N_10339,N_14368);
and U15580 (N_15580,N_12285,N_14574);
nor U15581 (N_15581,N_10930,N_11540);
xor U15582 (N_15582,N_12875,N_11753);
nand U15583 (N_15583,N_10318,N_13519);
nand U15584 (N_15584,N_12877,N_14727);
and U15585 (N_15585,N_10859,N_10321);
nand U15586 (N_15586,N_13194,N_12517);
nor U15587 (N_15587,N_13352,N_13123);
or U15588 (N_15588,N_13350,N_14069);
and U15589 (N_15589,N_13795,N_12749);
xor U15590 (N_15590,N_14800,N_12264);
nand U15591 (N_15591,N_14205,N_12113);
or U15592 (N_15592,N_11283,N_14779);
nor U15593 (N_15593,N_11175,N_10730);
and U15594 (N_15594,N_10323,N_14517);
nor U15595 (N_15595,N_11511,N_14060);
and U15596 (N_15596,N_13097,N_12539);
nor U15597 (N_15597,N_13289,N_14673);
xor U15598 (N_15598,N_13024,N_10531);
and U15599 (N_15599,N_11059,N_13332);
nor U15600 (N_15600,N_10523,N_14942);
nor U15601 (N_15601,N_12497,N_14272);
and U15602 (N_15602,N_11849,N_12073);
nor U15603 (N_15603,N_12472,N_12491);
nor U15604 (N_15604,N_14712,N_12102);
nor U15605 (N_15605,N_12734,N_13411);
and U15606 (N_15606,N_13313,N_10043);
or U15607 (N_15607,N_13985,N_13651);
nor U15608 (N_15608,N_10253,N_13525);
xor U15609 (N_15609,N_13558,N_12729);
nor U15610 (N_15610,N_10364,N_13726);
and U15611 (N_15611,N_11123,N_12195);
nand U15612 (N_15612,N_13053,N_14397);
and U15613 (N_15613,N_12895,N_10831);
and U15614 (N_15614,N_14222,N_12685);
nand U15615 (N_15615,N_14716,N_11362);
xnor U15616 (N_15616,N_10807,N_11486);
nand U15617 (N_15617,N_14631,N_10751);
nand U15618 (N_15618,N_14390,N_11134);
and U15619 (N_15619,N_12233,N_12606);
and U15620 (N_15620,N_13139,N_10444);
nand U15621 (N_15621,N_13331,N_14743);
nand U15622 (N_15622,N_12796,N_14648);
nor U15623 (N_15623,N_14444,N_11686);
nor U15624 (N_15624,N_10934,N_13689);
nand U15625 (N_15625,N_10282,N_10616);
xnor U15626 (N_15626,N_13380,N_11704);
and U15627 (N_15627,N_11223,N_10290);
and U15628 (N_15628,N_10349,N_13560);
or U15629 (N_15629,N_10170,N_14458);
nand U15630 (N_15630,N_14769,N_13205);
or U15631 (N_15631,N_14290,N_10853);
xnor U15632 (N_15632,N_12713,N_14816);
xor U15633 (N_15633,N_13000,N_10107);
nor U15634 (N_15634,N_14103,N_13701);
and U15635 (N_15635,N_12148,N_14588);
xor U15636 (N_15636,N_11584,N_14978);
and U15637 (N_15637,N_14924,N_11869);
xnor U15638 (N_15638,N_13218,N_10921);
xnor U15639 (N_15639,N_10498,N_12237);
nand U15640 (N_15640,N_13492,N_11630);
and U15641 (N_15641,N_11220,N_12461);
nor U15642 (N_15642,N_10271,N_13208);
xor U15643 (N_15643,N_11288,N_14405);
xor U15644 (N_15644,N_11319,N_13033);
xnor U15645 (N_15645,N_11209,N_10024);
xor U15646 (N_15646,N_13294,N_10634);
or U15647 (N_15647,N_12563,N_14360);
or U15648 (N_15648,N_14759,N_11927);
nand U15649 (N_15649,N_12027,N_14277);
and U15650 (N_15650,N_14776,N_10813);
nor U15651 (N_15651,N_13008,N_14315);
nor U15652 (N_15652,N_14100,N_11154);
nand U15653 (N_15653,N_14960,N_13140);
nand U15654 (N_15654,N_10347,N_14402);
nor U15655 (N_15655,N_11378,N_12882);
or U15656 (N_15656,N_11198,N_12725);
nor U15657 (N_15657,N_14426,N_14134);
xnor U15658 (N_15658,N_14987,N_11353);
xor U15659 (N_15659,N_10354,N_14620);
or U15660 (N_15660,N_14435,N_12088);
xor U15661 (N_15661,N_10557,N_10357);
nor U15662 (N_15662,N_13292,N_10480);
or U15663 (N_15663,N_10586,N_13173);
xnor U15664 (N_15664,N_13343,N_10599);
or U15665 (N_15665,N_12187,N_13043);
nand U15666 (N_15666,N_11497,N_12569);
nand U15667 (N_15667,N_14914,N_12985);
or U15668 (N_15668,N_11050,N_11640);
nor U15669 (N_15669,N_13354,N_13853);
or U15670 (N_15670,N_12391,N_12571);
or U15671 (N_15671,N_10875,N_13849);
and U15672 (N_15672,N_10100,N_10447);
xor U15673 (N_15673,N_14203,N_13233);
xnor U15674 (N_15674,N_14798,N_11720);
or U15675 (N_15675,N_13170,N_11255);
xor U15676 (N_15676,N_12383,N_13093);
nor U15677 (N_15677,N_10583,N_10267);
xnor U15678 (N_15678,N_12175,N_12762);
or U15679 (N_15679,N_11853,N_11816);
and U15680 (N_15680,N_11649,N_13296);
or U15681 (N_15681,N_11759,N_11594);
nand U15682 (N_15682,N_11328,N_10709);
or U15683 (N_15683,N_11280,N_14227);
or U15684 (N_15684,N_11164,N_12394);
nor U15685 (N_15685,N_11500,N_14586);
or U15686 (N_15686,N_12763,N_13537);
nor U15687 (N_15687,N_14029,N_13904);
xor U15688 (N_15688,N_13994,N_10704);
and U15689 (N_15689,N_11408,N_10098);
or U15690 (N_15690,N_13878,N_10182);
or U15691 (N_15691,N_10778,N_10733);
nor U15692 (N_15692,N_10915,N_13277);
nor U15693 (N_15693,N_12587,N_13201);
xor U15694 (N_15694,N_10195,N_10473);
xnor U15695 (N_15695,N_14316,N_14934);
or U15696 (N_15696,N_10052,N_10614);
xor U15697 (N_15697,N_13195,N_10548);
nand U15698 (N_15698,N_11258,N_14171);
nand U15699 (N_15699,N_11106,N_10332);
nand U15700 (N_15700,N_13457,N_13455);
and U15701 (N_15701,N_13861,N_13807);
xor U15702 (N_15702,N_10818,N_14076);
nor U15703 (N_15703,N_13465,N_11525);
xnor U15704 (N_15704,N_14651,N_11781);
or U15705 (N_15705,N_13974,N_14958);
nand U15706 (N_15706,N_10140,N_14369);
nand U15707 (N_15707,N_14156,N_12704);
and U15708 (N_15708,N_12364,N_13118);
and U15709 (N_15709,N_13912,N_13181);
nor U15710 (N_15710,N_12079,N_14578);
xnor U15711 (N_15711,N_11845,N_11833);
xnor U15712 (N_15712,N_14084,N_10275);
nor U15713 (N_15713,N_14869,N_11770);
or U15714 (N_15714,N_12646,N_10454);
xor U15715 (N_15715,N_10307,N_13102);
nand U15716 (N_15716,N_11375,N_14067);
or U15717 (N_15717,N_10682,N_13448);
nand U15718 (N_15718,N_13164,N_14662);
or U15719 (N_15719,N_13160,N_13211);
nor U15720 (N_15720,N_13739,N_10319);
nor U15721 (N_15721,N_13800,N_14729);
xnor U15722 (N_15722,N_13324,N_11263);
or U15723 (N_15723,N_12413,N_10784);
or U15724 (N_15724,N_14464,N_13874);
xor U15725 (N_15725,N_13022,N_11007);
nor U15726 (N_15726,N_11103,N_13433);
xor U15727 (N_15727,N_11327,N_10309);
xnor U15728 (N_15728,N_12898,N_10534);
nor U15729 (N_15729,N_12449,N_12523);
nand U15730 (N_15730,N_11291,N_10802);
and U15731 (N_15731,N_13004,N_11430);
or U15732 (N_15732,N_10826,N_13622);
and U15733 (N_15733,N_11181,N_14663);
and U15734 (N_15734,N_14158,N_11267);
nand U15735 (N_15735,N_13619,N_10499);
nand U15736 (N_15736,N_13526,N_13491);
nand U15737 (N_15737,N_11575,N_14117);
or U15738 (N_15738,N_14632,N_10379);
nand U15739 (N_15739,N_14020,N_10754);
nor U15740 (N_15740,N_11475,N_12614);
nand U15741 (N_15741,N_10436,N_10607);
xor U15742 (N_15742,N_12525,N_13171);
nor U15743 (N_15743,N_13088,N_12465);
nor U15744 (N_15744,N_14747,N_14874);
nor U15745 (N_15745,N_14062,N_11938);
nor U15746 (N_15746,N_10245,N_10736);
nand U15747 (N_15747,N_13036,N_11578);
or U15748 (N_15748,N_14876,N_12206);
xnor U15749 (N_15749,N_11413,N_14208);
nor U15750 (N_15750,N_10135,N_12688);
and U15751 (N_15751,N_13453,N_10111);
or U15752 (N_15752,N_11607,N_14093);
and U15753 (N_15753,N_14573,N_10939);
or U15754 (N_15754,N_10526,N_10739);
nand U15755 (N_15755,N_12076,N_12215);
nor U15756 (N_15756,N_10676,N_10546);
or U15757 (N_15757,N_12213,N_12304);
nand U15758 (N_15758,N_10948,N_11961);
or U15759 (N_15759,N_11429,N_13304);
nor U15760 (N_15760,N_11758,N_14073);
nand U15761 (N_15761,N_10983,N_10814);
nor U15762 (N_15762,N_14309,N_11192);
nand U15763 (N_15763,N_13426,N_12261);
and U15764 (N_15764,N_14610,N_11666);
nand U15765 (N_15765,N_12053,N_10997);
and U15766 (N_15766,N_14828,N_13715);
and U15767 (N_15767,N_12753,N_13454);
nand U15768 (N_15768,N_10431,N_14319);
and U15769 (N_15769,N_12697,N_10287);
nor U15770 (N_15770,N_11148,N_10125);
and U15771 (N_15771,N_14339,N_12524);
xor U15772 (N_15772,N_11137,N_12477);
xnor U15773 (N_15773,N_10322,N_10566);
xnor U15774 (N_15774,N_12538,N_12676);
nand U15775 (N_15775,N_11208,N_10016);
xor U15776 (N_15776,N_13842,N_14455);
nand U15777 (N_15777,N_14849,N_14652);
xnor U15778 (N_15778,N_13203,N_13145);
nor U15779 (N_15779,N_11743,N_10982);
nand U15780 (N_15780,N_13908,N_14889);
or U15781 (N_15781,N_13655,N_14098);
nand U15782 (N_15782,N_10760,N_12127);
xor U15783 (N_15783,N_13230,N_12368);
or U15784 (N_15784,N_10099,N_13754);
nor U15785 (N_15785,N_12188,N_11270);
nor U15786 (N_15786,N_11142,N_14975);
nand U15787 (N_15787,N_13395,N_10268);
xor U15788 (N_15788,N_13483,N_13348);
nor U15789 (N_15789,N_14507,N_12584);
or U15790 (N_15790,N_12290,N_13847);
or U15791 (N_15791,N_14492,N_14847);
xnor U15792 (N_15792,N_11302,N_14261);
and U15793 (N_15793,N_11412,N_12515);
nand U15794 (N_15794,N_14054,N_14774);
nand U15795 (N_15795,N_14655,N_11091);
nor U15796 (N_15796,N_10836,N_14240);
and U15797 (N_15797,N_10467,N_11622);
nor U15798 (N_15798,N_11459,N_10295);
nand U15799 (N_15799,N_10500,N_12740);
and U15800 (N_15800,N_12860,N_10151);
or U15801 (N_15801,N_11010,N_12049);
or U15802 (N_15802,N_14037,N_10958);
xnor U15803 (N_15803,N_13523,N_11110);
nor U15804 (N_15804,N_14113,N_11581);
or U15805 (N_15805,N_12031,N_13369);
nor U15806 (N_15806,N_12229,N_13733);
xnor U15807 (N_15807,N_10691,N_13295);
nand U15808 (N_15808,N_11477,N_11432);
and U15809 (N_15809,N_13184,N_14526);
xnor U15810 (N_15810,N_11893,N_14933);
nor U15811 (N_15811,N_13602,N_11308);
nor U15812 (N_15812,N_13383,N_12001);
and U15813 (N_15813,N_10401,N_11470);
xnor U15814 (N_15814,N_13447,N_13924);
nand U15815 (N_15815,N_12634,N_11911);
nand U15816 (N_15816,N_10074,N_14778);
nor U15817 (N_15817,N_14494,N_12997);
or U15818 (N_15818,N_14609,N_12151);
or U15819 (N_15819,N_11002,N_14970);
and U15820 (N_15820,N_13515,N_11125);
nand U15821 (N_15821,N_12374,N_10578);
nand U15822 (N_15822,N_14384,N_14378);
or U15823 (N_15823,N_10589,N_14549);
xor U15824 (N_15824,N_13397,N_11986);
xnor U15825 (N_15825,N_14299,N_10184);
xnor U15826 (N_15826,N_10327,N_12411);
nor U15827 (N_15827,N_12245,N_14988);
and U15828 (N_15828,N_12804,N_12097);
nand U15829 (N_15829,N_11804,N_12334);
nor U15830 (N_15830,N_12217,N_10412);
nor U15831 (N_15831,N_10946,N_10968);
or U15832 (N_15832,N_13784,N_13586);
nand U15833 (N_15833,N_12790,N_10705);
and U15834 (N_15834,N_13011,N_13497);
and U15835 (N_15835,N_14972,N_10721);
or U15836 (N_15836,N_13826,N_14348);
or U15837 (N_15837,N_14904,N_11454);
nand U15838 (N_15838,N_10230,N_11300);
and U15839 (N_15839,N_14591,N_14728);
and U15840 (N_15840,N_13385,N_10830);
and U15841 (N_15841,N_10911,N_13445);
nand U15842 (N_15842,N_13190,N_13656);
nor U15843 (N_15843,N_11948,N_14202);
nand U15844 (N_15844,N_14125,N_12949);
nor U15845 (N_15845,N_14257,N_10315);
nand U15846 (N_15846,N_10373,N_10622);
nand U15847 (N_15847,N_12315,N_11177);
or U15848 (N_15848,N_14077,N_11842);
and U15849 (N_15849,N_14939,N_12930);
xor U15850 (N_15850,N_10567,N_10097);
nand U15851 (N_15851,N_13615,N_10869);
xor U15852 (N_15852,N_14698,N_14500);
nor U15853 (N_15853,N_10937,N_10273);
nand U15854 (N_15854,N_10895,N_10805);
and U15855 (N_15855,N_14903,N_11878);
nand U15856 (N_15856,N_10272,N_10576);
nand U15857 (N_15857,N_11503,N_11621);
nor U15858 (N_15858,N_14977,N_12692);
and U15859 (N_15859,N_13528,N_14394);
xnor U15860 (N_15860,N_13410,N_12289);
and U15861 (N_15861,N_11820,N_12375);
or U15862 (N_15862,N_13925,N_10493);
nor U15863 (N_15863,N_14148,N_12010);
xor U15864 (N_15864,N_13349,N_10518);
xor U15865 (N_15865,N_14142,N_11563);
or U15866 (N_15866,N_13262,N_13516);
xor U15867 (N_15867,N_12083,N_13499);
and U15868 (N_15868,N_11631,N_14354);
xnor U15869 (N_15869,N_10217,N_10687);
nor U15870 (N_15870,N_10303,N_14355);
nor U15871 (N_15871,N_10019,N_10711);
nand U15872 (N_15872,N_14048,N_10198);
xor U15873 (N_15873,N_12760,N_12456);
nand U15874 (N_15874,N_12121,N_11410);
and U15875 (N_15875,N_14669,N_10259);
xor U15876 (N_15876,N_12018,N_10749);
nand U15877 (N_15877,N_13197,N_11746);
nand U15878 (N_15878,N_14780,N_14775);
nor U15879 (N_15879,N_12981,N_14502);
nand U15880 (N_15880,N_12055,N_11985);
xor U15881 (N_15881,N_12712,N_11084);
nor U15882 (N_15882,N_11796,N_10910);
xor U15883 (N_15883,N_12464,N_12544);
or U15884 (N_15884,N_13984,N_10785);
or U15885 (N_15885,N_10358,N_11202);
and U15886 (N_15886,N_12610,N_12890);
and U15887 (N_15887,N_14916,N_12116);
or U15888 (N_15888,N_14515,N_11954);
and U15889 (N_15889,N_14437,N_13612);
nand U15890 (N_15890,N_12303,N_14708);
or U15891 (N_15891,N_11426,N_12341);
xor U15892 (N_15892,N_12301,N_13127);
or U15893 (N_15893,N_12586,N_13898);
or U15894 (N_15894,N_12312,N_13479);
xnor U15895 (N_15895,N_13975,N_12994);
xor U15896 (N_15896,N_13281,N_10409);
nand U15897 (N_15897,N_13265,N_14310);
and U15898 (N_15898,N_14613,N_14630);
and U15899 (N_15899,N_13901,N_13957);
nor U15900 (N_15900,N_13017,N_10855);
xor U15901 (N_15901,N_14477,N_13377);
nor U15902 (N_15902,N_11023,N_14579);
xnor U15903 (N_15903,N_14340,N_14921);
xor U15904 (N_15904,N_13258,N_12070);
or U15905 (N_15905,N_12675,N_11155);
and U15906 (N_15906,N_10248,N_14932);
nor U15907 (N_15907,N_12040,N_13375);
nor U15908 (N_15908,N_11064,N_11887);
nand U15909 (N_15909,N_11794,N_10894);
nand U15910 (N_15910,N_10223,N_10962);
nand U15911 (N_15911,N_14764,N_11827);
xor U15912 (N_15912,N_13496,N_13923);
nor U15913 (N_15913,N_10624,N_12916);
and U15914 (N_15914,N_11958,N_14058);
or U15915 (N_15915,N_11529,N_11322);
nand U15916 (N_15916,N_11182,N_13583);
or U15917 (N_15917,N_11452,N_10753);
and U15918 (N_15918,N_13964,N_13960);
nand U15919 (N_15919,N_14448,N_12439);
nor U15920 (N_15920,N_12434,N_14057);
nand U15921 (N_15921,N_13461,N_12424);
xor U15922 (N_15922,N_13949,N_14556);
xor U15923 (N_15923,N_11641,N_12414);
nor U15924 (N_15924,N_11237,N_12271);
or U15925 (N_15925,N_10212,N_12128);
and U15926 (N_15926,N_14722,N_10122);
xor U15927 (N_15927,N_11075,N_14522);
xor U15928 (N_15928,N_12443,N_13805);
nand U15929 (N_15929,N_14749,N_13044);
xor U15930 (N_15930,N_10854,N_11304);
nor U15931 (N_15931,N_14491,N_13725);
xor U15932 (N_15932,N_10487,N_13192);
nand U15933 (N_15933,N_14347,N_13050);
nor U15934 (N_15934,N_12274,N_10692);
xnor U15935 (N_15935,N_13432,N_14690);
and U15936 (N_15936,N_11127,N_10356);
or U15937 (N_15937,N_13470,N_13503);
nand U15938 (N_15938,N_10767,N_10255);
nor U15939 (N_15939,N_13728,N_10745);
nand U15940 (N_15940,N_11532,N_13710);
xnor U15941 (N_15941,N_13948,N_11169);
and U15942 (N_15942,N_11179,N_10296);
nor U15943 (N_15943,N_14638,N_13885);
xnor U15944 (N_15944,N_12668,N_10655);
and U15945 (N_15945,N_12633,N_13721);
nor U15946 (N_15946,N_13552,N_13105);
nor U15947 (N_15947,N_13408,N_13361);
nand U15948 (N_15948,N_13286,N_13500);
nand U15949 (N_15949,N_13450,N_12978);
nor U15950 (N_15950,N_13020,N_13128);
nand U15951 (N_15951,N_10865,N_12064);
or U15952 (N_15952,N_11673,N_14639);
or U15953 (N_15953,N_12363,N_14329);
or U15954 (N_15954,N_11425,N_10411);
or U15955 (N_15955,N_13366,N_12335);
or U15956 (N_15956,N_13472,N_14256);
xor U15957 (N_15957,N_11981,N_13971);
nor U15958 (N_15958,N_13667,N_11589);
nand U15959 (N_15959,N_10398,N_10460);
nand U15960 (N_15960,N_12017,N_12581);
nand U15961 (N_15961,N_14576,N_12948);
xnor U15962 (N_15962,N_11795,N_11783);
and U15963 (N_15963,N_13449,N_11395);
xnor U15964 (N_15964,N_11632,N_10565);
xor U15965 (N_15965,N_12230,N_10712);
nand U15966 (N_15966,N_14236,N_14019);
and U15967 (N_15967,N_14243,N_10627);
and U15968 (N_15968,N_14184,N_10173);
and U15969 (N_15969,N_10700,N_13776);
or U15970 (N_15970,N_10799,N_11514);
or U15971 (N_15971,N_10089,N_12056);
nand U15972 (N_15972,N_12054,N_11230);
nand U15973 (N_15973,N_10870,N_10076);
and U15974 (N_15974,N_11268,N_14021);
xnor U15975 (N_15975,N_12258,N_14294);
and U15976 (N_15976,N_10776,N_14909);
nor U15977 (N_15977,N_14733,N_13633);
xor U15978 (N_15978,N_14274,N_12795);
xnor U15979 (N_15979,N_11974,N_11596);
xnor U15980 (N_15980,N_12032,N_10876);
or U15981 (N_15981,N_13274,N_13604);
xnor U15982 (N_15982,N_12039,N_10261);
nand U15983 (N_15983,N_10994,N_13830);
and U15984 (N_15984,N_12695,N_11730);
nor U15985 (N_15985,N_13783,N_14863);
xor U15986 (N_15986,N_11521,N_13567);
xor U15987 (N_15987,N_12784,N_13213);
nor U15988 (N_15988,N_11036,N_12298);
nand U15989 (N_15989,N_12767,N_11186);
nor U15990 (N_15990,N_14074,N_12846);
and U15991 (N_15991,N_13117,N_13996);
nand U15992 (N_15992,N_11693,N_10279);
nand U15993 (N_15993,N_13832,N_11292);
nor U15994 (N_15994,N_14865,N_13660);
xor U15995 (N_15995,N_12436,N_12060);
nor U15996 (N_15996,N_11627,N_13766);
xnor U15997 (N_15997,N_11643,N_11888);
and U15998 (N_15998,N_12108,N_13986);
xor U15999 (N_15999,N_13404,N_14420);
nor U16000 (N_16000,N_14540,N_13116);
or U16001 (N_16001,N_11806,N_10162);
or U16002 (N_16002,N_10901,N_11610);
nand U16003 (N_16003,N_12382,N_13269);
nor U16004 (N_16004,N_10015,N_12814);
or U16005 (N_16005,N_11560,N_11019);
and U16006 (N_16006,N_13779,N_14133);
and U16007 (N_16007,N_12510,N_10857);
xor U16008 (N_16008,N_13086,N_14018);
or U16009 (N_16009,N_12991,N_14411);
xor U16010 (N_16010,N_10220,N_14929);
nand U16011 (N_16011,N_10550,N_10892);
xnor U16012 (N_16012,N_12590,N_12837);
and U16013 (N_16013,N_11684,N_11994);
nand U16014 (N_16014,N_12159,N_14005);
xnor U16015 (N_16015,N_10117,N_14913);
and U16016 (N_16016,N_14232,N_10839);
nor U16017 (N_16017,N_11052,N_14330);
nand U16018 (N_16018,N_11374,N_11303);
or U16019 (N_16019,N_13774,N_10477);
or U16020 (N_16020,N_12968,N_10204);
nand U16021 (N_16021,N_14523,N_11603);
nand U16022 (N_16022,N_12388,N_10203);
and U16023 (N_16023,N_11279,N_10057);
or U16024 (N_16024,N_14263,N_12672);
and U16025 (N_16025,N_12632,N_13029);
or U16026 (N_16026,N_10504,N_11683);
and U16027 (N_16027,N_14637,N_11038);
xor U16028 (N_16028,N_12500,N_13468);
nand U16029 (N_16029,N_12429,N_13881);
and U16030 (N_16030,N_13541,N_12794);
nand U16031 (N_16031,N_10592,N_12899);
and U16032 (N_16032,N_11349,N_13748);
nor U16033 (N_16033,N_11301,N_11923);
or U16034 (N_16034,N_13637,N_10581);
or U16035 (N_16035,N_12081,N_12033);
or U16036 (N_16036,N_11491,N_13435);
and U16037 (N_16037,N_12047,N_14593);
nor U16038 (N_16038,N_11359,N_10113);
nand U16039 (N_16039,N_14209,N_11122);
nand U16040 (N_16040,N_12597,N_13588);
nor U16041 (N_16041,N_12030,N_13031);
and U16042 (N_16042,N_13654,N_10060);
nor U16043 (N_16043,N_14548,N_13831);
and U16044 (N_16044,N_11388,N_12866);
xnor U16045 (N_16045,N_11625,N_10375);
xnor U16046 (N_16046,N_12310,N_12469);
and U16047 (N_16047,N_12359,N_12147);
nor U16048 (N_16048,N_13507,N_14201);
nand U16049 (N_16049,N_14872,N_12327);
nor U16050 (N_16050,N_13566,N_13063);
nand U16051 (N_16051,N_14370,N_13359);
xnor U16052 (N_16052,N_11420,N_12705);
or U16053 (N_16053,N_13259,N_13587);
nor U16054 (N_16054,N_10445,N_12536);
xor U16055 (N_16055,N_13221,N_14542);
nor U16056 (N_16056,N_11022,N_10838);
and U16057 (N_16057,N_12800,N_13420);
nor U16058 (N_16058,N_12864,N_14899);
and U16059 (N_16059,N_10292,N_14831);
xnor U16060 (N_16060,N_13406,N_11107);
nor U16061 (N_16061,N_13486,N_10190);
and U16062 (N_16062,N_12319,N_10536);
nor U16063 (N_16063,N_11830,N_12722);
nand U16064 (N_16064,N_12869,N_11340);
nand U16065 (N_16065,N_11153,N_13720);
nor U16066 (N_16066,N_11814,N_14389);
nand U16067 (N_16067,N_14618,N_10418);
nor U16068 (N_16068,N_10954,N_13398);
xor U16069 (N_16069,N_12809,N_12601);
nand U16070 (N_16070,N_12112,N_14270);
nor U16071 (N_16071,N_14180,N_10175);
or U16072 (N_16072,N_12398,N_10972);
and U16073 (N_16073,N_13768,N_14080);
nand U16074 (N_16074,N_12062,N_10094);
or U16075 (N_16075,N_11480,N_12400);
xnor U16076 (N_16076,N_14010,N_12275);
or U16077 (N_16077,N_11638,N_13639);
and U16078 (N_16078,N_13154,N_12752);
and U16079 (N_16079,N_10631,N_14451);
nand U16080 (N_16080,N_14128,N_11026);
nor U16081 (N_16081,N_12494,N_13545);
and U16082 (N_16082,N_13246,N_10918);
or U16083 (N_16083,N_14323,N_14546);
and U16084 (N_16084,N_14928,N_13753);
xnor U16085 (N_16085,N_13722,N_14196);
nor U16086 (N_16086,N_13972,N_12821);
nor U16087 (N_16087,N_11495,N_10996);
nor U16088 (N_16088,N_10791,N_10363);
nand U16089 (N_16089,N_14470,N_14813);
or U16090 (N_16090,N_14717,N_13390);
nand U16091 (N_16091,N_11212,N_11711);
or U16092 (N_16092,N_13113,N_11077);
and U16093 (N_16093,N_12242,N_13143);
nor U16094 (N_16094,N_10515,N_10872);
nor U16095 (N_16095,N_11675,N_13522);
xnor U16096 (N_16096,N_13307,N_13328);
nor U16097 (N_16097,N_10145,N_10608);
and U16098 (N_16098,N_13034,N_13319);
or U16099 (N_16099,N_11734,N_13548);
xor U16100 (N_16100,N_12628,N_10242);
nor U16101 (N_16101,N_13469,N_14095);
xnor U16102 (N_16102,N_13466,N_12050);
xnor U16103 (N_16103,N_13995,N_10678);
nand U16104 (N_16104,N_10391,N_11694);
and U16105 (N_16105,N_10210,N_11760);
and U16106 (N_16106,N_10970,N_10606);
nand U16107 (N_16107,N_11669,N_14848);
or U16108 (N_16108,N_14344,N_12490);
nand U16109 (N_16109,N_14996,N_12914);
and U16110 (N_16110,N_12090,N_10058);
or U16111 (N_16111,N_12917,N_11929);
or U16112 (N_16112,N_13290,N_10903);
nand U16113 (N_16113,N_14359,N_10144);
xnor U16114 (N_16114,N_13323,N_13141);
nand U16115 (N_16115,N_10828,N_12085);
nand U16116 (N_16116,N_14115,N_12277);
or U16117 (N_16117,N_13627,N_13719);
xnor U16118 (N_16118,N_12284,N_12783);
nor U16119 (N_16119,N_12667,N_12306);
nor U16120 (N_16120,N_12024,N_12868);
nor U16121 (N_16121,N_13674,N_12988);
and U16122 (N_16122,N_13441,N_13506);
xnor U16123 (N_16123,N_13098,N_10366);
or U16124 (N_16124,N_13363,N_13076);
nor U16125 (N_16125,N_11916,N_14488);
nor U16126 (N_16126,N_13333,N_13539);
nor U16127 (N_16127,N_11069,N_13327);
or U16128 (N_16128,N_11379,N_13049);
xnor U16129 (N_16129,N_10200,N_12904);
nor U16130 (N_16130,N_10422,N_14056);
and U16131 (N_16131,N_10909,N_11389);
nand U16132 (N_16132,N_13045,N_10907);
nand U16133 (N_16133,N_12480,N_13886);
xor U16134 (N_16134,N_14303,N_13185);
nor U16135 (N_16135,N_12201,N_14527);
or U16136 (N_16136,N_10345,N_11618);
nand U16137 (N_16137,N_13175,N_10710);
xnor U16138 (N_16138,N_10949,N_12355);
xnor U16139 (N_16139,N_14785,N_14101);
nand U16140 (N_16140,N_14850,N_11341);
nor U16141 (N_16141,N_14738,N_13099);
nor U16142 (N_16142,N_13625,N_11574);
xnor U16143 (N_16143,N_13683,N_11057);
nor U16144 (N_16144,N_14830,N_13232);
and U16145 (N_16145,N_12990,N_14879);
nor U16146 (N_16146,N_12244,N_11639);
xnor U16147 (N_16147,N_10503,N_10437);
or U16148 (N_16148,N_12776,N_12094);
or U16149 (N_16149,N_13760,N_13846);
and U16150 (N_16150,N_13936,N_14952);
xnor U16151 (N_16151,N_10199,N_12329);
xnor U16152 (N_16152,N_14114,N_11606);
nand U16153 (N_16153,N_14877,N_14011);
xor U16154 (N_16154,N_10684,N_12501);
or U16155 (N_16155,N_10501,N_13144);
nor U16156 (N_16156,N_14823,N_11221);
nand U16157 (N_16157,N_12320,N_14172);
or U16158 (N_16158,N_14456,N_14518);
xnor U16159 (N_16159,N_12663,N_13142);
nand U16160 (N_16160,N_14999,N_11668);
or U16161 (N_16161,N_14428,N_10874);
and U16162 (N_16162,N_12718,N_11634);
nand U16163 (N_16163,N_11671,N_14366);
nor U16164 (N_16164,N_12835,N_10293);
or U16165 (N_16165,N_13594,N_12322);
or U16166 (N_16166,N_10320,N_10274);
or U16167 (N_16167,N_10653,N_10715);
xnor U16168 (N_16168,N_11964,N_10152);
xnor U16169 (N_16169,N_13306,N_14118);
nor U16170 (N_16170,N_11191,N_12308);
nand U16171 (N_16171,N_11567,N_10632);
xnor U16172 (N_16172,N_12309,N_12235);
nand U16173 (N_16173,N_14365,N_12416);
or U16174 (N_16174,N_14238,N_12564);
nand U16175 (N_16175,N_10146,N_12486);
xor U16176 (N_16176,N_11952,N_12164);
and U16177 (N_16177,N_12983,N_13813);
nand U16178 (N_16178,N_10530,N_11200);
or U16179 (N_16179,N_10574,N_14692);
and U16180 (N_16180,N_14349,N_14482);
and U16181 (N_16181,N_12724,N_11361);
xor U16182 (N_16182,N_10476,N_14353);
nor U16183 (N_16183,N_13367,N_11334);
xnor U16184 (N_16184,N_13089,N_14814);
xnor U16185 (N_16185,N_10675,N_12764);
nand U16186 (N_16186,N_13838,N_13636);
xor U16187 (N_16187,N_12323,N_10510);
nor U16188 (N_16188,N_14612,N_12011);
and U16189 (N_16189,N_12114,N_10947);
and U16190 (N_16190,N_14106,N_12214);
nand U16191 (N_16191,N_12471,N_11348);
and U16192 (N_16192,N_10280,N_14013);
xor U16193 (N_16193,N_13334,N_10216);
nor U16194 (N_16194,N_11053,N_12596);
and U16195 (N_16195,N_12283,N_14511);
nor U16196 (N_16196,N_13699,N_13770);
and U16197 (N_16197,N_14619,N_12174);
or U16198 (N_16198,N_14331,N_11446);
and U16199 (N_16199,N_10664,N_14015);
or U16200 (N_16200,N_12432,N_13804);
xnor U16201 (N_16201,N_11161,N_12234);
or U16202 (N_16202,N_14671,N_11336);
xnor U16203 (N_16203,N_11306,N_12813);
or U16204 (N_16204,N_11983,N_12892);
xnor U16205 (N_16205,N_11310,N_13913);
and U16206 (N_16206,N_14552,N_11213);
xnor U16207 (N_16207,N_11006,N_13283);
and U16208 (N_16208,N_12184,N_14539);
and U16209 (N_16209,N_14697,N_12854);
nand U16210 (N_16210,N_12550,N_12572);
or U16211 (N_16211,N_12812,N_14843);
or U16212 (N_16212,N_14108,N_14126);
and U16213 (N_16213,N_13867,N_13992);
xnor U16214 (N_16214,N_11855,N_11275);
nor U16215 (N_16215,N_13582,N_11928);
nor U16216 (N_16216,N_13330,N_13693);
and U16217 (N_16217,N_11484,N_13379);
and U16218 (N_16218,N_11416,N_12658);
and U16219 (N_16219,N_12227,N_12911);
xor U16220 (N_16220,N_14628,N_10054);
or U16221 (N_16221,N_11821,N_13509);
xnor U16222 (N_16222,N_12426,N_11254);
nand U16223 (N_16223,N_11966,N_12379);
nor U16224 (N_16224,N_10062,N_13864);
or U16225 (N_16225,N_13933,N_14750);
and U16226 (N_16226,N_14116,N_12463);
and U16227 (N_16227,N_11619,N_11650);
nand U16228 (N_16228,N_10971,N_14050);
nor U16229 (N_16229,N_10353,N_13075);
nor U16230 (N_16230,N_13429,N_12495);
and U16231 (N_16231,N_10612,N_12909);
or U16232 (N_16232,N_11058,N_12664);
nor U16233 (N_16233,N_11096,N_10017);
or U16234 (N_16234,N_10346,N_13773);
or U16235 (N_16235,N_12057,N_14408);
xor U16236 (N_16236,N_10611,N_11333);
nor U16237 (N_16237,N_12146,N_14852);
xor U16238 (N_16238,N_10850,N_10435);
xnor U16239 (N_16239,N_13430,N_10468);
and U16240 (N_16240,N_10642,N_12933);
and U16241 (N_16241,N_10986,N_11891);
nand U16242 (N_16242,N_11440,N_11370);
or U16243 (N_16243,N_12975,N_13255);
nand U16244 (N_16244,N_10243,N_13297);
or U16245 (N_16245,N_13928,N_12508);
xnor U16246 (N_16246,N_10888,N_10741);
and U16247 (N_16247,N_10866,N_11424);
nor U16248 (N_16248,N_14395,N_11602);
nor U16249 (N_16249,N_14603,N_10559);
nor U16250 (N_16250,N_12918,N_14467);
xnor U16251 (N_16251,N_11483,N_11469);
or U16252 (N_16252,N_14442,N_12240);
xor U16253 (N_16253,N_14956,N_14007);
nor U16254 (N_16254,N_13634,N_14267);
xor U16255 (N_16255,N_14401,N_13308);
nand U16256 (N_16256,N_13159,N_14110);
or U16257 (N_16257,N_14979,N_13961);
xor U16258 (N_16258,N_11073,N_13848);
and U16259 (N_16259,N_12958,N_13607);
nand U16260 (N_16260,N_10288,N_13915);
nor U16261 (N_16261,N_11592,N_10070);
or U16262 (N_16262,N_12078,N_14951);
nand U16263 (N_16263,N_12861,N_10679);
nand U16264 (N_16264,N_10868,N_12238);
and U16265 (N_16265,N_11873,N_14819);
xnor U16266 (N_16266,N_10474,N_12619);
nor U16267 (N_16267,N_13780,N_13225);
nor U16268 (N_16268,N_11448,N_13761);
or U16269 (N_16269,N_11716,N_12987);
or U16270 (N_16270,N_12279,N_10975);
nand U16271 (N_16271,N_14471,N_13489);
or U16272 (N_16272,N_10824,N_12451);
or U16273 (N_16273,N_11193,N_12236);
nand U16274 (N_16274,N_11553,N_11960);
nand U16275 (N_16275,N_10156,N_14183);
or U16276 (N_16276,N_12888,N_12842);
or U16277 (N_16277,N_12644,N_13371);
nor U16278 (N_16278,N_10400,N_12270);
nand U16279 (N_16279,N_10419,N_14512);
and U16280 (N_16280,N_10128,N_10491);
nand U16281 (N_16281,N_10665,N_10621);
nand U16282 (N_16282,N_12604,N_11046);
xor U16283 (N_16283,N_14014,N_13533);
and U16284 (N_16284,N_11897,N_11992);
nand U16285 (N_16285,N_12110,N_12332);
and U16286 (N_16286,N_11977,N_10178);
and U16287 (N_16287,N_11699,N_13019);
nand U16288 (N_16288,N_11854,N_11751);
xor U16289 (N_16289,N_12402,N_10469);
nand U16290 (N_16290,N_14821,N_10130);
nor U16291 (N_16291,N_11119,N_11320);
or U16292 (N_16292,N_10925,N_13162);
nor U16293 (N_16293,N_12527,N_12220);
nor U16294 (N_16294,N_13939,N_14079);
xnor U16295 (N_16295,N_12834,N_14152);
xor U16296 (N_16296,N_14550,N_11656);
and U16297 (N_16297,N_13714,N_13210);
or U16298 (N_16298,N_10049,N_12605);
nand U16299 (N_16299,N_11242,N_13325);
nand U16300 (N_16300,N_10542,N_11687);
or U16301 (N_16301,N_13464,N_13755);
nor U16302 (N_16302,N_11947,N_10941);
xor U16303 (N_16303,N_12041,N_14755);
nor U16304 (N_16304,N_11244,N_14901);
xor U16305 (N_16305,N_14168,N_14937);
or U16306 (N_16306,N_12761,N_11859);
and U16307 (N_16307,N_11318,N_14608);
or U16308 (N_16308,N_14589,N_11386);
or U16309 (N_16309,N_13691,N_10940);
nor U16310 (N_16310,N_13437,N_14683);
nor U16311 (N_16311,N_13082,N_12020);
or U16312 (N_16312,N_12935,N_11787);
nor U16313 (N_16313,N_14147,N_13514);
or U16314 (N_16314,N_11249,N_11943);
nand U16315 (N_16315,N_14725,N_11732);
or U16316 (N_16316,N_14204,N_10101);
nor U16317 (N_16317,N_11722,N_12069);
nor U16318 (N_16318,N_14127,N_11504);
xor U16319 (N_16319,N_13666,N_12537);
and U16320 (N_16320,N_10633,N_12380);
nand U16321 (N_16321,N_14302,N_11518);
or U16322 (N_16322,N_13498,N_14720);
nand U16323 (N_16323,N_12952,N_10719);
and U16324 (N_16324,N_10806,N_11707);
or U16325 (N_16325,N_14855,N_12492);
nor U16326 (N_16326,N_10310,N_13771);
or U16327 (N_16327,N_10981,N_12066);
xnor U16328 (N_16328,N_10408,N_12023);
nand U16329 (N_16329,N_12701,N_10810);
nor U16330 (N_16330,N_10724,N_13757);
nand U16331 (N_16331,N_13630,N_12992);
or U16332 (N_16332,N_10877,N_14842);
and U16333 (N_16333,N_11003,N_10202);
xnor U16334 (N_16334,N_11910,N_12203);
and U16335 (N_16335,N_10276,N_11239);
nand U16336 (N_16336,N_14528,N_13440);
nor U16337 (N_16337,N_14206,N_12950);
or U16338 (N_16338,N_11409,N_11519);
nor U16339 (N_16339,N_10525,N_11585);
nor U16340 (N_16340,N_14555,N_13750);
or U16341 (N_16341,N_12038,N_14317);
and U16342 (N_16342,N_14447,N_12684);
or U16343 (N_16343,N_14109,N_12803);
and U16344 (N_16344,N_13251,N_14188);
and U16345 (N_16345,N_12362,N_13243);
nand U16346 (N_16346,N_11577,N_13110);
or U16347 (N_16347,N_11879,N_13988);
nor U16348 (N_16348,N_10222,N_12543);
and U16349 (N_16349,N_14920,N_10943);
or U16350 (N_16350,N_14143,N_11236);
nor U16351 (N_16351,N_14145,N_14465);
and U16352 (N_16352,N_13606,N_14343);
or U16353 (N_16353,N_11642,N_13863);
nor U16354 (N_16354,N_14443,N_14372);
or U16355 (N_16355,N_11385,N_13216);
and U16356 (N_16356,N_12318,N_13072);
nand U16357 (N_16357,N_11990,N_13291);
nand U16358 (N_16358,N_14387,N_13877);
and U16359 (N_16359,N_13108,N_12280);
nor U16360 (N_16360,N_14562,N_11539);
and U16361 (N_16361,N_12210,N_10804);
nor U16362 (N_16362,N_10127,N_14803);
nor U16363 (N_16363,N_11097,N_14997);
or U16364 (N_16364,N_11824,N_14225);
nor U16365 (N_16365,N_13534,N_10787);
or U16366 (N_16366,N_14868,N_14873);
and U16367 (N_16367,N_10914,N_10330);
nor U16368 (N_16368,N_11789,N_13227);
and U16369 (N_16369,N_13058,N_10396);
or U16370 (N_16370,N_11554,N_12377);
and U16371 (N_16371,N_10979,N_14333);
and U16372 (N_16372,N_14276,N_10927);
nor U16373 (N_16373,N_11841,N_10848);
xor U16374 (N_16374,N_13342,N_10147);
xor U16375 (N_16375,N_14995,N_11792);
and U16376 (N_16376,N_14756,N_13713);
or U16377 (N_16377,N_14543,N_12071);
and U16378 (N_16378,N_13921,N_10584);
xor U16379 (N_16379,N_12021,N_13130);
or U16380 (N_16380,N_13860,N_11251);
nand U16381 (N_16381,N_14681,N_10138);
nor U16382 (N_16382,N_14833,N_10174);
or U16383 (N_16383,N_13413,N_13854);
nor U16384 (N_16384,N_12673,N_12161);
or U16385 (N_16385,N_13396,N_10386);
nor U16386 (N_16386,N_13550,N_10464);
xnor U16387 (N_16387,N_11524,N_11358);
nor U16388 (N_16388,N_13188,N_11968);
and U16389 (N_16389,N_11822,N_10334);
and U16390 (N_16390,N_14626,N_13261);
xor U16391 (N_16391,N_10126,N_12862);
nor U16392 (N_16392,N_12932,N_13811);
nor U16393 (N_16393,N_13009,N_10371);
nand U16394 (N_16394,N_14563,N_10110);
or U16395 (N_16395,N_12378,N_13119);
or U16396 (N_16396,N_10388,N_13841);
nor U16397 (N_16397,N_13505,N_11101);
xor U16398 (N_16398,N_13676,N_13355);
nor U16399 (N_16399,N_10617,N_14917);
and U16400 (N_16400,N_14969,N_11819);
nand U16401 (N_16401,N_14254,N_10610);
and U16402 (N_16402,N_11391,N_14091);
nand U16403 (N_16403,N_10131,N_12608);
xnor U16404 (N_16404,N_13788,N_10297);
nor U16405 (N_16405,N_11474,N_10088);
nor U16406 (N_16406,N_14861,N_13951);
xnor U16407 (N_16407,N_12894,N_13738);
nor U16408 (N_16408,N_13121,N_13927);
or U16409 (N_16409,N_12162,N_10648);
nor U16410 (N_16410,N_13790,N_11837);
or U16411 (N_16411,N_11189,N_12343);
and U16412 (N_16412,N_12186,N_11999);
xnor U16413 (N_16413,N_14306,N_12489);
nand U16414 (N_16414,N_10071,N_11112);
nor U16415 (N_16415,N_12009,N_13480);
nand U16416 (N_16416,N_12117,N_13929);
nor U16417 (N_16417,N_10055,N_12865);
nor U16418 (N_16418,N_11124,N_12082);
and U16419 (N_16419,N_10582,N_11373);
nand U16420 (N_16420,N_13758,N_12593);
or U16421 (N_16421,N_10305,N_10246);
nor U16422 (N_16422,N_14352,N_14902);
nand U16423 (N_16423,N_14312,N_11895);
or U16424 (N_16424,N_13547,N_11645);
nor U16425 (N_16425,N_11274,N_11690);
and U16426 (N_16426,N_11199,N_13301);
or U16427 (N_16427,N_14181,N_10969);
and U16428 (N_16428,N_10496,N_14525);
nand U16429 (N_16429,N_10861,N_12849);
or U16430 (N_16430,N_10461,N_13576);
nand U16431 (N_16431,N_13419,N_12540);
nor U16432 (N_16432,N_11762,N_14237);
or U16433 (N_16433,N_11467,N_11120);
and U16434 (N_16434,N_11146,N_12653);
nand U16435 (N_16435,N_12316,N_13032);
nand U16436 (N_16436,N_13229,N_13107);
nor U16437 (N_16437,N_12696,N_10809);
nor U16438 (N_16438,N_14981,N_14976);
nand U16439 (N_16439,N_11116,N_11682);
and U16440 (N_16440,N_13696,N_13882);
nand U16441 (N_16441,N_10051,N_13549);
xnor U16442 (N_16442,N_13236,N_13844);
and U16443 (N_16443,N_10341,N_14736);
and U16444 (N_16444,N_11100,N_11245);
or U16445 (N_16445,N_13234,N_10602);
or U16446 (N_16446,N_11940,N_11234);
and U16447 (N_16447,N_13135,N_10404);
or U16448 (N_16448,N_13601,N_11698);
or U16449 (N_16449,N_12974,N_14771);
and U16450 (N_16450,N_12488,N_13372);
nor U16451 (N_16451,N_10044,N_14955);
nand U16452 (N_16452,N_11697,N_14878);
nand U16453 (N_16453,N_10817,N_11406);
or U16454 (N_16454,N_10250,N_10669);
and U16455 (N_16455,N_11387,N_10458);
or U16456 (N_16456,N_12648,N_14793);
nand U16457 (N_16457,N_12092,N_12272);
or U16458 (N_16458,N_13193,N_11289);
and U16459 (N_16459,N_14466,N_14425);
nand U16460 (N_16460,N_12973,N_13436);
nand U16461 (N_16461,N_11726,N_10284);
and U16462 (N_16462,N_13869,N_11033);
nor U16463 (N_16463,N_11216,N_11271);
and U16464 (N_16464,N_11998,N_12134);
and U16465 (N_16465,N_13244,N_12680);
nor U16466 (N_16466,N_13911,N_11305);
nand U16467 (N_16467,N_10723,N_13129);
or U16468 (N_16468,N_12460,N_12522);
xor U16469 (N_16469,N_12766,N_13443);
xor U16470 (N_16470,N_11537,N_12155);
nor U16471 (N_16471,N_10438,N_11840);
nor U16472 (N_16472,N_14122,N_10158);
or U16473 (N_16473,N_12836,N_13644);
nor U16474 (N_16474,N_10772,N_14900);
nand U16475 (N_16475,N_13958,N_12084);
nand U16476 (N_16476,N_13462,N_10160);
xor U16477 (N_16477,N_12396,N_12765);
xnor U16478 (N_16478,N_12799,N_12282);
xor U16479 (N_16479,N_12415,N_10083);
nand U16480 (N_16480,N_10841,N_11590);
xor U16481 (N_16481,N_12847,N_10822);
nor U16482 (N_16482,N_13392,N_10998);
nand U16483 (N_16483,N_13400,N_11114);
nand U16484 (N_16484,N_13563,N_14481);
and U16485 (N_16485,N_13875,N_11513);
and U16486 (N_16486,N_14041,N_13962);
nor U16487 (N_16487,N_12115,N_13909);
nand U16488 (N_16488,N_12931,N_14918);
nand U16489 (N_16489,N_14810,N_12885);
and U16490 (N_16490,N_11496,N_14198);
nor U16491 (N_16491,N_10820,N_12297);
nor U16492 (N_16492,N_14102,N_11793);
nor U16493 (N_16493,N_10847,N_11740);
xor U16494 (N_16494,N_14600,N_12263);
nor U16495 (N_16495,N_11436,N_11976);
xor U16496 (N_16496,N_11332,N_14286);
or U16497 (N_16497,N_10765,N_14584);
nor U16498 (N_16498,N_13690,N_11901);
xor U16499 (N_16499,N_10081,N_13467);
xnor U16500 (N_16500,N_10834,N_13900);
xor U16501 (N_16501,N_11020,N_14027);
nor U16502 (N_16502,N_11065,N_14283);
and U16503 (N_16503,N_11653,N_13293);
xnor U16504 (N_16504,N_10591,N_11093);
and U16505 (N_16505,N_12473,N_12191);
and U16506 (N_16506,N_10453,N_12818);
xnor U16507 (N_16507,N_14075,N_13876);
and U16508 (N_16508,N_11404,N_12896);
xnor U16509 (N_16509,N_13668,N_10362);
or U16510 (N_16510,N_12848,N_13235);
nand U16511 (N_16511,N_13605,N_13284);
or U16512 (N_16512,N_10519,N_14450);
or U16513 (N_16513,N_14506,N_13675);
xnor U16514 (N_16514,N_14140,N_12158);
or U16515 (N_16515,N_10257,N_13207);
xnor U16516 (N_16516,N_12999,N_11725);
nand U16517 (N_16517,N_12340,N_12194);
nand U16518 (N_16518,N_10186,N_14253);
xnor U16519 (N_16519,N_11667,N_13239);
xnor U16520 (N_16520,N_11111,N_10640);
or U16521 (N_16521,N_11932,N_12616);
nand U16522 (N_16522,N_12579,N_14592);
and U16523 (N_16523,N_10463,N_11351);
xor U16524 (N_16524,N_12617,N_11252);
or U16525 (N_16525,N_13981,N_12305);
nand U16526 (N_16526,N_13855,N_13241);
xnor U16527 (N_16527,N_13727,N_14072);
nor U16528 (N_16528,N_10801,N_11219);
and U16529 (N_16529,N_10420,N_14055);
nand U16530 (N_16530,N_13809,N_13520);
and U16531 (N_16531,N_11764,N_11076);
and U16532 (N_16532,N_12462,N_13417);
or U16533 (N_16533,N_12660,N_12998);
nor U16534 (N_16534,N_14834,N_13950);
nor U16535 (N_16535,N_11788,N_10770);
nand U16536 (N_16536,N_12738,N_13322);
nand U16537 (N_16537,N_10685,N_11651);
or U16538 (N_16538,N_11366,N_11700);
xnor U16539 (N_16539,N_12635,N_10241);
and U16540 (N_16540,N_10898,N_14364);
nor U16541 (N_16541,N_11094,N_13376);
nor U16542 (N_16542,N_14284,N_13935);
nor U16543 (N_16543,N_11248,N_13134);
xor U16544 (N_16544,N_11705,N_12533);
nand U16545 (N_16545,N_14649,N_12855);
or U16546 (N_16546,N_14531,N_12551);
and U16547 (N_16547,N_13476,N_13577);
xnor U16548 (N_16548,N_12447,N_12346);
xnor U16549 (N_16549,N_12403,N_10006);
nand U16550 (N_16550,N_13955,N_13356);
and U16551 (N_16551,N_14544,N_11728);
nand U16552 (N_16552,N_12185,N_13442);
nand U16553 (N_16553,N_10359,N_10143);
xnor U16554 (N_16554,N_11238,N_14431);
nand U16555 (N_16555,N_11530,N_11779);
or U16556 (N_16556,N_14838,N_14674);
nand U16557 (N_16557,N_12819,N_14418);
nand U16558 (N_16558,N_12252,N_13481);
or U16559 (N_16559,N_10213,N_11629);
or U16560 (N_16560,N_13812,N_11445);
xor U16561 (N_16561,N_11456,N_10390);
xor U16562 (N_16562,N_11950,N_12333);
nor U16563 (N_16563,N_11321,N_10166);
and U16564 (N_16564,N_14452,N_13252);
nand U16565 (N_16565,N_12603,N_11665);
or U16566 (N_16566,N_10945,N_11276);
xor U16567 (N_16567,N_14258,N_11942);
and U16568 (N_16568,N_11118,N_13555);
nand U16569 (N_16569,N_12183,N_10766);
or U16570 (N_16570,N_14946,N_11231);
nand U16571 (N_16571,N_11570,N_13559);
and U16572 (N_16572,N_12145,N_13381);
or U16573 (N_16573,N_11168,N_12588);
xnor U16574 (N_16574,N_10201,N_11951);
or U16575 (N_16575,N_13336,N_12209);
xor U16576 (N_16576,N_11080,N_10952);
or U16577 (N_16577,N_14249,N_13180);
or U16578 (N_16578,N_13310,N_10644);
nand U16579 (N_16579,N_13148,N_11396);
or U16580 (N_16580,N_11517,N_14534);
or U16581 (N_16581,N_12351,N_11526);
and U16582 (N_16582,N_14462,N_12412);
nand U16583 (N_16583,N_14089,N_13493);
or U16584 (N_16584,N_13456,N_10036);
xor U16585 (N_16585,N_10013,N_11515);
or U16586 (N_16586,N_14191,N_13374);
nor U16587 (N_16587,N_12457,N_14679);
xnor U16588 (N_16588,N_11975,N_11613);
nor U16589 (N_16589,N_10326,N_12845);
nand U16590 (N_16590,N_13278,N_10680);
or U16591 (N_16591,N_11541,N_11926);
nor U16592 (N_16592,N_11836,N_14737);
or U16593 (N_16593,N_11883,N_13394);
nand U16594 (N_16594,N_12293,N_13591);
xnor U16595 (N_16595,N_13557,N_11843);
xor U16596 (N_16596,N_10695,N_14078);
nor U16597 (N_16597,N_10219,N_14726);
xor U16598 (N_16598,N_14676,N_12441);
xor U16599 (N_16599,N_11260,N_13529);
nor U16600 (N_16600,N_12509,N_10666);
or U16601 (N_16601,N_13112,N_14702);
nand U16602 (N_16602,N_12080,N_10905);
nor U16603 (N_16603,N_14693,N_14051);
xor U16604 (N_16604,N_12267,N_14179);
or U16605 (N_16605,N_14532,N_11904);
nor U16606 (N_16606,N_14884,N_11492);
or U16607 (N_16607,N_13382,N_14473);
nor U16608 (N_16608,N_14485,N_14604);
and U16609 (N_16609,N_13578,N_10867);
nand U16610 (N_16610,N_11194,N_13797);
xor U16611 (N_16611,N_11368,N_10507);
xor U16612 (N_16612,N_12620,N_13415);
nor U16613 (N_16613,N_12929,N_14730);
and U16614 (N_16614,N_11655,N_14320);
and U16615 (N_16615,N_13990,N_14357);
xnor U16616 (N_16616,N_14300,N_10471);
and U16617 (N_16617,N_11598,N_11648);
nand U16618 (N_16618,N_11316,N_11449);
and U16619 (N_16619,N_13222,N_10260);
and U16620 (N_16620,N_10572,N_13982);
xor U16621 (N_16621,N_10179,N_11703);
nor U16622 (N_16622,N_13926,N_13977);
nand U16623 (N_16623,N_10734,N_10917);
xnor U16624 (N_16624,N_14797,N_11004);
xor U16625 (N_16625,N_12956,N_13828);
xnor U16626 (N_16626,N_12612,N_13647);
and U16627 (N_16627,N_10079,N_11970);
xor U16628 (N_16628,N_14699,N_12565);
and U16629 (N_16629,N_10747,N_14434);
or U16630 (N_16630,N_12253,N_10352);
or U16631 (N_16631,N_11573,N_13568);
and U16632 (N_16632,N_10539,N_12726);
nor U16633 (N_16633,N_13762,N_12294);
xnor U16634 (N_16634,N_14064,N_13687);
nand U16635 (N_16635,N_14645,N_11072);
nand U16636 (N_16636,N_11933,N_12853);
or U16637 (N_16637,N_10092,N_10433);
nand U16638 (N_16638,N_12755,N_13151);
and U16639 (N_16639,N_13817,N_14949);
nor U16640 (N_16640,N_12528,N_10637);
or U16641 (N_16641,N_14350,N_14938);
and U16642 (N_16642,N_13438,N_12192);
and U16643 (N_16643,N_10858,N_10887);
xor U16644 (N_16644,N_10141,N_11068);
nand U16645 (N_16645,N_12980,N_10742);
or U16646 (N_16646,N_10344,N_12903);
nand U16647 (N_16647,N_14711,N_10891);
nor U16648 (N_16648,N_11092,N_11749);
and U16649 (N_16649,N_13257,N_10080);
or U16650 (N_16650,N_10595,N_14547);
nor U16651 (N_16651,N_13698,N_14991);
and U16652 (N_16652,N_14930,N_13628);
or U16653 (N_16653,N_12775,N_13916);
nand U16654 (N_16654,N_14594,N_10832);
xnor U16655 (N_16655,N_14163,N_12286);
nand U16656 (N_16656,N_12889,N_14176);
or U16657 (N_16657,N_10262,N_10740);
and U16658 (N_16658,N_11721,N_13482);
nand U16659 (N_16659,N_10995,N_13910);
or U16660 (N_16660,N_11180,N_11367);
nor U16661 (N_16661,N_10605,N_14881);
nor U16662 (N_16662,N_14941,N_10928);
nor U16663 (N_16663,N_11133,N_11543);
or U16664 (N_16664,N_14036,N_10424);
nor U16665 (N_16665,N_13565,N_12096);
nand U16666 (N_16666,N_12004,N_11892);
or U16667 (N_16667,N_11347,N_10104);
or U16668 (N_16668,N_12541,N_11345);
xor U16669 (N_16669,N_11433,N_11832);
xnor U16670 (N_16670,N_13288,N_11294);
xor U16671 (N_16671,N_12212,N_14751);
nand U16672 (N_16672,N_12883,N_12879);
nor U16673 (N_16673,N_13070,N_12321);
nor U16674 (N_16674,N_11147,N_10953);
xnor U16675 (N_16675,N_12331,N_13967);
or U16676 (N_16676,N_11054,N_14228);
and U16677 (N_16677,N_11393,N_10020);
nor U16678 (N_16678,N_13712,N_10625);
xor U16679 (N_16679,N_10812,N_10545);
nor U16680 (N_16680,N_12744,N_14919);
xnor U16681 (N_16681,N_10025,N_12498);
nor U16682 (N_16682,N_10935,N_11105);
or U16683 (N_16683,N_12255,N_11935);
xnor U16684 (N_16684,N_14313,N_11143);
or U16685 (N_16685,N_10782,N_13311);
xnor U16686 (N_16686,N_12636,N_13983);
nand U16687 (N_16687,N_12708,N_13884);
nand U16688 (N_16688,N_12058,N_10842);
xor U16689 (N_16689,N_12410,N_11241);
nand U16690 (N_16690,N_12381,N_14998);
xor U16691 (N_16691,N_10961,N_10224);
and U16692 (N_16692,N_12168,N_14380);
or U16693 (N_16693,N_12077,N_10650);
xnor U16694 (N_16694,N_11718,N_10365);
nand U16695 (N_16695,N_14016,N_10932);
nand U16696 (N_16696,N_11719,N_11108);
nor U16697 (N_16697,N_11965,N_14409);
nand U16698 (N_16698,N_13487,N_10864);
nor U16699 (N_16699,N_10376,N_11012);
or U16700 (N_16700,N_11501,N_11337);
xor U16701 (N_16701,N_10177,N_13746);
or U16702 (N_16702,N_10172,N_11095);
xor U16703 (N_16703,N_12197,N_14611);
and U16704 (N_16704,N_11848,N_10251);
or U16705 (N_16705,N_11799,N_13792);
nor U16706 (N_16706,N_12138,N_12807);
or U16707 (N_16707,N_12455,N_10450);
nand U16708 (N_16708,N_11750,N_10403);
or U16709 (N_16709,N_10416,N_11912);
or U16710 (N_16710,N_14980,N_11397);
xor U16711 (N_16711,N_11489,N_10792);
xnor U16712 (N_16712,N_10472,N_11863);
and U16713 (N_16713,N_11431,N_12840);
xnor U16714 (N_16714,N_12942,N_14026);
nand U16715 (N_16715,N_12288,N_14992);
xnor U16716 (N_16716,N_12831,N_13858);
nand U16717 (N_16717,N_13271,N_14862);
nand U16718 (N_16718,N_14229,N_14497);
nor U16719 (N_16719,N_14773,N_10277);
nand U16720 (N_16720,N_13414,N_10959);
nor U16721 (N_16721,N_10694,N_12170);
nand U16722 (N_16722,N_12513,N_14334);
nor U16723 (N_16723,N_13891,N_10002);
xnor U16724 (N_16724,N_14293,N_11995);
nand U16725 (N_16725,N_12142,N_14033);
nand U16726 (N_16726,N_14009,N_11865);
or U16727 (N_16727,N_11222,N_11689);
xnor U16728 (N_16728,N_12251,N_12556);
xnor U16729 (N_16729,N_11851,N_14022);
and U16730 (N_16730,N_11523,N_12369);
or U16731 (N_16731,N_13055,N_11502);
xor U16732 (N_16732,N_14910,N_14392);
and U16733 (N_16733,N_10490,N_11922);
nand U16734 (N_16734,N_13697,N_12124);
xor U16735 (N_16735,N_13922,N_14211);
or U16736 (N_16736,N_11583,N_14680);
nand U16737 (N_16737,N_10338,N_11079);
xor U16738 (N_16738,N_12816,N_14644);
xnor U16739 (N_16739,N_10938,N_12246);
or U16740 (N_16740,N_11415,N_11343);
xnor U16741 (N_16741,N_10923,N_12273);
xor U16742 (N_16742,N_11997,N_10999);
nor U16743 (N_16743,N_14739,N_11166);
or U16744 (N_16744,N_14657,N_10763);
nor U16745 (N_16745,N_14940,N_14675);
xnor U16746 (N_16746,N_10328,N_11394);
or U16747 (N_16747,N_13833,N_11670);
nand U16748 (N_16748,N_10823,N_10011);
xnor U16749 (N_16749,N_10774,N_12409);
or U16750 (N_16750,N_10672,N_13618);
xnor U16751 (N_16751,N_11281,N_12438);
nor U16752 (N_16752,N_14460,N_12265);
xor U16753 (N_16753,N_10026,N_10197);
xnor U16754 (N_16754,N_12721,N_13678);
nand U16755 (N_16755,N_11232,N_12797);
and U16756 (N_16756,N_13664,N_13025);
nor U16757 (N_16757,N_10881,N_13999);
xnor U16758 (N_16758,N_10004,N_11031);
and U16759 (N_16759,N_14499,N_14135);
nand U16760 (N_16760,N_14835,N_14583);
xor U16761 (N_16761,N_10299,N_12401);
nor U16762 (N_16762,N_10668,N_14974);
and U16763 (N_16763,N_11874,N_13989);
and U16764 (N_16764,N_13946,N_13952);
nor U16765 (N_16765,N_10816,N_14836);
nor U16766 (N_16766,N_11969,N_11937);
nor U16767 (N_16767,N_13896,N_10670);
nor U16768 (N_16768,N_12137,N_14104);
or U16769 (N_16769,N_13953,N_11427);
nand U16770 (N_16770,N_14248,N_12768);
nor U16771 (N_16771,N_13138,N_14647);
xnor U16772 (N_16772,N_14635,N_14811);
nand U16773 (N_16773,N_14440,N_10394);
nand U16774 (N_16774,N_10466,N_12022);
xor U16775 (N_16775,N_10193,N_12946);
or U16776 (N_16776,N_10977,N_13752);
or U16777 (N_16777,N_13870,N_13095);
and U16778 (N_16778,N_10764,N_14231);
and U16779 (N_16779,N_14841,N_10957);
or U16780 (N_16780,N_10846,N_10852);
or U16781 (N_16781,N_11401,N_11196);
nand U16782 (N_16782,N_11499,N_13149);
xor U16783 (N_16783,N_14386,N_13789);
nor U16784 (N_16784,N_10378,N_14190);
xnor U16785 (N_16785,N_10593,N_14002);
xnor U16786 (N_16786,N_10336,N_13825);
xor U16787 (N_16787,N_12984,N_12759);
nand U16788 (N_16788,N_14239,N_10720);
or U16789 (N_16789,N_10442,N_14475);
and U16790 (N_16790,N_11165,N_12732);
nor U16791 (N_16791,N_14099,N_14153);
nand U16792 (N_16792,N_10659,N_10521);
nand U16793 (N_16793,N_11662,N_11802);
or U16794 (N_16794,N_11402,N_14685);
or U16795 (N_16795,N_14599,N_11930);
nor U16796 (N_16796,N_13282,N_11355);
and U16797 (N_16797,N_10564,N_11599);
and U16798 (N_16798,N_14314,N_13564);
nand U16799 (N_16799,N_12798,N_11810);
nand U16800 (N_16800,N_13358,N_12872);
nor U16801 (N_16801,N_11041,N_11078);
or U16802 (N_16802,N_11061,N_14634);
nand U16803 (N_16803,N_12595,N_11657);
and U16804 (N_16804,N_14660,N_10372);
xnor U16805 (N_16805,N_12221,N_11224);
and U16806 (N_16806,N_12623,N_12228);
and U16807 (N_16807,N_12995,N_12833);
nor U16808 (N_16808,N_13378,N_11085);
and U16809 (N_16809,N_14990,N_13510);
nor U16810 (N_16810,N_14629,N_14700);
nor U16811 (N_16811,N_12278,N_12919);
and U16812 (N_16812,N_14684,N_11455);
xor U16813 (N_16813,N_12651,N_13187);
nand U16814 (N_16814,N_11551,N_10660);
xnor U16815 (N_16815,N_10441,N_12743);
and U16816 (N_16816,N_10651,N_12711);
or U16817 (N_16817,N_10351,N_13314);
and U16818 (N_16818,N_12008,N_12976);
nand U16819 (N_16819,N_14193,N_11807);
xor U16820 (N_16820,N_13611,N_11286);
and U16821 (N_16821,N_13150,N_11550);
xor U16822 (N_16822,N_12793,N_10773);
or U16823 (N_16823,N_13391,N_11680);
nand U16824 (N_16824,N_10007,N_14664);
and U16825 (N_16825,N_13165,N_11207);
or U16826 (N_16826,N_10413,N_10483);
nor U16827 (N_16827,N_12493,N_10482);
xor U16828 (N_16828,N_11042,N_14829);
nand U16829 (N_16829,N_11773,N_13880);
or U16830 (N_16830,N_14031,N_11739);
and U16831 (N_16831,N_10314,N_12700);
or U16832 (N_16832,N_14220,N_13169);
xnor U16833 (N_16833,N_11015,N_14607);
or U16834 (N_16834,N_11919,N_11595);
or U16835 (N_16835,N_14496,N_14070);
nor U16836 (N_16836,N_13598,N_14598);
xnor U16837 (N_16837,N_13206,N_13978);
xor U16838 (N_16838,N_14595,N_14615);
nor U16839 (N_16839,N_13513,N_12470);
or U16840 (N_16840,N_14107,N_12120);
xor U16841 (N_16841,N_11844,N_11163);
or U16842 (N_16842,N_12000,N_11812);
nor U16843 (N_16843,N_12993,N_12723);
xnor U16844 (N_16844,N_11712,N_12703);
nor U16845 (N_16845,N_12982,N_13692);
or U16846 (N_16846,N_10795,N_10066);
and U16847 (N_16847,N_13014,N_14682);
nor U16848 (N_16848,N_12714,N_12099);
or U16849 (N_16849,N_11443,N_12458);
and U16850 (N_16850,N_10649,N_14864);
xor U16851 (N_16851,N_11063,N_11235);
nor U16852 (N_16852,N_10556,N_13729);
xnor U16853 (N_16853,N_12647,N_11183);
or U16854 (N_16854,N_11104,N_10139);
nand U16855 (N_16855,N_13799,N_10737);
nand U16856 (N_16856,N_14377,N_10118);
nand U16857 (N_16857,N_10311,N_12939);
or U16858 (N_16858,N_13344,N_13326);
or U16859 (N_16859,N_14602,N_12757);
nand U16860 (N_16860,N_13287,N_11941);
or U16861 (N_16861,N_12468,N_10355);
xor U16862 (N_16862,N_14519,N_13973);
or U16863 (N_16863,N_11778,N_10046);
nor U16864 (N_16864,N_10335,N_10761);
and U16865 (N_16865,N_14412,N_14837);
xnor U16866 (N_16866,N_11688,N_12589);
nor U16867 (N_16867,N_10428,N_12781);
or U16868 (N_16868,N_11559,N_11681);
or U16869 (N_16869,N_12858,N_13893);
and U16870 (N_16870,N_10077,N_14931);
and U16871 (N_16871,N_11126,N_10157);
nand U16872 (N_16872,N_11786,N_14658);
xnor U16873 (N_16873,N_11293,N_10671);
xor U16874 (N_16874,N_14034,N_13906);
and U16875 (N_16875,N_11262,N_11829);
and U16876 (N_16876,N_13094,N_10758);
xor U16877 (N_16877,N_10553,N_13504);
or U16878 (N_16878,N_12035,N_12356);
nor U16879 (N_16879,N_12211,N_11899);
and U16880 (N_16880,N_10783,N_10662);
and U16881 (N_16881,N_10748,N_11660);
or U16882 (N_16882,N_12125,N_13027);
and U16883 (N_16883,N_12921,N_10643);
nor U16884 (N_16884,N_10196,N_11885);
nor U16885 (N_16885,N_10912,N_12224);
and U16886 (N_16886,N_14719,N_14536);
nand U16887 (N_16887,N_12656,N_13635);
xnor U16888 (N_16888,N_13688,N_11034);
and U16889 (N_16889,N_12682,N_12063);
nand U16890 (N_16890,N_14141,N_10645);
nor U16891 (N_16891,N_12727,N_14241);
nand U16892 (N_16892,N_13518,N_10095);
or U16893 (N_16893,N_11604,N_10727);
xnor U16894 (N_16894,N_13155,N_11299);
or U16895 (N_16895,N_11520,N_11971);
and U16896 (N_16896,N_12913,N_13659);
or U16897 (N_16897,N_10524,N_11214);
or U16898 (N_16898,N_13626,N_11365);
or U16899 (N_16899,N_12098,N_14535);
nor U16900 (N_16900,N_12219,N_12422);
and U16901 (N_16901,N_14763,N_11701);
nor U16902 (N_16902,N_14246,N_14686);
nor U16903 (N_16903,N_11284,N_12437);
and U16904 (N_16904,N_14338,N_14000);
nor U16905 (N_16905,N_13132,N_11307);
nor U16906 (N_16906,N_10427,N_11419);
nand U16907 (N_16907,N_11159,N_10797);
and U16908 (N_16908,N_13264,N_10283);
or U16909 (N_16909,N_12817,N_12440);
or U16910 (N_16910,N_10862,N_11369);
or U16911 (N_16911,N_14622,N_12141);
xnor U16912 (N_16912,N_14870,N_12013);
nand U16913 (N_16913,N_11752,N_14677);
nand U16914 (N_16914,N_14463,N_11246);
nor U16915 (N_16915,N_11738,N_13275);
xor U16916 (N_16916,N_14964,N_10781);
nand U16917 (N_16917,N_12583,N_13351);
xnor U16918 (N_16918,N_14794,N_13250);
and U16919 (N_16919,N_12748,N_12719);
nand U16920 (N_16920,N_12268,N_12167);
nor U16921 (N_16921,N_10991,N_12820);
nor U16922 (N_16922,N_14545,N_14419);
xnor U16923 (N_16923,N_13871,N_12649);
nand U16924 (N_16924,N_14346,N_13125);
and U16925 (N_16925,N_12792,N_11784);
or U16926 (N_16926,N_12576,N_10402);
xnor U16927 (N_16927,N_14882,N_12876);
and U16928 (N_16928,N_11190,N_14296);
and U16929 (N_16929,N_14189,N_11663);
xor U16930 (N_16930,N_11544,N_10342);
xor U16931 (N_16931,N_14501,N_10851);
or U16932 (N_16932,N_11418,N_10619);
or U16933 (N_16933,N_14905,N_10380);
nor U16934 (N_16934,N_13179,N_14963);
xnor U16935 (N_16935,N_14416,N_11277);
xnor U16936 (N_16936,N_14149,N_10698);
nand U16937 (N_16937,N_12045,N_10677);
nor U16938 (N_16938,N_10367,N_12754);
or U16939 (N_16939,N_10121,N_12208);
or U16940 (N_16940,N_11535,N_11088);
xor U16941 (N_16941,N_14400,N_13700);
and U16942 (N_16942,N_10844,N_14063);
nor U16943 (N_16943,N_12223,N_13131);
and U16944 (N_16944,N_10951,N_14493);
and U16945 (N_16945,N_12408,N_12552);
or U16946 (N_16946,N_13818,N_11049);
nand U16947 (N_16947,N_14087,N_11490);
nor U16948 (N_16948,N_13339,N_12674);
xor U16949 (N_16949,N_11861,N_14480);
nand U16950 (N_16950,N_12373,N_10426);
nor U16951 (N_16951,N_11013,N_13494);
nor U16952 (N_16952,N_13079,N_10031);
xor U16953 (N_16953,N_14789,N_11152);
and U16954 (N_16954,N_13196,N_11989);
nor U16955 (N_16955,N_11644,N_10615);
nor U16956 (N_16956,N_12609,N_14489);
nand U16957 (N_16957,N_13471,N_14820);
xor U16958 (N_16958,N_14966,N_11506);
nand U16959 (N_16959,N_13894,N_12689);
and U16960 (N_16960,N_10456,N_12969);
nor U16961 (N_16961,N_13166,N_10716);
or U16962 (N_16962,N_10451,N_10860);
nor U16963 (N_16963,N_10985,N_10845);
nand U16964 (N_16964,N_11508,N_14413);
or U16965 (N_16965,N_12637,N_12908);
or U16966 (N_16966,N_14654,N_10594);
or U16967 (N_16967,N_10752,N_10601);
nor U16968 (N_16968,N_11561,N_11188);
xor U16969 (N_16969,N_11774,N_13711);
and U16970 (N_16970,N_12016,N_14606);
nand U16971 (N_16971,N_10768,N_14006);
nor U16972 (N_16972,N_12900,N_14182);
and U16973 (N_16973,N_12591,N_11713);
nor U16974 (N_16974,N_12769,N_10037);
nor U16975 (N_16975,N_13940,N_13133);
xor U16976 (N_16976,N_12342,N_11150);
or U16977 (N_16977,N_11533,N_13393);
or U16978 (N_16978,N_12485,N_14804);
nand U16979 (N_16979,N_14311,N_12963);
or U16980 (N_16980,N_12299,N_13980);
and U16981 (N_16981,N_13836,N_12874);
nor U16982 (N_16982,N_11128,N_11417);
nand U16983 (N_16983,N_14740,N_11331);
nor U16984 (N_16984,N_13364,N_12172);
nand U16985 (N_16985,N_12928,N_10035);
xor U16986 (N_16986,N_10410,N_12745);
and U16987 (N_16987,N_14510,N_11815);
or U16988 (N_16988,N_12358,N_10103);
and U16989 (N_16989,N_10906,N_12655);
and U16990 (N_16990,N_14291,N_14788);
or U16991 (N_16991,N_10286,N_13919);
or U16992 (N_16992,N_13037,N_11867);
and U16993 (N_16993,N_14269,N_10209);
nor U16994 (N_16994,N_10059,N_13178);
or U16995 (N_16995,N_11141,N_11860);
nor U16996 (N_16996,N_10517,N_11616);
or U16997 (N_16997,N_12867,N_14356);
nor U16998 (N_16998,N_11601,N_10385);
nor U16999 (N_16999,N_13749,N_10229);
and U17000 (N_17000,N_10112,N_13966);
or U17001 (N_17001,N_14989,N_12376);
and U17002 (N_17002,N_12905,N_14441);
xnor U17003 (N_17003,N_12557,N_12871);
nand U17004 (N_17004,N_11884,N_14279);
nand U17005 (N_17005,N_12100,N_10072);
or U17006 (N_17006,N_12196,N_12287);
and U17007 (N_17007,N_12507,N_14484);
nor U17008 (N_17008,N_11803,N_13071);
or U17009 (N_17009,N_11329,N_10440);
nor U17010 (N_17010,N_10423,N_14560);
nor U17011 (N_17011,N_13182,N_14973);
xor U17012 (N_17012,N_14703,N_11171);
nor U17013 (N_17013,N_13530,N_11342);
or U17014 (N_17014,N_10093,N_12640);
and U17015 (N_17015,N_13866,N_14787);
nand U17016 (N_17016,N_10392,N_10630);
and U17017 (N_17017,N_10638,N_13360);
xor U17018 (N_17018,N_12996,N_10609);
nor U17019 (N_17019,N_11709,N_13247);
nand U17020 (N_17020,N_10028,N_10161);
and U17021 (N_17021,N_13484,N_13620);
nand U17022 (N_17022,N_14235,N_11534);
nor U17023 (N_17023,N_10078,N_12562);
nand U17024 (N_17024,N_10600,N_13767);
xor U17025 (N_17025,N_10936,N_11228);
nor U17026 (N_17026,N_14042,N_12925);
nor U17027 (N_17027,N_10798,N_11710);
nand U17028 (N_17028,N_11894,N_13584);
nor U17029 (N_17029,N_14672,N_13835);
nand U17030 (N_17030,N_14709,N_11407);
nor U17031 (N_17031,N_14721,N_10042);
or U17032 (N_17032,N_10124,N_13681);
xnor U17033 (N_17033,N_13763,N_11569);
or U17034 (N_17034,N_10048,N_11633);
or U17035 (N_17035,N_12421,N_13220);
or U17036 (N_17036,N_14571,N_10882);
and U17037 (N_17037,N_11905,N_12067);
nor U17038 (N_17038,N_13402,N_11218);
nor U17039 (N_17039,N_14173,N_12189);
nand U17040 (N_17040,N_11037,N_14731);
or U17041 (N_17041,N_12880,N_12778);
and U17042 (N_17042,N_12826,N_11265);
xor U17043 (N_17043,N_12248,N_11880);
nor U17044 (N_17044,N_12773,N_12856);
or U17045 (N_17045,N_12830,N_14752);
and U17046 (N_17046,N_13643,N_11597);
and U17047 (N_17047,N_11090,N_13993);
nand U17048 (N_17048,N_13745,N_13318);
xor U17049 (N_17049,N_13146,N_12389);
xnor U17050 (N_17050,N_10658,N_14410);
xnor U17051 (N_17051,N_11717,N_13542);
or U17052 (N_17052,N_13174,N_14278);
and U17053 (N_17053,N_14623,N_11775);
and U17054 (N_17054,N_11261,N_10819);
or U17055 (N_17055,N_10485,N_14894);
or U17056 (N_17056,N_14641,N_12806);
nor U17057 (N_17057,N_12736,N_14860);
xnor U17058 (N_17058,N_14840,N_13317);
nand U17059 (N_17059,N_13389,N_11398);
nand U17060 (N_17060,N_13309,N_13177);
and U17061 (N_17061,N_14943,N_11282);
and U17062 (N_17062,N_13511,N_12960);
nand U17063 (N_17063,N_12423,N_10096);
nor U17064 (N_17064,N_10965,N_14318);
and U17065 (N_17065,N_12737,N_10835);
xor U17066 (N_17066,N_14944,N_13460);
nand U17067 (N_17067,N_12786,N_12180);
and U17068 (N_17068,N_14088,N_10218);
nand U17069 (N_17069,N_13562,N_11444);
nor U17070 (N_17070,N_13735,N_11029);
and U17071 (N_17071,N_10397,N_11167);
or U17072 (N_17072,N_10786,N_12349);
and U17073 (N_17073,N_10003,N_14053);
or U17074 (N_17074,N_14617,N_12964);
and U17075 (N_17075,N_11098,N_12044);
xnor U17076 (N_17076,N_13340,N_10974);
nand U17077 (N_17077,N_11315,N_10191);
xnor U17078 (N_17078,N_12751,N_14817);
xnor U17079 (N_17079,N_14633,N_12741);
or U17080 (N_17080,N_11678,N_12104);
xnor U17081 (N_17081,N_14175,N_12823);
xnor U17082 (N_17082,N_13245,N_11312);
nor U17083 (N_17083,N_14885,N_12487);
or U17084 (N_17084,N_12239,N_10883);
nor U17085 (N_17085,N_12989,N_13081);
xor U17086 (N_17086,N_10481,N_14661);
nand U17087 (N_17087,N_11677,N_13791);
or U17088 (N_17088,N_10443,N_11605);
nand U17089 (N_17089,N_10623,N_12427);
nand U17090 (N_17090,N_10560,N_11018);
nor U17091 (N_17091,N_13204,N_14809);
nand U17092 (N_17092,N_10626,N_12679);
and U17093 (N_17093,N_14710,N_10580);
and U17094 (N_17094,N_14200,N_10728);
xnor U17095 (N_17095,N_14895,N_13862);
and U17096 (N_17096,N_14468,N_11907);
nor U17097 (N_17097,N_13662,N_14907);
and U17098 (N_17098,N_10547,N_13137);
and U17099 (N_17099,N_12986,N_14538);
and U17100 (N_17100,N_10102,N_13062);
nand U17101 (N_17101,N_13425,N_14783);
or U17102 (N_17102,N_10073,N_14753);
xor U17103 (N_17103,N_14806,N_12241);
xnor U17104 (N_17104,N_11944,N_11055);
nor U17105 (N_17105,N_14911,N_10873);
nor U17106 (N_17106,N_14207,N_13312);
or U17107 (N_17107,N_11729,N_12357);
or U17108 (N_17108,N_13695,N_10738);
nor U17109 (N_17109,N_11936,N_12399);
or U17110 (N_17110,N_10980,N_11801);
or U17111 (N_17111,N_12160,N_14083);
nand U17112 (N_17112,N_12119,N_14520);
xor U17113 (N_17113,N_10266,N_11582);
nand U17114 (N_17114,N_12344,N_13021);
nand U17115 (N_17115,N_14505,N_13401);
or U17116 (N_17116,N_10090,N_11962);
nand U17117 (N_17117,N_10374,N_10735);
and U17118 (N_17118,N_11360,N_12479);
nor U17119 (N_17119,N_14375,N_13917);
and U17120 (N_17120,N_13508,N_11466);
or U17121 (N_17121,N_10808,N_13595);
nor U17122 (N_17122,N_10187,N_11877);
nor U17123 (N_17123,N_12179,N_10446);
nand U17124 (N_17124,N_13941,N_13473);
and U17125 (N_17125,N_13249,N_10929);
or U17126 (N_17126,N_14234,N_11771);
nand U17127 (N_17127,N_13263,N_13879);
and U17128 (N_17128,N_12250,N_11047);
and U17129 (N_17129,N_13837,N_11434);
nor U17130 (N_17130,N_13517,N_10916);
or U17131 (N_17131,N_14177,N_13136);
or U17132 (N_17132,N_14845,N_10629);
nor U17133 (N_17133,N_14280,N_10302);
nand U17134 (N_17134,N_14045,N_14247);
and U17135 (N_17135,N_12666,N_10833);
and U17136 (N_17136,N_14131,N_11889);
or U17137 (N_17137,N_12516,N_13012);
xor U17138 (N_17138,N_13122,N_10084);
and U17139 (N_17139,N_14478,N_10214);
nor U17140 (N_17140,N_10588,N_12573);
xnor U17141 (N_17141,N_11083,N_12502);
nand U17142 (N_17142,N_13035,N_10744);
or U17143 (N_17143,N_13153,N_12979);
or U17144 (N_17144,N_14724,N_10596);
and U17145 (N_17145,N_12325,N_14337);
nand U17146 (N_17146,N_14210,N_11021);
xor U17147 (N_17147,N_14754,N_14212);
xor U17148 (N_17148,N_14092,N_13803);
nor U17149 (N_17149,N_14399,N_11115);
and U17150 (N_17150,N_14219,N_10731);
or U17151 (N_17151,N_12961,N_11442);
nor U17152 (N_17152,N_11696,N_10455);
nand U17153 (N_17153,N_10933,N_12311);
and U17154 (N_17154,N_10759,N_12226);
or U17155 (N_17155,N_10984,N_12345);
nand U17156 (N_17156,N_13101,N_10529);
nor U17157 (N_17157,N_12307,N_12691);
nand U17158 (N_17158,N_10587,N_12407);
and U17159 (N_17159,N_12716,N_14393);
xor U17160 (N_17160,N_10029,N_14959);
and U17161 (N_17161,N_12912,N_13217);
nor U17162 (N_17162,N_11138,N_10142);
xor U17163 (N_17163,N_14564,N_10988);
or U17164 (N_17164,N_13039,N_14185);
nand U17165 (N_17165,N_12962,N_11991);
nor U17166 (N_17166,N_13386,N_13741);
nor U17167 (N_17167,N_12476,N_11256);
xnor U17168 (N_17168,N_10383,N_14896);
and U17169 (N_17169,N_14476,N_13987);
or U17170 (N_17170,N_12555,N_10522);
and U17171 (N_17171,N_11350,N_12153);
nand U17172 (N_17172,N_13191,N_11772);
xnor U17173 (N_17173,N_11768,N_13815);
and U17174 (N_17174,N_13527,N_11229);
nand U17175 (N_17175,N_12859,N_12387);
or U17176 (N_17176,N_10045,N_10667);
nand U17177 (N_17177,N_11875,N_11600);
xor U17178 (N_17178,N_14590,N_11635);
xor U17179 (N_17179,N_11979,N_14786);
and U17180 (N_17180,N_12435,N_13798);
nand U17181 (N_17181,N_12296,N_10258);
nor U17182 (N_17182,N_10256,N_10169);
nor U17183 (N_17183,N_10154,N_13938);
nor U17184 (N_17184,N_13114,N_11176);
nor U17185 (N_17185,N_13596,N_10030);
and U17186 (N_17186,N_10068,N_14758);
nor U17187 (N_17187,N_14530,N_13540);
nand U17188 (N_17188,N_11311,N_10018);
or U17189 (N_17189,N_13046,N_14120);
nor U17190 (N_17190,N_11392,N_11135);
nor U17191 (N_17191,N_11399,N_14696);
or U17192 (N_17192,N_10194,N_14446);
nor U17193 (N_17193,N_13787,N_14097);
or U17194 (N_17194,N_13865,N_12046);
xnor U17195 (N_17195,N_11227,N_13490);
nand U17196 (N_17196,N_11898,N_14777);
or U17197 (N_17197,N_14807,N_10508);
or U17198 (N_17198,N_13240,N_12157);
nand U17199 (N_17199,N_13772,N_12292);
nand U17200 (N_17200,N_14994,N_12514);
nand U17201 (N_17201,N_12392,N_11136);
nand U17202 (N_17202,N_14948,N_13373);
xor U17203 (N_17203,N_14723,N_13092);
nand U17204 (N_17204,N_14765,N_11001);
nor U17205 (N_17205,N_11731,N_13495);
nor U17206 (N_17206,N_13944,N_12669);
nor U17207 (N_17207,N_13868,N_10429);
nand U17208 (N_17208,N_14886,N_12955);
nand U17209 (N_17209,N_14297,N_12386);
nand U17210 (N_17210,N_10885,N_14734);
nand U17211 (N_17211,N_14432,N_12089);
xor U17212 (N_17212,N_10908,N_13316);
or U17213 (N_17213,N_11089,N_10254);
nor U17214 (N_17214,N_10900,N_14601);
and U17215 (N_17215,N_11876,N_12143);
nor U17216 (N_17216,N_10533,N_14417);
nand U17217 (N_17217,N_14888,N_10032);
or U17218 (N_17218,N_11421,N_10897);
nor U17219 (N_17219,N_11081,N_12154);
or U17220 (N_17220,N_11149,N_13047);
or U17221 (N_17221,N_11390,N_11264);
xor U17222 (N_17222,N_13669,N_13005);
nor U17223 (N_17223,N_12630,N_14373);
and U17224 (N_17224,N_11654,N_10484);
or U17225 (N_17225,N_12715,N_10636);
nor U17226 (N_17226,N_13808,N_13759);
nand U17227 (N_17227,N_12621,N_11062);
xor U17228 (N_17228,N_13551,N_13001);
or U17229 (N_17229,N_11825,N_14461);
xor U17230 (N_17230,N_12746,N_14157);
xnor U17231 (N_17231,N_12205,N_10231);
nor U17232 (N_17232,N_11591,N_12887);
xnor U17233 (N_17233,N_11637,N_14326);
or U17234 (N_17234,N_14221,N_10119);
nand U17235 (N_17235,N_12574,N_12453);
xnor U17236 (N_17236,N_13685,N_11835);
nor U17237 (N_17237,N_12232,N_11959);
or U17238 (N_17238,N_12204,N_12007);
nor U17239 (N_17239,N_11330,N_10703);
xor U17240 (N_17240,N_13786,N_14052);
xnor U17241 (N_17241,N_11113,N_13474);
nor U17242 (N_17242,N_11536,N_10829);
nor U17243 (N_17243,N_14385,N_13589);
nor U17244 (N_17244,N_14151,N_10628);
and U17245 (N_17245,N_13889,N_10886);
and U17246 (N_17246,N_14281,N_10340);
nand U17247 (N_17247,N_10657,N_14383);
or U17248 (N_17248,N_11441,N_13345);
or U17249 (N_17249,N_10331,N_10532);
or U17250 (N_17250,N_10236,N_10221);
nand U17251 (N_17251,N_12360,N_10115);
nor U17252 (N_17252,N_11130,N_11512);
xor U17253 (N_17253,N_12048,N_11040);
nor U17254 (N_17254,N_11450,N_11896);
and U17255 (N_17255,N_13609,N_12163);
or U17256 (N_17256,N_12906,N_12547);
xor U17257 (N_17257,N_11043,N_12934);
or U17258 (N_17258,N_10896,N_10249);
nand U17259 (N_17259,N_10788,N_10164);
and U17260 (N_17260,N_10086,N_13431);
or U17261 (N_17261,N_14186,N_13903);
or U17262 (N_17262,N_14213,N_10683);
nand U17263 (N_17263,N_14001,N_14533);
nand U17264 (N_17264,N_12353,N_12531);
nand U17265 (N_17265,N_12474,N_11620);
xnor U17266 (N_17266,N_12580,N_14551);
nor U17267 (N_17267,N_11324,N_11587);
nand U17268 (N_17268,N_12677,N_10993);
xor U17269 (N_17269,N_11383,N_12467);
xnor U17270 (N_17270,N_12870,N_10235);
or U17271 (N_17271,N_12560,N_11809);
or U17272 (N_17272,N_12549,N_12101);
nand U17273 (N_17273,N_13883,N_12811);
or U17274 (N_17274,N_14666,N_11528);
nand U17275 (N_17275,N_14472,N_13299);
xnor U17276 (N_17276,N_12481,N_14427);
nand U17277 (N_17277,N_11233,N_10324);
nor U17278 (N_17278,N_10185,N_14421);
and U17279 (N_17279,N_12808,N_10008);
xnor U17280 (N_17280,N_12832,N_11011);
nand U17281 (N_17281,N_14361,N_12742);
xnor U17282 (N_17282,N_10956,N_10815);
or U17283 (N_17283,N_11172,N_11858);
xor U17284 (N_17284,N_12126,N_13242);
nor U17285 (N_17285,N_10878,N_12338);
nand U17286 (N_17286,N_13934,N_10646);
nor U17287 (N_17287,N_12881,N_14035);
nand U17288 (N_17288,N_14580,N_14012);
xor U17289 (N_17289,N_12131,N_13412);
and U17290 (N_17290,N_11659,N_10722);
nor U17291 (N_17291,N_11287,N_13816);
xor U17292 (N_17292,N_14223,N_10849);
and U17293 (N_17293,N_13189,N_14486);
or U17294 (N_17294,N_13744,N_12801);
nand U17295 (N_17295,N_13087,N_13061);
nand U17296 (N_17296,N_12805,N_14028);
nor U17297 (N_17297,N_13890,N_14024);
or U17298 (N_17298,N_14748,N_14742);
or U17299 (N_17299,N_14129,N_10056);
nand U17300 (N_17300,N_10926,N_11805);
nand U17301 (N_17301,N_10252,N_11674);
or U17302 (N_17302,N_13041,N_10291);
nand U17303 (N_17303,N_10992,N_11850);
and U17304 (N_17304,N_12065,N_10613);
nand U17305 (N_17305,N_11203,N_11797);
and U17306 (N_17306,N_10377,N_13834);
xor U17307 (N_17307,N_12971,N_12166);
nor U17308 (N_17308,N_12029,N_11498);
nand U17309 (N_17309,N_14965,N_11988);
and U17310 (N_17310,N_11996,N_11522);
nand U17311 (N_17311,N_12198,N_12361);
nand U17312 (N_17312,N_14162,N_14846);
and U17313 (N_17313,N_14880,N_13219);
nand U17314 (N_17314,N_10652,N_13553);
or U17315 (N_17315,N_10514,N_13571);
xnor U17316 (N_17316,N_14187,N_11886);
nor U17317 (N_17317,N_14701,N_10551);
and U17318 (N_17318,N_12136,N_12072);
or U17319 (N_17319,N_14744,N_13781);
nor U17320 (N_17320,N_11400,N_12526);
or U17321 (N_17321,N_13827,N_14275);
nand U17322 (N_17322,N_11566,N_13002);
nor U17323 (N_17323,N_10033,N_11847);
nor U17324 (N_17324,N_13597,N_11980);
nor U17325 (N_17325,N_12902,N_13892);
or U17326 (N_17326,N_10087,N_13186);
nand U17327 (N_17327,N_11290,N_14983);
xor U17328 (N_17328,N_10205,N_11906);
nor U17329 (N_17329,N_13080,N_10294);
nand U17330 (N_17330,N_14165,N_11082);
or U17331 (N_17331,N_11005,N_10486);
nor U17332 (N_17332,N_10237,N_11363);
xnor U17333 (N_17333,N_13248,N_13819);
xnor U17334 (N_17334,N_14741,N_12317);
nand U17335 (N_17335,N_11014,N_11568);
or U17336 (N_17336,N_14597,N_10871);
and U17337 (N_17337,N_14557,N_14689);
and U17338 (N_17338,N_11767,N_14137);
nor U17339 (N_17339,N_11460,N_12256);
xor U17340 (N_17340,N_10964,N_13126);
nand U17341 (N_17341,N_13052,N_14226);
and U17342 (N_17342,N_14195,N_11765);
nand U17343 (N_17343,N_10034,N_13423);
and U17344 (N_17344,N_14439,N_12965);
xnor U17345 (N_17345,N_14967,N_11527);
or U17346 (N_17346,N_13920,N_13463);
nand U17347 (N_17347,N_11915,N_11487);
xnor U17348 (N_17348,N_14328,N_10674);
or U17349 (N_17349,N_10393,N_10108);
nand U17350 (N_17350,N_12295,N_14327);
and U17351 (N_17351,N_14732,N_14345);
or U17352 (N_17352,N_13823,N_11215);
nand U17353 (N_17353,N_11987,N_14124);
xnor U17354 (N_17354,N_13593,N_10167);
nor U17355 (N_17355,N_12269,N_11405);
xor U17356 (N_17356,N_11571,N_10686);
nor U17357 (N_17357,N_10343,N_10067);
and U17358 (N_17358,N_14854,N_14259);
or U17359 (N_17359,N_14335,N_14438);
xor U17360 (N_17360,N_14503,N_14336);
xor U17361 (N_17361,N_13845,N_11465);
nor U17362 (N_17362,N_10743,N_13416);
nor U17363 (N_17363,N_11685,N_10681);
and U17364 (N_17364,N_11285,N_12758);
nand U17365 (N_17365,N_13969,N_13267);
nand U17366 (N_17366,N_13418,N_14766);
nand U17367 (N_17367,N_10479,N_11949);
nor U17368 (N_17368,N_11056,N_11817);
or U17369 (N_17369,N_11790,N_10165);
nor U17370 (N_17370,N_12504,N_13631);
or U17371 (N_17371,N_11967,N_10462);
and U17372 (N_17372,N_13718,N_11507);
or U17373 (N_17373,N_14627,N_13569);
nor U17374 (N_17374,N_10457,N_10211);
nor U17375 (N_17375,N_12529,N_13478);
nor U17376 (N_17376,N_12782,N_11909);
and U17377 (N_17377,N_12003,N_13650);
and U17378 (N_17378,N_14307,N_12681);
xnor U17379 (N_17379,N_12028,N_11626);
nand U17380 (N_17380,N_13399,N_11766);
xor U17381 (N_17381,N_11226,N_10538);
nand U17382 (N_17382,N_13905,N_10944);
nor U17383 (N_17383,N_14985,N_13018);
xor U17384 (N_17384,N_12582,N_11205);
or U17385 (N_17385,N_10133,N_10544);
nand U17386 (N_17386,N_12747,N_12512);
or U17387 (N_17387,N_12558,N_10285);
and U17388 (N_17388,N_13091,N_14159);
nand U17389 (N_17389,N_11266,N_13028);
and U17390 (N_17390,N_10528,N_14587);
or U17391 (N_17391,N_14457,N_11309);
and U17392 (N_17392,N_13353,N_13839);
nor U17393 (N_17393,N_14790,N_13723);
nor U17394 (N_17394,N_14925,N_14784);
or U17395 (N_17395,N_10661,N_10585);
nand U17396 (N_17396,N_13899,N_12367);
or U17397 (N_17397,N_10913,N_13907);
and U17398 (N_17398,N_12546,N_11204);
xnor U17399 (N_17399,N_11335,N_10597);
nand U17400 (N_17400,N_10105,N_14271);
xor U17401 (N_17401,N_14046,N_10579);
nand U17402 (N_17402,N_12393,N_13778);
nor U17403 (N_17403,N_12728,N_13538);
xor U17404 (N_17404,N_14746,N_10132);
nor U17405 (N_17405,N_13914,N_14541);
nor U17406 (N_17406,N_14694,N_10136);
xor U17407 (N_17407,N_13629,N_14487);
nor U17408 (N_17408,N_10189,N_13532);
or U17409 (N_17409,N_12683,N_13665);
nor U17410 (N_17410,N_12182,N_14524);
nor U17411 (N_17411,N_12787,N_11769);
or U17412 (N_17412,N_13521,N_14382);
nand U17413 (N_17413,N_12611,N_13346);
or U17414 (N_17414,N_11755,N_13459);
nand U17415 (N_17415,N_13298,N_10495);
nand U17416 (N_17416,N_12503,N_12371);
nor U17417 (N_17417,N_10009,N_13302);
nor U17418 (N_17418,N_13820,N_10693);
nor U17419 (N_17419,N_12720,N_12026);
and U17420 (N_17420,N_13026,N_13434);
and U17421 (N_17421,N_11881,N_12706);
xor U17422 (N_17422,N_11217,N_11691);
nor U17423 (N_17423,N_13793,N_14832);
and U17424 (N_17424,N_10967,N_11882);
nand U17425 (N_17425,N_13954,N_10325);
and U17426 (N_17426,N_11356,N_11439);
nor U17427 (N_17427,N_14321,N_11586);
nand U17428 (N_17428,N_13409,N_11326);
or U17429 (N_17429,N_11708,N_12225);
xnor U17430 (N_17430,N_11381,N_13543);
xor U17431 (N_17431,N_13895,N_14986);
and U17432 (N_17432,N_13090,N_10109);
nand U17433 (N_17433,N_14105,N_14561);
xnor U17434 (N_17434,N_12430,N_11195);
xor U17435 (N_17435,N_10329,N_10270);
nand U17436 (N_17436,N_11458,N_10000);
or U17437 (N_17437,N_14668,N_13918);
nand U17438 (N_17438,N_12750,N_13069);
xor U17439 (N_17439,N_12967,N_13764);
or U17440 (N_17440,N_13824,N_11278);
or U17441 (N_17441,N_11481,N_11225);
or U17442 (N_17442,N_13932,N_11371);
nand U17443 (N_17443,N_12511,N_10369);
and U17444 (N_17444,N_14642,N_13320);
nand U17445 (N_17445,N_11946,N_10570);
nand U17446 (N_17446,N_12372,N_11035);
nor U17447 (N_17447,N_12122,N_12852);
xor U17448 (N_17448,N_13579,N_13531);
nand U17449 (N_17449,N_11028,N_14367);
and U17450 (N_17450,N_12259,N_12336);
nand U17451 (N_17451,N_10106,N_11756);
nand U17452 (N_17452,N_13561,N_11715);
or U17453 (N_17453,N_10183,N_13887);
and U17454 (N_17454,N_13152,N_14802);
nor U17455 (N_17455,N_12123,N_14407);
and U17456 (N_17456,N_14665,N_13084);
xnor U17457 (N_17457,N_12694,N_11352);
xor U17458 (N_17458,N_12178,N_10027);
xnor U17459 (N_17459,N_12943,N_11737);
and U17460 (N_17460,N_12923,N_12851);
nor U17461 (N_17461,N_14169,N_12922);
or U17462 (N_17462,N_14230,N_10942);
and U17463 (N_17463,N_11000,N_11646);
nand U17464 (N_17464,N_13704,N_12926);
nand U17465 (N_17465,N_11364,N_12670);
and U17466 (N_17466,N_11482,N_10207);
xnor U17467 (N_17467,N_13592,N_12828);
nand U17468 (N_17468,N_10726,N_13796);
nand U17469 (N_17469,N_12785,N_13573);
and U17470 (N_17470,N_10226,N_14768);
xor U17471 (N_17471,N_13856,N_13775);
nand U17472 (N_17472,N_14292,N_14822);
or U17473 (N_17473,N_12891,N_14957);
nor U17474 (N_17474,N_13023,N_11457);
and U17475 (N_17475,N_14859,N_10793);
nand U17476 (N_17476,N_11510,N_13617);
xnor U17477 (N_17477,N_10790,N_13716);
nand U17478 (N_17478,N_12829,N_14926);
and U17479 (N_17479,N_11157,N_14282);
nor U17480 (N_17480,N_10713,N_14414);
nand U17481 (N_17481,N_14071,N_10879);
nor U17482 (N_17482,N_12548,N_11834);
xnor U17483 (N_17483,N_12951,N_11852);
or U17484 (N_17484,N_13806,N_11542);
nand U17485 (N_17485,N_13428,N_11479);
and U17486 (N_17486,N_13621,N_14264);
xor U17487 (N_17487,N_13124,N_10577);
or U17488 (N_17488,N_14892,N_14688);
nand U17489 (N_17489,N_14982,N_12521);
xor U17490 (N_17490,N_12483,N_12478);
nor U17491 (N_17491,N_13632,N_10762);
and U17492 (N_17492,N_10561,N_13010);
xor U17493 (N_17493,N_13888,N_12920);
xor U17494 (N_17494,N_13959,N_10021);
xor U17495 (N_17495,N_11615,N_12650);
and U17496 (N_17496,N_12036,N_10264);
and U17497 (N_17497,N_11826,N_14745);
nand U17498 (N_17498,N_12051,N_10569);
nor U17499 (N_17499,N_14049,N_12140);
and U17500 (N_17500,N_10784,N_14943);
xnor U17501 (N_17501,N_12013,N_13326);
nand U17502 (N_17502,N_14388,N_14346);
xnor U17503 (N_17503,N_11682,N_12931);
and U17504 (N_17504,N_12447,N_10911);
nor U17505 (N_17505,N_11183,N_10644);
or U17506 (N_17506,N_14298,N_12560);
and U17507 (N_17507,N_12033,N_10330);
nand U17508 (N_17508,N_14987,N_13105);
or U17509 (N_17509,N_13522,N_12773);
nand U17510 (N_17510,N_12313,N_11675);
xnor U17511 (N_17511,N_10893,N_12133);
xnor U17512 (N_17512,N_12888,N_12631);
nand U17513 (N_17513,N_10240,N_13596);
xor U17514 (N_17514,N_11953,N_13265);
xor U17515 (N_17515,N_14678,N_14201);
nand U17516 (N_17516,N_10758,N_10129);
or U17517 (N_17517,N_11701,N_13274);
xor U17518 (N_17518,N_10141,N_14470);
xor U17519 (N_17519,N_13907,N_11717);
xor U17520 (N_17520,N_10340,N_11418);
nand U17521 (N_17521,N_12111,N_11086);
xor U17522 (N_17522,N_13797,N_13869);
nand U17523 (N_17523,N_13246,N_10265);
nand U17524 (N_17524,N_11124,N_14560);
xnor U17525 (N_17525,N_11658,N_14960);
xor U17526 (N_17526,N_10831,N_13349);
and U17527 (N_17527,N_12004,N_14404);
xnor U17528 (N_17528,N_14007,N_10585);
or U17529 (N_17529,N_14768,N_11733);
nand U17530 (N_17530,N_13146,N_12351);
nor U17531 (N_17531,N_14928,N_14773);
nor U17532 (N_17532,N_10063,N_11999);
nor U17533 (N_17533,N_14924,N_11186);
nand U17534 (N_17534,N_13462,N_11224);
nor U17535 (N_17535,N_11331,N_13758);
nand U17536 (N_17536,N_14821,N_12754);
xnor U17537 (N_17537,N_10628,N_13557);
and U17538 (N_17538,N_10490,N_10560);
nand U17539 (N_17539,N_14721,N_10900);
or U17540 (N_17540,N_10070,N_10901);
nor U17541 (N_17541,N_13098,N_14368);
or U17542 (N_17542,N_12426,N_13444);
nor U17543 (N_17543,N_13393,N_10631);
or U17544 (N_17544,N_10815,N_13696);
xnor U17545 (N_17545,N_14043,N_13215);
or U17546 (N_17546,N_13673,N_10659);
nand U17547 (N_17547,N_11759,N_11737);
and U17548 (N_17548,N_13314,N_11922);
nand U17549 (N_17549,N_14380,N_11214);
and U17550 (N_17550,N_11219,N_10094);
xor U17551 (N_17551,N_11972,N_12585);
nand U17552 (N_17552,N_10167,N_10364);
nand U17553 (N_17553,N_12382,N_12619);
nor U17554 (N_17554,N_14435,N_11418);
or U17555 (N_17555,N_13960,N_11759);
xor U17556 (N_17556,N_14973,N_10721);
and U17557 (N_17557,N_12285,N_14575);
nand U17558 (N_17558,N_13781,N_13142);
and U17559 (N_17559,N_10642,N_14278);
nor U17560 (N_17560,N_12395,N_12235);
and U17561 (N_17561,N_14857,N_10957);
and U17562 (N_17562,N_12279,N_11449);
or U17563 (N_17563,N_14892,N_13462);
nand U17564 (N_17564,N_11069,N_14187);
nand U17565 (N_17565,N_10852,N_10073);
xor U17566 (N_17566,N_13913,N_14072);
xor U17567 (N_17567,N_11611,N_14780);
xor U17568 (N_17568,N_12769,N_11967);
or U17569 (N_17569,N_11616,N_11126);
nor U17570 (N_17570,N_12077,N_11966);
or U17571 (N_17571,N_14711,N_10086);
xor U17572 (N_17572,N_10009,N_14644);
nand U17573 (N_17573,N_11678,N_13030);
or U17574 (N_17574,N_12960,N_13076);
and U17575 (N_17575,N_10099,N_11326);
and U17576 (N_17576,N_12272,N_11050);
xor U17577 (N_17577,N_12932,N_10292);
or U17578 (N_17578,N_12195,N_14088);
or U17579 (N_17579,N_11856,N_10510);
nand U17580 (N_17580,N_11106,N_12940);
or U17581 (N_17581,N_12927,N_12708);
or U17582 (N_17582,N_11335,N_11326);
or U17583 (N_17583,N_11850,N_11573);
and U17584 (N_17584,N_10521,N_14784);
or U17585 (N_17585,N_11988,N_13128);
nand U17586 (N_17586,N_14887,N_13830);
and U17587 (N_17587,N_11536,N_12790);
xor U17588 (N_17588,N_10769,N_12859);
nor U17589 (N_17589,N_12975,N_14033);
nand U17590 (N_17590,N_13213,N_12063);
xnor U17591 (N_17591,N_11111,N_10842);
and U17592 (N_17592,N_14527,N_12900);
xnor U17593 (N_17593,N_12377,N_12985);
nor U17594 (N_17594,N_14767,N_11127);
xnor U17595 (N_17595,N_14434,N_10310);
nor U17596 (N_17596,N_11038,N_10257);
and U17597 (N_17597,N_13739,N_14895);
nor U17598 (N_17598,N_11087,N_11399);
or U17599 (N_17599,N_10928,N_14108);
and U17600 (N_17600,N_11869,N_10916);
nor U17601 (N_17601,N_10019,N_12734);
nor U17602 (N_17602,N_13185,N_12429);
or U17603 (N_17603,N_11836,N_11572);
nor U17604 (N_17604,N_12381,N_10319);
xor U17605 (N_17605,N_12783,N_14323);
or U17606 (N_17606,N_13071,N_11209);
nor U17607 (N_17607,N_13507,N_11932);
and U17608 (N_17608,N_11900,N_12265);
or U17609 (N_17609,N_12136,N_10482);
nor U17610 (N_17610,N_13002,N_11261);
xor U17611 (N_17611,N_13414,N_10760);
nor U17612 (N_17612,N_10699,N_11720);
or U17613 (N_17613,N_14609,N_12073);
and U17614 (N_17614,N_12449,N_10790);
xnor U17615 (N_17615,N_14653,N_14278);
and U17616 (N_17616,N_10212,N_12166);
xnor U17617 (N_17617,N_13681,N_10998);
xor U17618 (N_17618,N_13562,N_13268);
and U17619 (N_17619,N_13626,N_14634);
xor U17620 (N_17620,N_13857,N_10875);
or U17621 (N_17621,N_13464,N_12936);
nor U17622 (N_17622,N_14805,N_13098);
and U17623 (N_17623,N_13149,N_13131);
xnor U17624 (N_17624,N_14000,N_10794);
or U17625 (N_17625,N_10562,N_14736);
nand U17626 (N_17626,N_12584,N_12975);
xor U17627 (N_17627,N_10757,N_11706);
xor U17628 (N_17628,N_10911,N_13993);
xnor U17629 (N_17629,N_14376,N_12616);
or U17630 (N_17630,N_14535,N_11854);
nor U17631 (N_17631,N_12877,N_12976);
or U17632 (N_17632,N_12641,N_12940);
nand U17633 (N_17633,N_14726,N_14284);
or U17634 (N_17634,N_14945,N_11624);
nor U17635 (N_17635,N_13285,N_10052);
nand U17636 (N_17636,N_14766,N_11990);
and U17637 (N_17637,N_10360,N_13006);
xnor U17638 (N_17638,N_13550,N_14409);
or U17639 (N_17639,N_13867,N_14563);
and U17640 (N_17640,N_13560,N_10382);
or U17641 (N_17641,N_10527,N_14714);
xor U17642 (N_17642,N_14673,N_13636);
nor U17643 (N_17643,N_11253,N_11685);
and U17644 (N_17644,N_14514,N_14774);
or U17645 (N_17645,N_12069,N_13597);
and U17646 (N_17646,N_11474,N_10467);
nor U17647 (N_17647,N_14279,N_10474);
xnor U17648 (N_17648,N_13353,N_14630);
and U17649 (N_17649,N_10102,N_13847);
nor U17650 (N_17650,N_12828,N_12193);
nor U17651 (N_17651,N_13717,N_14365);
and U17652 (N_17652,N_14093,N_14371);
and U17653 (N_17653,N_11937,N_13767);
nand U17654 (N_17654,N_14292,N_12719);
nor U17655 (N_17655,N_11737,N_10314);
xor U17656 (N_17656,N_13821,N_12804);
xnor U17657 (N_17657,N_13428,N_11553);
nor U17658 (N_17658,N_11025,N_13001);
or U17659 (N_17659,N_12342,N_12515);
and U17660 (N_17660,N_12238,N_14682);
xnor U17661 (N_17661,N_13924,N_11895);
nand U17662 (N_17662,N_10214,N_11871);
nand U17663 (N_17663,N_11632,N_10385);
or U17664 (N_17664,N_13841,N_14407);
nand U17665 (N_17665,N_10382,N_10306);
and U17666 (N_17666,N_14837,N_12361);
nand U17667 (N_17667,N_14975,N_12037);
or U17668 (N_17668,N_12254,N_12090);
or U17669 (N_17669,N_11116,N_14697);
or U17670 (N_17670,N_14133,N_13555);
xor U17671 (N_17671,N_10371,N_14840);
and U17672 (N_17672,N_11142,N_11207);
xor U17673 (N_17673,N_10788,N_14391);
and U17674 (N_17674,N_12394,N_10885);
nand U17675 (N_17675,N_11783,N_13354);
and U17676 (N_17676,N_12263,N_10942);
nand U17677 (N_17677,N_10791,N_11358);
nand U17678 (N_17678,N_14924,N_13592);
or U17679 (N_17679,N_10057,N_12940);
xor U17680 (N_17680,N_11064,N_12879);
nand U17681 (N_17681,N_12000,N_13581);
and U17682 (N_17682,N_14068,N_13725);
nor U17683 (N_17683,N_12321,N_11966);
nand U17684 (N_17684,N_12857,N_11450);
and U17685 (N_17685,N_11800,N_10257);
nor U17686 (N_17686,N_10972,N_11288);
xor U17687 (N_17687,N_11756,N_14107);
or U17688 (N_17688,N_13542,N_13952);
nand U17689 (N_17689,N_13821,N_13493);
and U17690 (N_17690,N_11448,N_11939);
nor U17691 (N_17691,N_14785,N_10004);
nor U17692 (N_17692,N_12797,N_12241);
nand U17693 (N_17693,N_12811,N_14465);
xnor U17694 (N_17694,N_13679,N_10388);
xor U17695 (N_17695,N_11698,N_11693);
xnor U17696 (N_17696,N_10158,N_12839);
nand U17697 (N_17697,N_13592,N_13408);
nand U17698 (N_17698,N_14151,N_12340);
nand U17699 (N_17699,N_11749,N_13665);
xor U17700 (N_17700,N_14129,N_13055);
nor U17701 (N_17701,N_14032,N_13100);
nor U17702 (N_17702,N_11371,N_12302);
and U17703 (N_17703,N_12623,N_14643);
or U17704 (N_17704,N_11371,N_13995);
and U17705 (N_17705,N_10708,N_12636);
and U17706 (N_17706,N_12685,N_11019);
and U17707 (N_17707,N_10545,N_13029);
xor U17708 (N_17708,N_14792,N_14091);
xnor U17709 (N_17709,N_10241,N_10508);
nand U17710 (N_17710,N_14345,N_13429);
xor U17711 (N_17711,N_11730,N_12512);
xnor U17712 (N_17712,N_10468,N_14066);
or U17713 (N_17713,N_14878,N_10829);
nand U17714 (N_17714,N_10576,N_10948);
nand U17715 (N_17715,N_12510,N_12201);
xor U17716 (N_17716,N_12779,N_12652);
nor U17717 (N_17717,N_14796,N_14364);
nor U17718 (N_17718,N_12986,N_12166);
and U17719 (N_17719,N_13836,N_10195);
nand U17720 (N_17720,N_14816,N_11270);
or U17721 (N_17721,N_14370,N_13933);
or U17722 (N_17722,N_12457,N_14186);
and U17723 (N_17723,N_12313,N_13903);
or U17724 (N_17724,N_11388,N_12156);
or U17725 (N_17725,N_10628,N_11551);
or U17726 (N_17726,N_10414,N_14782);
and U17727 (N_17727,N_13001,N_10340);
xor U17728 (N_17728,N_10281,N_10928);
and U17729 (N_17729,N_10835,N_14193);
or U17730 (N_17730,N_12003,N_12915);
or U17731 (N_17731,N_11612,N_12426);
nand U17732 (N_17732,N_10706,N_10278);
or U17733 (N_17733,N_10364,N_12662);
nand U17734 (N_17734,N_11917,N_12982);
or U17735 (N_17735,N_12989,N_11106);
and U17736 (N_17736,N_11531,N_14040);
and U17737 (N_17737,N_14552,N_14078);
nor U17738 (N_17738,N_12107,N_11930);
nand U17739 (N_17739,N_12508,N_14029);
and U17740 (N_17740,N_10612,N_10054);
xor U17741 (N_17741,N_14139,N_13424);
nor U17742 (N_17742,N_12033,N_10555);
nand U17743 (N_17743,N_10304,N_14468);
nor U17744 (N_17744,N_12374,N_13102);
xnor U17745 (N_17745,N_10364,N_10362);
and U17746 (N_17746,N_10844,N_13016);
xor U17747 (N_17747,N_12669,N_13717);
nand U17748 (N_17748,N_10792,N_13368);
xor U17749 (N_17749,N_14590,N_10558);
or U17750 (N_17750,N_10741,N_11038);
xor U17751 (N_17751,N_10836,N_13714);
nor U17752 (N_17752,N_12949,N_13010);
and U17753 (N_17753,N_12874,N_14674);
nand U17754 (N_17754,N_11470,N_13255);
nand U17755 (N_17755,N_13732,N_11471);
or U17756 (N_17756,N_14865,N_13839);
nand U17757 (N_17757,N_14956,N_10993);
nor U17758 (N_17758,N_12495,N_13928);
nor U17759 (N_17759,N_12722,N_11056);
and U17760 (N_17760,N_13463,N_11301);
nor U17761 (N_17761,N_13131,N_10309);
nand U17762 (N_17762,N_10957,N_11972);
nand U17763 (N_17763,N_12869,N_11269);
xnor U17764 (N_17764,N_11463,N_14916);
and U17765 (N_17765,N_13172,N_13343);
xnor U17766 (N_17766,N_13883,N_13251);
xor U17767 (N_17767,N_11441,N_12197);
nand U17768 (N_17768,N_13478,N_14743);
and U17769 (N_17769,N_14198,N_14520);
or U17770 (N_17770,N_11473,N_13739);
or U17771 (N_17771,N_11140,N_11516);
nor U17772 (N_17772,N_11833,N_12075);
nand U17773 (N_17773,N_11511,N_13308);
nand U17774 (N_17774,N_10727,N_10692);
and U17775 (N_17775,N_12663,N_14647);
nor U17776 (N_17776,N_10550,N_14712);
nand U17777 (N_17777,N_12978,N_11876);
xor U17778 (N_17778,N_12976,N_10811);
nor U17779 (N_17779,N_13313,N_13457);
nor U17780 (N_17780,N_14482,N_10367);
nor U17781 (N_17781,N_10745,N_12585);
or U17782 (N_17782,N_11244,N_12511);
nand U17783 (N_17783,N_10407,N_13901);
or U17784 (N_17784,N_14294,N_14743);
nor U17785 (N_17785,N_11910,N_12472);
or U17786 (N_17786,N_14264,N_12801);
xnor U17787 (N_17787,N_12768,N_13777);
or U17788 (N_17788,N_12930,N_12996);
nor U17789 (N_17789,N_10259,N_14146);
or U17790 (N_17790,N_13085,N_10805);
nand U17791 (N_17791,N_13394,N_12967);
or U17792 (N_17792,N_14531,N_13719);
and U17793 (N_17793,N_13382,N_11590);
xnor U17794 (N_17794,N_10296,N_12668);
nand U17795 (N_17795,N_11741,N_12524);
xnor U17796 (N_17796,N_12498,N_11022);
nand U17797 (N_17797,N_11831,N_13308);
or U17798 (N_17798,N_12832,N_13645);
xnor U17799 (N_17799,N_10840,N_11885);
xnor U17800 (N_17800,N_11498,N_11451);
or U17801 (N_17801,N_10946,N_12776);
xnor U17802 (N_17802,N_12874,N_13404);
nand U17803 (N_17803,N_11151,N_13677);
and U17804 (N_17804,N_10427,N_10152);
nand U17805 (N_17805,N_14718,N_10511);
or U17806 (N_17806,N_13775,N_13091);
nand U17807 (N_17807,N_12361,N_12963);
nand U17808 (N_17808,N_12613,N_14137);
nand U17809 (N_17809,N_14070,N_10330);
xor U17810 (N_17810,N_10491,N_10838);
nand U17811 (N_17811,N_13637,N_13749);
xnor U17812 (N_17812,N_11466,N_10925);
and U17813 (N_17813,N_14282,N_13737);
or U17814 (N_17814,N_12223,N_14746);
nor U17815 (N_17815,N_13471,N_10619);
and U17816 (N_17816,N_13209,N_14409);
and U17817 (N_17817,N_14488,N_10896);
or U17818 (N_17818,N_10854,N_13207);
xnor U17819 (N_17819,N_13215,N_14178);
and U17820 (N_17820,N_12640,N_11412);
nand U17821 (N_17821,N_11758,N_11823);
xnor U17822 (N_17822,N_12417,N_14696);
xnor U17823 (N_17823,N_13039,N_14394);
or U17824 (N_17824,N_14133,N_11737);
nor U17825 (N_17825,N_10171,N_10705);
and U17826 (N_17826,N_13682,N_14640);
xnor U17827 (N_17827,N_14427,N_10059);
nor U17828 (N_17828,N_12898,N_11351);
and U17829 (N_17829,N_14114,N_12591);
nor U17830 (N_17830,N_10021,N_12783);
nor U17831 (N_17831,N_12123,N_14835);
and U17832 (N_17832,N_12064,N_14629);
xnor U17833 (N_17833,N_13551,N_10980);
and U17834 (N_17834,N_14815,N_13923);
and U17835 (N_17835,N_14900,N_12781);
nand U17836 (N_17836,N_12473,N_14113);
xnor U17837 (N_17837,N_10977,N_12840);
nor U17838 (N_17838,N_11311,N_12694);
and U17839 (N_17839,N_11749,N_10653);
and U17840 (N_17840,N_12592,N_10338);
or U17841 (N_17841,N_12948,N_14702);
xnor U17842 (N_17842,N_12976,N_13688);
nand U17843 (N_17843,N_13220,N_14853);
xnor U17844 (N_17844,N_11194,N_13478);
or U17845 (N_17845,N_11327,N_13539);
xnor U17846 (N_17846,N_10133,N_14402);
or U17847 (N_17847,N_10979,N_10498);
xor U17848 (N_17848,N_13754,N_11936);
nand U17849 (N_17849,N_11444,N_13876);
nor U17850 (N_17850,N_13738,N_13775);
nor U17851 (N_17851,N_13593,N_13936);
nor U17852 (N_17852,N_10199,N_14101);
and U17853 (N_17853,N_14625,N_11945);
or U17854 (N_17854,N_13018,N_12176);
xor U17855 (N_17855,N_13515,N_13966);
and U17856 (N_17856,N_14531,N_14468);
or U17857 (N_17857,N_10387,N_13839);
nor U17858 (N_17858,N_12444,N_12779);
nand U17859 (N_17859,N_12563,N_11154);
and U17860 (N_17860,N_11683,N_10097);
or U17861 (N_17861,N_13630,N_14775);
or U17862 (N_17862,N_11774,N_13399);
nor U17863 (N_17863,N_10638,N_11615);
nor U17864 (N_17864,N_11546,N_13711);
or U17865 (N_17865,N_13487,N_11957);
and U17866 (N_17866,N_10501,N_11829);
or U17867 (N_17867,N_10044,N_14881);
nand U17868 (N_17868,N_14462,N_10235);
or U17869 (N_17869,N_10702,N_12565);
or U17870 (N_17870,N_11587,N_14412);
or U17871 (N_17871,N_13567,N_10869);
nand U17872 (N_17872,N_10309,N_13975);
nand U17873 (N_17873,N_11539,N_14719);
nand U17874 (N_17874,N_14975,N_12336);
or U17875 (N_17875,N_13625,N_13352);
nor U17876 (N_17876,N_11944,N_11248);
nand U17877 (N_17877,N_14249,N_11928);
nand U17878 (N_17878,N_11389,N_13230);
and U17879 (N_17879,N_12238,N_13338);
nor U17880 (N_17880,N_10381,N_12792);
xnor U17881 (N_17881,N_11055,N_12381);
nand U17882 (N_17882,N_14174,N_12269);
nand U17883 (N_17883,N_14446,N_10502);
and U17884 (N_17884,N_11657,N_13786);
nor U17885 (N_17885,N_11726,N_10153);
or U17886 (N_17886,N_13478,N_14486);
and U17887 (N_17887,N_13328,N_13718);
nor U17888 (N_17888,N_12611,N_11368);
or U17889 (N_17889,N_13976,N_10782);
and U17890 (N_17890,N_11422,N_12940);
xor U17891 (N_17891,N_14457,N_10854);
or U17892 (N_17892,N_10262,N_13797);
or U17893 (N_17893,N_13710,N_14514);
and U17894 (N_17894,N_14437,N_11119);
and U17895 (N_17895,N_12823,N_12509);
nor U17896 (N_17896,N_13558,N_10703);
nand U17897 (N_17897,N_12916,N_14339);
nor U17898 (N_17898,N_10110,N_14567);
xor U17899 (N_17899,N_13501,N_13807);
or U17900 (N_17900,N_10419,N_13526);
xor U17901 (N_17901,N_12364,N_10574);
nor U17902 (N_17902,N_10744,N_14756);
or U17903 (N_17903,N_11729,N_13609);
or U17904 (N_17904,N_12153,N_11394);
nand U17905 (N_17905,N_10976,N_10177);
xnor U17906 (N_17906,N_10674,N_13147);
and U17907 (N_17907,N_14119,N_10088);
or U17908 (N_17908,N_11384,N_10442);
nand U17909 (N_17909,N_14103,N_12730);
nand U17910 (N_17910,N_13526,N_13097);
and U17911 (N_17911,N_10026,N_12880);
xnor U17912 (N_17912,N_12341,N_10028);
and U17913 (N_17913,N_10367,N_11325);
and U17914 (N_17914,N_12625,N_10316);
nand U17915 (N_17915,N_10094,N_13834);
xnor U17916 (N_17916,N_11795,N_11281);
nand U17917 (N_17917,N_13761,N_13110);
and U17918 (N_17918,N_13391,N_14519);
nand U17919 (N_17919,N_10410,N_14750);
and U17920 (N_17920,N_13693,N_13420);
nor U17921 (N_17921,N_14437,N_12078);
nand U17922 (N_17922,N_11828,N_14548);
and U17923 (N_17923,N_11234,N_11644);
xnor U17924 (N_17924,N_10321,N_14706);
nand U17925 (N_17925,N_13490,N_11194);
xor U17926 (N_17926,N_14770,N_10773);
nand U17927 (N_17927,N_10619,N_12485);
nand U17928 (N_17928,N_13623,N_12263);
xor U17929 (N_17929,N_12008,N_13114);
or U17930 (N_17930,N_10321,N_13980);
nand U17931 (N_17931,N_11055,N_10510);
nor U17932 (N_17932,N_13201,N_11285);
nand U17933 (N_17933,N_14657,N_10964);
nor U17934 (N_17934,N_10073,N_12846);
or U17935 (N_17935,N_10647,N_14873);
nor U17936 (N_17936,N_12142,N_14291);
and U17937 (N_17937,N_13594,N_10466);
and U17938 (N_17938,N_13602,N_12401);
xor U17939 (N_17939,N_11924,N_14860);
and U17940 (N_17940,N_13553,N_10296);
xnor U17941 (N_17941,N_13078,N_12039);
nor U17942 (N_17942,N_14320,N_10482);
nor U17943 (N_17943,N_11704,N_13713);
nand U17944 (N_17944,N_11827,N_11539);
and U17945 (N_17945,N_13325,N_10382);
and U17946 (N_17946,N_10285,N_13027);
and U17947 (N_17947,N_12845,N_12916);
or U17948 (N_17948,N_12154,N_13372);
nor U17949 (N_17949,N_10603,N_11034);
nor U17950 (N_17950,N_12298,N_14761);
and U17951 (N_17951,N_10501,N_13435);
xor U17952 (N_17952,N_13792,N_13645);
or U17953 (N_17953,N_12718,N_13341);
xnor U17954 (N_17954,N_11101,N_11334);
and U17955 (N_17955,N_14879,N_12907);
or U17956 (N_17956,N_12601,N_10311);
and U17957 (N_17957,N_13579,N_11219);
nor U17958 (N_17958,N_11010,N_14403);
nor U17959 (N_17959,N_10678,N_12972);
nor U17960 (N_17960,N_13740,N_11813);
and U17961 (N_17961,N_10584,N_14192);
xnor U17962 (N_17962,N_12170,N_14011);
nand U17963 (N_17963,N_14272,N_10680);
nand U17964 (N_17964,N_14578,N_10312);
and U17965 (N_17965,N_11856,N_14550);
and U17966 (N_17966,N_12339,N_13865);
or U17967 (N_17967,N_13778,N_11511);
nand U17968 (N_17968,N_12127,N_10739);
xnor U17969 (N_17969,N_12363,N_13730);
nor U17970 (N_17970,N_10539,N_11811);
nor U17971 (N_17971,N_13655,N_13300);
xor U17972 (N_17972,N_13957,N_13568);
and U17973 (N_17973,N_10055,N_14273);
nor U17974 (N_17974,N_10171,N_10473);
or U17975 (N_17975,N_14132,N_12499);
nand U17976 (N_17976,N_12201,N_13695);
nor U17977 (N_17977,N_11147,N_12659);
and U17978 (N_17978,N_10297,N_12777);
nor U17979 (N_17979,N_13690,N_12435);
nor U17980 (N_17980,N_13370,N_10939);
nor U17981 (N_17981,N_14777,N_14311);
xnor U17982 (N_17982,N_11092,N_11823);
nor U17983 (N_17983,N_13618,N_14314);
xor U17984 (N_17984,N_10252,N_12948);
xnor U17985 (N_17985,N_11133,N_10070);
and U17986 (N_17986,N_12634,N_14362);
or U17987 (N_17987,N_11651,N_10176);
and U17988 (N_17988,N_13980,N_12032);
nand U17989 (N_17989,N_13287,N_14441);
and U17990 (N_17990,N_12923,N_14797);
nand U17991 (N_17991,N_12425,N_14689);
xor U17992 (N_17992,N_12081,N_14018);
nor U17993 (N_17993,N_12219,N_11053);
nor U17994 (N_17994,N_12153,N_11560);
nand U17995 (N_17995,N_10579,N_12088);
xnor U17996 (N_17996,N_13840,N_12721);
or U17997 (N_17997,N_10154,N_10199);
nor U17998 (N_17998,N_13653,N_11540);
nand U17999 (N_17999,N_10645,N_14702);
xnor U18000 (N_18000,N_10705,N_11015);
nand U18001 (N_18001,N_10048,N_12926);
and U18002 (N_18002,N_11188,N_10675);
xnor U18003 (N_18003,N_12558,N_14645);
xnor U18004 (N_18004,N_11529,N_11595);
xnor U18005 (N_18005,N_13969,N_10703);
and U18006 (N_18006,N_14672,N_12322);
or U18007 (N_18007,N_10029,N_10503);
or U18008 (N_18008,N_10034,N_12788);
and U18009 (N_18009,N_11278,N_14458);
or U18010 (N_18010,N_13211,N_11146);
or U18011 (N_18011,N_12618,N_13836);
nand U18012 (N_18012,N_13483,N_11115);
xnor U18013 (N_18013,N_12700,N_11741);
and U18014 (N_18014,N_13241,N_10660);
or U18015 (N_18015,N_10309,N_13196);
nand U18016 (N_18016,N_11531,N_11412);
xor U18017 (N_18017,N_12779,N_14790);
nand U18018 (N_18018,N_12152,N_11598);
and U18019 (N_18019,N_13065,N_14028);
and U18020 (N_18020,N_10994,N_11737);
nand U18021 (N_18021,N_10541,N_13988);
or U18022 (N_18022,N_14066,N_13101);
or U18023 (N_18023,N_12472,N_13701);
xor U18024 (N_18024,N_10118,N_12637);
xor U18025 (N_18025,N_11072,N_12812);
nand U18026 (N_18026,N_12150,N_14298);
or U18027 (N_18027,N_11289,N_12748);
nand U18028 (N_18028,N_12636,N_13550);
or U18029 (N_18029,N_10219,N_12277);
and U18030 (N_18030,N_11390,N_13682);
nand U18031 (N_18031,N_13262,N_13027);
nor U18032 (N_18032,N_10226,N_11720);
xnor U18033 (N_18033,N_11797,N_12465);
xnor U18034 (N_18034,N_12699,N_10299);
and U18035 (N_18035,N_14275,N_12427);
or U18036 (N_18036,N_12862,N_13908);
and U18037 (N_18037,N_14559,N_14459);
nor U18038 (N_18038,N_14139,N_13945);
xnor U18039 (N_18039,N_10145,N_12706);
nor U18040 (N_18040,N_13673,N_14410);
nand U18041 (N_18041,N_14353,N_14692);
xor U18042 (N_18042,N_14196,N_12471);
or U18043 (N_18043,N_13158,N_12861);
or U18044 (N_18044,N_14356,N_14594);
nor U18045 (N_18045,N_10113,N_12700);
or U18046 (N_18046,N_11627,N_12512);
nand U18047 (N_18047,N_14426,N_11013);
nand U18048 (N_18048,N_12687,N_14969);
nor U18049 (N_18049,N_13996,N_10612);
xor U18050 (N_18050,N_11278,N_10522);
nor U18051 (N_18051,N_14889,N_11348);
or U18052 (N_18052,N_10429,N_12755);
nand U18053 (N_18053,N_11598,N_10764);
nor U18054 (N_18054,N_13839,N_13757);
xnor U18055 (N_18055,N_13368,N_14501);
xor U18056 (N_18056,N_14889,N_14355);
or U18057 (N_18057,N_11214,N_11141);
and U18058 (N_18058,N_10729,N_11593);
nand U18059 (N_18059,N_13128,N_14640);
xnor U18060 (N_18060,N_11472,N_11217);
nand U18061 (N_18061,N_12175,N_10683);
nand U18062 (N_18062,N_13257,N_13671);
nor U18063 (N_18063,N_14937,N_10108);
nor U18064 (N_18064,N_13223,N_10770);
xor U18065 (N_18065,N_14204,N_10252);
and U18066 (N_18066,N_13819,N_14338);
xor U18067 (N_18067,N_11341,N_10839);
xor U18068 (N_18068,N_12495,N_11746);
nor U18069 (N_18069,N_11871,N_14443);
and U18070 (N_18070,N_13745,N_11773);
or U18071 (N_18071,N_11987,N_11281);
nand U18072 (N_18072,N_12342,N_10897);
nand U18073 (N_18073,N_13055,N_10940);
nand U18074 (N_18074,N_12412,N_13348);
or U18075 (N_18075,N_13753,N_11898);
nand U18076 (N_18076,N_12270,N_14758);
or U18077 (N_18077,N_11968,N_11398);
nand U18078 (N_18078,N_12740,N_11883);
and U18079 (N_18079,N_13069,N_11428);
and U18080 (N_18080,N_14280,N_10357);
and U18081 (N_18081,N_11711,N_12279);
and U18082 (N_18082,N_10946,N_10133);
xnor U18083 (N_18083,N_13447,N_10218);
nand U18084 (N_18084,N_10721,N_12122);
or U18085 (N_18085,N_11681,N_12300);
and U18086 (N_18086,N_11684,N_10914);
nor U18087 (N_18087,N_14223,N_14270);
nand U18088 (N_18088,N_12596,N_11581);
and U18089 (N_18089,N_10965,N_10759);
xor U18090 (N_18090,N_10498,N_12387);
xnor U18091 (N_18091,N_13686,N_12720);
and U18092 (N_18092,N_10571,N_13712);
nand U18093 (N_18093,N_14033,N_10859);
xnor U18094 (N_18094,N_11635,N_10765);
xor U18095 (N_18095,N_10505,N_11667);
nor U18096 (N_18096,N_12057,N_12506);
xor U18097 (N_18097,N_14889,N_14201);
and U18098 (N_18098,N_10229,N_11698);
xnor U18099 (N_18099,N_11691,N_11509);
and U18100 (N_18100,N_14593,N_13036);
nor U18101 (N_18101,N_13881,N_11571);
or U18102 (N_18102,N_14609,N_14312);
xnor U18103 (N_18103,N_14080,N_11312);
and U18104 (N_18104,N_13271,N_13065);
nand U18105 (N_18105,N_10181,N_13966);
or U18106 (N_18106,N_13603,N_14810);
xor U18107 (N_18107,N_14894,N_10292);
and U18108 (N_18108,N_11100,N_14479);
nor U18109 (N_18109,N_13935,N_10250);
nor U18110 (N_18110,N_14023,N_14282);
xor U18111 (N_18111,N_13251,N_13716);
or U18112 (N_18112,N_10484,N_10490);
xor U18113 (N_18113,N_13077,N_12556);
xnor U18114 (N_18114,N_14032,N_13298);
xor U18115 (N_18115,N_10112,N_14282);
and U18116 (N_18116,N_11293,N_12561);
nor U18117 (N_18117,N_12470,N_12223);
nor U18118 (N_18118,N_10032,N_11653);
or U18119 (N_18119,N_10410,N_10933);
and U18120 (N_18120,N_12835,N_14800);
xnor U18121 (N_18121,N_14263,N_13774);
nor U18122 (N_18122,N_12214,N_13717);
xor U18123 (N_18123,N_10608,N_13974);
or U18124 (N_18124,N_12671,N_13711);
nor U18125 (N_18125,N_13195,N_12542);
xor U18126 (N_18126,N_14176,N_14202);
and U18127 (N_18127,N_14186,N_13757);
nor U18128 (N_18128,N_13096,N_12568);
nor U18129 (N_18129,N_11935,N_14292);
nand U18130 (N_18130,N_13359,N_13430);
and U18131 (N_18131,N_14323,N_11088);
and U18132 (N_18132,N_10629,N_13591);
xnor U18133 (N_18133,N_12072,N_11938);
and U18134 (N_18134,N_12934,N_14824);
nor U18135 (N_18135,N_10077,N_11866);
nand U18136 (N_18136,N_10688,N_12709);
and U18137 (N_18137,N_10800,N_13416);
or U18138 (N_18138,N_11870,N_13212);
xor U18139 (N_18139,N_12600,N_10785);
nor U18140 (N_18140,N_14473,N_10020);
nor U18141 (N_18141,N_13574,N_11037);
nor U18142 (N_18142,N_14271,N_13521);
nor U18143 (N_18143,N_11857,N_13083);
xor U18144 (N_18144,N_10895,N_14530);
nand U18145 (N_18145,N_14883,N_10631);
or U18146 (N_18146,N_12609,N_10347);
or U18147 (N_18147,N_14391,N_11110);
nor U18148 (N_18148,N_12377,N_13727);
nand U18149 (N_18149,N_14244,N_12685);
xnor U18150 (N_18150,N_11931,N_11364);
xnor U18151 (N_18151,N_13617,N_11253);
nor U18152 (N_18152,N_11369,N_10532);
nor U18153 (N_18153,N_12633,N_13235);
and U18154 (N_18154,N_10853,N_11471);
and U18155 (N_18155,N_13497,N_12535);
and U18156 (N_18156,N_10804,N_11773);
and U18157 (N_18157,N_14128,N_14459);
and U18158 (N_18158,N_11058,N_11673);
nor U18159 (N_18159,N_12168,N_10399);
or U18160 (N_18160,N_10644,N_13102);
nor U18161 (N_18161,N_10545,N_12971);
or U18162 (N_18162,N_12608,N_10354);
or U18163 (N_18163,N_12330,N_14248);
nor U18164 (N_18164,N_11729,N_12934);
or U18165 (N_18165,N_12626,N_10919);
and U18166 (N_18166,N_10561,N_14126);
or U18167 (N_18167,N_13531,N_10177);
xor U18168 (N_18168,N_12412,N_11220);
or U18169 (N_18169,N_10918,N_13665);
nand U18170 (N_18170,N_10556,N_10124);
and U18171 (N_18171,N_12966,N_10409);
and U18172 (N_18172,N_12255,N_10218);
nand U18173 (N_18173,N_10877,N_14515);
nor U18174 (N_18174,N_11925,N_12906);
nor U18175 (N_18175,N_14948,N_12957);
and U18176 (N_18176,N_13774,N_14284);
or U18177 (N_18177,N_14277,N_14214);
xor U18178 (N_18178,N_10835,N_10760);
xor U18179 (N_18179,N_10577,N_11654);
nand U18180 (N_18180,N_12244,N_10360);
nand U18181 (N_18181,N_11874,N_12708);
xnor U18182 (N_18182,N_14357,N_14781);
or U18183 (N_18183,N_13408,N_12137);
or U18184 (N_18184,N_14114,N_14409);
xnor U18185 (N_18185,N_12262,N_11270);
nand U18186 (N_18186,N_13113,N_13963);
xnor U18187 (N_18187,N_12093,N_13348);
nor U18188 (N_18188,N_10154,N_14249);
or U18189 (N_18189,N_10811,N_10963);
xnor U18190 (N_18190,N_10397,N_10941);
nand U18191 (N_18191,N_13884,N_11522);
xor U18192 (N_18192,N_11727,N_11415);
nor U18193 (N_18193,N_10317,N_11477);
or U18194 (N_18194,N_10509,N_11829);
xor U18195 (N_18195,N_11472,N_11581);
and U18196 (N_18196,N_11490,N_10575);
nand U18197 (N_18197,N_12605,N_10762);
and U18198 (N_18198,N_10738,N_12367);
and U18199 (N_18199,N_13925,N_12500);
xor U18200 (N_18200,N_14548,N_14049);
or U18201 (N_18201,N_13584,N_12562);
and U18202 (N_18202,N_13298,N_10544);
or U18203 (N_18203,N_14916,N_12211);
nor U18204 (N_18204,N_13976,N_11569);
nor U18205 (N_18205,N_12982,N_11019);
xnor U18206 (N_18206,N_12610,N_12202);
xnor U18207 (N_18207,N_14683,N_14389);
nand U18208 (N_18208,N_11447,N_14885);
nor U18209 (N_18209,N_11791,N_12748);
nand U18210 (N_18210,N_11402,N_13069);
nor U18211 (N_18211,N_13059,N_14915);
and U18212 (N_18212,N_14839,N_13668);
or U18213 (N_18213,N_10196,N_14076);
or U18214 (N_18214,N_13556,N_11386);
nand U18215 (N_18215,N_10206,N_10650);
xnor U18216 (N_18216,N_13797,N_12003);
nand U18217 (N_18217,N_14883,N_13834);
nor U18218 (N_18218,N_12751,N_12993);
xnor U18219 (N_18219,N_13220,N_12322);
nor U18220 (N_18220,N_13090,N_12964);
nor U18221 (N_18221,N_11258,N_13578);
nor U18222 (N_18222,N_12976,N_11127);
and U18223 (N_18223,N_13054,N_10671);
xor U18224 (N_18224,N_11002,N_13829);
xnor U18225 (N_18225,N_13502,N_12255);
nor U18226 (N_18226,N_12963,N_14715);
xor U18227 (N_18227,N_12914,N_11549);
nand U18228 (N_18228,N_12321,N_10066);
nor U18229 (N_18229,N_11074,N_11623);
nor U18230 (N_18230,N_11158,N_14783);
or U18231 (N_18231,N_14930,N_12125);
and U18232 (N_18232,N_13268,N_11712);
or U18233 (N_18233,N_10442,N_10347);
and U18234 (N_18234,N_12631,N_13894);
and U18235 (N_18235,N_14400,N_12290);
xor U18236 (N_18236,N_10363,N_12823);
nor U18237 (N_18237,N_10086,N_12828);
and U18238 (N_18238,N_13184,N_13711);
xor U18239 (N_18239,N_12277,N_11147);
nand U18240 (N_18240,N_11579,N_11640);
xnor U18241 (N_18241,N_10002,N_13330);
nand U18242 (N_18242,N_11762,N_11301);
and U18243 (N_18243,N_12673,N_12179);
and U18244 (N_18244,N_14312,N_14978);
xor U18245 (N_18245,N_12420,N_13909);
xnor U18246 (N_18246,N_10168,N_14630);
or U18247 (N_18247,N_13004,N_10399);
nand U18248 (N_18248,N_12152,N_13654);
nor U18249 (N_18249,N_13827,N_10146);
and U18250 (N_18250,N_11273,N_14058);
or U18251 (N_18251,N_14017,N_12312);
nor U18252 (N_18252,N_14516,N_11523);
nand U18253 (N_18253,N_13008,N_10674);
nor U18254 (N_18254,N_10238,N_11525);
xor U18255 (N_18255,N_12951,N_10378);
and U18256 (N_18256,N_12634,N_10288);
xor U18257 (N_18257,N_12818,N_10022);
and U18258 (N_18258,N_11017,N_14976);
or U18259 (N_18259,N_11285,N_13151);
and U18260 (N_18260,N_11585,N_12161);
or U18261 (N_18261,N_12570,N_12878);
nor U18262 (N_18262,N_14430,N_10082);
nor U18263 (N_18263,N_13984,N_11098);
nor U18264 (N_18264,N_13309,N_12268);
or U18265 (N_18265,N_12946,N_11574);
and U18266 (N_18266,N_14454,N_10582);
xor U18267 (N_18267,N_14042,N_14889);
xor U18268 (N_18268,N_10068,N_11987);
or U18269 (N_18269,N_14558,N_14053);
nand U18270 (N_18270,N_14032,N_13290);
and U18271 (N_18271,N_13311,N_11183);
nor U18272 (N_18272,N_10338,N_14098);
xor U18273 (N_18273,N_11918,N_11129);
nor U18274 (N_18274,N_14567,N_14969);
or U18275 (N_18275,N_12364,N_13143);
nor U18276 (N_18276,N_14129,N_10138);
or U18277 (N_18277,N_11335,N_11725);
nor U18278 (N_18278,N_12953,N_10996);
or U18279 (N_18279,N_12608,N_12496);
xnor U18280 (N_18280,N_13123,N_10822);
nor U18281 (N_18281,N_10944,N_13871);
nand U18282 (N_18282,N_11170,N_10782);
and U18283 (N_18283,N_12558,N_12317);
nand U18284 (N_18284,N_13843,N_11334);
nor U18285 (N_18285,N_10434,N_10847);
and U18286 (N_18286,N_14386,N_10911);
or U18287 (N_18287,N_10088,N_11562);
nand U18288 (N_18288,N_14900,N_10922);
or U18289 (N_18289,N_10044,N_10706);
nand U18290 (N_18290,N_12570,N_11273);
or U18291 (N_18291,N_14573,N_10184);
or U18292 (N_18292,N_14218,N_13895);
or U18293 (N_18293,N_10600,N_12610);
nor U18294 (N_18294,N_10375,N_12211);
nand U18295 (N_18295,N_10970,N_13836);
nor U18296 (N_18296,N_14312,N_11759);
nand U18297 (N_18297,N_10788,N_13673);
and U18298 (N_18298,N_12463,N_11313);
or U18299 (N_18299,N_12365,N_10959);
xor U18300 (N_18300,N_14244,N_10979);
xor U18301 (N_18301,N_12280,N_11587);
nor U18302 (N_18302,N_13278,N_12960);
nor U18303 (N_18303,N_14890,N_10347);
nor U18304 (N_18304,N_11487,N_14694);
or U18305 (N_18305,N_13988,N_13949);
nand U18306 (N_18306,N_14040,N_12942);
nor U18307 (N_18307,N_14293,N_14955);
nand U18308 (N_18308,N_11657,N_13924);
xnor U18309 (N_18309,N_11409,N_11972);
and U18310 (N_18310,N_11939,N_13401);
nand U18311 (N_18311,N_10429,N_12758);
nor U18312 (N_18312,N_13994,N_12294);
or U18313 (N_18313,N_14240,N_12866);
and U18314 (N_18314,N_11218,N_13366);
or U18315 (N_18315,N_14398,N_14090);
and U18316 (N_18316,N_13351,N_12155);
nor U18317 (N_18317,N_14066,N_14021);
xnor U18318 (N_18318,N_12990,N_13683);
or U18319 (N_18319,N_13884,N_14445);
xnor U18320 (N_18320,N_14608,N_13861);
nand U18321 (N_18321,N_11674,N_12216);
and U18322 (N_18322,N_14427,N_14502);
and U18323 (N_18323,N_11878,N_14217);
xor U18324 (N_18324,N_13966,N_13451);
or U18325 (N_18325,N_11596,N_10704);
nor U18326 (N_18326,N_14050,N_13831);
xnor U18327 (N_18327,N_12925,N_13347);
nand U18328 (N_18328,N_10613,N_14849);
and U18329 (N_18329,N_11342,N_12189);
and U18330 (N_18330,N_11159,N_10756);
nor U18331 (N_18331,N_13668,N_12329);
nor U18332 (N_18332,N_12287,N_14906);
or U18333 (N_18333,N_10137,N_10589);
nor U18334 (N_18334,N_13053,N_14268);
xnor U18335 (N_18335,N_10777,N_10734);
or U18336 (N_18336,N_11345,N_11005);
and U18337 (N_18337,N_13422,N_12127);
xor U18338 (N_18338,N_12146,N_10281);
xor U18339 (N_18339,N_13216,N_11899);
and U18340 (N_18340,N_11741,N_13089);
or U18341 (N_18341,N_13909,N_11799);
nor U18342 (N_18342,N_14907,N_10874);
and U18343 (N_18343,N_10706,N_12314);
nor U18344 (N_18344,N_13935,N_13618);
xor U18345 (N_18345,N_10656,N_14157);
or U18346 (N_18346,N_11398,N_11638);
nand U18347 (N_18347,N_12846,N_10034);
or U18348 (N_18348,N_13515,N_10328);
xnor U18349 (N_18349,N_10765,N_14922);
nand U18350 (N_18350,N_11217,N_14385);
and U18351 (N_18351,N_12007,N_10972);
xnor U18352 (N_18352,N_10782,N_11300);
xnor U18353 (N_18353,N_14334,N_12742);
nand U18354 (N_18354,N_10232,N_10281);
nand U18355 (N_18355,N_13571,N_12764);
and U18356 (N_18356,N_14156,N_12206);
and U18357 (N_18357,N_13538,N_12697);
nor U18358 (N_18358,N_10086,N_11421);
xor U18359 (N_18359,N_10967,N_13767);
or U18360 (N_18360,N_12098,N_14768);
xor U18361 (N_18361,N_12915,N_11294);
and U18362 (N_18362,N_13889,N_14220);
nor U18363 (N_18363,N_10258,N_10543);
nor U18364 (N_18364,N_14346,N_10693);
and U18365 (N_18365,N_11475,N_11252);
nand U18366 (N_18366,N_10179,N_12295);
or U18367 (N_18367,N_11913,N_11145);
and U18368 (N_18368,N_12005,N_14836);
nor U18369 (N_18369,N_14828,N_14265);
and U18370 (N_18370,N_14418,N_13453);
or U18371 (N_18371,N_10916,N_13084);
nand U18372 (N_18372,N_11456,N_10054);
nor U18373 (N_18373,N_12634,N_10873);
nand U18374 (N_18374,N_14815,N_14656);
xor U18375 (N_18375,N_13074,N_12780);
and U18376 (N_18376,N_14542,N_12883);
nand U18377 (N_18377,N_14392,N_14201);
nand U18378 (N_18378,N_14870,N_10522);
nand U18379 (N_18379,N_12408,N_13452);
and U18380 (N_18380,N_12960,N_12121);
nand U18381 (N_18381,N_12533,N_13452);
nor U18382 (N_18382,N_14565,N_14560);
nor U18383 (N_18383,N_13568,N_11763);
or U18384 (N_18384,N_12429,N_14162);
or U18385 (N_18385,N_12451,N_13248);
or U18386 (N_18386,N_12198,N_10358);
nand U18387 (N_18387,N_10853,N_14636);
nand U18388 (N_18388,N_11098,N_14098);
nor U18389 (N_18389,N_10279,N_10571);
xor U18390 (N_18390,N_11953,N_11890);
and U18391 (N_18391,N_14615,N_11388);
xnor U18392 (N_18392,N_14944,N_11972);
nand U18393 (N_18393,N_10157,N_13407);
xor U18394 (N_18394,N_11693,N_11384);
xor U18395 (N_18395,N_10617,N_11586);
nand U18396 (N_18396,N_13251,N_10071);
xor U18397 (N_18397,N_13571,N_14194);
nand U18398 (N_18398,N_14783,N_10501);
nor U18399 (N_18399,N_13917,N_10532);
and U18400 (N_18400,N_10665,N_11758);
nor U18401 (N_18401,N_12381,N_12909);
xor U18402 (N_18402,N_14906,N_14692);
and U18403 (N_18403,N_11863,N_14236);
nor U18404 (N_18404,N_14386,N_11246);
nand U18405 (N_18405,N_13896,N_12717);
nor U18406 (N_18406,N_10123,N_14924);
or U18407 (N_18407,N_11265,N_12199);
xnor U18408 (N_18408,N_10661,N_11289);
and U18409 (N_18409,N_13002,N_12075);
xnor U18410 (N_18410,N_12925,N_12870);
and U18411 (N_18411,N_12612,N_10179);
nor U18412 (N_18412,N_11024,N_14368);
xor U18413 (N_18413,N_11952,N_12659);
nand U18414 (N_18414,N_11890,N_12836);
nor U18415 (N_18415,N_10268,N_12481);
and U18416 (N_18416,N_11007,N_13657);
nand U18417 (N_18417,N_13629,N_12433);
or U18418 (N_18418,N_13765,N_12690);
nand U18419 (N_18419,N_11523,N_12683);
nand U18420 (N_18420,N_12463,N_11572);
or U18421 (N_18421,N_14533,N_10001);
or U18422 (N_18422,N_12723,N_12397);
xnor U18423 (N_18423,N_10697,N_10181);
or U18424 (N_18424,N_14975,N_12390);
or U18425 (N_18425,N_10809,N_11723);
and U18426 (N_18426,N_14347,N_10302);
or U18427 (N_18427,N_12787,N_10072);
nor U18428 (N_18428,N_11345,N_14770);
and U18429 (N_18429,N_10876,N_11875);
or U18430 (N_18430,N_10785,N_13080);
or U18431 (N_18431,N_13349,N_13005);
nand U18432 (N_18432,N_13376,N_11395);
nand U18433 (N_18433,N_14564,N_11513);
xor U18434 (N_18434,N_12920,N_12413);
and U18435 (N_18435,N_13241,N_13392);
nor U18436 (N_18436,N_11310,N_11221);
xor U18437 (N_18437,N_12426,N_10681);
nor U18438 (N_18438,N_11661,N_11251);
or U18439 (N_18439,N_11719,N_12988);
xor U18440 (N_18440,N_13266,N_13847);
xor U18441 (N_18441,N_13263,N_11387);
nand U18442 (N_18442,N_14833,N_11384);
or U18443 (N_18443,N_14340,N_14022);
xnor U18444 (N_18444,N_12566,N_10566);
or U18445 (N_18445,N_10641,N_12308);
nand U18446 (N_18446,N_12976,N_13299);
xor U18447 (N_18447,N_12997,N_10620);
and U18448 (N_18448,N_11977,N_12734);
or U18449 (N_18449,N_14817,N_11117);
nor U18450 (N_18450,N_13979,N_10507);
or U18451 (N_18451,N_11431,N_14840);
and U18452 (N_18452,N_12323,N_12222);
nand U18453 (N_18453,N_14136,N_14093);
nor U18454 (N_18454,N_10364,N_13664);
nor U18455 (N_18455,N_11163,N_12745);
and U18456 (N_18456,N_12187,N_13590);
nor U18457 (N_18457,N_13058,N_11241);
xnor U18458 (N_18458,N_14930,N_12709);
xor U18459 (N_18459,N_10268,N_11108);
or U18460 (N_18460,N_12705,N_14995);
and U18461 (N_18461,N_11273,N_12840);
and U18462 (N_18462,N_10264,N_12197);
nand U18463 (N_18463,N_13513,N_12639);
xnor U18464 (N_18464,N_10255,N_12259);
nor U18465 (N_18465,N_13097,N_10947);
or U18466 (N_18466,N_11093,N_13026);
or U18467 (N_18467,N_13757,N_10328);
or U18468 (N_18468,N_11285,N_11160);
nand U18469 (N_18469,N_11205,N_10137);
nor U18470 (N_18470,N_12083,N_14609);
or U18471 (N_18471,N_12701,N_10108);
nor U18472 (N_18472,N_12651,N_11601);
nand U18473 (N_18473,N_11444,N_14053);
nand U18474 (N_18474,N_14836,N_12276);
and U18475 (N_18475,N_13450,N_10576);
or U18476 (N_18476,N_12724,N_13607);
nor U18477 (N_18477,N_12556,N_13640);
nand U18478 (N_18478,N_13460,N_12464);
nand U18479 (N_18479,N_11536,N_11712);
nand U18480 (N_18480,N_14537,N_13600);
and U18481 (N_18481,N_10352,N_12147);
xor U18482 (N_18482,N_13752,N_11453);
and U18483 (N_18483,N_11823,N_13589);
nand U18484 (N_18484,N_13294,N_12473);
xnor U18485 (N_18485,N_14502,N_10043);
or U18486 (N_18486,N_13365,N_14638);
xnor U18487 (N_18487,N_12982,N_12918);
nand U18488 (N_18488,N_13502,N_11779);
xnor U18489 (N_18489,N_11058,N_13010);
and U18490 (N_18490,N_12119,N_12039);
nor U18491 (N_18491,N_12008,N_10784);
xor U18492 (N_18492,N_13444,N_14770);
xor U18493 (N_18493,N_10078,N_10430);
or U18494 (N_18494,N_11607,N_14906);
or U18495 (N_18495,N_11182,N_11368);
or U18496 (N_18496,N_14196,N_11363);
and U18497 (N_18497,N_10412,N_12730);
nor U18498 (N_18498,N_10631,N_14397);
and U18499 (N_18499,N_13243,N_10362);
xnor U18500 (N_18500,N_11834,N_13400);
and U18501 (N_18501,N_12956,N_14263);
xnor U18502 (N_18502,N_11220,N_10917);
and U18503 (N_18503,N_10248,N_10464);
xor U18504 (N_18504,N_10936,N_14537);
and U18505 (N_18505,N_14619,N_10668);
xnor U18506 (N_18506,N_12123,N_14730);
and U18507 (N_18507,N_14206,N_13167);
or U18508 (N_18508,N_11600,N_13692);
or U18509 (N_18509,N_13821,N_12639);
nor U18510 (N_18510,N_13281,N_13258);
or U18511 (N_18511,N_11847,N_11424);
or U18512 (N_18512,N_11649,N_10068);
nor U18513 (N_18513,N_13415,N_11513);
or U18514 (N_18514,N_14029,N_10437);
or U18515 (N_18515,N_12938,N_11958);
nor U18516 (N_18516,N_14262,N_14376);
nor U18517 (N_18517,N_10890,N_13970);
xnor U18518 (N_18518,N_11048,N_13902);
and U18519 (N_18519,N_11982,N_10650);
nand U18520 (N_18520,N_14921,N_11985);
and U18521 (N_18521,N_11360,N_10727);
or U18522 (N_18522,N_10684,N_11584);
nor U18523 (N_18523,N_14548,N_11066);
xnor U18524 (N_18524,N_10447,N_14735);
nand U18525 (N_18525,N_13057,N_12181);
or U18526 (N_18526,N_10922,N_14707);
nand U18527 (N_18527,N_12828,N_13744);
and U18528 (N_18528,N_13713,N_10549);
or U18529 (N_18529,N_14002,N_11251);
xor U18530 (N_18530,N_13626,N_11070);
nand U18531 (N_18531,N_10101,N_12337);
xnor U18532 (N_18532,N_14499,N_14303);
xor U18533 (N_18533,N_12704,N_13559);
xnor U18534 (N_18534,N_11347,N_14631);
xnor U18535 (N_18535,N_14210,N_12319);
or U18536 (N_18536,N_13336,N_12767);
nor U18537 (N_18537,N_13839,N_12894);
nor U18538 (N_18538,N_12382,N_13071);
nor U18539 (N_18539,N_14315,N_11891);
nor U18540 (N_18540,N_13387,N_10763);
nand U18541 (N_18541,N_13919,N_14064);
xor U18542 (N_18542,N_13030,N_13771);
and U18543 (N_18543,N_10924,N_12899);
xor U18544 (N_18544,N_10533,N_13298);
xnor U18545 (N_18545,N_12365,N_13054);
or U18546 (N_18546,N_12437,N_10060);
and U18547 (N_18547,N_10705,N_11382);
xnor U18548 (N_18548,N_13564,N_10869);
or U18549 (N_18549,N_14611,N_12596);
xor U18550 (N_18550,N_11510,N_11384);
xor U18551 (N_18551,N_12069,N_11657);
or U18552 (N_18552,N_12516,N_10673);
and U18553 (N_18553,N_12290,N_11516);
or U18554 (N_18554,N_10424,N_10825);
or U18555 (N_18555,N_10698,N_11639);
and U18556 (N_18556,N_13753,N_10038);
xnor U18557 (N_18557,N_14080,N_14960);
nand U18558 (N_18558,N_10445,N_12373);
xnor U18559 (N_18559,N_11470,N_13393);
nand U18560 (N_18560,N_14105,N_14766);
xnor U18561 (N_18561,N_11663,N_12751);
nor U18562 (N_18562,N_10367,N_12515);
and U18563 (N_18563,N_14515,N_13357);
and U18564 (N_18564,N_14153,N_12734);
nand U18565 (N_18565,N_14534,N_14927);
nor U18566 (N_18566,N_11692,N_14659);
xor U18567 (N_18567,N_14910,N_11874);
or U18568 (N_18568,N_13721,N_12073);
or U18569 (N_18569,N_12966,N_11344);
and U18570 (N_18570,N_13172,N_12591);
nand U18571 (N_18571,N_14241,N_10998);
or U18572 (N_18572,N_10961,N_13980);
xnor U18573 (N_18573,N_12536,N_11592);
xor U18574 (N_18574,N_12594,N_14536);
xor U18575 (N_18575,N_11889,N_13763);
xor U18576 (N_18576,N_11718,N_13701);
nand U18577 (N_18577,N_11926,N_14843);
and U18578 (N_18578,N_14627,N_10888);
xnor U18579 (N_18579,N_12500,N_12323);
and U18580 (N_18580,N_14265,N_10800);
nor U18581 (N_18581,N_12596,N_12742);
nand U18582 (N_18582,N_14330,N_13997);
or U18583 (N_18583,N_14683,N_14636);
xor U18584 (N_18584,N_12986,N_10891);
nand U18585 (N_18585,N_14661,N_10425);
xor U18586 (N_18586,N_10870,N_13463);
xnor U18587 (N_18587,N_14106,N_12767);
and U18588 (N_18588,N_10840,N_13045);
xnor U18589 (N_18589,N_14658,N_12007);
nor U18590 (N_18590,N_12848,N_14180);
or U18591 (N_18591,N_13046,N_10194);
xnor U18592 (N_18592,N_10414,N_10330);
or U18593 (N_18593,N_11739,N_11648);
nand U18594 (N_18594,N_11928,N_10213);
and U18595 (N_18595,N_13886,N_14499);
nor U18596 (N_18596,N_14440,N_11900);
nand U18597 (N_18597,N_12919,N_14099);
nor U18598 (N_18598,N_12272,N_14242);
nand U18599 (N_18599,N_14651,N_14064);
and U18600 (N_18600,N_10661,N_12370);
or U18601 (N_18601,N_14929,N_13754);
and U18602 (N_18602,N_12371,N_10911);
nand U18603 (N_18603,N_14954,N_10478);
xnor U18604 (N_18604,N_13842,N_11605);
xor U18605 (N_18605,N_10014,N_13497);
or U18606 (N_18606,N_10377,N_13413);
xor U18607 (N_18607,N_12266,N_10380);
or U18608 (N_18608,N_14199,N_12967);
nand U18609 (N_18609,N_12570,N_14943);
or U18610 (N_18610,N_13720,N_11617);
xnor U18611 (N_18611,N_14891,N_11005);
xnor U18612 (N_18612,N_13444,N_14818);
or U18613 (N_18613,N_11195,N_10885);
and U18614 (N_18614,N_11950,N_12631);
or U18615 (N_18615,N_13645,N_13850);
nand U18616 (N_18616,N_11811,N_14047);
nor U18617 (N_18617,N_12174,N_11452);
and U18618 (N_18618,N_14524,N_12356);
xor U18619 (N_18619,N_10046,N_13494);
nand U18620 (N_18620,N_10436,N_12354);
nor U18621 (N_18621,N_10588,N_13733);
and U18622 (N_18622,N_10649,N_11367);
nor U18623 (N_18623,N_12441,N_11348);
nor U18624 (N_18624,N_11626,N_13358);
or U18625 (N_18625,N_11259,N_14543);
nor U18626 (N_18626,N_10136,N_10332);
nor U18627 (N_18627,N_13922,N_10306);
or U18628 (N_18628,N_13668,N_14972);
nor U18629 (N_18629,N_13235,N_11708);
and U18630 (N_18630,N_14529,N_12130);
and U18631 (N_18631,N_13081,N_12060);
or U18632 (N_18632,N_10767,N_12669);
nand U18633 (N_18633,N_12242,N_10634);
nand U18634 (N_18634,N_13234,N_10035);
nor U18635 (N_18635,N_10513,N_11510);
and U18636 (N_18636,N_13672,N_12934);
nand U18637 (N_18637,N_12357,N_11534);
and U18638 (N_18638,N_11742,N_10338);
nor U18639 (N_18639,N_12400,N_14950);
nor U18640 (N_18640,N_10683,N_13875);
xor U18641 (N_18641,N_12380,N_11949);
and U18642 (N_18642,N_10434,N_10406);
and U18643 (N_18643,N_14470,N_13695);
nand U18644 (N_18644,N_10524,N_13820);
nor U18645 (N_18645,N_10396,N_10663);
nand U18646 (N_18646,N_10819,N_14007);
and U18647 (N_18647,N_11818,N_11150);
nor U18648 (N_18648,N_10148,N_13728);
xor U18649 (N_18649,N_12835,N_12882);
nand U18650 (N_18650,N_10244,N_10602);
nor U18651 (N_18651,N_10570,N_10959);
xor U18652 (N_18652,N_11894,N_10268);
nand U18653 (N_18653,N_14683,N_11452);
nand U18654 (N_18654,N_13858,N_12162);
and U18655 (N_18655,N_12502,N_12097);
xnor U18656 (N_18656,N_14097,N_13868);
nand U18657 (N_18657,N_11071,N_11869);
xnor U18658 (N_18658,N_10179,N_12610);
nor U18659 (N_18659,N_11056,N_10619);
or U18660 (N_18660,N_10327,N_10731);
or U18661 (N_18661,N_10820,N_12423);
xor U18662 (N_18662,N_14473,N_10670);
xor U18663 (N_18663,N_11322,N_11425);
nand U18664 (N_18664,N_10502,N_10791);
or U18665 (N_18665,N_11495,N_11440);
xor U18666 (N_18666,N_12426,N_13394);
xor U18667 (N_18667,N_10116,N_10169);
and U18668 (N_18668,N_11609,N_14946);
or U18669 (N_18669,N_13389,N_13424);
nand U18670 (N_18670,N_14811,N_13975);
xnor U18671 (N_18671,N_14874,N_12863);
nand U18672 (N_18672,N_11282,N_11356);
nand U18673 (N_18673,N_11837,N_13628);
and U18674 (N_18674,N_14148,N_12112);
xor U18675 (N_18675,N_14339,N_10615);
nand U18676 (N_18676,N_12762,N_14949);
nor U18677 (N_18677,N_13924,N_10226);
nor U18678 (N_18678,N_12835,N_14775);
xor U18679 (N_18679,N_11249,N_11804);
and U18680 (N_18680,N_13458,N_14688);
nor U18681 (N_18681,N_14781,N_13228);
xor U18682 (N_18682,N_10994,N_11689);
and U18683 (N_18683,N_10848,N_10971);
nor U18684 (N_18684,N_11636,N_13868);
nand U18685 (N_18685,N_11007,N_14444);
and U18686 (N_18686,N_10667,N_14524);
and U18687 (N_18687,N_10774,N_10100);
nand U18688 (N_18688,N_14051,N_13139);
xor U18689 (N_18689,N_12077,N_14330);
xor U18690 (N_18690,N_12785,N_13771);
and U18691 (N_18691,N_12615,N_12354);
nor U18692 (N_18692,N_10469,N_11912);
and U18693 (N_18693,N_10986,N_12441);
or U18694 (N_18694,N_10680,N_11359);
or U18695 (N_18695,N_12774,N_13115);
or U18696 (N_18696,N_11044,N_14077);
or U18697 (N_18697,N_14325,N_10258);
or U18698 (N_18698,N_12916,N_13448);
nand U18699 (N_18699,N_13423,N_12379);
nor U18700 (N_18700,N_12666,N_13274);
nor U18701 (N_18701,N_11922,N_14364);
and U18702 (N_18702,N_11241,N_12858);
xnor U18703 (N_18703,N_11011,N_11737);
or U18704 (N_18704,N_11182,N_11791);
and U18705 (N_18705,N_10540,N_10623);
and U18706 (N_18706,N_11355,N_14069);
nor U18707 (N_18707,N_10299,N_13591);
xor U18708 (N_18708,N_13569,N_11943);
and U18709 (N_18709,N_14427,N_10168);
nand U18710 (N_18710,N_13246,N_11059);
xnor U18711 (N_18711,N_11159,N_14708);
or U18712 (N_18712,N_14061,N_11367);
nand U18713 (N_18713,N_14256,N_13987);
xnor U18714 (N_18714,N_14314,N_14990);
and U18715 (N_18715,N_12900,N_14272);
and U18716 (N_18716,N_13196,N_14957);
xnor U18717 (N_18717,N_12768,N_12138);
xnor U18718 (N_18718,N_14623,N_13364);
nor U18719 (N_18719,N_11617,N_13916);
nand U18720 (N_18720,N_13391,N_14754);
or U18721 (N_18721,N_10728,N_13613);
nand U18722 (N_18722,N_12243,N_12085);
nor U18723 (N_18723,N_11795,N_12609);
xnor U18724 (N_18724,N_12517,N_10150);
nand U18725 (N_18725,N_12773,N_10330);
and U18726 (N_18726,N_12231,N_14419);
nand U18727 (N_18727,N_10857,N_12776);
nor U18728 (N_18728,N_11777,N_13826);
and U18729 (N_18729,N_13483,N_14499);
and U18730 (N_18730,N_10790,N_12341);
xnor U18731 (N_18731,N_11203,N_10087);
and U18732 (N_18732,N_13561,N_11451);
nor U18733 (N_18733,N_12978,N_12030);
and U18734 (N_18734,N_11201,N_14865);
nor U18735 (N_18735,N_14093,N_13000);
xor U18736 (N_18736,N_10457,N_10200);
nor U18737 (N_18737,N_14474,N_10977);
or U18738 (N_18738,N_10676,N_10852);
xnor U18739 (N_18739,N_11897,N_14053);
xor U18740 (N_18740,N_12870,N_11344);
xnor U18741 (N_18741,N_13960,N_13447);
xnor U18742 (N_18742,N_12047,N_14287);
xnor U18743 (N_18743,N_12053,N_12220);
xnor U18744 (N_18744,N_12552,N_12407);
nand U18745 (N_18745,N_10749,N_10898);
nand U18746 (N_18746,N_12102,N_12730);
nor U18747 (N_18747,N_12256,N_12090);
nand U18748 (N_18748,N_10342,N_14663);
or U18749 (N_18749,N_12715,N_13658);
or U18750 (N_18750,N_14434,N_12625);
or U18751 (N_18751,N_13322,N_11557);
and U18752 (N_18752,N_10200,N_12069);
or U18753 (N_18753,N_14820,N_13903);
and U18754 (N_18754,N_14283,N_12535);
nand U18755 (N_18755,N_12396,N_12624);
nand U18756 (N_18756,N_14457,N_14312);
and U18757 (N_18757,N_12584,N_11840);
nand U18758 (N_18758,N_10169,N_10726);
xor U18759 (N_18759,N_13709,N_13207);
xnor U18760 (N_18760,N_13050,N_13042);
or U18761 (N_18761,N_10920,N_10855);
or U18762 (N_18762,N_14698,N_10695);
nor U18763 (N_18763,N_14395,N_13754);
and U18764 (N_18764,N_11219,N_13613);
nand U18765 (N_18765,N_11318,N_13619);
nor U18766 (N_18766,N_10393,N_11960);
or U18767 (N_18767,N_11487,N_12112);
or U18768 (N_18768,N_10775,N_13875);
xor U18769 (N_18769,N_11297,N_11739);
nor U18770 (N_18770,N_13245,N_11152);
nand U18771 (N_18771,N_11216,N_11252);
nor U18772 (N_18772,N_11163,N_13844);
xnor U18773 (N_18773,N_13545,N_14133);
nor U18774 (N_18774,N_14746,N_10757);
nand U18775 (N_18775,N_12350,N_13431);
nor U18776 (N_18776,N_13292,N_12971);
nand U18777 (N_18777,N_14941,N_11538);
xor U18778 (N_18778,N_13815,N_10321);
nand U18779 (N_18779,N_11590,N_11025);
xor U18780 (N_18780,N_14136,N_12256);
xnor U18781 (N_18781,N_10003,N_10653);
or U18782 (N_18782,N_14556,N_13534);
nand U18783 (N_18783,N_13230,N_12323);
and U18784 (N_18784,N_12306,N_10750);
nand U18785 (N_18785,N_10067,N_14816);
xnor U18786 (N_18786,N_14394,N_14835);
and U18787 (N_18787,N_10661,N_14746);
nor U18788 (N_18788,N_13269,N_10478);
nor U18789 (N_18789,N_13532,N_10698);
nand U18790 (N_18790,N_14027,N_11487);
or U18791 (N_18791,N_12842,N_12732);
nand U18792 (N_18792,N_12439,N_10664);
nand U18793 (N_18793,N_12675,N_11705);
nor U18794 (N_18794,N_10560,N_14042);
and U18795 (N_18795,N_14430,N_11074);
nor U18796 (N_18796,N_10904,N_10964);
or U18797 (N_18797,N_12595,N_14806);
nand U18798 (N_18798,N_11717,N_11521);
or U18799 (N_18799,N_14662,N_14818);
xnor U18800 (N_18800,N_10701,N_11834);
nor U18801 (N_18801,N_13361,N_13321);
and U18802 (N_18802,N_14473,N_13611);
or U18803 (N_18803,N_10605,N_11968);
or U18804 (N_18804,N_11244,N_14715);
and U18805 (N_18805,N_11565,N_13389);
nor U18806 (N_18806,N_12666,N_14039);
or U18807 (N_18807,N_14417,N_11279);
and U18808 (N_18808,N_11405,N_13069);
and U18809 (N_18809,N_12519,N_12438);
nor U18810 (N_18810,N_12961,N_13314);
nor U18811 (N_18811,N_10974,N_10930);
or U18812 (N_18812,N_13054,N_10754);
and U18813 (N_18813,N_10587,N_10398);
or U18814 (N_18814,N_10586,N_12500);
nor U18815 (N_18815,N_12419,N_11892);
xor U18816 (N_18816,N_10577,N_11099);
and U18817 (N_18817,N_14278,N_13863);
and U18818 (N_18818,N_10747,N_12570);
or U18819 (N_18819,N_13284,N_12157);
nor U18820 (N_18820,N_13560,N_11503);
nor U18821 (N_18821,N_14805,N_12698);
nor U18822 (N_18822,N_14442,N_11829);
and U18823 (N_18823,N_12475,N_14405);
and U18824 (N_18824,N_10043,N_12080);
nand U18825 (N_18825,N_10307,N_10793);
nand U18826 (N_18826,N_14402,N_12921);
or U18827 (N_18827,N_12448,N_14668);
nor U18828 (N_18828,N_12195,N_10815);
or U18829 (N_18829,N_12728,N_14198);
nor U18830 (N_18830,N_11312,N_10375);
nand U18831 (N_18831,N_13442,N_13970);
and U18832 (N_18832,N_11258,N_14764);
nand U18833 (N_18833,N_11660,N_11079);
nand U18834 (N_18834,N_13320,N_12993);
xor U18835 (N_18835,N_11496,N_14024);
nor U18836 (N_18836,N_13230,N_10186);
and U18837 (N_18837,N_11711,N_13047);
and U18838 (N_18838,N_12371,N_13335);
or U18839 (N_18839,N_13197,N_13397);
or U18840 (N_18840,N_10214,N_11514);
nand U18841 (N_18841,N_12506,N_13091);
nand U18842 (N_18842,N_14720,N_13492);
or U18843 (N_18843,N_14734,N_13113);
or U18844 (N_18844,N_13287,N_14889);
nor U18845 (N_18845,N_14307,N_14587);
xnor U18846 (N_18846,N_11442,N_11195);
or U18847 (N_18847,N_11086,N_12440);
xor U18848 (N_18848,N_11425,N_12742);
nand U18849 (N_18849,N_14301,N_14375);
and U18850 (N_18850,N_13428,N_12821);
nand U18851 (N_18851,N_12897,N_10307);
and U18852 (N_18852,N_12920,N_13174);
nor U18853 (N_18853,N_13237,N_10729);
xnor U18854 (N_18854,N_14389,N_11377);
or U18855 (N_18855,N_11887,N_12571);
and U18856 (N_18856,N_10565,N_10662);
nand U18857 (N_18857,N_11469,N_10468);
and U18858 (N_18858,N_13713,N_14464);
xnor U18859 (N_18859,N_11919,N_14494);
nand U18860 (N_18860,N_13605,N_14787);
or U18861 (N_18861,N_13321,N_11382);
nor U18862 (N_18862,N_14997,N_13162);
or U18863 (N_18863,N_12311,N_14984);
nor U18864 (N_18864,N_12749,N_12252);
or U18865 (N_18865,N_11789,N_12841);
xnor U18866 (N_18866,N_12466,N_10399);
nor U18867 (N_18867,N_10613,N_10848);
and U18868 (N_18868,N_11612,N_10877);
or U18869 (N_18869,N_13596,N_14944);
or U18870 (N_18870,N_11018,N_14312);
nor U18871 (N_18871,N_12476,N_11651);
nand U18872 (N_18872,N_11012,N_11492);
xnor U18873 (N_18873,N_11615,N_14268);
nor U18874 (N_18874,N_10331,N_14689);
xor U18875 (N_18875,N_12546,N_13703);
nor U18876 (N_18876,N_10235,N_13957);
nand U18877 (N_18877,N_13274,N_11638);
xnor U18878 (N_18878,N_10104,N_13994);
xnor U18879 (N_18879,N_10409,N_13883);
and U18880 (N_18880,N_11962,N_10961);
xnor U18881 (N_18881,N_11335,N_12590);
xnor U18882 (N_18882,N_14146,N_12534);
or U18883 (N_18883,N_12864,N_10911);
nor U18884 (N_18884,N_13783,N_10603);
or U18885 (N_18885,N_11791,N_13803);
and U18886 (N_18886,N_11992,N_10590);
nand U18887 (N_18887,N_14847,N_10029);
and U18888 (N_18888,N_11058,N_10847);
and U18889 (N_18889,N_14258,N_12137);
nand U18890 (N_18890,N_14987,N_11294);
nand U18891 (N_18891,N_14099,N_14881);
or U18892 (N_18892,N_12675,N_13733);
or U18893 (N_18893,N_14477,N_13730);
or U18894 (N_18894,N_10078,N_12874);
nor U18895 (N_18895,N_13674,N_12915);
and U18896 (N_18896,N_12864,N_13190);
nor U18897 (N_18897,N_10626,N_13964);
nor U18898 (N_18898,N_10586,N_12784);
xor U18899 (N_18899,N_11787,N_12826);
and U18900 (N_18900,N_12023,N_11975);
and U18901 (N_18901,N_10188,N_12000);
or U18902 (N_18902,N_12139,N_14759);
xor U18903 (N_18903,N_11604,N_10950);
or U18904 (N_18904,N_13599,N_13486);
nand U18905 (N_18905,N_14782,N_13598);
and U18906 (N_18906,N_14614,N_14603);
or U18907 (N_18907,N_13087,N_14351);
xnor U18908 (N_18908,N_12562,N_14799);
and U18909 (N_18909,N_11843,N_14381);
nor U18910 (N_18910,N_13078,N_12243);
or U18911 (N_18911,N_12253,N_14488);
xnor U18912 (N_18912,N_13932,N_10823);
nand U18913 (N_18913,N_11476,N_14643);
nor U18914 (N_18914,N_13237,N_10857);
or U18915 (N_18915,N_12975,N_13410);
or U18916 (N_18916,N_10721,N_10203);
and U18917 (N_18917,N_13856,N_10260);
nor U18918 (N_18918,N_13953,N_10048);
nor U18919 (N_18919,N_13197,N_14253);
or U18920 (N_18920,N_11918,N_11188);
or U18921 (N_18921,N_12326,N_14189);
and U18922 (N_18922,N_11996,N_14610);
xor U18923 (N_18923,N_13222,N_10986);
or U18924 (N_18924,N_11030,N_10409);
nand U18925 (N_18925,N_14158,N_14226);
nand U18926 (N_18926,N_12541,N_14619);
nor U18927 (N_18927,N_12290,N_11879);
nor U18928 (N_18928,N_12108,N_11049);
nor U18929 (N_18929,N_10902,N_12213);
nand U18930 (N_18930,N_14707,N_13667);
and U18931 (N_18931,N_12442,N_11315);
xnor U18932 (N_18932,N_11418,N_12667);
or U18933 (N_18933,N_11666,N_13546);
xor U18934 (N_18934,N_12080,N_10707);
xor U18935 (N_18935,N_11192,N_13943);
xnor U18936 (N_18936,N_13247,N_12193);
xor U18937 (N_18937,N_12817,N_12085);
or U18938 (N_18938,N_14752,N_11951);
nand U18939 (N_18939,N_10136,N_13685);
nor U18940 (N_18940,N_12651,N_12621);
nor U18941 (N_18941,N_12342,N_14048);
and U18942 (N_18942,N_14176,N_13673);
and U18943 (N_18943,N_10774,N_13666);
and U18944 (N_18944,N_10751,N_14463);
xor U18945 (N_18945,N_13127,N_10416);
nand U18946 (N_18946,N_13614,N_13264);
and U18947 (N_18947,N_14129,N_13483);
nor U18948 (N_18948,N_12834,N_12571);
nand U18949 (N_18949,N_14506,N_11551);
nor U18950 (N_18950,N_12804,N_12919);
or U18951 (N_18951,N_12222,N_11494);
or U18952 (N_18952,N_12446,N_14434);
and U18953 (N_18953,N_10608,N_13417);
and U18954 (N_18954,N_11371,N_13049);
and U18955 (N_18955,N_12325,N_12683);
xnor U18956 (N_18956,N_14301,N_13654);
nor U18957 (N_18957,N_11648,N_11322);
nand U18958 (N_18958,N_14295,N_12531);
and U18959 (N_18959,N_11987,N_10034);
xnor U18960 (N_18960,N_14401,N_10209);
xor U18961 (N_18961,N_12807,N_14628);
and U18962 (N_18962,N_12865,N_10654);
or U18963 (N_18963,N_12919,N_12922);
or U18964 (N_18964,N_11133,N_14045);
nand U18965 (N_18965,N_10789,N_11813);
nor U18966 (N_18966,N_14880,N_10603);
or U18967 (N_18967,N_14404,N_14139);
and U18968 (N_18968,N_11224,N_14127);
nand U18969 (N_18969,N_13734,N_10250);
xor U18970 (N_18970,N_12726,N_13591);
nor U18971 (N_18971,N_14794,N_14634);
and U18972 (N_18972,N_13824,N_14516);
nor U18973 (N_18973,N_11203,N_10601);
nor U18974 (N_18974,N_11660,N_14449);
and U18975 (N_18975,N_14124,N_11510);
xnor U18976 (N_18976,N_14764,N_12006);
xor U18977 (N_18977,N_10669,N_12477);
nor U18978 (N_18978,N_14118,N_13328);
nand U18979 (N_18979,N_12417,N_10276);
xor U18980 (N_18980,N_11215,N_11306);
or U18981 (N_18981,N_14091,N_14574);
or U18982 (N_18982,N_13377,N_14928);
or U18983 (N_18983,N_12265,N_10168);
xor U18984 (N_18984,N_11930,N_10525);
nand U18985 (N_18985,N_10687,N_12744);
xnor U18986 (N_18986,N_14400,N_10065);
xnor U18987 (N_18987,N_14263,N_14206);
xor U18988 (N_18988,N_13279,N_13489);
or U18989 (N_18989,N_12441,N_11489);
or U18990 (N_18990,N_11496,N_14246);
xor U18991 (N_18991,N_13409,N_11270);
xnor U18992 (N_18992,N_13705,N_10422);
nand U18993 (N_18993,N_11412,N_13065);
nor U18994 (N_18994,N_10498,N_11164);
or U18995 (N_18995,N_11696,N_14296);
or U18996 (N_18996,N_10008,N_11568);
or U18997 (N_18997,N_14936,N_10203);
nand U18998 (N_18998,N_14453,N_13747);
and U18999 (N_18999,N_11058,N_10160);
nand U19000 (N_19000,N_10994,N_10785);
or U19001 (N_19001,N_11866,N_10247);
nor U19002 (N_19002,N_14279,N_14435);
or U19003 (N_19003,N_13744,N_10607);
nand U19004 (N_19004,N_13585,N_10140);
or U19005 (N_19005,N_12438,N_13556);
xor U19006 (N_19006,N_12016,N_14514);
nor U19007 (N_19007,N_13306,N_12762);
and U19008 (N_19008,N_13698,N_14351);
xor U19009 (N_19009,N_10996,N_14401);
nor U19010 (N_19010,N_12714,N_13598);
nand U19011 (N_19011,N_14089,N_14295);
nor U19012 (N_19012,N_10035,N_10892);
xnor U19013 (N_19013,N_12904,N_10550);
nand U19014 (N_19014,N_13585,N_11074);
or U19015 (N_19015,N_11217,N_14451);
nand U19016 (N_19016,N_13737,N_12738);
nand U19017 (N_19017,N_11822,N_11666);
or U19018 (N_19018,N_13407,N_12759);
and U19019 (N_19019,N_12783,N_13512);
nor U19020 (N_19020,N_11242,N_10193);
or U19021 (N_19021,N_11090,N_13683);
xor U19022 (N_19022,N_10437,N_10851);
and U19023 (N_19023,N_13215,N_12188);
nand U19024 (N_19024,N_14940,N_12744);
xnor U19025 (N_19025,N_10840,N_12607);
nor U19026 (N_19026,N_14674,N_14364);
and U19027 (N_19027,N_14307,N_10028);
nand U19028 (N_19028,N_11154,N_13102);
and U19029 (N_19029,N_10528,N_10858);
and U19030 (N_19030,N_14502,N_11384);
and U19031 (N_19031,N_13639,N_11488);
or U19032 (N_19032,N_12394,N_14097);
nand U19033 (N_19033,N_12752,N_10647);
nand U19034 (N_19034,N_14447,N_12559);
nand U19035 (N_19035,N_11164,N_10571);
and U19036 (N_19036,N_11872,N_12732);
nor U19037 (N_19037,N_12499,N_13111);
xor U19038 (N_19038,N_12038,N_11146);
nor U19039 (N_19039,N_13625,N_13330);
nand U19040 (N_19040,N_10886,N_13761);
nand U19041 (N_19041,N_13949,N_10200);
xnor U19042 (N_19042,N_14200,N_13251);
nand U19043 (N_19043,N_13441,N_12136);
or U19044 (N_19044,N_11009,N_14048);
and U19045 (N_19045,N_11845,N_12557);
or U19046 (N_19046,N_14631,N_10844);
or U19047 (N_19047,N_13748,N_13321);
nand U19048 (N_19048,N_13854,N_11363);
or U19049 (N_19049,N_10233,N_10880);
nand U19050 (N_19050,N_11787,N_12580);
xor U19051 (N_19051,N_11208,N_11555);
and U19052 (N_19052,N_13152,N_13206);
and U19053 (N_19053,N_14010,N_10474);
xnor U19054 (N_19054,N_10985,N_10199);
and U19055 (N_19055,N_12674,N_10775);
or U19056 (N_19056,N_10267,N_14435);
xor U19057 (N_19057,N_13177,N_11554);
nor U19058 (N_19058,N_13393,N_10801);
nor U19059 (N_19059,N_14375,N_12098);
nor U19060 (N_19060,N_11327,N_10157);
nor U19061 (N_19061,N_10827,N_11613);
nor U19062 (N_19062,N_10562,N_14955);
or U19063 (N_19063,N_14106,N_12234);
xor U19064 (N_19064,N_10132,N_14816);
xnor U19065 (N_19065,N_14063,N_14688);
nand U19066 (N_19066,N_10125,N_12925);
nor U19067 (N_19067,N_11828,N_10371);
nor U19068 (N_19068,N_10393,N_14244);
and U19069 (N_19069,N_12343,N_10372);
xor U19070 (N_19070,N_11569,N_12867);
nor U19071 (N_19071,N_13431,N_13427);
xor U19072 (N_19072,N_12210,N_12054);
and U19073 (N_19073,N_13503,N_13076);
nand U19074 (N_19074,N_12418,N_11391);
and U19075 (N_19075,N_10445,N_12559);
or U19076 (N_19076,N_11463,N_14631);
xnor U19077 (N_19077,N_13886,N_14258);
or U19078 (N_19078,N_11568,N_12516);
nor U19079 (N_19079,N_12884,N_14616);
nand U19080 (N_19080,N_12766,N_13130);
nand U19081 (N_19081,N_11068,N_10951);
nand U19082 (N_19082,N_13830,N_10710);
nand U19083 (N_19083,N_14993,N_10896);
nor U19084 (N_19084,N_14895,N_11872);
or U19085 (N_19085,N_14479,N_11651);
xor U19086 (N_19086,N_11473,N_11095);
nor U19087 (N_19087,N_14639,N_14675);
and U19088 (N_19088,N_10818,N_10584);
and U19089 (N_19089,N_14586,N_11503);
nand U19090 (N_19090,N_14802,N_14007);
xnor U19091 (N_19091,N_14052,N_11869);
or U19092 (N_19092,N_12322,N_12600);
nor U19093 (N_19093,N_14912,N_14411);
xor U19094 (N_19094,N_13471,N_14431);
or U19095 (N_19095,N_13060,N_12768);
nor U19096 (N_19096,N_10021,N_11170);
or U19097 (N_19097,N_10978,N_13394);
and U19098 (N_19098,N_13265,N_10550);
nand U19099 (N_19099,N_10064,N_12931);
nor U19100 (N_19100,N_13517,N_10509);
nor U19101 (N_19101,N_12324,N_11453);
xor U19102 (N_19102,N_13600,N_13270);
or U19103 (N_19103,N_13310,N_12894);
nand U19104 (N_19104,N_12322,N_13051);
or U19105 (N_19105,N_11239,N_11892);
nor U19106 (N_19106,N_14400,N_13393);
xnor U19107 (N_19107,N_13487,N_14862);
or U19108 (N_19108,N_14521,N_11543);
xor U19109 (N_19109,N_11208,N_13110);
nor U19110 (N_19110,N_14302,N_10874);
nor U19111 (N_19111,N_10814,N_14696);
and U19112 (N_19112,N_11816,N_11929);
nor U19113 (N_19113,N_13565,N_11005);
xnor U19114 (N_19114,N_11320,N_13491);
and U19115 (N_19115,N_11285,N_12188);
or U19116 (N_19116,N_13565,N_11889);
or U19117 (N_19117,N_12621,N_13148);
nand U19118 (N_19118,N_13876,N_11834);
and U19119 (N_19119,N_14777,N_11792);
and U19120 (N_19120,N_14058,N_14522);
nand U19121 (N_19121,N_11945,N_11418);
or U19122 (N_19122,N_12314,N_14532);
xor U19123 (N_19123,N_13030,N_14837);
nand U19124 (N_19124,N_14060,N_13069);
and U19125 (N_19125,N_13396,N_14977);
nand U19126 (N_19126,N_12144,N_11784);
xnor U19127 (N_19127,N_10603,N_11072);
nor U19128 (N_19128,N_14403,N_14357);
xnor U19129 (N_19129,N_11464,N_14299);
xor U19130 (N_19130,N_14920,N_14900);
nand U19131 (N_19131,N_11927,N_12044);
xnor U19132 (N_19132,N_13742,N_10742);
nor U19133 (N_19133,N_10532,N_11154);
nand U19134 (N_19134,N_13364,N_10892);
nor U19135 (N_19135,N_13364,N_12510);
xor U19136 (N_19136,N_12715,N_14889);
and U19137 (N_19137,N_10835,N_12660);
nand U19138 (N_19138,N_12466,N_13365);
xnor U19139 (N_19139,N_12550,N_11646);
xor U19140 (N_19140,N_14435,N_14454);
nand U19141 (N_19141,N_10542,N_11720);
nand U19142 (N_19142,N_13669,N_13895);
nand U19143 (N_19143,N_12767,N_12530);
xor U19144 (N_19144,N_13035,N_11265);
or U19145 (N_19145,N_11543,N_13238);
or U19146 (N_19146,N_10614,N_13329);
nand U19147 (N_19147,N_11835,N_14359);
nor U19148 (N_19148,N_14054,N_10892);
or U19149 (N_19149,N_13468,N_10697);
xnor U19150 (N_19150,N_11306,N_12104);
nand U19151 (N_19151,N_11360,N_14449);
xnor U19152 (N_19152,N_10867,N_13036);
or U19153 (N_19153,N_11349,N_14533);
and U19154 (N_19154,N_13257,N_10513);
nor U19155 (N_19155,N_12309,N_10629);
nand U19156 (N_19156,N_14194,N_14753);
and U19157 (N_19157,N_12651,N_14279);
and U19158 (N_19158,N_12772,N_10111);
and U19159 (N_19159,N_12462,N_12810);
nand U19160 (N_19160,N_10750,N_14811);
or U19161 (N_19161,N_10891,N_12408);
and U19162 (N_19162,N_14970,N_10078);
or U19163 (N_19163,N_13763,N_14973);
or U19164 (N_19164,N_14774,N_14599);
xnor U19165 (N_19165,N_13063,N_12092);
or U19166 (N_19166,N_10671,N_11947);
or U19167 (N_19167,N_13241,N_11996);
or U19168 (N_19168,N_14668,N_14831);
xnor U19169 (N_19169,N_14060,N_10386);
nand U19170 (N_19170,N_12517,N_10360);
nor U19171 (N_19171,N_14530,N_10554);
or U19172 (N_19172,N_12153,N_12201);
nor U19173 (N_19173,N_13269,N_14255);
nor U19174 (N_19174,N_12951,N_13170);
nor U19175 (N_19175,N_14880,N_11977);
or U19176 (N_19176,N_14056,N_10713);
and U19177 (N_19177,N_12813,N_10456);
nor U19178 (N_19178,N_14801,N_10760);
nor U19179 (N_19179,N_12639,N_14635);
nand U19180 (N_19180,N_14147,N_13842);
or U19181 (N_19181,N_11608,N_11487);
nand U19182 (N_19182,N_11032,N_10309);
nand U19183 (N_19183,N_13611,N_10374);
and U19184 (N_19184,N_12843,N_14135);
nor U19185 (N_19185,N_10802,N_13026);
nand U19186 (N_19186,N_11212,N_10043);
nand U19187 (N_19187,N_10144,N_11982);
and U19188 (N_19188,N_10436,N_11843);
nor U19189 (N_19189,N_11047,N_10297);
xor U19190 (N_19190,N_14901,N_11436);
xor U19191 (N_19191,N_10781,N_13264);
nand U19192 (N_19192,N_10982,N_10321);
nand U19193 (N_19193,N_11587,N_14949);
or U19194 (N_19194,N_11074,N_10387);
xnor U19195 (N_19195,N_12386,N_14824);
nor U19196 (N_19196,N_13886,N_10974);
nor U19197 (N_19197,N_13333,N_13367);
nand U19198 (N_19198,N_10534,N_11152);
nand U19199 (N_19199,N_11050,N_14201);
or U19200 (N_19200,N_10140,N_13181);
and U19201 (N_19201,N_11392,N_13404);
and U19202 (N_19202,N_12243,N_12338);
or U19203 (N_19203,N_13010,N_12161);
nor U19204 (N_19204,N_12318,N_11203);
nand U19205 (N_19205,N_12865,N_10553);
nand U19206 (N_19206,N_13926,N_10616);
or U19207 (N_19207,N_14993,N_13204);
nand U19208 (N_19208,N_13556,N_10265);
nor U19209 (N_19209,N_12787,N_14905);
or U19210 (N_19210,N_10854,N_11398);
and U19211 (N_19211,N_12261,N_13409);
and U19212 (N_19212,N_14196,N_10752);
and U19213 (N_19213,N_11442,N_14074);
nor U19214 (N_19214,N_12169,N_12128);
nand U19215 (N_19215,N_12436,N_13330);
and U19216 (N_19216,N_14040,N_14317);
nand U19217 (N_19217,N_13980,N_11470);
and U19218 (N_19218,N_13983,N_10878);
nor U19219 (N_19219,N_12492,N_10144);
xor U19220 (N_19220,N_14355,N_11788);
xor U19221 (N_19221,N_10208,N_12653);
nor U19222 (N_19222,N_11798,N_10100);
nand U19223 (N_19223,N_10944,N_12061);
nand U19224 (N_19224,N_11183,N_11729);
or U19225 (N_19225,N_11665,N_11818);
nand U19226 (N_19226,N_14137,N_14314);
nand U19227 (N_19227,N_12190,N_13302);
and U19228 (N_19228,N_13974,N_11943);
or U19229 (N_19229,N_13770,N_11181);
xnor U19230 (N_19230,N_11297,N_10937);
or U19231 (N_19231,N_11308,N_14390);
nor U19232 (N_19232,N_14955,N_12149);
and U19233 (N_19233,N_14925,N_13860);
nand U19234 (N_19234,N_14830,N_10375);
xnor U19235 (N_19235,N_10385,N_13525);
or U19236 (N_19236,N_10797,N_11686);
nor U19237 (N_19237,N_14574,N_13985);
or U19238 (N_19238,N_12703,N_14732);
or U19239 (N_19239,N_13323,N_13703);
nor U19240 (N_19240,N_11055,N_14157);
xor U19241 (N_19241,N_12432,N_12057);
or U19242 (N_19242,N_13127,N_10648);
and U19243 (N_19243,N_14081,N_11760);
or U19244 (N_19244,N_12768,N_11826);
nor U19245 (N_19245,N_12934,N_13484);
and U19246 (N_19246,N_12400,N_13489);
nor U19247 (N_19247,N_11227,N_14880);
xnor U19248 (N_19248,N_12437,N_14565);
nand U19249 (N_19249,N_12326,N_14618);
nand U19250 (N_19250,N_13340,N_12199);
or U19251 (N_19251,N_10731,N_12168);
nand U19252 (N_19252,N_11115,N_12249);
nand U19253 (N_19253,N_12313,N_11563);
and U19254 (N_19254,N_12213,N_14758);
xor U19255 (N_19255,N_11839,N_12356);
nand U19256 (N_19256,N_13534,N_12735);
nor U19257 (N_19257,N_13096,N_11263);
nand U19258 (N_19258,N_11219,N_14368);
nand U19259 (N_19259,N_11062,N_14266);
or U19260 (N_19260,N_10859,N_11236);
and U19261 (N_19261,N_11449,N_10025);
nor U19262 (N_19262,N_11631,N_10894);
xor U19263 (N_19263,N_13469,N_13819);
xor U19264 (N_19264,N_13302,N_11009);
and U19265 (N_19265,N_11261,N_12904);
nor U19266 (N_19266,N_11837,N_12647);
nor U19267 (N_19267,N_14560,N_12809);
and U19268 (N_19268,N_13203,N_12806);
and U19269 (N_19269,N_10566,N_11391);
nand U19270 (N_19270,N_11693,N_14966);
nand U19271 (N_19271,N_10195,N_10223);
nor U19272 (N_19272,N_13306,N_12388);
xor U19273 (N_19273,N_10470,N_10375);
or U19274 (N_19274,N_10117,N_11411);
or U19275 (N_19275,N_13676,N_14576);
xor U19276 (N_19276,N_10103,N_14062);
nand U19277 (N_19277,N_14258,N_12608);
and U19278 (N_19278,N_12217,N_11124);
xor U19279 (N_19279,N_12351,N_14270);
xnor U19280 (N_19280,N_13532,N_10647);
xor U19281 (N_19281,N_11674,N_11586);
nor U19282 (N_19282,N_13328,N_11582);
and U19283 (N_19283,N_11196,N_10974);
nor U19284 (N_19284,N_10963,N_13376);
and U19285 (N_19285,N_12996,N_13366);
and U19286 (N_19286,N_14984,N_13462);
and U19287 (N_19287,N_11364,N_13712);
nor U19288 (N_19288,N_13939,N_10207);
and U19289 (N_19289,N_14118,N_12706);
xnor U19290 (N_19290,N_12203,N_10116);
xnor U19291 (N_19291,N_11369,N_11871);
and U19292 (N_19292,N_11744,N_10977);
nor U19293 (N_19293,N_10727,N_12070);
xor U19294 (N_19294,N_12150,N_13462);
nor U19295 (N_19295,N_11509,N_10001);
nor U19296 (N_19296,N_11803,N_12099);
nand U19297 (N_19297,N_13796,N_12421);
and U19298 (N_19298,N_11018,N_12484);
or U19299 (N_19299,N_13443,N_13192);
nand U19300 (N_19300,N_14797,N_14039);
nor U19301 (N_19301,N_10045,N_14981);
nand U19302 (N_19302,N_11652,N_12181);
and U19303 (N_19303,N_12733,N_12190);
nand U19304 (N_19304,N_10284,N_11086);
and U19305 (N_19305,N_14982,N_12132);
nor U19306 (N_19306,N_11844,N_14870);
nor U19307 (N_19307,N_13888,N_10115);
xor U19308 (N_19308,N_14066,N_13008);
or U19309 (N_19309,N_11156,N_10330);
and U19310 (N_19310,N_12493,N_14237);
nand U19311 (N_19311,N_10365,N_13512);
nor U19312 (N_19312,N_11529,N_14848);
or U19313 (N_19313,N_10334,N_10314);
and U19314 (N_19314,N_12287,N_12065);
nand U19315 (N_19315,N_12300,N_13904);
nand U19316 (N_19316,N_10358,N_14586);
and U19317 (N_19317,N_14134,N_14276);
xnor U19318 (N_19318,N_12805,N_12091);
and U19319 (N_19319,N_10686,N_10339);
nand U19320 (N_19320,N_11564,N_10207);
xnor U19321 (N_19321,N_10550,N_11489);
and U19322 (N_19322,N_13291,N_11466);
xor U19323 (N_19323,N_10503,N_13946);
and U19324 (N_19324,N_10681,N_10560);
or U19325 (N_19325,N_11201,N_14636);
and U19326 (N_19326,N_11251,N_13640);
or U19327 (N_19327,N_10745,N_13358);
and U19328 (N_19328,N_12091,N_10276);
or U19329 (N_19329,N_12931,N_12991);
xor U19330 (N_19330,N_11137,N_12808);
xor U19331 (N_19331,N_12773,N_10091);
or U19332 (N_19332,N_12119,N_14117);
and U19333 (N_19333,N_12907,N_13792);
and U19334 (N_19334,N_13879,N_13663);
xor U19335 (N_19335,N_12608,N_12584);
nor U19336 (N_19336,N_14419,N_12379);
nor U19337 (N_19337,N_11270,N_14961);
or U19338 (N_19338,N_10421,N_14879);
or U19339 (N_19339,N_13744,N_14448);
or U19340 (N_19340,N_10308,N_14519);
or U19341 (N_19341,N_13234,N_11413);
and U19342 (N_19342,N_10327,N_11472);
nand U19343 (N_19343,N_10408,N_10333);
xor U19344 (N_19344,N_12639,N_12899);
nand U19345 (N_19345,N_11785,N_11584);
nand U19346 (N_19346,N_12364,N_10737);
or U19347 (N_19347,N_10643,N_11147);
nor U19348 (N_19348,N_13558,N_13537);
nor U19349 (N_19349,N_10361,N_10939);
or U19350 (N_19350,N_13420,N_10152);
xnor U19351 (N_19351,N_12222,N_13726);
xnor U19352 (N_19352,N_11833,N_11674);
nand U19353 (N_19353,N_10422,N_12557);
xor U19354 (N_19354,N_11775,N_13566);
nor U19355 (N_19355,N_10434,N_12066);
and U19356 (N_19356,N_11461,N_14417);
nor U19357 (N_19357,N_12758,N_13557);
nor U19358 (N_19358,N_12471,N_10207);
and U19359 (N_19359,N_12955,N_10579);
or U19360 (N_19360,N_12635,N_11399);
nor U19361 (N_19361,N_10214,N_10643);
and U19362 (N_19362,N_11497,N_14121);
nand U19363 (N_19363,N_11488,N_12840);
xnor U19364 (N_19364,N_11580,N_13844);
nor U19365 (N_19365,N_11756,N_14438);
nand U19366 (N_19366,N_10665,N_10067);
nand U19367 (N_19367,N_14047,N_11825);
or U19368 (N_19368,N_13200,N_13164);
nor U19369 (N_19369,N_11054,N_14375);
or U19370 (N_19370,N_14028,N_10656);
xor U19371 (N_19371,N_13624,N_11713);
and U19372 (N_19372,N_14297,N_13897);
or U19373 (N_19373,N_12600,N_10252);
nand U19374 (N_19374,N_11646,N_13774);
and U19375 (N_19375,N_14896,N_13046);
or U19376 (N_19376,N_10455,N_13546);
or U19377 (N_19377,N_10905,N_14672);
and U19378 (N_19378,N_13006,N_13960);
nor U19379 (N_19379,N_14820,N_12564);
nand U19380 (N_19380,N_13829,N_10506);
xor U19381 (N_19381,N_10246,N_14259);
nor U19382 (N_19382,N_11886,N_10698);
or U19383 (N_19383,N_11721,N_14894);
and U19384 (N_19384,N_14893,N_12614);
or U19385 (N_19385,N_11715,N_11995);
xnor U19386 (N_19386,N_10855,N_10701);
nor U19387 (N_19387,N_12767,N_10817);
or U19388 (N_19388,N_12385,N_12347);
nand U19389 (N_19389,N_10737,N_13734);
nand U19390 (N_19390,N_11053,N_12597);
nand U19391 (N_19391,N_12365,N_12219);
nor U19392 (N_19392,N_14045,N_14173);
xor U19393 (N_19393,N_11190,N_10980);
nand U19394 (N_19394,N_14988,N_10929);
nand U19395 (N_19395,N_12421,N_13061);
nor U19396 (N_19396,N_11360,N_14323);
xnor U19397 (N_19397,N_10730,N_11008);
nand U19398 (N_19398,N_14226,N_11810);
and U19399 (N_19399,N_10084,N_12078);
nor U19400 (N_19400,N_13363,N_11169);
xnor U19401 (N_19401,N_13656,N_10540);
and U19402 (N_19402,N_10677,N_11398);
nor U19403 (N_19403,N_10202,N_11401);
nand U19404 (N_19404,N_10528,N_14667);
or U19405 (N_19405,N_13051,N_14015);
nor U19406 (N_19406,N_11623,N_11884);
and U19407 (N_19407,N_14751,N_13510);
nor U19408 (N_19408,N_12483,N_12235);
xnor U19409 (N_19409,N_11982,N_11080);
nand U19410 (N_19410,N_12523,N_13407);
nand U19411 (N_19411,N_10987,N_14689);
nor U19412 (N_19412,N_14690,N_12213);
and U19413 (N_19413,N_11225,N_12521);
and U19414 (N_19414,N_11937,N_10396);
or U19415 (N_19415,N_11133,N_10925);
xor U19416 (N_19416,N_14096,N_12780);
nor U19417 (N_19417,N_12926,N_12472);
nor U19418 (N_19418,N_10245,N_14988);
nand U19419 (N_19419,N_12744,N_10033);
xnor U19420 (N_19420,N_14938,N_14523);
or U19421 (N_19421,N_13666,N_13919);
or U19422 (N_19422,N_11464,N_11940);
and U19423 (N_19423,N_14895,N_10422);
xor U19424 (N_19424,N_14199,N_12731);
or U19425 (N_19425,N_11432,N_12343);
and U19426 (N_19426,N_12857,N_10036);
nor U19427 (N_19427,N_14655,N_12062);
nand U19428 (N_19428,N_11280,N_14793);
nand U19429 (N_19429,N_14100,N_11752);
and U19430 (N_19430,N_10299,N_13446);
nand U19431 (N_19431,N_10606,N_10130);
nand U19432 (N_19432,N_12373,N_14241);
and U19433 (N_19433,N_10769,N_11834);
or U19434 (N_19434,N_14804,N_11067);
xor U19435 (N_19435,N_14320,N_13721);
nand U19436 (N_19436,N_13280,N_11501);
nand U19437 (N_19437,N_12992,N_12633);
and U19438 (N_19438,N_12479,N_10781);
and U19439 (N_19439,N_10754,N_11592);
and U19440 (N_19440,N_14215,N_12466);
and U19441 (N_19441,N_11394,N_11684);
nor U19442 (N_19442,N_12182,N_13905);
xor U19443 (N_19443,N_13361,N_11971);
xnor U19444 (N_19444,N_10810,N_14810);
xnor U19445 (N_19445,N_14419,N_14979);
nand U19446 (N_19446,N_10693,N_10389);
nor U19447 (N_19447,N_13254,N_13732);
or U19448 (N_19448,N_13143,N_10331);
xor U19449 (N_19449,N_10964,N_12134);
xnor U19450 (N_19450,N_11296,N_12061);
or U19451 (N_19451,N_14810,N_13259);
nor U19452 (N_19452,N_13020,N_10595);
nor U19453 (N_19453,N_14497,N_14717);
nor U19454 (N_19454,N_11269,N_12635);
nor U19455 (N_19455,N_11860,N_10967);
xor U19456 (N_19456,N_11056,N_11833);
xor U19457 (N_19457,N_11730,N_14773);
xnor U19458 (N_19458,N_12552,N_11092);
nand U19459 (N_19459,N_10784,N_12045);
nand U19460 (N_19460,N_13177,N_11248);
nand U19461 (N_19461,N_13425,N_14728);
nand U19462 (N_19462,N_11312,N_10977);
xnor U19463 (N_19463,N_10328,N_12803);
and U19464 (N_19464,N_11863,N_13542);
or U19465 (N_19465,N_10487,N_12546);
and U19466 (N_19466,N_14721,N_10807);
or U19467 (N_19467,N_10149,N_13987);
nor U19468 (N_19468,N_11606,N_14846);
nand U19469 (N_19469,N_11635,N_11417);
nor U19470 (N_19470,N_12534,N_10636);
and U19471 (N_19471,N_14099,N_13458);
xor U19472 (N_19472,N_12140,N_12532);
and U19473 (N_19473,N_12416,N_10719);
and U19474 (N_19474,N_10664,N_11884);
xnor U19475 (N_19475,N_12780,N_10824);
xor U19476 (N_19476,N_10053,N_12302);
xor U19477 (N_19477,N_10906,N_13960);
nand U19478 (N_19478,N_13227,N_12719);
nor U19479 (N_19479,N_12839,N_11228);
and U19480 (N_19480,N_13863,N_13853);
nor U19481 (N_19481,N_11132,N_11795);
nand U19482 (N_19482,N_10230,N_12076);
nand U19483 (N_19483,N_10554,N_14001);
or U19484 (N_19484,N_14118,N_12419);
nand U19485 (N_19485,N_12633,N_10166);
nand U19486 (N_19486,N_13334,N_12826);
xnor U19487 (N_19487,N_10242,N_10034);
and U19488 (N_19488,N_14813,N_11335);
or U19489 (N_19489,N_14626,N_11392);
or U19490 (N_19490,N_14395,N_13552);
or U19491 (N_19491,N_13148,N_14209);
xnor U19492 (N_19492,N_13680,N_13790);
and U19493 (N_19493,N_12513,N_10336);
xnor U19494 (N_19494,N_10446,N_13879);
or U19495 (N_19495,N_10515,N_13418);
xnor U19496 (N_19496,N_11833,N_12634);
or U19497 (N_19497,N_11143,N_13347);
nand U19498 (N_19498,N_13220,N_11199);
and U19499 (N_19499,N_12766,N_10549);
xnor U19500 (N_19500,N_13196,N_10686);
or U19501 (N_19501,N_13904,N_14754);
xnor U19502 (N_19502,N_14818,N_11995);
xnor U19503 (N_19503,N_12115,N_10249);
nor U19504 (N_19504,N_11668,N_10103);
nor U19505 (N_19505,N_13507,N_12540);
nor U19506 (N_19506,N_11430,N_12814);
nand U19507 (N_19507,N_14042,N_11053);
nand U19508 (N_19508,N_12001,N_13328);
nand U19509 (N_19509,N_14868,N_12645);
xor U19510 (N_19510,N_11393,N_14837);
nand U19511 (N_19511,N_14245,N_12030);
and U19512 (N_19512,N_14088,N_10518);
xnor U19513 (N_19513,N_12576,N_14013);
or U19514 (N_19514,N_14759,N_14023);
or U19515 (N_19515,N_13848,N_12436);
xor U19516 (N_19516,N_13407,N_12262);
nand U19517 (N_19517,N_13555,N_14558);
and U19518 (N_19518,N_12465,N_10713);
xor U19519 (N_19519,N_10186,N_12258);
or U19520 (N_19520,N_14440,N_13732);
nor U19521 (N_19521,N_11160,N_12145);
and U19522 (N_19522,N_14618,N_14907);
nor U19523 (N_19523,N_10318,N_11236);
nand U19524 (N_19524,N_12763,N_10344);
xnor U19525 (N_19525,N_10749,N_13442);
nand U19526 (N_19526,N_14392,N_13566);
and U19527 (N_19527,N_10876,N_13421);
xor U19528 (N_19528,N_12329,N_13660);
and U19529 (N_19529,N_11762,N_13110);
xor U19530 (N_19530,N_12054,N_14533);
xor U19531 (N_19531,N_14320,N_13307);
or U19532 (N_19532,N_13122,N_10620);
or U19533 (N_19533,N_12651,N_13993);
nand U19534 (N_19534,N_10322,N_12390);
nand U19535 (N_19535,N_12549,N_10365);
or U19536 (N_19536,N_10289,N_14585);
or U19537 (N_19537,N_10631,N_12863);
xnor U19538 (N_19538,N_12780,N_12124);
or U19539 (N_19539,N_10461,N_10578);
xnor U19540 (N_19540,N_11338,N_10240);
and U19541 (N_19541,N_13461,N_14451);
nand U19542 (N_19542,N_11389,N_10035);
xor U19543 (N_19543,N_12877,N_10952);
nor U19544 (N_19544,N_14309,N_13869);
or U19545 (N_19545,N_12948,N_14330);
nor U19546 (N_19546,N_11315,N_10024);
xor U19547 (N_19547,N_11284,N_13203);
xor U19548 (N_19548,N_10103,N_13873);
nand U19549 (N_19549,N_11452,N_14640);
and U19550 (N_19550,N_12456,N_10973);
nand U19551 (N_19551,N_10863,N_14959);
nor U19552 (N_19552,N_13470,N_11082);
or U19553 (N_19553,N_13969,N_10492);
xnor U19554 (N_19554,N_13697,N_14867);
xor U19555 (N_19555,N_10876,N_14245);
and U19556 (N_19556,N_11250,N_12317);
nand U19557 (N_19557,N_12905,N_11341);
nand U19558 (N_19558,N_14396,N_12181);
xnor U19559 (N_19559,N_12973,N_10458);
xnor U19560 (N_19560,N_11317,N_10830);
and U19561 (N_19561,N_11223,N_13058);
xnor U19562 (N_19562,N_11380,N_13803);
xor U19563 (N_19563,N_10475,N_13769);
xor U19564 (N_19564,N_10981,N_12098);
and U19565 (N_19565,N_12347,N_13094);
nor U19566 (N_19566,N_10230,N_12290);
nor U19567 (N_19567,N_10911,N_10033);
nor U19568 (N_19568,N_10908,N_14931);
xor U19569 (N_19569,N_14670,N_10289);
or U19570 (N_19570,N_12235,N_11925);
and U19571 (N_19571,N_12642,N_12388);
or U19572 (N_19572,N_14468,N_13590);
and U19573 (N_19573,N_13882,N_11312);
nor U19574 (N_19574,N_12231,N_11952);
and U19575 (N_19575,N_12218,N_10921);
or U19576 (N_19576,N_13774,N_13230);
nand U19577 (N_19577,N_12185,N_14025);
or U19578 (N_19578,N_14867,N_14959);
and U19579 (N_19579,N_10031,N_13434);
nor U19580 (N_19580,N_14155,N_14141);
or U19581 (N_19581,N_10106,N_11046);
and U19582 (N_19582,N_10418,N_14640);
xor U19583 (N_19583,N_14876,N_12544);
or U19584 (N_19584,N_11334,N_10294);
xnor U19585 (N_19585,N_11901,N_10452);
nor U19586 (N_19586,N_12886,N_11809);
or U19587 (N_19587,N_14542,N_11901);
nand U19588 (N_19588,N_13061,N_13930);
and U19589 (N_19589,N_11655,N_13526);
nand U19590 (N_19590,N_13868,N_12295);
nor U19591 (N_19591,N_11913,N_13594);
or U19592 (N_19592,N_13163,N_11284);
nor U19593 (N_19593,N_14934,N_12946);
xor U19594 (N_19594,N_14467,N_11238);
nand U19595 (N_19595,N_10204,N_11477);
nand U19596 (N_19596,N_11677,N_14344);
and U19597 (N_19597,N_14984,N_10675);
xor U19598 (N_19598,N_12995,N_13323);
nor U19599 (N_19599,N_13668,N_13602);
xor U19600 (N_19600,N_14551,N_14956);
nand U19601 (N_19601,N_10380,N_11186);
xor U19602 (N_19602,N_14998,N_10322);
nor U19603 (N_19603,N_13721,N_10839);
and U19604 (N_19604,N_11550,N_12391);
or U19605 (N_19605,N_11342,N_14686);
nor U19606 (N_19606,N_13312,N_11347);
or U19607 (N_19607,N_10960,N_13094);
and U19608 (N_19608,N_11319,N_11985);
xor U19609 (N_19609,N_10536,N_12274);
xnor U19610 (N_19610,N_10383,N_11519);
or U19611 (N_19611,N_13809,N_13718);
nor U19612 (N_19612,N_11416,N_10658);
nand U19613 (N_19613,N_14098,N_14264);
xor U19614 (N_19614,N_10733,N_10330);
and U19615 (N_19615,N_10475,N_14388);
or U19616 (N_19616,N_12678,N_12101);
xor U19617 (N_19617,N_14040,N_14930);
xnor U19618 (N_19618,N_12870,N_11693);
nand U19619 (N_19619,N_11155,N_10597);
xor U19620 (N_19620,N_11708,N_13413);
and U19621 (N_19621,N_14077,N_13138);
xor U19622 (N_19622,N_12690,N_12673);
nor U19623 (N_19623,N_14285,N_14221);
nand U19624 (N_19624,N_13612,N_14275);
or U19625 (N_19625,N_11857,N_11139);
xor U19626 (N_19626,N_14702,N_14908);
xor U19627 (N_19627,N_13713,N_12462);
or U19628 (N_19628,N_12304,N_11820);
nand U19629 (N_19629,N_10860,N_12812);
or U19630 (N_19630,N_14739,N_13408);
and U19631 (N_19631,N_14206,N_11025);
or U19632 (N_19632,N_13065,N_11002);
nor U19633 (N_19633,N_13964,N_10917);
nor U19634 (N_19634,N_14020,N_10328);
xnor U19635 (N_19635,N_14847,N_13851);
nand U19636 (N_19636,N_14341,N_10610);
and U19637 (N_19637,N_14723,N_10179);
nor U19638 (N_19638,N_10050,N_10727);
and U19639 (N_19639,N_14029,N_14673);
xor U19640 (N_19640,N_13339,N_13242);
or U19641 (N_19641,N_13017,N_13163);
xor U19642 (N_19642,N_10065,N_11171);
nor U19643 (N_19643,N_11079,N_11603);
nor U19644 (N_19644,N_12397,N_10765);
and U19645 (N_19645,N_10943,N_14816);
or U19646 (N_19646,N_14419,N_10402);
nand U19647 (N_19647,N_13499,N_12119);
or U19648 (N_19648,N_12546,N_13295);
or U19649 (N_19649,N_14588,N_11935);
xnor U19650 (N_19650,N_11095,N_11242);
and U19651 (N_19651,N_14803,N_14259);
and U19652 (N_19652,N_10325,N_14129);
and U19653 (N_19653,N_13122,N_12362);
and U19654 (N_19654,N_13080,N_14444);
xnor U19655 (N_19655,N_13619,N_10811);
nand U19656 (N_19656,N_10106,N_13050);
or U19657 (N_19657,N_11380,N_14878);
or U19658 (N_19658,N_10566,N_12515);
nand U19659 (N_19659,N_12316,N_13465);
nor U19660 (N_19660,N_12073,N_11896);
nand U19661 (N_19661,N_13704,N_12001);
nor U19662 (N_19662,N_10707,N_12131);
xor U19663 (N_19663,N_10874,N_14851);
or U19664 (N_19664,N_12641,N_14950);
nor U19665 (N_19665,N_10973,N_10930);
and U19666 (N_19666,N_12511,N_11452);
and U19667 (N_19667,N_14086,N_14754);
and U19668 (N_19668,N_13283,N_14604);
xnor U19669 (N_19669,N_13785,N_10340);
nor U19670 (N_19670,N_10255,N_13508);
xnor U19671 (N_19671,N_12883,N_11657);
xnor U19672 (N_19672,N_12870,N_11363);
or U19673 (N_19673,N_13048,N_10390);
xnor U19674 (N_19674,N_11029,N_14831);
nand U19675 (N_19675,N_13216,N_10900);
or U19676 (N_19676,N_13325,N_10627);
or U19677 (N_19677,N_13714,N_12910);
nand U19678 (N_19678,N_14547,N_11331);
and U19679 (N_19679,N_11508,N_11728);
nor U19680 (N_19680,N_13729,N_11140);
nand U19681 (N_19681,N_14010,N_10887);
xnor U19682 (N_19682,N_13942,N_14513);
xor U19683 (N_19683,N_11062,N_12345);
nor U19684 (N_19684,N_11652,N_11611);
and U19685 (N_19685,N_10629,N_14426);
nand U19686 (N_19686,N_14203,N_14370);
nor U19687 (N_19687,N_10768,N_12787);
nand U19688 (N_19688,N_10565,N_10536);
nand U19689 (N_19689,N_12131,N_11937);
nor U19690 (N_19690,N_11444,N_12749);
nand U19691 (N_19691,N_13217,N_12490);
and U19692 (N_19692,N_10692,N_11996);
or U19693 (N_19693,N_11060,N_10673);
or U19694 (N_19694,N_12444,N_13512);
or U19695 (N_19695,N_12308,N_14200);
and U19696 (N_19696,N_11006,N_13383);
or U19697 (N_19697,N_11773,N_10816);
and U19698 (N_19698,N_11589,N_12898);
nor U19699 (N_19699,N_14139,N_11841);
nand U19700 (N_19700,N_12886,N_14096);
nor U19701 (N_19701,N_11125,N_13703);
xnor U19702 (N_19702,N_14179,N_10864);
and U19703 (N_19703,N_11650,N_13912);
xnor U19704 (N_19704,N_12817,N_12652);
or U19705 (N_19705,N_12499,N_14737);
and U19706 (N_19706,N_13133,N_10754);
or U19707 (N_19707,N_11649,N_10573);
nor U19708 (N_19708,N_11298,N_11553);
and U19709 (N_19709,N_14804,N_14813);
nor U19710 (N_19710,N_11289,N_11816);
nand U19711 (N_19711,N_13097,N_13583);
and U19712 (N_19712,N_14144,N_11281);
nor U19713 (N_19713,N_10187,N_11712);
and U19714 (N_19714,N_10118,N_14020);
nand U19715 (N_19715,N_11654,N_11374);
nand U19716 (N_19716,N_13876,N_11318);
or U19717 (N_19717,N_13629,N_10893);
xor U19718 (N_19718,N_10707,N_12192);
or U19719 (N_19719,N_14306,N_12839);
and U19720 (N_19720,N_11638,N_10624);
or U19721 (N_19721,N_13329,N_13455);
or U19722 (N_19722,N_12043,N_13202);
nor U19723 (N_19723,N_12460,N_12002);
or U19724 (N_19724,N_10117,N_11241);
nor U19725 (N_19725,N_10317,N_12711);
nand U19726 (N_19726,N_13081,N_13205);
nand U19727 (N_19727,N_12106,N_10471);
and U19728 (N_19728,N_10219,N_10531);
and U19729 (N_19729,N_13834,N_12739);
and U19730 (N_19730,N_14840,N_12794);
or U19731 (N_19731,N_11153,N_14382);
or U19732 (N_19732,N_12409,N_13007);
or U19733 (N_19733,N_11973,N_14311);
or U19734 (N_19734,N_11880,N_11791);
nand U19735 (N_19735,N_10480,N_10926);
or U19736 (N_19736,N_11957,N_10601);
or U19737 (N_19737,N_12760,N_12673);
nor U19738 (N_19738,N_11994,N_13698);
and U19739 (N_19739,N_11989,N_14097);
and U19740 (N_19740,N_14374,N_13042);
nand U19741 (N_19741,N_13466,N_14693);
nor U19742 (N_19742,N_12178,N_14495);
nand U19743 (N_19743,N_11552,N_12473);
and U19744 (N_19744,N_11187,N_11774);
nand U19745 (N_19745,N_10766,N_12844);
xor U19746 (N_19746,N_14502,N_14332);
xor U19747 (N_19747,N_11814,N_10281);
xnor U19748 (N_19748,N_13626,N_14148);
or U19749 (N_19749,N_14864,N_12580);
and U19750 (N_19750,N_12595,N_10863);
nand U19751 (N_19751,N_10271,N_13797);
or U19752 (N_19752,N_14476,N_11624);
xor U19753 (N_19753,N_13726,N_11888);
xnor U19754 (N_19754,N_12179,N_11597);
xor U19755 (N_19755,N_10039,N_14369);
nand U19756 (N_19756,N_12661,N_14372);
nand U19757 (N_19757,N_11382,N_10651);
nor U19758 (N_19758,N_12987,N_13243);
or U19759 (N_19759,N_10556,N_12521);
or U19760 (N_19760,N_10324,N_10331);
nand U19761 (N_19761,N_12799,N_14374);
nor U19762 (N_19762,N_11206,N_10930);
xnor U19763 (N_19763,N_11267,N_11113);
nor U19764 (N_19764,N_10948,N_11878);
xor U19765 (N_19765,N_12221,N_10742);
and U19766 (N_19766,N_10450,N_14990);
or U19767 (N_19767,N_12579,N_10896);
and U19768 (N_19768,N_13224,N_12251);
nor U19769 (N_19769,N_14702,N_11243);
nor U19770 (N_19770,N_13481,N_14098);
nor U19771 (N_19771,N_14850,N_13859);
xor U19772 (N_19772,N_13098,N_14538);
and U19773 (N_19773,N_10782,N_13774);
nor U19774 (N_19774,N_14473,N_13150);
nand U19775 (N_19775,N_14046,N_10079);
or U19776 (N_19776,N_13576,N_10941);
nand U19777 (N_19777,N_13451,N_11382);
nand U19778 (N_19778,N_10604,N_14537);
and U19779 (N_19779,N_12085,N_13161);
or U19780 (N_19780,N_14958,N_11511);
xor U19781 (N_19781,N_10010,N_11251);
or U19782 (N_19782,N_11764,N_13297);
nor U19783 (N_19783,N_14225,N_13226);
or U19784 (N_19784,N_12445,N_14868);
and U19785 (N_19785,N_10853,N_11476);
nor U19786 (N_19786,N_14191,N_12406);
or U19787 (N_19787,N_10428,N_10726);
xnor U19788 (N_19788,N_13940,N_10525);
nor U19789 (N_19789,N_10222,N_11402);
and U19790 (N_19790,N_10037,N_14241);
nand U19791 (N_19791,N_14504,N_14975);
nand U19792 (N_19792,N_12224,N_14498);
xor U19793 (N_19793,N_14717,N_10861);
or U19794 (N_19794,N_12323,N_13306);
and U19795 (N_19795,N_11643,N_13523);
or U19796 (N_19796,N_12935,N_10730);
nand U19797 (N_19797,N_11880,N_13524);
nor U19798 (N_19798,N_14877,N_14026);
and U19799 (N_19799,N_10316,N_13990);
and U19800 (N_19800,N_14493,N_11239);
nor U19801 (N_19801,N_10282,N_12729);
xnor U19802 (N_19802,N_14762,N_13588);
nand U19803 (N_19803,N_13200,N_10598);
nor U19804 (N_19804,N_12701,N_10404);
xnor U19805 (N_19805,N_10361,N_14413);
or U19806 (N_19806,N_13960,N_10785);
nor U19807 (N_19807,N_12947,N_14873);
nand U19808 (N_19808,N_10222,N_10338);
nand U19809 (N_19809,N_12094,N_13935);
or U19810 (N_19810,N_13031,N_12393);
xnor U19811 (N_19811,N_11083,N_11060);
and U19812 (N_19812,N_10372,N_13325);
xnor U19813 (N_19813,N_13058,N_13558);
xor U19814 (N_19814,N_13341,N_14266);
xnor U19815 (N_19815,N_12866,N_14371);
nand U19816 (N_19816,N_14156,N_12784);
or U19817 (N_19817,N_12425,N_13570);
nand U19818 (N_19818,N_10792,N_10221);
nand U19819 (N_19819,N_14676,N_11789);
and U19820 (N_19820,N_10941,N_14402);
and U19821 (N_19821,N_14392,N_14255);
or U19822 (N_19822,N_10994,N_13787);
nand U19823 (N_19823,N_11265,N_13222);
nand U19824 (N_19824,N_12515,N_10152);
or U19825 (N_19825,N_14603,N_13055);
or U19826 (N_19826,N_14437,N_14230);
nand U19827 (N_19827,N_14498,N_13964);
and U19828 (N_19828,N_14566,N_13792);
nand U19829 (N_19829,N_11220,N_11164);
or U19830 (N_19830,N_12732,N_14140);
xor U19831 (N_19831,N_12554,N_11900);
or U19832 (N_19832,N_12270,N_12404);
nand U19833 (N_19833,N_10269,N_14065);
nand U19834 (N_19834,N_12328,N_13080);
nand U19835 (N_19835,N_13188,N_11379);
nor U19836 (N_19836,N_10717,N_10939);
and U19837 (N_19837,N_11460,N_13504);
nor U19838 (N_19838,N_12465,N_14749);
xor U19839 (N_19839,N_13183,N_10470);
nand U19840 (N_19840,N_12626,N_11096);
xor U19841 (N_19841,N_14806,N_14864);
nand U19842 (N_19842,N_12951,N_14354);
nor U19843 (N_19843,N_14163,N_12025);
and U19844 (N_19844,N_11764,N_14656);
or U19845 (N_19845,N_13959,N_10972);
xor U19846 (N_19846,N_11056,N_11018);
or U19847 (N_19847,N_12935,N_14630);
and U19848 (N_19848,N_13328,N_12772);
and U19849 (N_19849,N_12434,N_11773);
nor U19850 (N_19850,N_11306,N_14871);
nand U19851 (N_19851,N_13126,N_12875);
or U19852 (N_19852,N_10233,N_14470);
and U19853 (N_19853,N_14110,N_13698);
xnor U19854 (N_19854,N_10675,N_14199);
nor U19855 (N_19855,N_10853,N_13917);
or U19856 (N_19856,N_10918,N_14244);
and U19857 (N_19857,N_14031,N_11406);
and U19858 (N_19858,N_10296,N_14601);
nor U19859 (N_19859,N_12477,N_13056);
or U19860 (N_19860,N_11892,N_11390);
nand U19861 (N_19861,N_12074,N_14190);
and U19862 (N_19862,N_14600,N_10553);
and U19863 (N_19863,N_12434,N_10948);
or U19864 (N_19864,N_10668,N_10276);
xor U19865 (N_19865,N_13709,N_12370);
nand U19866 (N_19866,N_12534,N_13015);
or U19867 (N_19867,N_11153,N_10282);
nor U19868 (N_19868,N_14181,N_10514);
nor U19869 (N_19869,N_13320,N_10897);
or U19870 (N_19870,N_10466,N_12130);
nor U19871 (N_19871,N_13876,N_10747);
nor U19872 (N_19872,N_10366,N_13381);
or U19873 (N_19873,N_14147,N_13560);
or U19874 (N_19874,N_14797,N_14758);
nor U19875 (N_19875,N_12480,N_11794);
nor U19876 (N_19876,N_12152,N_10786);
nor U19877 (N_19877,N_11926,N_14519);
and U19878 (N_19878,N_13712,N_12928);
xnor U19879 (N_19879,N_14157,N_13307);
nand U19880 (N_19880,N_12857,N_14795);
xor U19881 (N_19881,N_14762,N_13160);
and U19882 (N_19882,N_11426,N_14431);
and U19883 (N_19883,N_14023,N_10138);
xor U19884 (N_19884,N_14870,N_10725);
or U19885 (N_19885,N_10486,N_14362);
nor U19886 (N_19886,N_13091,N_12736);
xor U19887 (N_19887,N_14290,N_10204);
or U19888 (N_19888,N_12219,N_11761);
nand U19889 (N_19889,N_10845,N_13930);
nor U19890 (N_19890,N_11070,N_14968);
nor U19891 (N_19891,N_11879,N_12795);
xor U19892 (N_19892,N_14305,N_10794);
nand U19893 (N_19893,N_13144,N_14146);
nand U19894 (N_19894,N_14687,N_10284);
nor U19895 (N_19895,N_14760,N_14698);
xnor U19896 (N_19896,N_12858,N_11288);
xor U19897 (N_19897,N_13519,N_13058);
and U19898 (N_19898,N_14704,N_12041);
nand U19899 (N_19899,N_14174,N_10407);
nand U19900 (N_19900,N_12830,N_13410);
nand U19901 (N_19901,N_11727,N_10559);
nor U19902 (N_19902,N_11905,N_11854);
or U19903 (N_19903,N_10364,N_14169);
nand U19904 (N_19904,N_14069,N_13551);
and U19905 (N_19905,N_13274,N_14990);
and U19906 (N_19906,N_12895,N_10044);
or U19907 (N_19907,N_12138,N_11986);
nor U19908 (N_19908,N_12077,N_13209);
xnor U19909 (N_19909,N_11809,N_14141);
nand U19910 (N_19910,N_10693,N_13111);
or U19911 (N_19911,N_13779,N_10448);
xor U19912 (N_19912,N_10871,N_11645);
xnor U19913 (N_19913,N_14784,N_14824);
and U19914 (N_19914,N_12916,N_10744);
or U19915 (N_19915,N_13157,N_14159);
nand U19916 (N_19916,N_13982,N_14516);
nand U19917 (N_19917,N_11037,N_12882);
xnor U19918 (N_19918,N_14231,N_11073);
or U19919 (N_19919,N_14842,N_10636);
nor U19920 (N_19920,N_12512,N_11648);
nand U19921 (N_19921,N_11130,N_11181);
nor U19922 (N_19922,N_13183,N_12535);
nor U19923 (N_19923,N_13147,N_13683);
or U19924 (N_19924,N_14658,N_14317);
or U19925 (N_19925,N_12052,N_10805);
and U19926 (N_19926,N_10552,N_13279);
nor U19927 (N_19927,N_10430,N_10090);
xnor U19928 (N_19928,N_11086,N_11324);
and U19929 (N_19929,N_12294,N_10603);
xor U19930 (N_19930,N_13361,N_13884);
and U19931 (N_19931,N_11704,N_10246);
and U19932 (N_19932,N_14406,N_12073);
or U19933 (N_19933,N_13096,N_14125);
nand U19934 (N_19934,N_10997,N_10243);
or U19935 (N_19935,N_11457,N_11473);
xor U19936 (N_19936,N_12645,N_13138);
xnor U19937 (N_19937,N_13234,N_14112);
nand U19938 (N_19938,N_10525,N_10761);
and U19939 (N_19939,N_12437,N_14369);
nand U19940 (N_19940,N_12817,N_12273);
nand U19941 (N_19941,N_14799,N_10420);
xnor U19942 (N_19942,N_10723,N_13489);
or U19943 (N_19943,N_14009,N_12552);
xor U19944 (N_19944,N_10508,N_11127);
and U19945 (N_19945,N_13495,N_10190);
nand U19946 (N_19946,N_13216,N_10925);
and U19947 (N_19947,N_10230,N_14066);
nor U19948 (N_19948,N_14960,N_13695);
xor U19949 (N_19949,N_11700,N_12133);
nor U19950 (N_19950,N_13935,N_10690);
nor U19951 (N_19951,N_11483,N_13756);
nand U19952 (N_19952,N_11913,N_11706);
xor U19953 (N_19953,N_13675,N_12178);
nand U19954 (N_19954,N_13605,N_13255);
xor U19955 (N_19955,N_11468,N_14918);
nand U19956 (N_19956,N_13569,N_11543);
and U19957 (N_19957,N_14295,N_10050);
or U19958 (N_19958,N_13707,N_14362);
and U19959 (N_19959,N_10734,N_14767);
and U19960 (N_19960,N_14844,N_12401);
or U19961 (N_19961,N_12449,N_13687);
xor U19962 (N_19962,N_12477,N_12940);
xor U19963 (N_19963,N_10373,N_12605);
xor U19964 (N_19964,N_13285,N_14456);
xnor U19965 (N_19965,N_14282,N_13565);
nand U19966 (N_19966,N_11622,N_13253);
and U19967 (N_19967,N_13093,N_14961);
nor U19968 (N_19968,N_13818,N_11938);
nor U19969 (N_19969,N_13848,N_10899);
or U19970 (N_19970,N_13440,N_12906);
xor U19971 (N_19971,N_12510,N_13620);
xnor U19972 (N_19972,N_11627,N_12306);
or U19973 (N_19973,N_11943,N_11109);
xnor U19974 (N_19974,N_13969,N_13057);
xnor U19975 (N_19975,N_11061,N_12173);
and U19976 (N_19976,N_11097,N_13299);
or U19977 (N_19977,N_13041,N_14198);
nor U19978 (N_19978,N_14208,N_11678);
and U19979 (N_19979,N_13667,N_11394);
and U19980 (N_19980,N_12338,N_12823);
or U19981 (N_19981,N_14034,N_13458);
nand U19982 (N_19982,N_13052,N_12165);
nor U19983 (N_19983,N_11764,N_13180);
and U19984 (N_19984,N_14432,N_12083);
xor U19985 (N_19985,N_10093,N_10698);
and U19986 (N_19986,N_13915,N_14824);
and U19987 (N_19987,N_12367,N_11838);
or U19988 (N_19988,N_13473,N_14263);
and U19989 (N_19989,N_11432,N_13997);
or U19990 (N_19990,N_12526,N_12295);
or U19991 (N_19991,N_10304,N_12090);
nor U19992 (N_19992,N_14846,N_10269);
or U19993 (N_19993,N_11295,N_10993);
nor U19994 (N_19994,N_12902,N_10141);
and U19995 (N_19995,N_12143,N_10210);
or U19996 (N_19996,N_13508,N_11005);
nand U19997 (N_19997,N_10369,N_11200);
xnor U19998 (N_19998,N_13348,N_12230);
or U19999 (N_19999,N_10182,N_13675);
and U20000 (N_20000,N_15267,N_15001);
or U20001 (N_20001,N_16202,N_15137);
nand U20002 (N_20002,N_15477,N_16181);
nand U20003 (N_20003,N_18836,N_16365);
xor U20004 (N_20004,N_17894,N_19086);
and U20005 (N_20005,N_17769,N_18464);
xor U20006 (N_20006,N_16186,N_17158);
and U20007 (N_20007,N_16423,N_19710);
and U20008 (N_20008,N_19879,N_16306);
nand U20009 (N_20009,N_17658,N_17906);
or U20010 (N_20010,N_19126,N_19929);
and U20011 (N_20011,N_18174,N_17618);
or U20012 (N_20012,N_17100,N_16744);
nand U20013 (N_20013,N_15718,N_19186);
xor U20014 (N_20014,N_16161,N_18095);
nand U20015 (N_20015,N_19627,N_17346);
xor U20016 (N_20016,N_15869,N_19258);
nor U20017 (N_20017,N_18722,N_17814);
nor U20018 (N_20018,N_17675,N_17933);
xnor U20019 (N_20019,N_17930,N_18092);
nor U20020 (N_20020,N_15060,N_17430);
nor U20021 (N_20021,N_19550,N_19094);
xor U20022 (N_20022,N_18142,N_16973);
and U20023 (N_20023,N_19776,N_15032);
nor U20024 (N_20024,N_15812,N_15949);
and U20025 (N_20025,N_16840,N_19051);
and U20026 (N_20026,N_15849,N_19592);
nor U20027 (N_20027,N_16948,N_19682);
and U20028 (N_20028,N_19208,N_17680);
nor U20029 (N_20029,N_19343,N_18735);
and U20030 (N_20030,N_15094,N_18505);
and U20031 (N_20031,N_18356,N_17195);
nand U20032 (N_20032,N_19523,N_18377);
or U20033 (N_20033,N_15815,N_18892);
and U20034 (N_20034,N_17247,N_17535);
nand U20035 (N_20035,N_17795,N_19254);
nand U20036 (N_20036,N_16382,N_19031);
and U20037 (N_20037,N_18342,N_15454);
xor U20038 (N_20038,N_16061,N_19000);
or U20039 (N_20039,N_17156,N_15133);
or U20040 (N_20040,N_15028,N_17250);
and U20041 (N_20041,N_19836,N_18711);
nor U20042 (N_20042,N_15316,N_16733);
and U20043 (N_20043,N_18762,N_16248);
xor U20044 (N_20044,N_17077,N_17687);
nor U20045 (N_20045,N_18900,N_18153);
nand U20046 (N_20046,N_19350,N_18058);
nand U20047 (N_20047,N_16172,N_18015);
xnor U20048 (N_20048,N_15994,N_17827);
and U20049 (N_20049,N_17872,N_18164);
or U20050 (N_20050,N_15836,N_19146);
nor U20051 (N_20051,N_19464,N_19145);
nor U20052 (N_20052,N_15546,N_15455);
xor U20053 (N_20053,N_17556,N_16588);
and U20054 (N_20054,N_18558,N_16038);
nor U20055 (N_20055,N_18929,N_16045);
nor U20056 (N_20056,N_16338,N_19573);
and U20057 (N_20057,N_17537,N_16701);
nand U20058 (N_20058,N_18828,N_17673);
nand U20059 (N_20059,N_15225,N_16342);
nand U20060 (N_20060,N_15453,N_16796);
xnor U20061 (N_20061,N_17981,N_16768);
nor U20062 (N_20062,N_16516,N_19124);
nand U20063 (N_20063,N_17748,N_19590);
nand U20064 (N_20064,N_17938,N_18884);
or U20065 (N_20065,N_17108,N_16280);
xnor U20066 (N_20066,N_16138,N_15073);
nor U20067 (N_20067,N_17330,N_17541);
or U20068 (N_20068,N_17759,N_16039);
nand U20069 (N_20069,N_16228,N_19117);
nand U20070 (N_20070,N_16509,N_17649);
or U20071 (N_20071,N_16388,N_19794);
nor U20072 (N_20072,N_18849,N_19948);
or U20073 (N_20073,N_15369,N_17338);
and U20074 (N_20074,N_15261,N_15727);
nor U20075 (N_20075,N_16513,N_15941);
nor U20076 (N_20076,N_17820,N_18835);
xor U20077 (N_20077,N_15173,N_19452);
nor U20078 (N_20078,N_18056,N_19528);
xnor U20079 (N_20079,N_15750,N_16488);
xor U20080 (N_20080,N_16400,N_15380);
and U20081 (N_20081,N_18724,N_16854);
nor U20082 (N_20082,N_18120,N_19930);
nand U20083 (N_20083,N_19974,N_17481);
and U20084 (N_20084,N_17390,N_16308);
nand U20085 (N_20085,N_15731,N_15931);
and U20086 (N_20086,N_19395,N_18664);
nor U20087 (N_20087,N_19058,N_18500);
xnor U20088 (N_20088,N_19656,N_18380);
or U20089 (N_20089,N_16037,N_18732);
xor U20090 (N_20090,N_16372,N_18744);
and U20091 (N_20091,N_16902,N_16102);
and U20092 (N_20092,N_16072,N_17695);
nor U20093 (N_20093,N_19471,N_17813);
nand U20094 (N_20094,N_16587,N_16196);
or U20095 (N_20095,N_19845,N_16195);
nand U20096 (N_20096,N_19808,N_15273);
or U20097 (N_20097,N_17446,N_19064);
or U20098 (N_20098,N_19455,N_18277);
nand U20099 (N_20099,N_15648,N_19993);
or U20100 (N_20100,N_17187,N_18230);
nor U20101 (N_20101,N_17357,N_18879);
nand U20102 (N_20102,N_15395,N_18938);
xnor U20103 (N_20103,N_16297,N_19480);
and U20104 (N_20104,N_19147,N_18333);
xnor U20105 (N_20105,N_18738,N_16781);
and U20106 (N_20106,N_17320,N_17552);
and U20107 (N_20107,N_15431,N_19504);
nand U20108 (N_20108,N_15972,N_15515);
xor U20109 (N_20109,N_17178,N_15258);
or U20110 (N_20110,N_15697,N_17570);
nor U20111 (N_20111,N_18872,N_15639);
nor U20112 (N_20112,N_16511,N_17788);
nor U20113 (N_20113,N_19494,N_18287);
xnor U20114 (N_20114,N_16101,N_19221);
nand U20115 (N_20115,N_19894,N_18376);
nand U20116 (N_20116,N_15976,N_18680);
nor U20117 (N_20117,N_17878,N_17644);
and U20118 (N_20118,N_15699,N_18981);
xor U20119 (N_20119,N_19474,N_18031);
nand U20120 (N_20120,N_18317,N_19834);
and U20121 (N_20121,N_16237,N_17198);
or U20122 (N_20122,N_18456,N_16075);
or U20123 (N_20123,N_15097,N_17163);
nand U20124 (N_20124,N_15143,N_16932);
nor U20125 (N_20125,N_16950,N_17661);
nand U20126 (N_20126,N_17309,N_15356);
xnor U20127 (N_20127,N_19493,N_19330);
and U20128 (N_20128,N_17274,N_17251);
xor U20129 (N_20129,N_16491,N_19373);
and U20130 (N_20130,N_17116,N_19810);
nor U20131 (N_20131,N_18304,N_17278);
xor U20132 (N_20132,N_19134,N_16141);
or U20133 (N_20133,N_17177,N_17526);
or U20134 (N_20134,N_16536,N_17600);
and U20135 (N_20135,N_19713,N_16864);
and U20136 (N_20136,N_19637,N_15277);
xor U20137 (N_20137,N_15478,N_17857);
xor U20138 (N_20138,N_17170,N_18799);
nand U20139 (N_20139,N_19998,N_17080);
xnor U20140 (N_20140,N_18394,N_16789);
nor U20141 (N_20141,N_19295,N_18370);
or U20142 (N_20142,N_15857,N_16656);
or U20143 (N_20143,N_18992,N_17034);
and U20144 (N_20144,N_18134,N_19040);
xnor U20145 (N_20145,N_16940,N_15989);
or U20146 (N_20146,N_15985,N_16259);
nand U20147 (N_20147,N_17733,N_16882);
and U20148 (N_20148,N_16352,N_17594);
nor U20149 (N_20149,N_18552,N_17019);
nor U20150 (N_20150,N_19203,N_19250);
xor U20151 (N_20151,N_16766,N_16152);
or U20152 (N_20152,N_17778,N_19061);
xnor U20153 (N_20153,N_15604,N_15285);
xnor U20154 (N_20154,N_16124,N_17962);
and U20155 (N_20155,N_17628,N_19874);
and U20156 (N_20156,N_17222,N_16569);
and U20157 (N_20157,N_16445,N_15338);
or U20158 (N_20158,N_16938,N_17207);
or U20159 (N_20159,N_18475,N_19537);
or U20160 (N_20160,N_18474,N_16020);
nand U20161 (N_20161,N_18989,N_16630);
nand U20162 (N_20162,N_17147,N_15191);
xor U20163 (N_20163,N_15992,N_17755);
or U20164 (N_20164,N_15096,N_15663);
xnor U20165 (N_20165,N_19082,N_15980);
nand U20166 (N_20166,N_15443,N_19322);
nand U20167 (N_20167,N_18877,N_16408);
nand U20168 (N_20168,N_19187,N_15091);
nand U20169 (N_20169,N_16679,N_18224);
xnor U20170 (N_20170,N_17284,N_19987);
and U20171 (N_20171,N_16390,N_16553);
nor U20172 (N_20172,N_19852,N_17070);
xnor U20173 (N_20173,N_17521,N_17886);
or U20174 (N_20174,N_16510,N_19230);
and U20175 (N_20175,N_19212,N_19819);
xor U20176 (N_20176,N_16374,N_17752);
nor U20177 (N_20177,N_17352,N_16953);
and U20178 (N_20178,N_16809,N_17035);
nand U20179 (N_20179,N_16058,N_18297);
nor U20180 (N_20180,N_17924,N_19160);
xnor U20181 (N_20181,N_19601,N_17418);
and U20182 (N_20182,N_15152,N_16606);
xor U20183 (N_20183,N_16193,N_15637);
nor U20184 (N_20184,N_15221,N_17779);
nor U20185 (N_20185,N_18649,N_15929);
or U20186 (N_20186,N_17692,N_19597);
and U20187 (N_20187,N_17515,N_15514);
xnor U20188 (N_20188,N_15297,N_17519);
and U20189 (N_20189,N_18005,N_15418);
and U20190 (N_20190,N_15935,N_17460);
nand U20191 (N_20191,N_19361,N_17956);
nand U20192 (N_20192,N_15232,N_18737);
nand U20193 (N_20193,N_18826,N_17561);
xor U20194 (N_20194,N_18368,N_17508);
and U20195 (N_20195,N_16512,N_16095);
or U20196 (N_20196,N_19267,N_15621);
nand U20197 (N_20197,N_15964,N_15831);
or U20198 (N_20198,N_17206,N_16718);
and U20199 (N_20199,N_15622,N_16219);
nor U20200 (N_20200,N_19880,N_15948);
or U20201 (N_20201,N_19437,N_15555);
or U20202 (N_20202,N_16357,N_18837);
or U20203 (N_20203,N_19642,N_16395);
xor U20204 (N_20204,N_17260,N_19060);
nand U20205 (N_20205,N_18655,N_19139);
nand U20206 (N_20206,N_17382,N_15315);
xor U20207 (N_20207,N_18227,N_17849);
nand U20208 (N_20208,N_16810,N_19435);
nand U20209 (N_20209,N_17232,N_16110);
nand U20210 (N_20210,N_15927,N_16986);
nor U20211 (N_20211,N_16201,N_17351);
nor U20212 (N_20212,N_19216,N_19584);
or U20213 (N_20213,N_16273,N_16769);
nor U20214 (N_20214,N_18741,N_19740);
and U20215 (N_20215,N_15673,N_18866);
nand U20216 (N_20216,N_17360,N_15124);
xnor U20217 (N_20217,N_15100,N_19189);
nor U20218 (N_20218,N_16534,N_19386);
xor U20219 (N_20219,N_15066,N_18736);
xnor U20220 (N_20220,N_16353,N_15151);
nand U20221 (N_20221,N_19300,N_19122);
nor U20222 (N_20222,N_18260,N_18650);
and U20223 (N_20223,N_18748,N_15585);
nor U20224 (N_20224,N_17533,N_18496);
xnor U20225 (N_20225,N_19917,N_17593);
xnor U20226 (N_20226,N_18413,N_19681);
xnor U20227 (N_20227,N_16318,N_19370);
or U20228 (N_20228,N_16296,N_15391);
nand U20229 (N_20229,N_16003,N_18118);
and U20230 (N_20230,N_19882,N_16485);
xor U20231 (N_20231,N_17441,N_19979);
xnor U20232 (N_20232,N_19037,N_16669);
or U20233 (N_20233,N_16078,N_18696);
or U20234 (N_20234,N_16617,N_16265);
nand U20235 (N_20235,N_18171,N_17907);
nand U20236 (N_20236,N_17489,N_17918);
xor U20237 (N_20237,N_15855,N_17058);
xor U20238 (N_20238,N_15282,N_18341);
nor U20239 (N_20239,N_15287,N_19706);
xor U20240 (N_20240,N_16339,N_16815);
xnor U20241 (N_20241,N_19772,N_19744);
nor U20242 (N_20242,N_16088,N_17806);
xor U20243 (N_20243,N_15237,N_16397);
nand U20244 (N_20244,N_16593,N_17427);
or U20245 (N_20245,N_15878,N_15002);
nand U20246 (N_20246,N_16852,N_15600);
and U20247 (N_20247,N_15756,N_17818);
or U20248 (N_20248,N_19308,N_19339);
or U20249 (N_20249,N_19498,N_15827);
xor U20250 (N_20250,N_17065,N_16988);
nand U20251 (N_20251,N_15298,N_18463);
xor U20252 (N_20252,N_16770,N_18555);
nand U20253 (N_20253,N_16419,N_18358);
xor U20254 (N_20254,N_17729,N_16584);
or U20255 (N_20255,N_17710,N_16793);
nand U20256 (N_20256,N_17588,N_18886);
nor U20257 (N_20257,N_15531,N_19833);
and U20258 (N_20258,N_16633,N_19021);
nor U20259 (N_20259,N_16916,N_16906);
nor U20260 (N_20260,N_18176,N_16239);
xnor U20261 (N_20261,N_19198,N_15306);
nand U20262 (N_20262,N_18339,N_16263);
or U20263 (N_20263,N_17409,N_18324);
and U20264 (N_20264,N_15130,N_15970);
xnor U20265 (N_20265,N_19415,N_17904);
nor U20266 (N_20266,N_15241,N_16571);
or U20267 (N_20267,N_17478,N_16984);
nand U20268 (N_20268,N_18852,N_17339);
or U20269 (N_20269,N_18298,N_19521);
nor U20270 (N_20270,N_17209,N_17839);
or U20271 (N_20271,N_15720,N_18674);
xnor U20272 (N_20272,N_18593,N_19408);
nand U20273 (N_20273,N_15871,N_19867);
nand U20274 (N_20274,N_19734,N_15185);
nand U20275 (N_20275,N_16247,N_17885);
or U20276 (N_20276,N_19196,N_17293);
xor U20277 (N_20277,N_19835,N_17799);
or U20278 (N_20278,N_18430,N_17610);
xnor U20279 (N_20279,N_17739,N_18041);
and U20280 (N_20280,N_15265,N_15414);
nor U20281 (N_20281,N_16505,N_17134);
or U20282 (N_20282,N_15072,N_18690);
nand U20283 (N_20283,N_16723,N_19104);
and U20284 (N_20284,N_15824,N_16689);
xor U20285 (N_20285,N_17109,N_18175);
or U20286 (N_20286,N_18986,N_19416);
nand U20287 (N_20287,N_17888,N_17234);
nand U20288 (N_20288,N_18961,N_15296);
xor U20289 (N_20289,N_16379,N_16478);
and U20290 (N_20290,N_17936,N_17525);
or U20291 (N_20291,N_18121,N_18200);
xnor U20292 (N_20292,N_17204,N_18661);
xor U20293 (N_20293,N_17679,N_19443);
and U20294 (N_20294,N_19508,N_18487);
nor U20295 (N_20295,N_19422,N_16346);
xor U20296 (N_20296,N_15921,N_15665);
nor U20297 (N_20297,N_16646,N_15219);
nand U20298 (N_20298,N_16700,N_16116);
or U20299 (N_20299,N_18600,N_17879);
nor U20300 (N_20300,N_19610,N_18228);
xor U20301 (N_20301,N_17201,N_16684);
nor U20302 (N_20302,N_15343,N_18767);
xor U20303 (N_20303,N_18479,N_18515);
xnor U20304 (N_20304,N_17974,N_19215);
and U20305 (N_20305,N_15489,N_17982);
or U20306 (N_20306,N_19354,N_17076);
or U20307 (N_20307,N_18679,N_19605);
nand U20308 (N_20308,N_17221,N_17828);
xor U20309 (N_20309,N_18660,N_18063);
nor U20310 (N_20310,N_17380,N_19210);
xor U20311 (N_20311,N_19421,N_16949);
and U20312 (N_20312,N_15164,N_18936);
and U20313 (N_20313,N_16891,N_15876);
or U20314 (N_20314,N_16272,N_15320);
xnor U20315 (N_20315,N_19136,N_16994);
or U20316 (N_20316,N_17868,N_18393);
nor U20317 (N_20317,N_15472,N_19684);
nor U20318 (N_20318,N_19892,N_16294);
nand U20319 (N_20319,N_16359,N_19385);
nor U20320 (N_20320,N_19305,N_15424);
or U20321 (N_20321,N_19956,N_15888);
or U20322 (N_20322,N_18784,N_16214);
nor U20323 (N_20323,N_17756,N_15597);
nor U20324 (N_20324,N_19320,N_15147);
and U20325 (N_20325,N_16585,N_16304);
nor U20326 (N_20326,N_18329,N_18335);
or U20327 (N_20327,N_16433,N_18256);
nand U20328 (N_20328,N_19281,N_16667);
xor U20329 (N_20329,N_19513,N_18863);
nand U20330 (N_20330,N_16113,N_16066);
or U20331 (N_20331,N_15202,N_16861);
nand U20332 (N_20332,N_18559,N_17388);
and U20333 (N_20333,N_16728,N_17738);
xor U20334 (N_20334,N_15760,N_18702);
nand U20335 (N_20335,N_16048,N_18445);
nand U20336 (N_20336,N_19673,N_19162);
nand U20337 (N_20337,N_18291,N_19854);
xor U20338 (N_20338,N_19658,N_15101);
or U20339 (N_20339,N_17870,N_17822);
xnor U20340 (N_20340,N_18124,N_15930);
nor U20341 (N_20341,N_16111,N_18853);
nor U20342 (N_20342,N_19377,N_16474);
and U20343 (N_20343,N_17713,N_17838);
xor U20344 (N_20344,N_19664,N_16576);
and U20345 (N_20345,N_17988,N_19752);
and U20346 (N_20346,N_18930,N_18804);
nor U20347 (N_20347,N_17215,N_19663);
nor U20348 (N_20348,N_16097,N_18055);
nor U20349 (N_20349,N_15695,N_16207);
or U20350 (N_20350,N_17744,N_16417);
nor U20351 (N_20351,N_18315,N_16441);
xor U20352 (N_20352,N_16976,N_18067);
or U20353 (N_20353,N_17291,N_18193);
nand U20354 (N_20354,N_16305,N_16911);
xnor U20355 (N_20355,N_18328,N_18446);
and U20356 (N_20356,N_17771,N_18369);
or U20357 (N_20357,N_18127,N_16862);
or U20358 (N_20358,N_19009,N_19355);
or U20359 (N_20359,N_18502,N_19755);
and U20360 (N_20360,N_19838,N_17671);
nor U20361 (N_20361,N_15601,N_19697);
xnor U20362 (N_20362,N_18848,N_16640);
nand U20363 (N_20363,N_16254,N_15868);
or U20364 (N_20364,N_17614,N_18421);
and U20365 (N_20365,N_16473,N_17750);
nor U20366 (N_20366,N_17362,N_17623);
or U20367 (N_20367,N_19075,N_17977);
nor U20368 (N_20368,N_16767,N_16454);
and U20369 (N_20369,N_16772,N_15245);
and U20370 (N_20370,N_17704,N_15607);
nand U20371 (N_20371,N_17727,N_19232);
nand U20372 (N_20372,N_15946,N_19848);
and U20373 (N_20373,N_15575,N_16847);
nor U20374 (N_20374,N_15016,N_17431);
nor U20375 (N_20375,N_15393,N_16914);
nor U20376 (N_20376,N_18211,N_18195);
nor U20377 (N_20377,N_17536,N_19516);
and U20378 (N_20378,N_15040,N_18082);
nand U20379 (N_20379,N_18905,N_18541);
or U20380 (N_20380,N_15795,N_16083);
nor U20381 (N_20381,N_15179,N_16626);
nand U20382 (N_20382,N_18371,N_15490);
nand U20383 (N_20383,N_15441,N_18987);
xnor U20384 (N_20384,N_15952,N_15262);
and U20385 (N_20385,N_17182,N_18202);
xor U20386 (N_20386,N_19759,N_18829);
and U20387 (N_20387,N_17627,N_19932);
and U20388 (N_20388,N_19054,N_16523);
or U20389 (N_20389,N_16910,N_15439);
xnor U20390 (N_20390,N_17851,N_17161);
nand U20391 (N_20391,N_15082,N_19680);
xor U20392 (N_20392,N_16165,N_19717);
xnor U20393 (N_20393,N_16295,N_19071);
nor U20394 (N_20394,N_19859,N_19259);
nand U20395 (N_20395,N_18128,N_19913);
xnor U20396 (N_20396,N_15198,N_15389);
and U20397 (N_20397,N_19985,N_16236);
nor U20398 (N_20398,N_18428,N_19241);
or U20399 (N_20399,N_17244,N_16170);
nand U20400 (N_20400,N_19309,N_18361);
or U20401 (N_20401,N_18654,N_16302);
xor U20402 (N_20402,N_18528,N_17368);
nor U20403 (N_20403,N_16846,N_16177);
nand U20404 (N_20404,N_16481,N_18873);
nand U20405 (N_20405,N_19600,N_16905);
nor U20406 (N_20406,N_15303,N_15543);
and U20407 (N_20407,N_15764,N_19935);
nor U20408 (N_20408,N_16637,N_19280);
or U20409 (N_20409,N_17509,N_16677);
and U20410 (N_20410,N_18347,N_15859);
xnor U20411 (N_20411,N_15728,N_18816);
or U20412 (N_20412,N_16583,N_15031);
nand U20413 (N_20413,N_16997,N_19293);
nor U20414 (N_20414,N_19840,N_19918);
or U20415 (N_20415,N_19766,N_18932);
and U20416 (N_20416,N_15561,N_19180);
nand U20417 (N_20417,N_15978,N_17117);
nand U20418 (N_20418,N_15005,N_17344);
nor U20419 (N_20419,N_19553,N_16120);
or U20420 (N_20420,N_19131,N_19798);
xnor U20421 (N_20421,N_15520,N_15612);
nand U20422 (N_20422,N_18433,N_17267);
nand U20423 (N_20423,N_15521,N_16205);
xor U20424 (N_20424,N_17630,N_17012);
and U20425 (N_20425,N_16238,N_15483);
or U20426 (N_20426,N_16006,N_18950);
xnor U20427 (N_20427,N_16154,N_15177);
nor U20428 (N_20428,N_16021,N_16612);
or U20429 (N_20429,N_16025,N_18151);
or U20430 (N_20430,N_15843,N_16314);
or U20431 (N_20431,N_15996,N_15884);
and U20432 (N_20432,N_15702,N_19316);
nor U20433 (N_20433,N_18018,N_17753);
nor U20434 (N_20434,N_17061,N_15215);
or U20435 (N_20435,N_19200,N_16760);
xor U20436 (N_20436,N_16887,N_19465);
xor U20437 (N_20437,N_17356,N_18706);
and U20438 (N_20438,N_19388,N_16705);
xor U20439 (N_20439,N_18024,N_16409);
nand U20440 (N_20440,N_15025,N_19624);
or U20441 (N_20441,N_17993,N_19331);
or U20442 (N_20442,N_15250,N_15973);
nand U20443 (N_20443,N_15430,N_17921);
xor U20444 (N_20444,N_17008,N_15474);
and U20445 (N_20445,N_18543,N_17681);
and U20446 (N_20446,N_18068,N_17167);
nand U20447 (N_20447,N_16197,N_15882);
and U20448 (N_20448,N_17017,N_19003);
nor U20449 (N_20449,N_18533,N_19512);
nand U20450 (N_20450,N_18726,N_15517);
and U20451 (N_20451,N_16027,N_16387);
and U20452 (N_20452,N_19453,N_16613);
or U20453 (N_20453,N_15349,N_18652);
xor U20454 (N_20454,N_18144,N_15162);
and U20455 (N_20455,N_17624,N_19988);
nor U20456 (N_20456,N_18613,N_16160);
nand U20457 (N_20457,N_17319,N_15360);
and U20458 (N_20458,N_15008,N_16620);
xnor U20459 (N_20459,N_16915,N_16839);
and U20460 (N_20460,N_17826,N_19356);
or U20461 (N_20461,N_16034,N_16759);
or U20462 (N_20462,N_16721,N_15144);
nand U20463 (N_20463,N_19286,N_19675);
or U20464 (N_20464,N_18903,N_19518);
xnor U20465 (N_20465,N_16127,N_15294);
or U20466 (N_20466,N_17792,N_19261);
nor U20467 (N_20467,N_17433,N_19016);
xnor U20468 (N_20468,N_19420,N_19263);
nand U20469 (N_20469,N_15381,N_17269);
nand U20470 (N_20470,N_17696,N_19378);
nor U20471 (N_20471,N_19662,N_16140);
or U20472 (N_20472,N_15830,N_16464);
xnor U20473 (N_20473,N_19581,N_16596);
or U20474 (N_20474,N_18130,N_18862);
nor U20475 (N_20475,N_18054,N_19118);
or U20476 (N_20476,N_18110,N_19721);
or U20477 (N_20477,N_19876,N_19202);
nand U20478 (N_20478,N_17550,N_15704);
nor U20479 (N_20479,N_19757,N_15504);
nor U20480 (N_20480,N_15866,N_17002);
or U20481 (N_20481,N_17554,N_19125);
nor U20482 (N_20482,N_17263,N_17176);
xor U20483 (N_20483,N_16217,N_17669);
nor U20484 (N_20484,N_16059,N_15022);
and U20485 (N_20485,N_18093,N_16266);
nor U20486 (N_20486,N_16444,N_17266);
or U20487 (N_20487,N_16675,N_18294);
nor U20488 (N_20488,N_18468,N_17208);
nor U20489 (N_20489,N_15451,N_16347);
xor U20490 (N_20490,N_15705,N_16643);
xor U20491 (N_20491,N_19526,N_19817);
and U20492 (N_20492,N_18458,N_17316);
nor U20493 (N_20493,N_18531,N_19864);
and U20494 (N_20494,N_17415,N_16876);
nor U20495 (N_20495,N_15708,N_17691);
nand U20496 (N_20496,N_17690,N_15317);
and U20497 (N_20497,N_17425,N_19842);
and U20498 (N_20498,N_18089,N_15684);
nor U20499 (N_20499,N_18278,N_19400);
nand U20500 (N_20500,N_18520,N_15918);
or U20501 (N_20501,N_16702,N_15467);
xor U20502 (N_20502,N_18440,N_16337);
nor U20503 (N_20503,N_19288,N_18630);
xnor U20504 (N_20504,N_19806,N_16665);
nor U20505 (N_20505,N_18460,N_15769);
nor U20506 (N_20506,N_18815,N_18285);
and U20507 (N_20507,N_19730,N_17439);
xor U20508 (N_20508,N_16753,N_15751);
and U20509 (N_20509,N_19358,N_17890);
nand U20510 (N_20510,N_18299,N_19121);
xor U20511 (N_20511,N_17620,N_15797);
nor U20512 (N_20512,N_17835,N_16851);
xnor U20513 (N_20513,N_15596,N_18366);
or U20514 (N_20514,N_18563,N_15926);
xnor U20515 (N_20515,N_15700,N_16913);
nand U20516 (N_20516,N_19901,N_19851);
nand U20517 (N_20517,N_15401,N_17531);
nand U20518 (N_20518,N_19344,N_19903);
xor U20519 (N_20519,N_16224,N_19256);
xnor U20520 (N_20520,N_17023,N_17423);
nand U20521 (N_20521,N_15093,N_18551);
or U20522 (N_20522,N_17773,N_16211);
xor U20523 (N_20523,N_19830,N_16747);
xnor U20524 (N_20524,N_18761,N_19499);
nand U20525 (N_20525,N_17859,N_19269);
or U20526 (N_20526,N_18167,N_15448);
nand U20527 (N_20527,N_18034,N_17928);
xnor U20528 (N_20528,N_15766,N_16220);
and U20529 (N_20529,N_17210,N_17392);
nor U20530 (N_20530,N_19831,N_19704);
nor U20531 (N_20531,N_17854,N_19635);
nor U20532 (N_20532,N_15506,N_18113);
nor U20533 (N_20533,N_17609,N_19371);
xor U20534 (N_20534,N_18478,N_17625);
or U20535 (N_20535,N_18148,N_15363);
and U20536 (N_20536,N_17995,N_18119);
and U20537 (N_20537,N_15800,N_19579);
nand U20538 (N_20538,N_15635,N_15524);
nand U20539 (N_20539,N_17777,N_15872);
and U20540 (N_20540,N_18997,N_17989);
and U20541 (N_20541,N_18300,N_19634);
xnor U20542 (N_20542,N_15677,N_17013);
xnor U20543 (N_20543,N_16797,N_16834);
nand U20544 (N_20544,N_17463,N_17470);
nand U20545 (N_20545,N_15461,N_17544);
or U20546 (N_20546,N_19243,N_17659);
and U20547 (N_20547,N_17367,N_19423);
nand U20548 (N_20548,N_16493,N_18514);
or U20549 (N_20549,N_17240,N_19073);
xor U20550 (N_20550,N_19133,N_17650);
and U20551 (N_20551,N_16043,N_18104);
nor U20552 (N_20552,N_19727,N_17285);
nor U20553 (N_20553,N_17566,N_19463);
xnor U20554 (N_20554,N_18688,N_15592);
xor U20555 (N_20555,N_16830,N_16460);
or U20556 (N_20556,N_15562,N_18639);
nand U20557 (N_20557,N_19018,N_18898);
nor U20558 (N_20558,N_15773,N_17584);
or U20559 (N_20559,N_18156,N_18576);
and U20560 (N_20560,N_18044,N_16108);
nand U20561 (N_20561,N_16865,N_15593);
nor U20562 (N_20562,N_17567,N_19689);
or U20563 (N_20563,N_19793,N_16627);
or U20564 (N_20564,N_16345,N_17036);
xnor U20565 (N_20565,N_18345,N_17484);
or U20566 (N_20566,N_17202,N_16398);
and U20567 (N_20567,N_17312,N_15302);
nand U20568 (N_20568,N_15491,N_18869);
and U20569 (N_20569,N_18605,N_18709);
and U20570 (N_20570,N_17965,N_16787);
xor U20571 (N_20571,N_17214,N_17639);
or U20572 (N_20572,N_15685,N_17075);
xor U20573 (N_20573,N_17272,N_17532);
xor U20574 (N_20574,N_19519,N_19151);
nand U20575 (N_20575,N_16099,N_16028);
nand U20576 (N_20576,N_18634,N_16002);
nor U20577 (N_20577,N_16972,N_18647);
nand U20578 (N_20578,N_17909,N_17925);
or U20579 (N_20579,N_18398,N_15383);
nor U20580 (N_20580,N_15190,N_18894);
nor U20581 (N_20581,N_18165,N_16706);
and U20582 (N_20582,N_19008,N_19116);
nand U20583 (N_20583,N_15588,N_17861);
or U20584 (N_20584,N_16442,N_16685);
or U20585 (N_20585,N_18046,N_15118);
and U20586 (N_20586,N_16968,N_19034);
and U20587 (N_20587,N_17832,N_17217);
or U20588 (N_20588,N_19657,N_16309);
nor U20589 (N_20589,N_16106,N_15175);
nor U20590 (N_20590,N_18901,N_19984);
and U20591 (N_20591,N_15488,N_17457);
or U20592 (N_20592,N_19185,N_17505);
nand U20593 (N_20593,N_18813,N_15233);
nand U20594 (N_20594,N_16699,N_17040);
or U20595 (N_20595,N_16198,N_18109);
nor U20596 (N_20596,N_15605,N_15382);
nand U20597 (N_20597,N_19595,N_18306);
nor U20598 (N_20598,N_16996,N_17749);
and U20599 (N_20599,N_15460,N_17960);
or U20600 (N_20600,N_19920,N_17412);
nor U20601 (N_20601,N_17128,N_17734);
and U20602 (N_20602,N_19460,N_15642);
and U20603 (N_20603,N_18662,N_18793);
xnor U20604 (N_20604,N_19391,N_18472);
nor U20605 (N_20605,N_15386,N_19353);
nand U20606 (N_20606,N_17770,N_18638);
nand U20607 (N_20607,N_15907,N_17829);
and U20608 (N_20608,N_18867,N_16350);
xor U20609 (N_20609,N_16383,N_15803);
xor U20610 (N_20610,N_15052,N_17689);
xnor U20611 (N_20611,N_15739,N_18597);
and U20612 (N_20612,N_18401,N_16162);
or U20613 (N_20613,N_18080,N_17447);
xnor U20614 (N_20614,N_16331,N_19801);
or U20615 (N_20615,N_17243,N_18521);
xnor U20616 (N_20616,N_18948,N_17518);
xnor U20617 (N_20617,N_19324,N_18143);
and U20618 (N_20618,N_19603,N_17112);
and U20619 (N_20619,N_18117,N_16438);
or U20620 (N_20620,N_15576,N_17099);
nor U20621 (N_20621,N_18577,N_16784);
nor U20622 (N_20622,N_16222,N_18141);
nor U20623 (N_20623,N_18447,N_19837);
nand U20624 (N_20624,N_16991,N_18170);
xnor U20625 (N_20625,N_19803,N_15056);
xnor U20626 (N_20626,N_19036,N_19724);
and U20627 (N_20627,N_18079,N_18822);
nor U20628 (N_20628,N_18883,N_19418);
or U20629 (N_20629,N_19213,N_15703);
nand U20630 (N_20630,N_17259,N_17046);
or U20631 (N_20631,N_15628,N_16935);
and U20632 (N_20632,N_17083,N_17155);
xor U20633 (N_20633,N_15452,N_19958);
or U20634 (N_20634,N_19352,N_19698);
or U20635 (N_20635,N_19781,N_17657);
and U20636 (N_20636,N_16880,N_17910);
or U20637 (N_20637,N_17699,N_15048);
nand U20638 (N_20638,N_19555,N_17621);
nor U20639 (N_20639,N_19080,N_16944);
and U20640 (N_20640,N_18296,N_17224);
or U20641 (N_20641,N_19621,N_15257);
nand U20642 (N_20642,N_17016,N_19092);
nor U20643 (N_20643,N_16341,N_15557);
or U20644 (N_20644,N_17922,N_17709);
or U20645 (N_20645,N_17617,N_16591);
or U20646 (N_20646,N_19175,N_15058);
xor U20647 (N_20647,N_16877,N_16241);
and U20648 (N_20648,N_16056,N_17523);
or U20649 (N_20649,N_15345,N_17118);
nand U20650 (N_20650,N_17539,N_17426);
xor U20651 (N_20651,N_17563,N_19271);
and U20652 (N_20652,N_15848,N_15893);
nand U20653 (N_20653,N_19608,N_16368);
nand U20654 (N_20654,N_18833,N_17629);
xnor U20655 (N_20655,N_17789,N_19454);
or U20656 (N_20656,N_18216,N_18069);
xor U20657 (N_20657,N_16187,N_16693);
nand U20658 (N_20658,N_19141,N_15388);
or U20659 (N_20659,N_19708,N_15323);
nor U20660 (N_20660,N_18071,N_15446);
or U20661 (N_20661,N_17581,N_16199);
and U20662 (N_20662,N_17211,N_17641);
nor U20663 (N_20663,N_16502,N_15281);
and U20664 (N_20664,N_15125,N_16933);
xnor U20665 (N_20665,N_19821,N_17632);
nor U20666 (N_20666,N_17308,N_19001);
nand U20667 (N_20667,N_18857,N_16496);
nand U20668 (N_20668,N_17969,N_17282);
nand U20669 (N_20669,N_16661,N_19679);
nor U20670 (N_20670,N_18953,N_15624);
xor U20671 (N_20671,N_17542,N_17591);
and U20672 (N_20672,N_15318,N_16719);
and U20673 (N_20673,N_19237,N_15721);
nor U20674 (N_20674,N_17672,N_19629);
xor U20675 (N_20675,N_17929,N_16157);
xor U20676 (N_20676,N_19085,N_18087);
nand U20677 (N_20677,N_15794,N_16000);
and U20678 (N_20678,N_17697,N_16896);
nand U20679 (N_20679,N_15877,N_15274);
or U20680 (N_20680,N_17502,N_15280);
and U20681 (N_20681,N_19614,N_16868);
nand U20682 (N_20682,N_18890,N_16094);
nor U20683 (N_20683,N_16325,N_15951);
and U20684 (N_20684,N_18166,N_15229);
or U20685 (N_20685,N_17985,N_19055);
xor U20686 (N_20686,N_16126,N_19960);
nor U20687 (N_20687,N_16149,N_16663);
nand U20688 (N_20688,N_16377,N_19789);
or U20689 (N_20689,N_15319,N_17768);
xor U20690 (N_20690,N_18441,N_15898);
or U20691 (N_20691,N_16889,N_17007);
xor U20692 (N_20692,N_17842,N_18564);
nand U20693 (N_20693,N_18016,N_15536);
xnor U20694 (N_20694,N_18565,N_16955);
xor U20695 (N_20695,N_18746,N_18740);
nor U20696 (N_20696,N_19915,N_16307);
and U20697 (N_20697,N_17703,N_15347);
and U20698 (N_20698,N_15765,N_15904);
or U20699 (N_20699,N_17808,N_16035);
xor U20700 (N_20700,N_19211,N_15355);
nor U20701 (N_20701,N_15442,N_18439);
nand U20702 (N_20702,N_15336,N_17972);
nor U20703 (N_20703,N_17162,N_18534);
and U20704 (N_20704,N_18396,N_17648);
or U20705 (N_20705,N_15107,N_18527);
and U20706 (N_20706,N_16091,N_16954);
or U20707 (N_20707,N_15435,N_17310);
nor U20708 (N_20708,N_17054,N_16282);
and U20709 (N_20709,N_15136,N_17175);
xnor U20710 (N_20710,N_17652,N_17595);
nor U20711 (N_20711,N_19501,N_19357);
or U20712 (N_20712,N_16327,N_17408);
and U20713 (N_20713,N_15095,N_16600);
nor U20714 (N_20714,N_15916,N_15771);
or U20715 (N_20715,N_19938,N_16326);
or U20716 (N_20716,N_18659,N_17559);
nor U20717 (N_20717,N_19559,N_16920);
nand U20718 (N_20718,N_18974,N_18451);
or U20719 (N_20719,N_15953,N_18231);
nor U20720 (N_20720,N_16081,N_16123);
or U20721 (N_20721,N_18498,N_16145);
and U20722 (N_20722,N_17227,N_15598);
and U20723 (N_20723,N_16416,N_19074);
xnor U20724 (N_20724,N_19561,N_16841);
xor U20725 (N_20725,N_17361,N_19802);
and U20726 (N_20726,N_15818,N_18425);
xnor U20727 (N_20727,N_17785,N_18169);
nor U20728 (N_20728,N_17616,N_16270);
or U20729 (N_20729,N_17762,N_17653);
and U20730 (N_20730,N_19364,N_19390);
and U20731 (N_20731,N_19873,N_18805);
nor U20732 (N_20732,N_17355,N_19883);
nor U20733 (N_20733,N_18179,N_17288);
nand U20734 (N_20734,N_16011,N_17238);
or U20735 (N_20735,N_16279,N_19888);
nand U20736 (N_20736,N_15286,N_19476);
xor U20737 (N_20737,N_15559,N_16057);
nand U20738 (N_20738,N_19688,N_17643);
nand U20739 (N_20739,N_17919,N_19220);
and U20740 (N_20740,N_15613,N_17287);
nor U20741 (N_20741,N_17436,N_17169);
nor U20742 (N_20742,N_17664,N_17725);
or U20743 (N_20743,N_17545,N_16216);
nand U20744 (N_20744,N_16828,N_19540);
nand U20745 (N_20745,N_15943,N_17670);
nor U20746 (N_20746,N_17350,N_15957);
and U20747 (N_20747,N_16166,N_16427);
nand U20748 (N_20748,N_18155,N_17486);
nor U20749 (N_20749,N_16826,N_15735);
and U20750 (N_20750,N_19265,N_18250);
and U20751 (N_20751,N_17875,N_19500);
xnor U20752 (N_20752,N_15573,N_18571);
nand U20753 (N_20753,N_16589,N_15207);
nor U20754 (N_20754,N_17406,N_16215);
nor U20755 (N_20755,N_15590,N_17817);
or U20756 (N_20756,N_16651,N_19329);
nor U20757 (N_20757,N_16812,N_17149);
and U20758 (N_20758,N_16808,N_19161);
and U20759 (N_20759,N_16129,N_19604);
nor U20760 (N_20760,N_16825,N_15404);
xor U20761 (N_20761,N_19996,N_18790);
and U20762 (N_20762,N_19229,N_16594);
or U20763 (N_20763,N_15870,N_15204);
xor U20764 (N_20764,N_18686,N_18586);
nor U20765 (N_20765,N_17429,N_17407);
xor U20766 (N_20766,N_16421,N_16184);
nor U20767 (N_20767,N_16014,N_18039);
nand U20768 (N_20768,N_17766,N_16785);
xor U20769 (N_20769,N_15791,N_15780);
nor U20770 (N_20770,N_19780,N_17674);
and U20771 (N_20771,N_16628,N_18979);
or U20772 (N_20772,N_16683,N_18184);
or U20773 (N_20773,N_17847,N_18778);
nor U20774 (N_20774,N_17970,N_19858);
nand U20775 (N_20775,N_15411,N_16979);
nand U20776 (N_20776,N_17438,N_18692);
nand U20777 (N_20777,N_17959,N_17622);
xor U20778 (N_20778,N_15024,N_17393);
nand U20779 (N_20779,N_19038,N_18934);
and U20780 (N_20780,N_18269,N_15903);
xnor U20781 (N_20781,N_18823,N_16635);
xnor U20782 (N_20782,N_15662,N_16064);
nand U20783 (N_20783,N_16873,N_15566);
or U20784 (N_20784,N_17840,N_18213);
and U20785 (N_20785,N_15594,N_16001);
or U20786 (N_20786,N_19583,N_19166);
xnor U20787 (N_20787,N_17558,N_19761);
xor U20788 (N_20788,N_15647,N_15465);
or U20789 (N_20789,N_17119,N_16668);
or U20790 (N_20790,N_15326,N_17242);
nor U20791 (N_20791,N_15309,N_17419);
xnor U20792 (N_20792,N_15819,N_17708);
nor U20793 (N_20793,N_17474,N_15146);
or U20794 (N_20794,N_18223,N_17135);
and U20795 (N_20795,N_19233,N_18841);
or U20796 (N_20796,N_15044,N_17500);
xor U20797 (N_20797,N_18365,N_17146);
and U20798 (N_20798,N_19014,N_17871);
or U20799 (N_20799,N_15180,N_17271);
and U20800 (N_20800,N_15579,N_16632);
and U20801 (N_20801,N_17978,N_18510);
nor U20802 (N_20802,N_19787,N_17520);
or U20803 (N_20803,N_19111,N_15860);
and U20804 (N_20804,N_16525,N_19775);
nand U20805 (N_20805,N_16928,N_18011);
or U20806 (N_20806,N_18509,N_18537);
nor U20807 (N_20807,N_15088,N_18190);
nor U20808 (N_20808,N_18830,N_19514);
or U20809 (N_20809,N_19194,N_19193);
nor U20810 (N_20810,N_17855,N_18601);
nor U20811 (N_20811,N_17501,N_18303);
xnor U20812 (N_20812,N_18919,N_18337);
or U20813 (N_20813,N_16614,N_18727);
or U20814 (N_20814,N_16053,N_18160);
and U20815 (N_20815,N_18665,N_17265);
nand U20816 (N_20816,N_16023,N_15141);
or U20817 (N_20817,N_18392,N_19811);
nand U20818 (N_20818,N_15947,N_18999);
xor U20819 (N_20819,N_16117,N_18234);
nor U20820 (N_20820,N_18859,N_15962);
xor U20821 (N_20821,N_19598,N_15484);
nand U20822 (N_20822,N_19433,N_18701);
and U20823 (N_20823,N_16167,N_17078);
and U20824 (N_20824,N_15670,N_17359);
nand U20825 (N_20825,N_16200,N_19692);
or U20826 (N_20826,N_18635,N_17587);
or U20827 (N_20827,N_18561,N_17724);
xnor U20828 (N_20828,N_17189,N_17084);
nor U20829 (N_20829,N_16696,N_15079);
nor U20830 (N_20830,N_15413,N_16471);
xnor U20831 (N_20831,N_17807,N_17903);
nand U20832 (N_20832,N_16260,N_16137);
nor U20833 (N_20833,N_18698,N_18860);
nand U20834 (N_20834,N_15422,N_17853);
or U20835 (N_20835,N_15899,N_19363);
or U20836 (N_20836,N_16030,N_18235);
xnor U20837 (N_20837,N_17354,N_15726);
and U20838 (N_20838,N_19995,N_16253);
and U20839 (N_20839,N_16565,N_15801);
nor U20840 (N_20840,N_17286,N_18242);
nor U20841 (N_20841,N_17923,N_18026);
xor U20842 (N_20842,N_16771,N_17754);
xnor U20843 (N_20843,N_15806,N_19132);
nor U20844 (N_20844,N_18910,N_18524);
nand U20845 (N_20845,N_16153,N_18771);
nor U20846 (N_20846,N_17767,N_15027);
or U20847 (N_20847,N_16918,N_15372);
nor U20848 (N_20848,N_16144,N_18266);
xor U20849 (N_20849,N_18824,N_17711);
and U20850 (N_20850,N_18273,N_15646);
xnor U20851 (N_20851,N_16192,N_18570);
nor U20852 (N_20852,N_19289,N_15892);
nand U20853 (N_20853,N_15944,N_15425);
nor U20854 (N_20854,N_18625,N_16818);
nand U20855 (N_20855,N_15006,N_19906);
xor U20856 (N_20856,N_15550,N_15875);
nor U20857 (N_20857,N_19505,N_16435);
nand U20858 (N_20858,N_15098,N_18483);
or U20859 (N_20859,N_18794,N_18889);
xnor U20860 (N_20860,N_15887,N_16054);
nand U20861 (N_20861,N_18684,N_17800);
and U20862 (N_20862,N_17665,N_18641);
xor U20863 (N_20863,N_15938,N_19007);
xor U20864 (N_20864,N_19594,N_15255);
or U20865 (N_20865,N_16621,N_19921);
or U20866 (N_20866,N_18075,N_17369);
or U20867 (N_20867,N_17548,N_18594);
xor U20868 (N_20868,N_15402,N_19456);
xnor U20869 (N_20869,N_19115,N_18747);
nor U20870 (N_20870,N_16963,N_18409);
nand U20871 (N_20871,N_19696,N_17004);
nand U20872 (N_20872,N_15981,N_15603);
nor U20873 (N_20873,N_15057,N_15427);
nand U20874 (N_20874,N_18751,N_18730);
nor U20875 (N_20875,N_15121,N_19284);
and U20876 (N_20876,N_19367,N_18453);
or U20877 (N_20877,N_18391,N_19942);
nor U20878 (N_20878,N_18003,N_15666);
nor U20879 (N_20879,N_18518,N_19412);
or U20880 (N_20880,N_17812,N_17546);
nand U20881 (N_20881,N_17253,N_19568);
nand U20882 (N_20882,N_19027,N_17772);
nand U20883 (N_20883,N_18875,N_17555);
and U20884 (N_20884,N_17504,N_17173);
or U20885 (N_20885,N_15782,N_19169);
xor U20886 (N_20886,N_18244,N_17728);
nor U20887 (N_20887,N_17947,N_17129);
nor U20888 (N_20888,N_17899,N_18319);
xor U20889 (N_20889,N_19515,N_18185);
nand U20890 (N_20890,N_15492,N_15437);
and U20891 (N_20891,N_17498,N_17245);
and U20892 (N_20892,N_19778,N_18501);
xor U20893 (N_20893,N_19703,N_19805);
xor U20894 (N_20894,N_18100,N_15761);
and U20895 (N_20895,N_18631,N_18508);
nand U20896 (N_20896,N_18247,N_17472);
nand U20897 (N_20897,N_18598,N_15291);
xnor U20898 (N_20898,N_15571,N_16952);
or U20899 (N_20899,N_18530,N_19641);
and U20900 (N_20900,N_19279,N_15919);
and U20901 (N_20901,N_18796,N_16517);
or U20902 (N_20902,N_19066,N_16562);
nand U20903 (N_20903,N_17102,N_18139);
and U20904 (N_20904,N_16364,N_16682);
or U20905 (N_20905,N_19099,N_19959);
nand U20906 (N_20906,N_16470,N_18927);
xnor U20907 (N_20907,N_16659,N_19646);
or U20908 (N_20908,N_18331,N_15227);
nor U20909 (N_20909,N_17396,N_19326);
nand U20910 (N_20910,N_15883,N_18320);
or U20911 (N_20911,N_18777,N_18418);
or U20912 (N_20912,N_18843,N_17896);
xnor U20913 (N_20913,N_17931,N_15676);
or U20914 (N_20914,N_19414,N_15631);
nand U20915 (N_20915,N_19076,N_16136);
or U20916 (N_20916,N_16418,N_18851);
or U20917 (N_20917,N_18773,N_16658);
nor U20918 (N_20918,N_19890,N_18708);
or U20919 (N_20919,N_19720,N_15160);
nor U20920 (N_20920,N_15378,N_17949);
nor U20921 (N_20921,N_17142,N_15587);
and U20922 (N_20922,N_15745,N_16431);
nand U20923 (N_20923,N_19963,N_19593);
and U20924 (N_20924,N_17005,N_19088);
nor U20925 (N_20925,N_18305,N_15967);
nor U20926 (N_20926,N_18970,N_19005);
xnor U20927 (N_20927,N_15426,N_16544);
nand U20928 (N_20928,N_19328,N_16577);
or U20929 (N_20929,N_19527,N_16173);
and U20930 (N_20930,N_17819,N_18756);
nand U20931 (N_20931,N_16776,N_15367);
xor U20932 (N_20932,N_15560,N_15746);
xor U20933 (N_20933,N_16183,N_15954);
or U20934 (N_20934,N_19255,N_17140);
nor U20935 (N_20935,N_15725,N_18924);
or U20936 (N_20936,N_17994,N_16756);
nor U20937 (N_20937,N_16519,N_16829);
or U20938 (N_20938,N_19939,N_19447);
xnor U20939 (N_20939,N_16504,N_15923);
nand U20940 (N_20940,N_18759,N_16412);
or U20941 (N_20941,N_17377,N_18098);
or U20942 (N_20942,N_17057,N_15120);
xnor U20943 (N_20943,N_15163,N_18181);
xnor U20944 (N_20944,N_18573,N_15462);
nand U20945 (N_20945,N_18891,N_16262);
and U20946 (N_20946,N_18271,N_16720);
and U20947 (N_20947,N_15853,N_19911);
or U20948 (N_20948,N_16114,N_15790);
xnor U20949 (N_20949,N_15737,N_19841);
and U20950 (N_20950,N_18572,N_16069);
nand U20951 (N_20951,N_18621,N_19690);
xnor U20952 (N_20952,N_16597,N_19792);
and U20953 (N_20953,N_15548,N_15445);
and U20954 (N_20954,N_18902,N_18752);
or U20955 (N_20955,N_15862,N_19419);
xor U20956 (N_20956,N_15111,N_18158);
and U20957 (N_20957,N_16369,N_15046);
nand U20958 (N_20958,N_18261,N_15632);
nor U20959 (N_20959,N_17512,N_18255);
nand U20960 (N_20960,N_17249,N_19401);
nand U20961 (N_20961,N_19517,N_19174);
or U20962 (N_20962,N_17301,N_18783);
and U20963 (N_20963,N_19725,N_16601);
nand U20964 (N_20964,N_19487,N_15334);
nand U20965 (N_20965,N_19954,N_19674);
nor U20966 (N_20966,N_16942,N_18387);
or U20967 (N_20967,N_15055,N_19541);
and U20968 (N_20968,N_17651,N_16281);
and U20969 (N_20969,N_15200,N_18348);
nand U20970 (N_20970,N_15251,N_15570);
nor U20971 (N_20971,N_18993,N_17435);
xnor U20972 (N_20972,N_15264,N_19002);
or U20973 (N_20973,N_16378,N_19816);
and U20974 (N_20974,N_16623,N_18622);
nor U20975 (N_20975,N_15686,N_15833);
or U20976 (N_20976,N_19321,N_17416);
and U20977 (N_20977,N_17940,N_17264);
nand U20978 (N_20978,N_17815,N_18241);
or U20979 (N_20979,N_16749,N_19033);
nor U20980 (N_20980,N_19260,N_16508);
and U20981 (N_20981,N_19825,N_17952);
and U20982 (N_20982,N_17041,N_16486);
xor U20983 (N_20983,N_17325,N_16610);
nor U20984 (N_20984,N_16052,N_19257);
or U20985 (N_20985,N_15529,N_15896);
nor U20986 (N_20986,N_15004,N_18906);
nand U20987 (N_20987,N_18785,N_15471);
nand U20988 (N_20988,N_17453,N_17414);
or U20989 (N_20989,N_15945,N_16730);
nor U20990 (N_20990,N_19591,N_17020);
and U20991 (N_20991,N_16618,N_18078);
nand U20992 (N_20992,N_15614,N_15440);
nand U20993 (N_20993,N_19451,N_19556);
and U20994 (N_20994,N_19149,N_18946);
nor U20995 (N_20995,N_17562,N_19262);
nor U20996 (N_20996,N_17185,N_15224);
nor U20997 (N_20997,N_18028,N_18163);
or U20998 (N_20998,N_16962,N_15582);
or U20999 (N_20999,N_15879,N_17138);
nor U21000 (N_21000,N_16194,N_17212);
nor U21001 (N_21001,N_15385,N_19726);
nor U21002 (N_21002,N_19891,N_16366);
and U21003 (N_21003,N_19105,N_18619);
nand U21004 (N_21004,N_17862,N_15788);
and U21005 (N_21005,N_18713,N_17893);
xnor U21006 (N_21006,N_15132,N_17986);
nand U21007 (N_21007,N_17860,N_19382);
and U21008 (N_21008,N_18210,N_19479);
nand U21009 (N_21009,N_18963,N_17280);
nand U21010 (N_21010,N_19264,N_16930);
xor U21011 (N_21011,N_16343,N_18233);
nand U21012 (N_21012,N_18725,N_17976);
xor U21013 (N_21013,N_15734,N_19588);
xor U21014 (N_21014,N_19908,N_15230);
nor U21015 (N_21015,N_19387,N_16466);
nand U21016 (N_21016,N_16526,N_19298);
nand U21017 (N_21017,N_15936,N_16537);
nand U21018 (N_21018,N_17033,N_16542);
nor U21019 (N_21019,N_17469,N_18653);
nor U21020 (N_21020,N_17141,N_18010);
nor U21021 (N_21021,N_15889,N_15167);
xor U21022 (N_21022,N_15150,N_18922);
nand U21023 (N_21023,N_19878,N_18257);
or U21024 (N_21024,N_17039,N_17613);
nor U21025 (N_21025,N_16634,N_16921);
and U21026 (N_21026,N_15186,N_17216);
xnor U21027 (N_21027,N_18338,N_19434);
nor U21028 (N_21028,N_17467,N_15153);
or U21029 (N_21029,N_17332,N_18834);
or U21030 (N_21030,N_18592,N_16782);
nand U21031 (N_21031,N_19109,N_16875);
and U21032 (N_21032,N_18683,N_16016);
nand U21033 (N_21033,N_16119,N_19093);
xor U21034 (N_21034,N_18957,N_16615);
nor U21035 (N_21035,N_19622,N_18469);
or U21036 (N_21036,N_17764,N_18135);
or U21037 (N_21037,N_15449,N_18422);
and U21038 (N_21038,N_17655,N_16269);
or U21039 (N_21039,N_19488,N_15249);
nand U21040 (N_21040,N_17205,N_17823);
nand U21041 (N_21041,N_18695,N_15508);
xnor U21042 (N_21042,N_15134,N_15748);
and U21043 (N_21043,N_15330,N_19564);
nand U21044 (N_21044,N_18798,N_15796);
or U21045 (N_21045,N_19032,N_18236);
nor U21046 (N_21046,N_19217,N_17529);
nand U21047 (N_21047,N_19643,N_16552);
nor U21048 (N_21048,N_18633,N_19670);
and U21049 (N_21049,N_15021,N_18249);
or U21050 (N_21050,N_18535,N_16133);
xor U21051 (N_21051,N_18268,N_16631);
or U21052 (N_21052,N_16231,N_19546);
or U21053 (N_21053,N_16085,N_17299);
and U21054 (N_21054,N_17402,N_18310);
or U21055 (N_21055,N_15358,N_15730);
nor U21056 (N_21056,N_15236,N_17192);
and U21057 (N_21057,N_16695,N_17948);
and U21058 (N_21058,N_19691,N_18644);
and U21059 (N_21059,N_16482,N_18239);
and U21060 (N_21060,N_16312,N_19439);
and U21061 (N_21061,N_19585,N_18351);
nand U21062 (N_21062,N_17939,N_16507);
xnor U21063 (N_21063,N_18177,N_18000);
nand U21064 (N_21064,N_17663,N_18465);
xnor U21065 (N_21065,N_15495,N_19228);
and U21066 (N_21066,N_16578,N_19458);
nor U21067 (N_21067,N_16104,N_16096);
nor U21068 (N_21068,N_19337,N_16549);
nand U21069 (N_21069,N_19013,N_19898);
or U21070 (N_21070,N_15636,N_19304);
nor U21071 (N_21071,N_19461,N_16082);
nor U21072 (N_21072,N_15295,N_18471);
nand U21073 (N_21073,N_19910,N_18648);
nand U21074 (N_21074,N_17700,N_18861);
xor U21075 (N_21075,N_15634,N_19087);
xnor U21076 (N_21076,N_16244,N_17902);
or U21077 (N_21077,N_17751,N_16572);
or U21078 (N_21078,N_18363,N_16335);
and U21079 (N_21079,N_16724,N_15611);
and U21080 (N_21080,N_18477,N_18292);
or U21081 (N_21081,N_18491,N_16535);
and U21082 (N_21082,N_17306,N_16556);
and U21083 (N_21083,N_15268,N_15643);
or U21084 (N_21084,N_18222,N_17916);
or U21085 (N_21085,N_19165,N_16761);
and U21086 (N_21086,N_19042,N_16897);
nor U21087 (N_21087,N_18243,N_15243);
and U21088 (N_21088,N_17450,N_18435);
xnor U21089 (N_21089,N_16734,N_19716);
xor U21090 (N_21090,N_19970,N_19912);
nand U21091 (N_21091,N_18322,N_16967);
nor U21092 (N_21092,N_17136,N_16547);
nor U21093 (N_21093,N_15373,N_16816);
or U21094 (N_21094,N_18053,N_18764);
and U21095 (N_21095,N_18051,N_17682);
nor U21096 (N_21096,N_16143,N_19914);
nand U21097 (N_21097,N_16278,N_19335);
or U21098 (N_21098,N_16538,N_16277);
nand U21099 (N_21099,N_19026,N_18855);
or U21100 (N_21100,N_15656,N_19853);
nand U21101 (N_21101,N_18803,N_15784);
and U21102 (N_21102,N_19846,N_15271);
and U21103 (N_21103,N_17166,N_19885);
or U21104 (N_21104,N_18772,N_15412);
nand U21105 (N_21105,N_17935,N_17874);
or U21106 (N_21106,N_19773,N_18937);
and U21107 (N_21107,N_18766,N_17290);
nand U21108 (N_21108,N_19403,N_19509);
or U21109 (N_21109,N_19826,N_19359);
nand U21110 (N_21110,N_15558,N_15423);
nor U21111 (N_21111,N_18897,N_18008);
xor U21112 (N_21112,N_16580,N_15564);
and U21113 (N_21113,N_18995,N_16664);
nand U21114 (N_21114,N_16349,N_19695);
nand U21115 (N_21115,N_19477,N_17790);
or U21116 (N_21116,N_17549,N_16886);
nor U21117 (N_21117,N_16255,N_18728);
nand U21118 (N_21118,N_17213,N_15192);
nor U21119 (N_21119,N_16959,N_16204);
nand U21120 (N_21120,N_16731,N_15410);
or U21121 (N_21121,N_16655,N_19068);
nand U21122 (N_21122,N_19219,N_16005);
or U21123 (N_21123,N_18657,N_19582);
nand U21124 (N_21124,N_19986,N_17333);
nand U21125 (N_21125,N_16567,N_18150);
xor U21126 (N_21126,N_16898,N_17884);
nand U21127 (N_21127,N_19236,N_19481);
nor U21128 (N_21128,N_15409,N_15178);
and U21129 (N_21129,N_16795,N_15609);
nand U21130 (N_21130,N_17220,N_17957);
nand U21131 (N_21131,N_19020,N_18703);
nor U21132 (N_21132,N_17656,N_19551);
or U21133 (N_21133,N_19290,N_19168);
nor U21134 (N_21134,N_18885,N_16070);
nand U21135 (N_21135,N_18896,N_17801);
or U21136 (N_21136,N_16859,N_19743);
and U21137 (N_21137,N_18951,N_19729);
nand U21138 (N_21138,N_15897,N_15240);
or U21139 (N_21139,N_17254,N_15902);
or U21140 (N_21140,N_18971,N_17079);
nor U21141 (N_21141,N_15687,N_18925);
or U21142 (N_21142,N_16459,N_16697);
nand U21143 (N_21143,N_19580,N_15181);
nand U21144 (N_21144,N_19292,N_16046);
nand U21145 (N_21145,N_15661,N_15105);
or U21146 (N_21146,N_15683,N_19790);
nand U21147 (N_21147,N_17398,N_15503);
or U21148 (N_21148,N_18959,N_17324);
or U21149 (N_21149,N_17413,N_16912);
and U21150 (N_21150,N_19562,N_15061);
xnor U21151 (N_21151,N_17506,N_18203);
nor U21152 (N_21152,N_15886,N_19409);
nor U21153 (N_21153,N_16212,N_18111);
and U21154 (N_21154,N_15327,N_17761);
and U21155 (N_21155,N_16843,N_15839);
and U21156 (N_21156,N_16936,N_18513);
xnor U21157 (N_21157,N_16344,N_18282);
nor U21158 (N_21158,N_15015,N_17069);
and U21159 (N_21159,N_17685,N_15392);
nor U21160 (N_21160,N_17113,N_19283);
nor U21161 (N_21161,N_15783,N_15370);
or U21162 (N_21162,N_18626,N_19771);
xor U21163 (N_21163,N_15626,N_17315);
xor U21164 (N_21164,N_18517,N_19226);
and U21165 (N_21165,N_17730,N_16607);
nor U21166 (N_21166,N_17171,N_19928);
nor U21167 (N_21167,N_17640,N_17693);
nor U21168 (N_21168,N_16029,N_16159);
nor U21169 (N_21169,N_17461,N_17908);
nand U21170 (N_21170,N_16922,N_19041);
or U21171 (N_21171,N_18809,N_18289);
or U21172 (N_21172,N_17666,N_18909);
nor U21173 (N_21173,N_16283,N_18264);
xnor U21174 (N_21174,N_18749,N_18191);
and U21175 (N_21175,N_15799,N_15881);
and U21176 (N_21176,N_16704,N_15109);
and U21177 (N_21177,N_19602,N_16155);
and U21178 (N_21178,N_15675,N_19677);
nand U21179 (N_21179,N_18220,N_19128);
or U21180 (N_21180,N_17258,N_19884);
or U21181 (N_21181,N_15569,N_17226);
nor U21182 (N_21182,N_16867,N_18229);
nor U21183 (N_21183,N_16449,N_19711);
nor U21184 (N_21184,N_16805,N_19017);
xnor U21185 (N_21185,N_16890,N_17151);
nor U21186 (N_21186,N_15201,N_19277);
nand U21187 (N_21187,N_17592,N_19968);
nor U21188 (N_21188,N_17499,N_17281);
or U21189 (N_21189,N_17270,N_19472);
and U21190 (N_21190,N_18019,N_19492);
and U21191 (N_21191,N_17980,N_16463);
nand U21192 (N_21192,N_15131,N_16135);
nand U21193 (N_21193,N_17574,N_18383);
and U21194 (N_21194,N_19895,N_17451);
and U21195 (N_21195,N_16590,N_18012);
xor U21196 (N_21196,N_18839,N_19577);
xnor U21197 (N_21197,N_16334,N_18646);
nand U21198 (N_21198,N_15420,N_15104);
nand U21199 (N_21199,N_17294,N_18494);
and U21200 (N_21200,N_16333,N_15156);
nand U21201 (N_21201,N_15793,N_17300);
nor U21202 (N_21202,N_16290,N_16146);
xnor U21203 (N_21203,N_15473,N_19231);
nand U21204 (N_21204,N_15394,N_19098);
nor U21205 (N_21205,N_18591,N_16943);
and U21206 (N_21206,N_19345,N_16084);
or U21207 (N_21207,N_16026,N_18022);
nand U21208 (N_21208,N_16109,N_17737);
xnor U21209 (N_21209,N_19181,N_15530);
nor U21210 (N_21210,N_18427,N_18640);
or U21211 (N_21211,N_16156,N_15523);
nor U21212 (N_21212,N_15778,N_17780);
xor U21213 (N_21213,N_17231,N_18821);
nor U21214 (N_21214,N_19982,N_18526);
nand U21215 (N_21215,N_18707,N_16592);
nand U21216 (N_21216,N_19144,N_15482);
or U21217 (N_21217,N_17071,N_17383);
nor U21218 (N_21218,N_18146,N_18308);
nor U21219 (N_21219,N_16024,N_19120);
nand U21220 (N_21220,N_15549,N_19015);
nand U21221 (N_21221,N_17912,N_18546);
xnor U21222 (N_21222,N_16745,N_15689);
xnor U21223 (N_21223,N_17719,N_15772);
or U21224 (N_21224,N_17443,N_16727);
nor U21225 (N_21225,N_15244,N_15083);
xnor U21226 (N_21226,N_17975,N_16773);
nand U21227 (N_21227,N_18914,N_19234);
and U21228 (N_21228,N_15682,N_18507);
nor U21229 (N_21229,N_16233,N_19676);
nand U21230 (N_21230,N_18878,N_15577);
nor U21231 (N_21231,N_17973,N_19589);
and U21232 (N_21232,N_16210,N_18499);
or U21233 (N_21233,N_18825,N_19770);
or U21234 (N_21234,N_17596,N_19897);
nand U21235 (N_21235,N_19889,N_16428);
and U21236 (N_21236,N_17228,N_15998);
nor U21237 (N_21237,N_16060,N_16310);
nor U21238 (N_21238,N_17064,N_17698);
and U21239 (N_21239,N_16540,N_19524);
and U21240 (N_21240,N_17740,N_16321);
and U21241 (N_21241,N_16358,N_16603);
and U21242 (N_21242,N_18522,N_15161);
xnor U21243 (N_21243,N_15817,N_15811);
nor U21244 (N_21244,N_18693,N_18988);
nand U21245 (N_21245,N_15974,N_17006);
nand U21246 (N_21246,N_18627,N_16073);
or U21247 (N_21247,N_17830,N_15293);
xnor U21248 (N_21248,N_19990,N_16545);
nor U21249 (N_21249,N_17381,N_16758);
or U21250 (N_21250,N_19712,N_16995);
nor U21251 (N_21251,N_15479,N_18059);
nand U21252 (N_21252,N_18699,N_16457);
nor U21253 (N_21253,N_16229,N_18154);
and U21254 (N_21254,N_17296,N_19924);
or U21255 (N_21255,N_19048,N_16833);
or U21256 (N_21256,N_15991,N_19089);
or U21257 (N_21257,N_19705,N_17345);
nand U21258 (N_21258,N_17745,N_19633);
and U21259 (N_21259,N_18001,N_17510);
nor U21260 (N_21260,N_17047,N_19860);
nor U21261 (N_21261,N_16490,N_18488);
nor U21262 (N_21262,N_19625,N_15519);
or U21263 (N_21263,N_18912,N_17934);
nand U21264 (N_21264,N_16792,N_18705);
or U21265 (N_21265,N_17678,N_19529);
nor U21266 (N_21266,N_16855,N_18114);
and U21267 (N_21267,N_15279,N_17488);
nor U21268 (N_21268,N_19178,N_19788);
nand U21269 (N_21269,N_19926,N_19011);
xor U21270 (N_21270,N_18206,N_18697);
nor U21271 (N_21271,N_18107,N_15842);
nand U21272 (N_21272,N_15214,N_19448);
or U21273 (N_21273,N_19558,N_18188);
nor U21274 (N_21274,N_17530,N_16670);
xor U21275 (N_21275,N_19952,N_16476);
xor U21276 (N_21276,N_18354,N_19737);
nand U21277 (N_21277,N_19489,N_16871);
nand U21278 (N_21278,N_19769,N_17364);
nand U21279 (N_21279,N_16227,N_19156);
xor U21280 (N_21280,N_19576,N_19266);
xnor U21281 (N_21281,N_19444,N_17370);
xnor U21282 (N_21282,N_16960,N_18750);
and U21283 (N_21283,N_16853,N_19379);
and U21284 (N_21284,N_19362,N_19554);
or U21285 (N_21285,N_16666,N_15059);
and U21286 (N_21286,N_15203,N_16561);
nand U21287 (N_21287,N_19374,N_19369);
xnor U21288 (N_21288,N_16122,N_19407);
and U21289 (N_21289,N_17144,N_19574);
nor U21290 (N_21290,N_18768,N_16520);
nor U21291 (N_21291,N_15007,N_15074);
nor U21292 (N_21292,N_17159,N_16402);
or U21293 (N_21293,N_18237,N_15518);
and U21294 (N_21294,N_19768,N_15660);
and U21295 (N_21295,N_15939,N_15568);
xor U21296 (N_21296,N_19774,N_18276);
or U21297 (N_21297,N_16735,N_15851);
or U21298 (N_21298,N_19973,N_15716);
nor U21299 (N_21299,N_19164,N_16909);
xor U21300 (N_21300,N_17327,N_17534);
xor U21301 (N_21301,N_17901,N_17358);
and U21302 (N_21302,N_15835,N_15873);
nand U21303 (N_21303,N_16256,N_17701);
nand U21304 (N_21304,N_19782,N_18311);
or U21305 (N_21305,N_17056,N_19341);
or U21306 (N_21306,N_15362,N_16799);
nand U21307 (N_21307,N_16844,N_16285);
or U21308 (N_21308,N_19006,N_17987);
xnor U21309 (N_21309,N_18888,N_18084);
xor U21310 (N_21310,N_16673,N_18168);
nand U21311 (N_21311,N_19392,N_17405);
nand U21312 (N_21312,N_15470,N_18581);
and U21313 (N_21313,N_16982,N_17816);
nor U21314 (N_21314,N_15248,N_17059);
nor U21315 (N_21315,N_15211,N_18275);
and U21316 (N_21316,N_17953,N_15466);
and U21317 (N_21317,N_17055,N_15965);
xor U21318 (N_21318,N_16188,N_17516);
and U21319 (N_21319,N_19947,N_16447);
and U21320 (N_21320,N_18149,N_15103);
or U21321 (N_21321,N_15763,N_18907);
or U21322 (N_21322,N_16676,N_16252);
nand U21323 (N_21323,N_17573,N_19389);
xnor U21324 (N_21324,N_19235,N_19102);
nand U21325 (N_21325,N_17184,N_18199);
nand U21326 (N_21326,N_15108,N_15069);
xor U21327 (N_21327,N_18020,N_15658);
nor U21328 (N_21328,N_16007,N_15854);
or U21329 (N_21329,N_15496,N_16313);
nor U21330 (N_21330,N_15493,N_17148);
nand U21331 (N_21331,N_19640,N_18467);
nor U21332 (N_21332,N_19665,N_17582);
and U21333 (N_21333,N_18353,N_19964);
nand U21334 (N_21334,N_16391,N_16729);
nand U21335 (N_21335,N_18416,N_15208);
nand U21336 (N_21336,N_16715,N_17598);
nand U21337 (N_21337,N_18145,N_16249);
and U21338 (N_21338,N_18550,N_18402);
xnor U21339 (N_21339,N_16977,N_15464);
xnor U21340 (N_21340,N_18429,N_15433);
xnor U21341 (N_21341,N_17298,N_18032);
or U21342 (N_21342,N_15499,N_16692);
and U21343 (N_21343,N_15743,N_15528);
nand U21344 (N_21344,N_17086,N_15733);
xnor U21345 (N_21345,N_18470,N_15619);
nand U21346 (N_21346,N_15602,N_16907);
nand U21347 (N_21347,N_16743,N_15651);
or U21348 (N_21348,N_18091,N_16458);
nand U21349 (N_21349,N_18424,N_16221);
and U21350 (N_21350,N_16998,N_17943);
nand U21351 (N_21351,N_17037,N_15864);
or U21352 (N_21352,N_19535,N_16604);
nor U21353 (N_21353,N_17601,N_19946);
nand U21354 (N_21354,N_19157,N_18106);
and U21355 (N_21355,N_16065,N_19127);
xor U21356 (N_21356,N_17349,N_17022);
nand U21357 (N_21357,N_16716,N_19919);
and U21358 (N_21358,N_17183,N_16838);
xor U21359 (N_21359,N_16531,N_17417);
xor U21360 (N_21360,N_16801,N_18076);
nand U21361 (N_21361,N_19383,N_19192);
and U21362 (N_21362,N_19565,N_15223);
or U21363 (N_21363,N_18323,N_15076);
and U21364 (N_21364,N_16403,N_19678);
or U21365 (N_21365,N_19025,N_16559);
nand U21366 (N_21366,N_17631,N_15266);
xnor U21367 (N_21367,N_15610,N_18567);
and U21368 (N_21368,N_19899,N_18610);
or U21369 (N_21369,N_17111,N_18007);
nand U21370 (N_21370,N_15847,N_15966);
xnor U21371 (N_21371,N_17900,N_17735);
nor U21372 (N_21372,N_18850,N_18714);
xnor U21373 (N_21373,N_16492,N_17314);
or U21374 (N_21374,N_16118,N_19916);
and U21375 (N_21375,N_17898,N_15113);
or U21376 (N_21376,N_15969,N_16257);
and U21377 (N_21377,N_17353,N_17602);
xor U21378 (N_21378,N_18663,N_15583);
nand U21379 (N_21379,N_18140,N_19784);
xor U21380 (N_21380,N_19129,N_15436);
or U21381 (N_21381,N_16599,N_15089);
xnor U21382 (N_21382,N_19902,N_18316);
xnor U21383 (N_21383,N_19348,N_15390);
nor U21384 (N_21384,N_17612,N_16381);
and U21385 (N_21385,N_17736,N_19191);
nor U21386 (N_21386,N_15102,N_15925);
xnor U21387 (N_21387,N_17191,N_15029);
nor U21388 (N_21388,N_15696,N_19997);
nor U21389 (N_21389,N_15578,N_15754);
and U21390 (N_21390,N_17329,N_18629);
nand U21391 (N_21391,N_19091,N_19467);
and U21392 (N_21392,N_17926,N_17917);
nor U21393 (N_21393,N_17165,N_17645);
nor U21394 (N_21394,N_17992,N_18716);
and U21395 (N_21395,N_17524,N_19285);
or U21396 (N_21396,N_16303,N_15432);
xor U21397 (N_21397,N_19072,N_15641);
or U21398 (N_21398,N_15335,N_15459);
and U21399 (N_21399,N_16008,N_16966);
and U21400 (N_21400,N_15253,N_16074);
nand U21401 (N_21401,N_16823,N_19334);
or U21402 (N_21402,N_15767,N_19429);
or U21403 (N_21403,N_17961,N_18049);
nand U21404 (N_21404,N_15584,N_15171);
and U21405 (N_21405,N_15554,N_16783);
xor U21406 (N_21406,N_18904,N_15804);
and U21407 (N_21407,N_15009,N_19722);
or U21408 (N_21408,N_18590,N_17440);
nand U21409 (N_21409,N_19466,N_17072);
and U21410 (N_21410,N_19586,N_19506);
nand U21411 (N_21411,N_19896,N_16654);
or U21412 (N_21412,N_19044,N_18603);
nand U21413 (N_21413,N_17105,N_15119);
and U21414 (N_21414,N_19522,N_19750);
nand U21415 (N_21415,N_17081,N_15655);
nand U21416 (N_21416,N_18854,N_17496);
xnor U21417 (N_21417,N_16978,N_18004);
and U21418 (N_21418,N_17576,N_15387);
xor U21419 (N_21419,N_19459,N_18327);
nand U21420 (N_21420,N_15532,N_15155);
or U21421 (N_21421,N_16093,N_17580);
xor U21422 (N_21422,N_19783,N_17052);
and U21423 (N_21423,N_16740,N_16992);
nor U21424 (N_21424,N_18786,N_18523);
or U21425 (N_21425,N_18562,N_18426);
and U21426 (N_21426,N_15544,N_18941);
nand U21427 (N_21427,N_16821,N_16213);
or U21428 (N_21428,N_17230,N_19981);
nor U21429 (N_21429,N_15715,N_18795);
or U21430 (N_21430,N_18739,N_17458);
nor U21431 (N_21431,N_18133,N_17095);
nor U21432 (N_21432,N_19777,N_19360);
and U21433 (N_21433,N_19273,N_19153);
and U21434 (N_21434,N_16462,N_15510);
and U21435 (N_21435,N_19314,N_19539);
nand U21436 (N_21436,N_15254,N_15379);
xnor U21437 (N_21437,N_17261,N_17950);
xor U21438 (N_21438,N_19425,N_16373);
nand U21439 (N_21439,N_17044,N_17793);
or U21440 (N_21440,N_16737,N_16090);
nor U21441 (N_21441,N_16134,N_19065);
nor U21442 (N_21442,N_19617,N_18623);
nor U21443 (N_21443,N_15922,N_16707);
or U21444 (N_21444,N_16386,N_16746);
nor U21445 (N_21445,N_19137,N_18052);
nand U21446 (N_21446,N_18077,N_18397);
nor U21447 (N_21447,N_19338,N_16824);
and U21448 (N_21448,N_18152,N_17517);
or U21449 (N_21449,N_17275,N_16103);
nor U21450 (N_21450,N_17194,N_15062);
or U21451 (N_21451,N_19626,N_18090);
nor U21452 (N_21452,N_18274,N_19270);
or U21453 (N_21453,N_15494,N_18017);
or U21454 (N_21454,N_17608,N_17605);
and U21455 (N_21455,N_17589,N_15757);
and U21456 (N_21456,N_17025,N_15187);
and U21457 (N_21457,N_15955,N_18246);
or U21458 (N_21458,N_15509,N_16185);
nand U21459 (N_21459,N_18404,N_18723);
nor U21460 (N_21460,N_15288,N_16465);
or U21461 (N_21461,N_16405,N_15629);
and U21462 (N_21462,N_18511,N_19745);
nand U21463 (N_21463,N_15913,N_15891);
nor U21464 (N_21464,N_16376,N_15498);
xnor U21465 (N_21465,N_16245,N_16533);
nor U21466 (N_21466,N_17837,N_17984);
nor U21467 (N_21467,N_16524,N_16732);
and U21468 (N_21468,N_19396,N_16301);
nor U21469 (N_21469,N_15507,N_18895);
xor U21470 (N_21470,N_17237,N_19503);
nand U21471 (N_21471,N_16860,N_15270);
xnor U21472 (N_21472,N_19393,N_19944);
xnor U21473 (N_21473,N_15915,N_19468);
or U21474 (N_21474,N_19630,N_15174);
or U21475 (N_21475,N_16107,N_18265);
xnor U21476 (N_21476,N_17125,N_16261);
and U21477 (N_21477,N_19795,N_17482);
nor U21478 (N_21478,N_17611,N_19639);
and U21479 (N_21479,N_15867,N_18215);
nor U21480 (N_21480,N_17090,N_19927);
xor U21481 (N_21481,N_15744,N_18344);
nor U21482 (N_21482,N_18868,N_19741);
and U21483 (N_21483,N_15300,N_16750);
and U21484 (N_21484,N_18998,N_18187);
and U21485 (N_21485,N_19103,N_17880);
or U21486 (N_21486,N_17432,N_18108);
or U21487 (N_21487,N_15858,N_18539);
or U21488 (N_21488,N_15950,N_19110);
nor U21489 (N_21489,N_18939,N_18975);
xnor U21490 (N_21490,N_15789,N_16394);
nand U21491 (N_21491,N_19599,N_17223);
xor U21492 (N_21492,N_19272,N_17660);
and U21493 (N_21493,N_19218,N_16234);
nor U21494 (N_21494,N_19957,N_15042);
or U21495 (N_21495,N_16208,N_19544);
or U21496 (N_21496,N_19427,N_16475);
nand U21497 (N_21497,N_16328,N_15589);
nand U21498 (N_21498,N_18681,N_19311);
xor U21499 (N_21499,N_16946,N_19651);
xnor U21500 (N_21500,N_18717,N_19949);
nand U21501 (N_21501,N_15774,N_19779);
xnor U21502 (N_21502,N_15312,N_15366);
nand U21503 (N_21503,N_19941,N_16845);
or U21504 (N_21504,N_19751,N_16320);
or U21505 (N_21505,N_16888,N_17400);
xnor U21506 (N_21506,N_18642,N_16570);
nand U21507 (N_21507,N_18921,N_19278);
nor U21508 (N_21508,N_17376,N_17179);
nand U21509 (N_21509,N_15779,N_19575);
nand U21510 (N_21510,N_18057,N_17276);
nor U21511 (N_21511,N_16393,N_16964);
nand U21512 (N_21512,N_18484,N_16317);
or U21513 (N_21513,N_18556,N_17883);
xnor U21514 (N_21514,N_16521,N_15880);
nor U21515 (N_21515,N_18584,N_15630);
nand U21516 (N_21516,N_15305,N_18964);
nand U21517 (N_21517,N_17082,N_18116);
or U21518 (N_21518,N_18192,N_19950);
nor U21519 (N_21519,N_17334,N_18408);
and U21520 (N_21520,N_16392,N_15822);
xnor U21521 (N_21521,N_19975,N_17074);
nand U21522 (N_21522,N_16939,N_17540);
or U21523 (N_21523,N_16885,N_16717);
and U21524 (N_21524,N_15979,N_18991);
nor U21525 (N_21525,N_19636,N_19863);
xnor U21526 (N_21526,N_15340,N_18687);
nand U21527 (N_21527,N_16452,N_18574);
nor U21528 (N_21528,N_16158,N_15501);
xnor U21529 (N_21529,N_19404,N_15776);
xor U21530 (N_21530,N_15595,N_18103);
nor U21531 (N_21531,N_16710,N_18858);
nand U21532 (N_21532,N_17866,N_18378);
and U21533 (N_21533,N_17686,N_15724);
or U21534 (N_21534,N_18913,N_15328);
and U21535 (N_21535,N_15917,N_18493);
xnor U21536 (N_21536,N_18411,N_18131);
xor U21537 (N_21537,N_18290,N_15908);
nor U21538 (N_21538,N_18710,N_16448);
nor U21539 (N_21539,N_17188,N_15064);
and U21540 (N_21540,N_19980,N_19440);
nor U21541 (N_21541,N_19728,N_15475);
nand U21542 (N_21542,N_18611,N_19715);
xor U21543 (N_21543,N_18595,N_17103);
and U21544 (N_21544,N_18326,N_18844);
nor U21545 (N_21545,N_16130,N_19829);
nor U21546 (N_21546,N_18672,N_17667);
xnor U21547 (N_21547,N_18731,N_15786);
nor U21548 (N_21548,N_17098,N_16414);
and U21549 (N_21549,N_18549,N_18183);
nor U21550 (N_21550,N_19114,N_18540);
or U21551 (N_21551,N_19719,N_19563);
or U21552 (N_21552,N_15199,N_16163);
nand U21553 (N_21553,N_17634,N_15551);
or U21554 (N_21554,N_16527,N_15444);
or U21555 (N_21555,N_19965,N_16856);
nor U21556 (N_21556,N_17401,N_19871);
xnor U21557 (N_21557,N_19442,N_18658);
and U21558 (N_21558,N_19062,N_15707);
xor U21559 (N_21559,N_16774,N_19207);
nand U21560 (N_21560,N_18083,N_18423);
nor U21561 (N_21561,N_18618,N_15397);
xor U21562 (N_21562,N_18817,N_19332);
nor U21563 (N_21563,N_18473,N_18245);
xnor U21564 (N_21564,N_18532,N_18434);
nand U21565 (N_21565,N_18548,N_19694);
and U21566 (N_21566,N_19922,N_17877);
nand U21567 (N_21567,N_19312,N_16086);
nand U21568 (N_21568,N_18037,N_16439);
and U21569 (N_21569,N_15468,N_15310);
or U21570 (N_21570,N_15540,N_19424);
or U21571 (N_21571,N_16566,N_16100);
or U21572 (N_21572,N_15959,N_15115);
nand U21573 (N_21573,N_17599,N_18870);
nor U21574 (N_21574,N_16738,N_17646);
or U21575 (N_21575,N_19814,N_17920);
xor U21576 (N_21576,N_18685,N_17003);
and U21577 (N_21577,N_15640,N_18589);
nor U21578 (N_21578,N_16330,N_18412);
nor U21579 (N_21579,N_19628,N_16467);
nand U21580 (N_21580,N_18173,N_17944);
nor U21581 (N_21581,N_19862,N_18162);
xor U21582 (N_21582,N_16863,N_16067);
nor U21583 (N_21583,N_19893,N_17514);
and U21584 (N_21584,N_16780,N_15712);
nor U21585 (N_21585,N_18691,N_16713);
nor U21586 (N_21586,N_16575,N_19756);
nand U21587 (N_21587,N_15299,N_18789);
xor U21588 (N_21588,N_15283,N_18968);
nand U21589 (N_21589,N_15206,N_17043);
or U21590 (N_21590,N_16605,N_15552);
xor U21591 (N_21591,N_15606,N_16323);
nand U21592 (N_21592,N_18238,N_19672);
and U21593 (N_21593,N_17389,N_17297);
or U21594 (N_21594,N_17848,N_19872);
nand U21595 (N_21595,N_17087,N_16690);
and U21596 (N_21596,N_16223,N_18669);
and U21597 (N_21597,N_16751,N_15139);
and U21598 (N_21598,N_18745,N_15117);
nand U21599 (N_21599,N_19707,N_19760);
or U21600 (N_21600,N_16736,N_15313);
or U21601 (N_21601,N_18088,N_15350);
and U21602 (N_21602,N_18334,N_17565);
or U21603 (N_21603,N_16077,N_19661);
xor U21604 (N_21604,N_19638,N_15193);
or U21605 (N_21605,N_19767,N_19204);
nand U21606 (N_21606,N_17121,N_16518);
nor U21607 (N_21607,N_19397,N_17527);
nand U21608 (N_21608,N_18620,N_16468);
xnor U21609 (N_21609,N_16709,N_15650);
or U21610 (N_21610,N_19333,N_17032);
xor U21611 (N_21611,N_19747,N_19214);
and U21612 (N_21612,N_15276,N_19560);
nor U21613 (N_21613,N_18776,N_15228);
and U21614 (N_21614,N_15762,N_18212);
and U21615 (N_21615,N_18346,N_17705);
and U21616 (N_21616,N_15234,N_16189);
or U21617 (N_21617,N_15127,N_18030);
xnor U21618 (N_21618,N_15099,N_16754);
nand U21619 (N_21619,N_18721,N_17824);
or U21620 (N_21620,N_15874,N_16648);
and U21621 (N_21621,N_18399,N_15077);
nand U21622 (N_21622,N_18916,N_15408);
nand U21623 (N_21623,N_16794,N_17262);
nor U21624 (N_21624,N_18272,N_17475);
xor U21625 (N_21625,N_19869,N_15940);
xnor U21626 (N_21626,N_16698,N_18137);
nor U21627 (N_21627,N_19748,N_15894);
xor U21628 (N_21628,N_16822,N_16595);
nand U21629 (N_21629,N_15246,N_18529);
and U21630 (N_21630,N_17114,N_19989);
nand U21631 (N_21631,N_15026,N_15086);
nand U21632 (N_21632,N_17107,N_17712);
nand U21633 (N_21633,N_17027,N_19875);
nor U21634 (N_21634,N_19754,N_15344);
xnor U21635 (N_21635,N_15403,N_16894);
and U21636 (N_21636,N_18349,N_15325);
nor U21637 (N_21637,N_19142,N_17092);
nand U21638 (N_21638,N_18994,N_16528);
nor U21639 (N_21639,N_17326,N_18720);
nand U21640 (N_21640,N_17911,N_16892);
or U21641 (N_21641,N_15339,N_15406);
xor U21642 (N_21642,N_17420,N_15986);
nor U21643 (N_21643,N_17304,N_18400);
nand U21644 (N_21644,N_15037,N_16814);
or U21645 (N_21645,N_17375,N_18050);
and U21646 (N_21646,N_16506,N_18021);
xnor U21647 (N_21647,N_15033,N_15599);
nand U21648 (N_21648,N_15885,N_17836);
nand U21649 (N_21649,N_19578,N_19632);
xor U21650 (N_21650,N_15463,N_18381);
nand U21651 (N_21651,N_17726,N_17490);
xnor U21652 (N_21652,N_19813,N_18607);
nand U21653 (N_21653,N_16883,N_18712);
and U21654 (N_21654,N_16176,N_16396);
xor U21655 (N_21655,N_15659,N_18996);
or U21656 (N_21656,N_19861,N_19197);
or U21657 (N_21657,N_18312,N_15834);
nor U21658 (N_21658,N_16622,N_18579);
or U21659 (N_21659,N_17821,N_16924);
xnor U21660 (N_21660,N_19446,N_17998);
nor U21661 (N_21661,N_15758,N_16644);
or U21662 (N_21662,N_17723,N_19473);
and U21663 (N_21663,N_18608,N_16274);
xnor U21664 (N_21664,N_17889,N_19731);
nor U21665 (N_21665,N_16849,N_17647);
nand U21666 (N_21666,N_18675,N_16179);
and U21667 (N_21667,N_19649,N_18757);
xnor U21668 (N_21668,N_19693,N_18480);
nor U21669 (N_21669,N_15003,N_19402);
xor U21670 (N_21670,N_15616,N_18536);
nand U21671 (N_21671,N_17743,N_15679);
and U21672 (N_21672,N_15256,N_19667);
xor U21673 (N_21673,N_19525,N_19945);
xnor U21674 (N_21674,N_15292,N_16662);
and U21675 (N_21675,N_16477,N_16835);
nand U21676 (N_21676,N_17434,N_19545);
and U21677 (N_21677,N_17741,N_16363);
or U21678 (N_21678,N_15314,N_16276);
xor U21679 (N_21679,N_15196,N_19252);
or U21680 (N_21680,N_15023,N_16788);
or U21681 (N_21681,N_18159,N_17583);
and U21682 (N_21682,N_19557,N_19179);
and U21683 (N_21683,N_17522,N_19799);
xnor U21684 (N_21684,N_19978,N_18676);
and U21685 (N_21685,N_15563,N_15138);
and U21686 (N_21686,N_17341,N_17863);
nand U21687 (N_21687,N_17233,N_15135);
nor U21688 (N_21688,N_17607,N_18047);
nand U21689 (N_21689,N_15035,N_15212);
nor U21690 (N_21690,N_18045,N_18972);
nand U21691 (N_21691,N_16712,N_16971);
nor U21692 (N_21692,N_15184,N_16360);
nand U21693 (N_21693,N_15222,N_19881);
and U21694 (N_21694,N_15043,N_17445);
or U21695 (N_21695,N_18985,N_16958);
and U21696 (N_21696,N_16125,N_18283);
xnor U21697 (N_21697,N_17106,N_19059);
or U21698 (N_21698,N_18029,N_16413);
and U21699 (N_21699,N_18928,N_16356);
and U21700 (N_21700,N_18765,N_16803);
xor U21701 (N_21701,N_16582,N_19538);
or U21702 (N_21702,N_18832,N_15513);
and U21703 (N_21703,N_16636,N_19648);
nor U21704 (N_21704,N_16827,N_16267);
xor U21705 (N_21705,N_15398,N_18094);
nor U21706 (N_21706,N_19096,N_15713);
xor U21707 (N_21707,N_17018,N_19937);
nand U21708 (N_21708,N_19249,N_15993);
nor U21709 (N_21709,N_15252,N_18700);
and U21710 (N_21710,N_17373,N_16765);
and U21711 (N_21711,N_18466,N_17283);
or U21712 (N_21712,N_15752,N_18295);
nor U21713 (N_21713,N_18390,N_15050);
or U21714 (N_21714,N_19548,N_18624);
and U21715 (N_21715,N_19699,N_18384);
xnor U21716 (N_21716,N_16711,N_19936);
or U21717 (N_21717,N_16190,N_19796);
nor U21718 (N_21718,N_18893,N_19247);
nand U21719 (N_21719,N_19083,N_17575);
nor U21720 (N_21720,N_18060,N_18455);
or U21721 (N_21721,N_18819,N_16925);
nor U21722 (N_21722,N_19496,N_15188);
or U21723 (N_21723,N_17307,N_17133);
nor U21724 (N_21724,N_16240,N_19010);
and U21725 (N_21725,N_19856,N_15505);
nor U21726 (N_21726,N_15983,N_19844);
or U21727 (N_21727,N_15982,N_15516);
xor U21728 (N_21728,N_18407,N_15011);
nor U21729 (N_21729,N_16175,N_16638);
nand U21730 (N_21730,N_17615,N_15159);
nand U21731 (N_21731,N_19470,N_17462);
and U21732 (N_21732,N_18557,N_18942);
nand U21733 (N_21733,N_17131,N_19301);
and U21734 (N_21734,N_18497,N_18279);
nand U21735 (N_21735,N_15664,N_19043);
xor U21736 (N_21736,N_19107,N_15740);
or U21737 (N_21737,N_18033,N_18960);
and U21738 (N_21738,N_18887,N_17257);
nor U21739 (N_21739,N_19190,N_15781);
xnor U21740 (N_21740,N_16055,N_18575);
nor U21741 (N_21741,N_16497,N_19753);
xor U21742 (N_21742,N_15798,N_19809);
nor U21743 (N_21743,N_15846,N_16779);
nand U21744 (N_21744,N_15361,N_19406);
nand U21745 (N_21745,N_17181,N_18882);
nor U21746 (N_21746,N_19552,N_19925);
and U21747 (N_21747,N_19123,N_15036);
nor U21748 (N_21748,N_15975,N_16226);
and U21749 (N_21749,N_18254,N_18614);
xnor U21750 (N_21750,N_16351,N_15371);
xnor U21751 (N_21751,N_17160,N_15114);
xnor U21752 (N_21752,N_19482,N_17015);
nor U21753 (N_21753,N_17914,N_18389);
nand U21754 (N_21754,N_15525,N_16443);
nor U21755 (N_21755,N_17473,N_16422);
nor U21756 (N_21756,N_18792,N_15260);
nand U21757 (N_21757,N_18431,N_17869);
nand U21758 (N_21758,N_16128,N_18253);
xnor U21759 (N_21759,N_17026,N_19057);
nand U21760 (N_21760,N_17028,N_16009);
nor U21761 (N_21761,N_17491,N_15961);
or U21762 (N_21762,N_18944,N_18457);
or U21763 (N_21763,N_16191,N_18544);
or U21764 (N_21764,N_18908,N_18637);
or U21765 (N_21765,N_19668,N_17913);
xnor U21766 (N_21766,N_17422,N_17279);
nor U21767 (N_21767,N_16813,N_16872);
nor U21768 (N_21768,N_17378,N_15078);
nor U21769 (N_21769,N_15691,N_16837);
or U21770 (N_21770,N_17292,N_17511);
xor U21771 (N_21771,N_16040,N_19940);
and U21772 (N_21772,N_17891,N_15770);
nand U21773 (N_21773,N_19618,N_17466);
and U21774 (N_21774,N_19195,N_17528);
nand U21775 (N_21775,N_18840,N_16483);
or U21776 (N_21776,N_19495,N_17363);
and U21777 (N_21777,N_15618,N_16098);
xnor U21778 (N_21778,N_16869,N_18779);
nand U21779 (N_21779,N_15065,N_19242);
xor U21780 (N_21780,N_15625,N_18512);
nor U21781 (N_21781,N_15681,N_19764);
nor U21782 (N_21782,N_15538,N_17085);
and U21783 (N_21783,N_18769,N_16050);
nor U21784 (N_21784,N_15140,N_19994);
or U21785 (N_21785,N_19177,N_16182);
nor U21786 (N_21786,N_15112,N_16714);
nand U21787 (N_21787,N_18388,N_16401);
nor U21788 (N_21788,N_18374,N_15054);
nand U21789 (N_21789,N_16209,N_17485);
nand U21790 (N_21790,N_17867,N_16042);
or U21791 (N_21791,N_17746,N_17011);
nor U21792 (N_21792,N_17336,N_16866);
nand U21793 (N_21793,N_15068,N_19491);
and U21794 (N_21794,N_19507,N_17295);
nor U21795 (N_21795,N_15116,N_16674);
nor U21796 (N_21796,N_15792,N_16641);
or U21797 (N_21797,N_19645,N_17154);
or U21798 (N_21798,N_17858,N_17180);
nor U21799 (N_21799,N_15840,N_19951);
nand U21800 (N_21800,N_17455,N_17089);
nand U21801 (N_21801,N_19274,N_16775);
and U21802 (N_21802,N_16436,N_17399);
or U21803 (N_21803,N_16501,N_16164);
nand U21804 (N_21804,N_16609,N_18806);
nor U21805 (N_21805,N_17798,N_17468);
xnor U21806 (N_21806,N_16022,N_15823);
and U21807 (N_21807,N_19732,N_19606);
or U21808 (N_21808,N_19268,N_19907);
xor U21809 (N_21809,N_17229,N_15694);
xnor U21810 (N_21810,N_17564,N_15481);
nand U21811 (N_21811,N_16884,N_18449);
nand U21812 (N_21812,N_17172,N_18811);
and U21813 (N_21813,N_16250,N_15844);
or U21814 (N_21814,N_18874,N_19431);
nor U21815 (N_21815,N_18876,N_16484);
nand U21816 (N_21816,N_15429,N_17497);
nand U21817 (N_21817,N_18454,N_18797);
xor U21818 (N_21818,N_18667,N_17067);
or U21819 (N_21819,N_19478,N_15182);
and U21820 (N_21820,N_16289,N_15706);
nor U21821 (N_21821,N_17543,N_16268);
or U21822 (N_21822,N_15717,N_18755);
xor U21823 (N_21823,N_19611,N_15895);
xnor U21824 (N_21824,N_19143,N_18205);
nand U21825 (N_21825,N_19307,N_17557);
xnor U21826 (N_21826,N_17104,N_19850);
nand U21827 (N_21827,N_17955,N_15968);
or U21828 (N_21828,N_15997,N_18742);
nand U21829 (N_21829,N_18102,N_15145);
nor U21830 (N_21830,N_17465,N_19534);
nor U21831 (N_21831,N_16079,N_15633);
nor U21832 (N_21832,N_19436,N_16551);
nand U21833 (N_21833,N_15669,N_18286);
or U21834 (N_21834,N_17538,N_18615);
nor U21835 (N_21835,N_19227,N_15321);
nor U21836 (N_21836,N_17635,N_18481);
and U21837 (N_21837,N_17954,N_18132);
nand U21838 (N_21838,N_16739,N_17782);
nand U21839 (N_21839,N_15216,N_18486);
and U21840 (N_21840,N_17717,N_18186);
or U21841 (N_21841,N_16657,N_15547);
and U21842 (N_21842,N_17864,N_19340);
xor U21843 (N_21843,N_19966,N_18596);
or U21844 (N_21844,N_19167,N_17865);
nor U21845 (N_21845,N_16616,N_17841);
or U21846 (N_21846,N_18976,N_19097);
nor U21847 (N_21847,N_18800,N_17387);
nand U21848 (N_21848,N_17783,N_18585);
or U21849 (N_21849,N_18490,N_19644);
nand U21850 (N_21850,N_16947,N_17572);
or U21851 (N_21851,N_16857,N_17442);
or U21852 (N_21852,N_17963,N_18064);
and U21853 (N_21853,N_16370,N_15809);
nand U21854 (N_21854,N_18704,N_15239);
nor U21855 (N_21855,N_17464,N_15051);
nand U21856 (N_21856,N_19812,N_18554);
nor U21857 (N_21857,N_17747,N_18432);
nand U21858 (N_21858,N_18990,N_16284);
nor U21859 (N_21859,N_19991,N_15289);
nor U21860 (N_21860,N_19886,N_15209);
or U21861 (N_21861,N_18314,N_17174);
nand U21862 (N_21862,N_18632,N_18616);
nor U21863 (N_21863,N_15487,N_19469);
and U21864 (N_21864,N_19302,N_18362);
and U21865 (N_21865,N_15987,N_17219);
or U21866 (N_21866,N_18267,N_15553);
nand U21867 (N_21867,N_16017,N_17881);
or U21868 (N_21868,N_19543,N_15591);
xnor U21869 (N_21869,N_15971,N_16817);
nand U21870 (N_21870,N_19785,N_15617);
and U21871 (N_21871,N_19225,N_19758);
or U21872 (N_21872,N_17603,N_17424);
and U21873 (N_21873,N_18666,N_18820);
nor U21874 (N_21874,N_18636,N_18074);
nand U21875 (N_21875,N_18489,N_15000);
or U21876 (N_21876,N_15235,N_15960);
xor U21877 (N_21877,N_17404,N_17732);
or U21878 (N_21878,N_15527,N_15063);
and U21879 (N_21879,N_18602,N_15012);
xor U21880 (N_21880,N_16235,N_17203);
and U21881 (N_21881,N_17317,N_17328);
and U21882 (N_21882,N_18065,N_16722);
and U21883 (N_21883,N_15272,N_17683);
and U21884 (N_21884,N_18410,N_17722);
and U21885 (N_21885,N_15307,N_18760);
or U21886 (N_21886,N_17200,N_19441);
nor U21887 (N_21887,N_17365,N_16804);
nor U21888 (N_21888,N_17760,N_18656);
nor U21889 (N_21889,N_18969,N_15526);
xor U21890 (N_21890,N_16332,N_17395);
xor U21891 (N_21891,N_17248,N_17444);
xnor U21892 (N_21892,N_15537,N_19807);
nor U21893 (N_21893,N_19426,N_15247);
nand U21894 (N_21894,N_15123,N_15533);
nand U21895 (N_21895,N_18196,N_18578);
nor U21896 (N_21896,N_17479,N_19532);
nor U21897 (N_21897,N_19182,N_15357);
nand U21898 (N_21898,N_19718,N_16324);
nor U21899 (N_21899,N_17856,N_16748);
nor U21900 (N_21900,N_15829,N_17781);
nand U21901 (N_21901,N_15688,N_15220);
and U21902 (N_21902,N_19253,N_19318);
xor U21903 (N_21903,N_15841,N_19244);
xor U21904 (N_21904,N_15447,N_19206);
nor U21905 (N_21905,N_17127,N_16742);
nor U21906 (N_21906,N_19905,N_19547);
and U21907 (N_21907,N_15157,N_17239);
xor U21908 (N_21908,N_15901,N_19457);
nand U21909 (N_21909,N_18689,N_18321);
nor U21910 (N_21910,N_16558,N_17053);
xor U21911 (N_21911,N_18406,N_19430);
nor U21912 (N_21912,N_18129,N_17471);
and U21913 (N_21913,N_18207,N_16802);
or U21914 (N_21914,N_19069,N_15331);
xor U21915 (N_21915,N_16985,N_15565);
and U21916 (N_21916,N_17372,N_17876);
nor U21917 (N_21917,N_17063,N_18395);
nand U21918 (N_21918,N_19342,N_16895);
nor U21919 (N_21919,N_19023,N_15755);
xnor U21920 (N_21920,N_19405,N_19035);
and U21921 (N_21921,N_18382,N_15469);
xnor U21922 (N_21922,N_19714,N_16987);
xor U21923 (N_21923,N_18259,N_19818);
xor U21924 (N_21924,N_17967,N_16581);
or U21925 (N_21925,N_16203,N_15376);
nor U21926 (N_21926,N_15667,N_16850);
nand U21927 (N_21927,N_15351,N_19742);
nand U21928 (N_21928,N_18161,N_15984);
nand U21929 (N_21929,N_19723,N_18670);
nor U21930 (N_21930,N_16568,N_16494);
and U21931 (N_21931,N_17196,N_15195);
and U21932 (N_21932,N_17720,N_19310);
nor U21933 (N_21933,N_17411,N_17255);
nor U21934 (N_21934,N_15278,N_16671);
and U21935 (N_21935,N_16965,N_16678);
or U21936 (N_21936,N_17895,N_16319);
or U21937 (N_21937,N_19569,N_15210);
and U21938 (N_21938,N_15914,N_15346);
xnor U21939 (N_21939,N_19347,N_15084);
and U21940 (N_21940,N_16406,N_18178);
or U21941 (N_21941,N_18476,N_16218);
xor U21942 (N_21942,N_15308,N_18318);
or U21943 (N_21943,N_15129,N_18036);
xnor U21944 (N_21944,N_16990,N_19839);
or U21945 (N_21945,N_19351,N_19746);
xor U21946 (N_21946,N_17456,N_18545);
nor U21947 (N_21947,N_16983,N_18462);
or U21948 (N_21948,N_19587,N_19163);
nand U21949 (N_21949,N_18599,N_16645);
nor U21950 (N_21950,N_15837,N_16681);
and U21951 (N_21951,N_18780,N_19022);
nand U21952 (N_21952,N_19319,N_16848);
nand U21953 (N_21953,N_18438,N_18013);
nand U21954 (N_21954,N_19449,N_15259);
and U21955 (N_21955,N_16112,N_15838);
and U21956 (N_21956,N_17225,N_17946);
and U21957 (N_21957,N_15217,N_17437);
nor U21958 (N_21958,N_19090,N_15231);
xnor U21959 (N_21959,N_17302,N_15999);
or U21960 (N_21960,N_19375,N_18385);
and U21961 (N_21961,N_17199,N_15863);
nor U21962 (N_21962,N_17758,N_16560);
and U21963 (N_21963,N_19652,N_16174);
xnor U21964 (N_21964,N_15126,N_16602);
nor U21965 (N_21965,N_19108,N_18734);
nor U21966 (N_21966,N_18096,N_17476);
xor U21967 (N_21967,N_18856,N_16489);
xor U21968 (N_21968,N_16032,N_17757);
nand U21969 (N_21969,N_16015,N_16726);
or U21970 (N_21970,N_15400,N_15785);
nor U21971 (N_21971,N_18405,N_15092);
and U21972 (N_21972,N_19004,N_16842);
xnor U21973 (N_21973,N_17385,N_19797);
xor U21974 (N_21974,N_15047,N_18198);
and U21975 (N_21975,N_15711,N_15480);
or U21976 (N_21976,N_15586,N_18180);
xor U21977 (N_21977,N_16881,N_16811);
nor U21978 (N_21978,N_19571,N_19384);
xor U21979 (N_21979,N_19171,N_15500);
nand U21980 (N_21980,N_18945,N_17124);
nand U21981 (N_21981,N_19654,N_15821);
or U21982 (N_21982,N_18204,N_15539);
nor U21983 (N_21983,N_18415,N_17654);
nand U21984 (N_21984,N_15324,N_18258);
and U21985 (N_21985,N_17809,N_17042);
nand U21986 (N_21986,N_16672,N_17021);
xnor U21987 (N_21987,N_19865,N_16232);
nand U21988 (N_21988,N_15912,N_16532);
nand U21989 (N_21989,N_18973,N_15364);
or U21990 (N_21990,N_17915,N_16934);
nor U21991 (N_21991,N_15942,N_18081);
or U21992 (N_21992,N_19176,N_19323);
nand U21993 (N_21993,N_17784,N_15645);
and U21994 (N_21994,N_17966,N_16778);
and U21995 (N_21995,N_19101,N_17348);
xor U21996 (N_21996,N_17991,N_17694);
nand U21997 (N_21997,N_19735,N_15623);
or U21998 (N_21998,N_16879,N_16639);
nand U21999 (N_21999,N_15678,N_19870);
or U22000 (N_22000,N_17619,N_16355);
and U22001 (N_22001,N_15671,N_18977);
xor U22002 (N_22002,N_18417,N_15826);
and U22003 (N_22003,N_16999,N_16206);
xor U22004 (N_22004,N_17765,N_17038);
xnor U22005 (N_22005,N_18420,N_19800);
and U22006 (N_22006,N_15353,N_15825);
xnor U22007 (N_22007,N_17305,N_16287);
and U22008 (N_22008,N_17153,N_18678);
and U22009 (N_22009,N_18966,N_16642);
xor U22010 (N_22010,N_18485,N_17775);
and U22011 (N_22011,N_16415,N_18444);
nor U22012 (N_22012,N_16242,N_15457);
nand U22013 (N_22013,N_17945,N_19349);
xor U22014 (N_22014,N_16089,N_16514);
nand U22015 (N_22015,N_18880,N_17101);
nand U22016 (N_22016,N_16080,N_16440);
nor U22017 (N_22017,N_18587,N_15301);
xnor U22018 (N_22018,N_15511,N_17834);
and U22019 (N_22019,N_18729,N_17742);
xor U22020 (N_22020,N_15690,N_17571);
xor U22021 (N_22021,N_19613,N_18157);
nand U22022 (N_22022,N_15407,N_16688);
nand U22023 (N_22023,N_17009,N_19130);
and U22024 (N_22024,N_19183,N_15189);
nand U22025 (N_22025,N_19607,N_16049);
and U22026 (N_22026,N_17246,N_17110);
nand U22027 (N_22027,N_19399,N_19428);
xnor U22028 (N_22028,N_16298,N_16018);
xnor U22029 (N_22029,N_19815,N_19765);
nor U22030 (N_22030,N_16586,N_15759);
nand U22031 (N_22031,N_19299,N_19832);
and U22032 (N_22032,N_17094,N_17313);
or U22033 (N_22033,N_17999,N_19152);
xor U22034 (N_22034,N_15541,N_19616);
or U22035 (N_22035,N_18209,N_16316);
nor U22036 (N_22036,N_17152,N_18956);
nor U22037 (N_22037,N_15719,N_17979);
nor U22038 (N_22038,N_15736,N_17513);
nor U22039 (N_22039,N_18218,N_15169);
or U22040 (N_22040,N_17774,N_17590);
nor U22041 (N_22041,N_16487,N_17637);
or U22042 (N_22042,N_15434,N_15165);
or U22043 (N_22043,N_18293,N_17049);
xnor U22044 (N_22044,N_17311,N_18375);
or U22045 (N_22045,N_17937,N_19962);
nor U22046 (N_22046,N_17941,N_17662);
or U22047 (N_22047,N_17676,N_19660);
xor U22048 (N_22048,N_19619,N_18566);
or U22049 (N_22049,N_17971,N_17340);
nor U22050 (N_22050,N_19510,N_17493);
xor U22051 (N_22051,N_16044,N_16981);
nand U22052 (N_22052,N_17507,N_17403);
and U22053 (N_22053,N_19240,N_18580);
or U22054 (N_22054,N_17029,N_19567);
or U22055 (N_22055,N_15396,N_17803);
or U22056 (N_22056,N_16499,N_15668);
or U22057 (N_22057,N_19475,N_16426);
xor U22058 (N_22058,N_19877,N_16624);
xnor U22059 (N_22059,N_18802,N_16031);
or U22060 (N_22060,N_18386,N_19631);
or U22061 (N_22061,N_17122,N_19887);
xnor U22062 (N_22062,N_19398,N_18086);
or U22063 (N_22063,N_15415,N_15322);
xnor U22064 (N_22064,N_15672,N_15106);
nand U22065 (N_22065,N_19820,N_15458);
nor U22066 (N_22066,N_18072,N_17636);
or U22067 (N_22067,N_19052,N_16131);
and U22068 (N_22068,N_16500,N_19170);
nand U22069 (N_22069,N_15722,N_19155);
nand U22070 (N_22070,N_19536,N_19317);
xnor U22071 (N_22071,N_18343,N_17366);
xnor U22072 (N_22072,N_19450,N_16275);
nor U22073 (N_22073,N_15657,N_19209);
or U22074 (N_22074,N_18980,N_17371);
and U22075 (N_22075,N_15158,N_18983);
nor U22076 (N_22076,N_18677,N_16180);
xor U22077 (N_22077,N_16092,N_18251);
nand U22078 (N_22078,N_18673,N_16411);
xor U22079 (N_22079,N_17831,N_16019);
or U22080 (N_22080,N_15450,N_17477);
nand U22081 (N_22081,N_17810,N_16010);
and U22082 (N_22082,N_17942,N_19868);
nand U22083 (N_22083,N_16437,N_18847);
or U22084 (N_22084,N_18194,N_16404);
or U22085 (N_22085,N_15852,N_19019);
or U22086 (N_22086,N_16498,N_19497);
or U22087 (N_22087,N_16139,N_15183);
nor U22088 (N_22088,N_16741,N_17715);
nand U22089 (N_22089,N_18753,N_16763);
or U22090 (N_22090,N_17062,N_19502);
or U22091 (N_22091,N_18221,N_18775);
nor U22092 (N_22092,N_19511,N_15534);
nor U22093 (N_22093,N_18360,N_19438);
nand U22094 (N_22094,N_17164,N_19119);
nand U22095 (N_22095,N_19368,N_18838);
xor U22096 (N_22096,N_18027,N_15486);
and U22097 (N_22097,N_17000,N_15205);
or U22098 (N_22098,N_18367,N_17668);
nand U22099 (N_22099,N_19201,N_18940);
or U22100 (N_22100,N_16340,N_18965);
nor U22101 (N_22101,N_18359,N_19849);
nand U22102 (N_22102,N_17448,N_19063);
or U22103 (N_22103,N_18352,N_19106);
nand U22104 (N_22104,N_17322,N_18147);
and U22105 (N_22105,N_15365,N_16293);
nand U22106 (N_22106,N_17932,N_15122);
or U22107 (N_22107,N_16013,N_18754);
nand U22108 (N_22108,N_18628,N_18947);
or U22109 (N_22109,N_15574,N_16300);
and U22110 (N_22110,N_19112,N_15732);
xnor U22111 (N_22111,N_16764,N_18126);
xnor U22112 (N_22112,N_19485,N_19824);
and U22113 (N_22113,N_15932,N_19972);
nand U22114 (N_22114,N_15749,N_16951);
xnor U22115 (N_22115,N_19205,N_19184);
xor U22116 (N_22116,N_16563,N_17218);
and U22117 (N_22117,N_17483,N_18845);
xor U22118 (N_22118,N_16169,N_19154);
nand U22119 (N_22119,N_19077,N_16870);
and U22120 (N_22120,N_15341,N_18284);
xor U22121 (N_22121,N_18009,N_18807);
and U22122 (N_22122,N_15080,N_15741);
and U22123 (N_22123,N_17882,N_17045);
or U22124 (N_22124,N_17852,N_15142);
nand U22125 (N_22125,N_19173,N_17804);
nand U22126 (N_22126,N_19297,N_15476);
and U22127 (N_22127,N_15802,N_19702);
xor U22128 (N_22128,N_16836,N_15226);
nor U22129 (N_22129,N_16945,N_19135);
nor U22130 (N_22130,N_17050,N_16063);
xor U22131 (N_22131,N_15832,N_17927);
and U22132 (N_22132,N_18788,N_15807);
and U22133 (N_22133,N_16243,N_19070);
nand U22134 (N_22134,N_16652,N_16258);
nor U22135 (N_22135,N_18949,N_16434);
xor U22136 (N_22136,N_18048,N_15910);
and U22137 (N_22137,N_17721,N_16047);
nor U22138 (N_22138,N_16522,N_17323);
xnor U22139 (N_22139,N_17303,N_16919);
xnor U22140 (N_22140,N_16033,N_19961);
or U22141 (N_22141,N_16472,N_18718);
and U22142 (N_22142,N_15087,N_15777);
or U22143 (N_22143,N_17990,N_17157);
nand U22144 (N_22144,N_17495,N_18232);
or U22145 (N_22145,N_18801,N_19763);
nor U22146 (N_22146,N_19325,N_18097);
nand U22147 (N_22147,N_17585,N_19248);
and U22148 (N_22148,N_17983,N_17794);
xnor U22149 (N_22149,N_17386,N_19943);
and U22150 (N_22150,N_19411,N_18617);
xnor U22151 (N_22151,N_19246,N_19239);
and U22152 (N_22152,N_19056,N_17379);
or U22153 (N_22153,N_17186,N_16937);
nand U22154 (N_22154,N_19843,N_16432);
xor U22155 (N_22155,N_17802,N_17277);
xor U22156 (N_22156,N_17449,N_18035);
xor U22157 (N_22157,N_17014,N_16543);
and U22158 (N_22158,N_19303,N_18448);
and U22159 (N_22159,N_15723,N_17145);
or U22160 (N_22160,N_18791,N_19804);
xnor U22161 (N_22161,N_15701,N_18252);
nand U22162 (N_22162,N_15710,N_16969);
or U22163 (N_22163,N_15937,N_19992);
nor U22164 (N_22164,N_17073,N_19615);
nor U22165 (N_22165,N_16798,N_15018);
or U22166 (N_22166,N_19282,N_15456);
nand U22167 (N_22167,N_16899,N_18450);
nand U22168 (N_22168,N_16115,N_16230);
nor U22169 (N_22169,N_17256,N_16041);
xor U22170 (N_22170,N_18379,N_16980);
xnor U22171 (N_22171,N_18182,N_19686);
nor U22172 (N_22172,N_16629,N_15075);
nor U22173 (N_22173,N_18812,N_16926);
nand U22174 (N_22174,N_15850,N_17066);
or U22175 (N_22175,N_16453,N_15375);
nand U22176 (N_22176,N_19666,N_17577);
nor U22177 (N_22177,N_16546,N_16874);
nand U22178 (N_22178,N_19045,N_15071);
nand U22179 (N_22179,N_16858,N_16539);
nand U22180 (N_22180,N_15081,N_17024);
or U22181 (N_22181,N_17397,N_16806);
nand U22182 (N_22182,N_17343,N_17051);
nor U22183 (N_22183,N_15988,N_16929);
and U22184 (N_22184,N_19847,N_18782);
nor U22185 (N_22185,N_18982,N_17139);
xor U22186 (N_22186,N_16291,N_19138);
or U22187 (N_22187,N_16322,N_15580);
nand U22188 (N_22188,N_15269,N_15890);
and U22189 (N_22189,N_18105,N_16878);
xor U22190 (N_22190,N_15417,N_19855);
nor U22191 (N_22191,N_19786,N_16430);
xor U22192 (N_22192,N_16554,N_15911);
or U22193 (N_22193,N_17547,N_19669);
nor U22194 (N_22194,N_19647,N_19739);
or U22195 (N_22195,N_15522,N_19251);
xnor U22196 (N_22196,N_16299,N_17001);
and U22197 (N_22197,N_19012,N_16791);
and U22198 (N_22198,N_18138,N_16399);
nor U22199 (N_22199,N_15090,N_18962);
and U22200 (N_22200,N_17335,N_16927);
and U22201 (N_22201,N_17897,N_15242);
xnor U22202 (N_22202,N_16923,N_17068);
xnor U22203 (N_22203,N_19078,N_16548);
or U22204 (N_22204,N_19923,N_18309);
xor U22205 (N_22205,N_15213,N_15497);
nand U22206 (N_22206,N_18332,N_16703);
nand U22207 (N_22207,N_18553,N_16062);
and U22208 (N_22208,N_19687,N_17060);
or U22209 (N_22209,N_15014,N_19983);
or U22210 (N_22210,N_15176,N_16515);
xnor U22211 (N_22211,N_15154,N_15275);
or U22212 (N_22212,N_17586,N_15861);
nor U22213 (N_22213,N_19365,N_16461);
xnor U22214 (N_22214,N_15928,N_15421);
xnor U22215 (N_22215,N_15284,N_18588);
or U22216 (N_22216,N_16555,N_18061);
or U22217 (N_22217,N_19490,N_18112);
and U22218 (N_22218,N_19659,N_18952);
nand U22219 (N_22219,N_19327,N_15170);
nand U22220 (N_22220,N_18002,N_19158);
nand U22221 (N_22221,N_15384,N_18774);
or U22222 (N_22222,N_16455,N_19432);
and U22223 (N_22223,N_19224,N_15039);
nor U22224 (N_22224,N_16649,N_19079);
or U22225 (N_22225,N_18719,N_19762);
and U22226 (N_22226,N_17964,N_15168);
and U22227 (N_22227,N_17347,N_19394);
nand U22228 (N_22228,N_19736,N_15644);
nand U22229 (N_22229,N_18954,N_18920);
and U22230 (N_22230,N_17797,N_15808);
xnor U22231 (N_22231,N_19159,N_19024);
or U22232 (N_22232,N_19566,N_16725);
nand U22233 (N_22233,N_19904,N_16625);
and U22234 (N_22234,N_16975,N_15070);
or U22235 (N_22235,N_17642,N_18073);
nor U22236 (N_22236,N_18787,N_15680);
nor U22237 (N_22237,N_18671,N_19623);
or U22238 (N_22238,N_15820,N_16687);
xor U22239 (N_22239,N_16450,N_17569);
xor U22240 (N_22240,N_15787,N_16900);
or U22241 (N_22241,N_18504,N_19900);
nand U22242 (N_22242,N_18984,N_16429);
xnor U22243 (N_22243,N_16380,N_19100);
nor U22244 (N_22244,N_18459,N_17494);
nor U22245 (N_22245,N_18437,N_17030);
and U22246 (N_22246,N_17845,N_18814);
or U22247 (N_22247,N_19857,N_15828);
or U22248 (N_22248,N_19140,N_17374);
nand U22249 (N_22249,N_15352,N_17048);
xor U22250 (N_22250,N_16903,N_15148);
and U22251 (N_22251,N_16389,N_17604);
nand U22252 (N_22252,N_17951,N_18978);
or U22253 (N_22253,N_18038,N_16132);
nand U22254 (N_22254,N_17568,N_18443);
or U22255 (N_22255,N_18715,N_16647);
xnor U22256 (N_22256,N_16329,N_17844);
and U22257 (N_22257,N_16410,N_16608);
and U22258 (N_22258,N_15924,N_19749);
or U22259 (N_22259,N_15654,N_15149);
nand U22260 (N_22260,N_19650,N_19969);
xor U22261 (N_22261,N_18225,N_16456);
nor U22262 (N_22262,N_18340,N_15816);
nand U22263 (N_22263,N_16288,N_16087);
nand U22264 (N_22264,N_18967,N_17252);
nor U22265 (N_22265,N_17289,N_17428);
or U22266 (N_22266,N_17123,N_19410);
xor U22267 (N_22267,N_18307,N_17597);
nor U22268 (N_22268,N_17454,N_19095);
or U22269 (N_22269,N_18758,N_18582);
and U22270 (N_22270,N_18612,N_18006);
xnor U22271 (N_22271,N_16292,N_17168);
and U22272 (N_22272,N_18062,N_17342);
or U22273 (N_22273,N_15653,N_18248);
xor U22274 (N_22274,N_18280,N_17551);
nor U22275 (N_22275,N_16246,N_16961);
nor U22276 (N_22276,N_16957,N_19039);
xor U22277 (N_22277,N_18373,N_18560);
or U22278 (N_22278,N_15627,N_17503);
or U22279 (N_22279,N_17633,N_18682);
nor U22280 (N_22280,N_19685,N_15608);
xnor U22281 (N_22281,N_16286,N_19306);
xor U22282 (N_22282,N_16271,N_18403);
nor U22283 (N_22283,N_19520,N_17268);
nor U22284 (N_22284,N_16142,N_16653);
nand U22285 (N_22285,N_15615,N_17873);
or U22286 (N_22286,N_15263,N_15814);
or U22287 (N_22287,N_17626,N_15172);
nand U22288 (N_22288,N_18503,N_18827);
and U22289 (N_22289,N_15753,N_18301);
or U22290 (N_22290,N_19287,N_17010);
xnor U22291 (N_22291,N_18101,N_19199);
and U22292 (N_22292,N_16503,N_19671);
xor U22293 (N_22293,N_16564,N_15304);
xnor U22294 (N_22294,N_18043,N_17091);
nand U22295 (N_22295,N_17132,N_15041);
nand U22296 (N_22296,N_16956,N_16529);
or U22297 (N_22297,N_17714,N_18357);
nor U22298 (N_22298,N_16557,N_18808);
nand U22299 (N_22299,N_16541,N_15845);
and U22300 (N_22300,N_18547,N_19977);
nor U22301 (N_22301,N_16686,N_15995);
or U22302 (N_22302,N_17843,N_15020);
nor U22303 (N_22303,N_15010,N_19572);
and U22304 (N_22304,N_18123,N_17805);
nor U22305 (N_22305,N_16225,N_16650);
nand U22306 (N_22306,N_17684,N_16151);
nand U22307 (N_22307,N_18915,N_15067);
nand U22308 (N_22308,N_18842,N_18042);
and U22309 (N_22309,N_15775,N_18542);
and U22310 (N_22310,N_18197,N_16105);
nor U22311 (N_22311,N_16832,N_15977);
nand U22312 (N_22312,N_16264,N_17996);
or U22313 (N_22313,N_18364,N_15342);
nor U22314 (N_22314,N_15438,N_16446);
nor U22315 (N_22315,N_17236,N_18568);
and U22316 (N_22316,N_16168,N_18302);
nand U22317 (N_22317,N_18270,N_16917);
nor U22318 (N_22318,N_15909,N_18694);
xor U22319 (N_22319,N_15348,N_17776);
nand U22320 (N_22320,N_16371,N_18733);
nand U22321 (N_22321,N_19315,N_17337);
and U22322 (N_22322,N_15572,N_19653);
nand U22323 (N_22323,N_18070,N_16931);
and U22324 (N_22324,N_16451,N_19376);
xor U22325 (N_22325,N_17606,N_17391);
xor U22326 (N_22326,N_15333,N_19296);
nand U22327 (N_22327,N_18014,N_16619);
xor U22328 (N_22328,N_18864,N_16150);
or U22329 (N_22329,N_17088,N_19971);
xnor U22330 (N_22330,N_15485,N_17791);
nor U22331 (N_22331,N_17421,N_17452);
and U22332 (N_22332,N_18770,N_19549);
nand U22333 (N_22333,N_19934,N_17384);
xor U22334 (N_22334,N_16790,N_16800);
nand U22335 (N_22335,N_17707,N_19483);
or U22336 (N_22336,N_16752,N_19028);
and U22337 (N_22337,N_15038,N_17331);
and U22338 (N_22338,N_15810,N_17892);
or U22339 (N_22339,N_18923,N_15045);
or U22340 (N_22340,N_19999,N_18219);
xnor U22341 (N_22341,N_18419,N_17492);
nand U22342 (N_22342,N_16036,N_15128);
nand U22343 (N_22343,N_19828,N_17787);
or U22344 (N_22344,N_16424,N_15674);
nand U22345 (N_22345,N_17850,N_19084);
nor U22346 (N_22346,N_19372,N_15290);
xnor U22347 (N_22347,N_18189,N_19530);
or U22348 (N_22348,N_16757,N_15542);
nor U22349 (N_22349,N_18846,N_15377);
xor U22350 (N_22350,N_16367,N_18313);
nand U22351 (N_22351,N_18226,N_18436);
and U22352 (N_22352,N_18781,N_17796);
nand U22353 (N_22353,N_19222,N_15545);
nor U22354 (N_22354,N_16071,N_16384);
or U22355 (N_22355,N_16820,N_19150);
xnor U22356 (N_22356,N_19701,N_17958);
nand U22357 (N_22357,N_18606,N_15638);
xor U22358 (N_22358,N_19531,N_16336);
nor U22359 (N_22359,N_17846,N_19953);
xnor U22360 (N_22360,N_16148,N_15428);
nor U22361 (N_22361,N_15693,N_17093);
and U22362 (N_22362,N_17578,N_18262);
or U22363 (N_22363,N_18525,N_19822);
and U22364 (N_22364,N_19570,N_16941);
or U22365 (N_22365,N_19081,N_18763);
and U22366 (N_22366,N_18651,N_16171);
or U22367 (N_22367,N_19791,N_16354);
xor U22368 (N_22368,N_19612,N_17273);
xnor U22369 (N_22369,N_15030,N_17702);
or U22370 (N_22370,N_17579,N_17150);
nand U22371 (N_22371,N_19683,N_19029);
nor U22372 (N_22372,N_15768,N_16076);
nand U22373 (N_22373,N_18645,N_16694);
nand U22374 (N_22374,N_18136,N_18931);
and U22375 (N_22375,N_19709,N_16348);
nor U22376 (N_22376,N_15956,N_16004);
and U22377 (N_22377,N_15311,N_15865);
nor U22378 (N_22378,N_19030,N_15963);
nand U22379 (N_22379,N_16550,N_17394);
and U22380 (N_22380,N_15581,N_17321);
and U22381 (N_22381,N_18492,N_16777);
xor U22382 (N_22382,N_15399,N_15652);
or U22383 (N_22383,N_16251,N_16051);
nand U22384 (N_22384,N_17887,N_19596);
nand U22385 (N_22385,N_19049,N_18201);
or U22386 (N_22386,N_15958,N_18099);
xnor U22387 (N_22387,N_19113,N_18604);
or U22388 (N_22388,N_18609,N_18288);
nor U22389 (N_22389,N_17193,N_15166);
nand U22390 (N_22390,N_18743,N_17905);
nand U22391 (N_22391,N_17638,N_15374);
or U22392 (N_22392,N_18214,N_19827);
or U22393 (N_22393,N_16989,N_17143);
or U22394 (N_22394,N_18355,N_18263);
and U22395 (N_22395,N_18519,N_15085);
and U22396 (N_22396,N_16974,N_19866);
or U22397 (N_22397,N_16807,N_18933);
nand U22398 (N_22398,N_19542,N_19445);
xnor U22399 (N_22399,N_19823,N_19245);
xor U22400 (N_22400,N_18911,N_19733);
and U22401 (N_22401,N_15017,N_18217);
or U22402 (N_22402,N_18172,N_16530);
nand U22403 (N_22403,N_17731,N_16425);
and U22404 (N_22404,N_15019,N_15567);
or U22405 (N_22405,N_16831,N_15329);
or U22406 (N_22406,N_18865,N_15110);
xnor U22407 (N_22407,N_17318,N_15218);
xnor U22408 (N_22408,N_19276,N_18336);
xor U22409 (N_22409,N_16819,N_19484);
or U22410 (N_22410,N_19486,N_15053);
xor U22411 (N_22411,N_17763,N_17235);
xor U22412 (N_22412,N_18871,N_16691);
or U22413 (N_22413,N_19413,N_19047);
xnor U22414 (N_22414,N_17833,N_18482);
nor U22415 (N_22415,N_18917,N_19291);
nor U22416 (N_22416,N_15512,N_18538);
xor U22417 (N_22417,N_19046,N_16970);
nand U22418 (N_22418,N_17688,N_19172);
nand U22419 (N_22419,N_17120,N_15419);
xnor U22420 (N_22420,N_19346,N_18452);
and U22421 (N_22421,N_19700,N_16573);
or U22422 (N_22422,N_15049,N_17718);
nor U22423 (N_22423,N_18040,N_15738);
xnor U22424 (N_22424,N_18208,N_19294);
and U22425 (N_22425,N_16611,N_18414);
nand U22426 (N_22426,N_17410,N_16375);
nor U22427 (N_22427,N_17459,N_15194);
or U22428 (N_22428,N_19053,N_19976);
or U22429 (N_22429,N_18115,N_19967);
nor U22430 (N_22430,N_16469,N_16574);
xor U22431 (N_22431,N_16680,N_18025);
nand U22432 (N_22432,N_17241,N_18899);
and U22433 (N_22433,N_19933,N_16901);
xor U22434 (N_22434,N_19381,N_18240);
and U22435 (N_22435,N_19609,N_15856);
xor U22436 (N_22436,N_15990,N_16068);
xor U22437 (N_22437,N_16420,N_19909);
or U22438 (N_22438,N_18958,N_19313);
xnor U22439 (N_22439,N_19336,N_19655);
nor U22440 (N_22440,N_16598,N_18926);
xnor U22441 (N_22441,N_16762,N_16147);
xor U22442 (N_22442,N_19462,N_17480);
and U22443 (N_22443,N_17553,N_15368);
or U22444 (N_22444,N_19620,N_16178);
xor U22445 (N_22445,N_18281,N_16904);
xnor U22446 (N_22446,N_15416,N_18372);
xor U22447 (N_22447,N_18955,N_15359);
nand U22448 (N_22448,N_17137,N_15337);
xor U22449 (N_22449,N_16385,N_15692);
nor U22450 (N_22450,N_15934,N_17126);
nor U22451 (N_22451,N_17031,N_15698);
and U22452 (N_22452,N_18810,N_18085);
xor U22453 (N_22453,N_19050,N_17716);
xnor U22454 (N_22454,N_16708,N_19238);
or U22455 (N_22455,N_16362,N_16480);
and U22456 (N_22456,N_15034,N_18569);
or U22457 (N_22457,N_18506,N_16121);
nand U22458 (N_22458,N_15900,N_17560);
nor U22459 (N_22459,N_17115,N_15747);
nor U22460 (N_22460,N_15354,N_16407);
xor U22461 (N_22461,N_18583,N_15197);
nand U22462 (N_22462,N_16893,N_17096);
or U22463 (N_22463,N_15709,N_19380);
or U22464 (N_22464,N_17997,N_19275);
nand U22465 (N_22465,N_17197,N_18330);
and U22466 (N_22466,N_15920,N_15556);
xnor U22467 (N_22467,N_16908,N_16315);
nand U22468 (N_22468,N_18125,N_15742);
or U22469 (N_22469,N_19417,N_16993);
or U22470 (N_22470,N_16579,N_15729);
xnor U22471 (N_22471,N_17968,N_18350);
or U22472 (N_22472,N_17097,N_15905);
xnor U22473 (N_22473,N_16311,N_18818);
nand U22474 (N_22474,N_18023,N_15013);
and U22475 (N_22475,N_18831,N_18643);
nand U22476 (N_22476,N_19931,N_15933);
and U22477 (N_22477,N_19188,N_15620);
and U22478 (N_22478,N_16495,N_19067);
nand U22479 (N_22479,N_18668,N_18935);
nand U22480 (N_22480,N_18918,N_15813);
nand U22481 (N_22481,N_17811,N_18461);
xnor U22482 (N_22482,N_18066,N_15535);
nor U22483 (N_22483,N_17677,N_15405);
or U22484 (N_22484,N_16786,N_18495);
and U22485 (N_22485,N_19955,N_17786);
or U22486 (N_22486,N_19366,N_15502);
and U22487 (N_22487,N_15238,N_16755);
nor U22488 (N_22488,N_17130,N_18325);
xor U22489 (N_22489,N_19148,N_19533);
or U22490 (N_22490,N_17706,N_15332);
and U22491 (N_22491,N_18442,N_18516);
xor U22492 (N_22492,N_18881,N_16479);
nand U22493 (N_22493,N_16012,N_17487);
or U22494 (N_22494,N_19738,N_19223);
xnor U22495 (N_22495,N_15714,N_16361);
and U22496 (N_22496,N_16660,N_15805);
xnor U22497 (N_22497,N_15649,N_18122);
and U22498 (N_22498,N_17825,N_17190);
nand U22499 (N_22499,N_18943,N_15906);
nor U22500 (N_22500,N_18135,N_19577);
nand U22501 (N_22501,N_15452,N_17891);
and U22502 (N_22502,N_16145,N_17837);
xnor U22503 (N_22503,N_16834,N_18590);
xnor U22504 (N_22504,N_16988,N_15922);
xnor U22505 (N_22505,N_17605,N_15647);
and U22506 (N_22506,N_15899,N_18332);
nor U22507 (N_22507,N_16564,N_18420);
nor U22508 (N_22508,N_15260,N_17243);
or U22509 (N_22509,N_19646,N_15929);
nand U22510 (N_22510,N_16869,N_15823);
nor U22511 (N_22511,N_17863,N_16363);
nor U22512 (N_22512,N_19056,N_15772);
xnor U22513 (N_22513,N_16856,N_16453);
or U22514 (N_22514,N_18896,N_17593);
and U22515 (N_22515,N_16674,N_17983);
and U22516 (N_22516,N_15929,N_17300);
xnor U22517 (N_22517,N_16705,N_16513);
nor U22518 (N_22518,N_18833,N_17636);
or U22519 (N_22519,N_17959,N_17166);
xnor U22520 (N_22520,N_17540,N_16231);
or U22521 (N_22521,N_15657,N_19241);
or U22522 (N_22522,N_15160,N_16861);
xor U22523 (N_22523,N_19864,N_16226);
nor U22524 (N_22524,N_18315,N_18395);
and U22525 (N_22525,N_18520,N_16928);
xnor U22526 (N_22526,N_17527,N_16972);
nand U22527 (N_22527,N_15460,N_17086);
nor U22528 (N_22528,N_18452,N_15460);
nand U22529 (N_22529,N_18706,N_18350);
xnor U22530 (N_22530,N_15167,N_15414);
nor U22531 (N_22531,N_16885,N_16692);
nor U22532 (N_22532,N_19244,N_19130);
nor U22533 (N_22533,N_17232,N_16790);
and U22534 (N_22534,N_15193,N_18634);
or U22535 (N_22535,N_18922,N_15492);
and U22536 (N_22536,N_17127,N_19422);
and U22537 (N_22537,N_18585,N_15120);
nand U22538 (N_22538,N_15154,N_17094);
xor U22539 (N_22539,N_16666,N_18869);
nand U22540 (N_22540,N_18456,N_18126);
nor U22541 (N_22541,N_16877,N_16163);
nor U22542 (N_22542,N_15882,N_19576);
or U22543 (N_22543,N_16575,N_19509);
and U22544 (N_22544,N_17243,N_16241);
or U22545 (N_22545,N_15041,N_19511);
nor U22546 (N_22546,N_15437,N_15636);
or U22547 (N_22547,N_19887,N_19440);
nand U22548 (N_22548,N_17286,N_16797);
nor U22549 (N_22549,N_17611,N_17852);
nor U22550 (N_22550,N_17057,N_19924);
nor U22551 (N_22551,N_18877,N_16705);
nor U22552 (N_22552,N_19285,N_19443);
nor U22553 (N_22553,N_19969,N_16035);
nor U22554 (N_22554,N_17501,N_15450);
or U22555 (N_22555,N_16176,N_16038);
nor U22556 (N_22556,N_18576,N_18196);
nand U22557 (N_22557,N_16997,N_16656);
or U22558 (N_22558,N_17440,N_18593);
nor U22559 (N_22559,N_17609,N_15578);
nor U22560 (N_22560,N_16503,N_15756);
or U22561 (N_22561,N_15644,N_17843);
nor U22562 (N_22562,N_15685,N_16949);
nand U22563 (N_22563,N_19848,N_19656);
nand U22564 (N_22564,N_15649,N_16262);
nand U22565 (N_22565,N_19374,N_16799);
xor U22566 (N_22566,N_15220,N_15430);
xnor U22567 (N_22567,N_17308,N_16530);
or U22568 (N_22568,N_15713,N_18418);
and U22569 (N_22569,N_19802,N_19116);
nor U22570 (N_22570,N_15640,N_15538);
nand U22571 (N_22571,N_18658,N_15137);
xor U22572 (N_22572,N_15610,N_17010);
nor U22573 (N_22573,N_19120,N_16479);
nor U22574 (N_22574,N_17237,N_17649);
xor U22575 (N_22575,N_19303,N_17188);
nand U22576 (N_22576,N_19448,N_16769);
xnor U22577 (N_22577,N_17116,N_18573);
and U22578 (N_22578,N_18007,N_18416);
nor U22579 (N_22579,N_18564,N_16904);
and U22580 (N_22580,N_19208,N_17561);
and U22581 (N_22581,N_17959,N_19137);
or U22582 (N_22582,N_15062,N_18047);
or U22583 (N_22583,N_17765,N_18591);
nand U22584 (N_22584,N_19920,N_16189);
nand U22585 (N_22585,N_16923,N_15108);
nand U22586 (N_22586,N_16392,N_17241);
or U22587 (N_22587,N_15671,N_16511);
or U22588 (N_22588,N_18855,N_15821);
and U22589 (N_22589,N_16878,N_19785);
or U22590 (N_22590,N_18214,N_17619);
nor U22591 (N_22591,N_15134,N_19006);
xnor U22592 (N_22592,N_18550,N_17212);
nand U22593 (N_22593,N_16892,N_16833);
nand U22594 (N_22594,N_18026,N_17553);
nand U22595 (N_22595,N_16415,N_16632);
or U22596 (N_22596,N_16971,N_16111);
nand U22597 (N_22597,N_19356,N_16046);
or U22598 (N_22598,N_18854,N_15170);
nand U22599 (N_22599,N_19096,N_17965);
nor U22600 (N_22600,N_17786,N_18842);
xnor U22601 (N_22601,N_15236,N_19318);
nand U22602 (N_22602,N_19541,N_16729);
nor U22603 (N_22603,N_18663,N_17906);
nor U22604 (N_22604,N_19406,N_17542);
or U22605 (N_22605,N_17665,N_17093);
and U22606 (N_22606,N_18221,N_15689);
nor U22607 (N_22607,N_17965,N_19676);
nand U22608 (N_22608,N_19136,N_16195);
nor U22609 (N_22609,N_15003,N_18507);
nand U22610 (N_22610,N_16125,N_16051);
nand U22611 (N_22611,N_16597,N_15518);
nand U22612 (N_22612,N_17539,N_15774);
nand U22613 (N_22613,N_19795,N_19025);
nand U22614 (N_22614,N_18051,N_16575);
or U22615 (N_22615,N_18030,N_18322);
nor U22616 (N_22616,N_18347,N_18628);
nand U22617 (N_22617,N_15837,N_18192);
xnor U22618 (N_22618,N_19972,N_16253);
xnor U22619 (N_22619,N_16775,N_19514);
or U22620 (N_22620,N_17737,N_17293);
xor U22621 (N_22621,N_15178,N_15093);
nor U22622 (N_22622,N_17475,N_16847);
or U22623 (N_22623,N_15108,N_19535);
and U22624 (N_22624,N_18557,N_17919);
xor U22625 (N_22625,N_16914,N_17192);
xnor U22626 (N_22626,N_16560,N_16716);
and U22627 (N_22627,N_18417,N_16504);
nor U22628 (N_22628,N_18404,N_15726);
xnor U22629 (N_22629,N_17214,N_16244);
nand U22630 (N_22630,N_15184,N_19147);
and U22631 (N_22631,N_16818,N_19836);
or U22632 (N_22632,N_18131,N_17230);
or U22633 (N_22633,N_17292,N_15989);
nand U22634 (N_22634,N_17626,N_15555);
xor U22635 (N_22635,N_16961,N_18504);
and U22636 (N_22636,N_18166,N_18559);
and U22637 (N_22637,N_17478,N_15378);
xor U22638 (N_22638,N_16112,N_15936);
and U22639 (N_22639,N_19245,N_15658);
nor U22640 (N_22640,N_16313,N_15470);
xor U22641 (N_22641,N_19229,N_19456);
or U22642 (N_22642,N_17663,N_15190);
and U22643 (N_22643,N_18810,N_18430);
and U22644 (N_22644,N_17824,N_17110);
nand U22645 (N_22645,N_15359,N_15806);
nor U22646 (N_22646,N_19224,N_19931);
or U22647 (N_22647,N_19071,N_17332);
nand U22648 (N_22648,N_15659,N_19212);
and U22649 (N_22649,N_19641,N_19210);
or U22650 (N_22650,N_17807,N_17061);
xnor U22651 (N_22651,N_19841,N_15900);
or U22652 (N_22652,N_19052,N_18654);
and U22653 (N_22653,N_19640,N_15267);
and U22654 (N_22654,N_18458,N_18887);
and U22655 (N_22655,N_19706,N_18746);
nor U22656 (N_22656,N_18575,N_15603);
nor U22657 (N_22657,N_18400,N_16649);
or U22658 (N_22658,N_18687,N_17494);
or U22659 (N_22659,N_19952,N_15080);
nand U22660 (N_22660,N_15767,N_19090);
and U22661 (N_22661,N_15191,N_18889);
nand U22662 (N_22662,N_16801,N_16436);
and U22663 (N_22663,N_19582,N_16017);
nand U22664 (N_22664,N_17864,N_18078);
xnor U22665 (N_22665,N_15251,N_17445);
nand U22666 (N_22666,N_16468,N_15841);
or U22667 (N_22667,N_18047,N_17984);
nor U22668 (N_22668,N_19311,N_17634);
and U22669 (N_22669,N_18393,N_15636);
nor U22670 (N_22670,N_15774,N_19527);
or U22671 (N_22671,N_15367,N_19097);
nand U22672 (N_22672,N_18621,N_15271);
nor U22673 (N_22673,N_16720,N_16784);
or U22674 (N_22674,N_15506,N_15554);
nor U22675 (N_22675,N_16797,N_19229);
or U22676 (N_22676,N_15638,N_15518);
and U22677 (N_22677,N_17148,N_16098);
or U22678 (N_22678,N_16391,N_19040);
nor U22679 (N_22679,N_16844,N_15772);
or U22680 (N_22680,N_17644,N_16326);
xnor U22681 (N_22681,N_17202,N_16580);
xor U22682 (N_22682,N_17743,N_15876);
nand U22683 (N_22683,N_16192,N_18335);
xor U22684 (N_22684,N_17967,N_17300);
nor U22685 (N_22685,N_17545,N_18183);
or U22686 (N_22686,N_17142,N_16531);
xnor U22687 (N_22687,N_15751,N_19273);
xor U22688 (N_22688,N_15143,N_18752);
nor U22689 (N_22689,N_16852,N_17431);
nor U22690 (N_22690,N_17665,N_19226);
and U22691 (N_22691,N_17696,N_18641);
and U22692 (N_22692,N_16550,N_17251);
and U22693 (N_22693,N_16604,N_18804);
and U22694 (N_22694,N_16275,N_18584);
nor U22695 (N_22695,N_19062,N_17908);
xor U22696 (N_22696,N_18241,N_15782);
nor U22697 (N_22697,N_16023,N_17594);
xor U22698 (N_22698,N_15281,N_18182);
or U22699 (N_22699,N_17864,N_19853);
nor U22700 (N_22700,N_19168,N_19512);
and U22701 (N_22701,N_15568,N_19133);
and U22702 (N_22702,N_19633,N_15110);
nand U22703 (N_22703,N_19656,N_15391);
or U22704 (N_22704,N_19501,N_16741);
or U22705 (N_22705,N_16660,N_19821);
or U22706 (N_22706,N_16388,N_18276);
or U22707 (N_22707,N_19827,N_16668);
and U22708 (N_22708,N_16684,N_15528);
nand U22709 (N_22709,N_15559,N_19340);
or U22710 (N_22710,N_17388,N_18183);
nor U22711 (N_22711,N_15004,N_15715);
and U22712 (N_22712,N_19367,N_16398);
or U22713 (N_22713,N_19460,N_15040);
or U22714 (N_22714,N_17495,N_19050);
and U22715 (N_22715,N_19640,N_16266);
and U22716 (N_22716,N_18791,N_16102);
or U22717 (N_22717,N_15392,N_15493);
xor U22718 (N_22718,N_18312,N_17369);
nand U22719 (N_22719,N_19796,N_19477);
and U22720 (N_22720,N_19924,N_19701);
nor U22721 (N_22721,N_15376,N_18659);
xor U22722 (N_22722,N_19382,N_16617);
xnor U22723 (N_22723,N_18491,N_17888);
or U22724 (N_22724,N_18230,N_15729);
xor U22725 (N_22725,N_15608,N_17096);
xnor U22726 (N_22726,N_16483,N_18758);
nor U22727 (N_22727,N_19313,N_19618);
and U22728 (N_22728,N_17712,N_16773);
nand U22729 (N_22729,N_15206,N_19632);
and U22730 (N_22730,N_18194,N_18011);
nand U22731 (N_22731,N_19980,N_16445);
nand U22732 (N_22732,N_17095,N_19424);
nor U22733 (N_22733,N_18303,N_15990);
or U22734 (N_22734,N_18901,N_18596);
or U22735 (N_22735,N_19322,N_15195);
and U22736 (N_22736,N_19122,N_15547);
or U22737 (N_22737,N_19332,N_18870);
or U22738 (N_22738,N_15320,N_17489);
xnor U22739 (N_22739,N_17071,N_16191);
and U22740 (N_22740,N_15899,N_19289);
xnor U22741 (N_22741,N_17939,N_17359);
and U22742 (N_22742,N_17087,N_17289);
or U22743 (N_22743,N_16428,N_18056);
xor U22744 (N_22744,N_18455,N_15324);
and U22745 (N_22745,N_18756,N_17019);
and U22746 (N_22746,N_18851,N_16477);
or U22747 (N_22747,N_15579,N_17763);
and U22748 (N_22748,N_18334,N_17918);
nor U22749 (N_22749,N_19860,N_16719);
xor U22750 (N_22750,N_15862,N_17533);
or U22751 (N_22751,N_17318,N_16088);
and U22752 (N_22752,N_19685,N_19496);
nand U22753 (N_22753,N_17778,N_19579);
and U22754 (N_22754,N_16041,N_18636);
or U22755 (N_22755,N_17373,N_18949);
nand U22756 (N_22756,N_19848,N_16740);
and U22757 (N_22757,N_17960,N_17704);
xor U22758 (N_22758,N_19360,N_19377);
xnor U22759 (N_22759,N_15736,N_19918);
and U22760 (N_22760,N_17751,N_19950);
xnor U22761 (N_22761,N_18064,N_19543);
nor U22762 (N_22762,N_18154,N_18648);
xnor U22763 (N_22763,N_17445,N_17813);
and U22764 (N_22764,N_18147,N_16784);
nand U22765 (N_22765,N_19678,N_16971);
or U22766 (N_22766,N_18678,N_19572);
xnor U22767 (N_22767,N_17638,N_17955);
xor U22768 (N_22768,N_17118,N_18973);
xnor U22769 (N_22769,N_18189,N_17966);
or U22770 (N_22770,N_15345,N_19475);
and U22771 (N_22771,N_15323,N_16614);
nand U22772 (N_22772,N_18580,N_17529);
xor U22773 (N_22773,N_15455,N_17008);
or U22774 (N_22774,N_17558,N_15398);
or U22775 (N_22775,N_19358,N_19854);
nor U22776 (N_22776,N_15034,N_17788);
and U22777 (N_22777,N_17880,N_18307);
xor U22778 (N_22778,N_16715,N_17956);
xor U22779 (N_22779,N_18218,N_18311);
nand U22780 (N_22780,N_15705,N_17857);
and U22781 (N_22781,N_16969,N_16048);
xor U22782 (N_22782,N_18432,N_17587);
xor U22783 (N_22783,N_15124,N_17168);
or U22784 (N_22784,N_18791,N_18596);
xor U22785 (N_22785,N_16249,N_15082);
nor U22786 (N_22786,N_15099,N_18480);
and U22787 (N_22787,N_19419,N_16117);
nand U22788 (N_22788,N_18893,N_16033);
or U22789 (N_22789,N_19960,N_19142);
nand U22790 (N_22790,N_15333,N_17590);
nand U22791 (N_22791,N_15445,N_16617);
nor U22792 (N_22792,N_15461,N_19336);
xnor U22793 (N_22793,N_15601,N_16610);
and U22794 (N_22794,N_17283,N_17657);
nor U22795 (N_22795,N_19086,N_17580);
nor U22796 (N_22796,N_18415,N_17012);
or U22797 (N_22797,N_18653,N_17341);
nand U22798 (N_22798,N_18493,N_18495);
xnor U22799 (N_22799,N_18571,N_16890);
or U22800 (N_22800,N_18739,N_15942);
and U22801 (N_22801,N_15183,N_15081);
and U22802 (N_22802,N_18078,N_17379);
or U22803 (N_22803,N_18129,N_16069);
nor U22804 (N_22804,N_15969,N_17910);
nor U22805 (N_22805,N_18789,N_15736);
nand U22806 (N_22806,N_17375,N_16795);
nor U22807 (N_22807,N_19589,N_17814);
nand U22808 (N_22808,N_15942,N_18369);
and U22809 (N_22809,N_17069,N_15718);
nand U22810 (N_22810,N_19371,N_15652);
nand U22811 (N_22811,N_15887,N_16026);
and U22812 (N_22812,N_17622,N_18670);
xnor U22813 (N_22813,N_15295,N_18342);
nor U22814 (N_22814,N_18252,N_17846);
and U22815 (N_22815,N_17097,N_15360);
and U22816 (N_22816,N_16240,N_15476);
and U22817 (N_22817,N_17401,N_19032);
nor U22818 (N_22818,N_18261,N_17563);
nor U22819 (N_22819,N_17944,N_15486);
xnor U22820 (N_22820,N_15565,N_19440);
or U22821 (N_22821,N_15414,N_18035);
and U22822 (N_22822,N_17783,N_16017);
nand U22823 (N_22823,N_18033,N_19647);
xor U22824 (N_22824,N_15193,N_15286);
nor U22825 (N_22825,N_17866,N_17491);
nor U22826 (N_22826,N_16875,N_17479);
nand U22827 (N_22827,N_19049,N_19034);
or U22828 (N_22828,N_16892,N_15000);
nor U22829 (N_22829,N_15138,N_18432);
xor U22830 (N_22830,N_15503,N_17648);
and U22831 (N_22831,N_15589,N_17679);
nand U22832 (N_22832,N_16370,N_18665);
xnor U22833 (N_22833,N_18267,N_19697);
or U22834 (N_22834,N_17829,N_16022);
xor U22835 (N_22835,N_17154,N_15661);
or U22836 (N_22836,N_18590,N_18454);
or U22837 (N_22837,N_19745,N_17408);
nor U22838 (N_22838,N_17198,N_16866);
xnor U22839 (N_22839,N_15121,N_15973);
xnor U22840 (N_22840,N_17484,N_18531);
or U22841 (N_22841,N_16106,N_18560);
nand U22842 (N_22842,N_19928,N_18656);
or U22843 (N_22843,N_16362,N_19158);
and U22844 (N_22844,N_18759,N_16685);
and U22845 (N_22845,N_18493,N_19251);
and U22846 (N_22846,N_18229,N_16062);
or U22847 (N_22847,N_15628,N_18561);
xnor U22848 (N_22848,N_16720,N_17857);
or U22849 (N_22849,N_17015,N_17771);
xor U22850 (N_22850,N_16075,N_16929);
xor U22851 (N_22851,N_19271,N_16676);
nor U22852 (N_22852,N_17870,N_18433);
nand U22853 (N_22853,N_16936,N_15386);
nand U22854 (N_22854,N_15179,N_18144);
and U22855 (N_22855,N_18344,N_15595);
xor U22856 (N_22856,N_17704,N_15565);
and U22857 (N_22857,N_16445,N_15642);
nand U22858 (N_22858,N_15986,N_15864);
xnor U22859 (N_22859,N_17336,N_19451);
or U22860 (N_22860,N_19462,N_17216);
nand U22861 (N_22861,N_16284,N_16098);
and U22862 (N_22862,N_18207,N_15350);
xor U22863 (N_22863,N_17762,N_15441);
xor U22864 (N_22864,N_17809,N_16144);
and U22865 (N_22865,N_19385,N_18563);
xor U22866 (N_22866,N_16068,N_16829);
or U22867 (N_22867,N_16088,N_15316);
and U22868 (N_22868,N_16917,N_18913);
or U22869 (N_22869,N_18196,N_19041);
nand U22870 (N_22870,N_15460,N_15986);
and U22871 (N_22871,N_16828,N_18576);
or U22872 (N_22872,N_17508,N_16628);
or U22873 (N_22873,N_17778,N_19598);
nor U22874 (N_22874,N_18363,N_17165);
nor U22875 (N_22875,N_18366,N_15715);
and U22876 (N_22876,N_15948,N_16798);
nor U22877 (N_22877,N_18573,N_16567);
and U22878 (N_22878,N_15188,N_16079);
xnor U22879 (N_22879,N_19263,N_15473);
nor U22880 (N_22880,N_17294,N_17524);
nand U22881 (N_22881,N_19413,N_15643);
xnor U22882 (N_22882,N_16143,N_18122);
nor U22883 (N_22883,N_17705,N_18775);
or U22884 (N_22884,N_16642,N_16984);
and U22885 (N_22885,N_19954,N_16209);
xor U22886 (N_22886,N_17021,N_18030);
xor U22887 (N_22887,N_15339,N_15837);
and U22888 (N_22888,N_16979,N_19020);
nand U22889 (N_22889,N_19940,N_17706);
or U22890 (N_22890,N_17502,N_18671);
nand U22891 (N_22891,N_16196,N_17407);
or U22892 (N_22892,N_19624,N_16082);
or U22893 (N_22893,N_19125,N_15695);
nand U22894 (N_22894,N_16044,N_17659);
or U22895 (N_22895,N_15792,N_18772);
or U22896 (N_22896,N_15416,N_18147);
nand U22897 (N_22897,N_19353,N_16000);
or U22898 (N_22898,N_17487,N_16868);
nand U22899 (N_22899,N_19546,N_19036);
nand U22900 (N_22900,N_17019,N_17757);
nand U22901 (N_22901,N_17910,N_16874);
xnor U22902 (N_22902,N_18366,N_17665);
nand U22903 (N_22903,N_18249,N_18981);
xnor U22904 (N_22904,N_19861,N_17533);
and U22905 (N_22905,N_18208,N_19248);
xnor U22906 (N_22906,N_15879,N_19997);
xor U22907 (N_22907,N_15088,N_18502);
nand U22908 (N_22908,N_17792,N_16615);
and U22909 (N_22909,N_16144,N_17869);
nor U22910 (N_22910,N_17994,N_17837);
and U22911 (N_22911,N_17154,N_17531);
or U22912 (N_22912,N_15079,N_16396);
nand U22913 (N_22913,N_15711,N_18719);
nor U22914 (N_22914,N_18348,N_19957);
nor U22915 (N_22915,N_19493,N_15857);
xor U22916 (N_22916,N_17226,N_17049);
xnor U22917 (N_22917,N_15986,N_19103);
and U22918 (N_22918,N_18115,N_16914);
nor U22919 (N_22919,N_18739,N_15817);
nand U22920 (N_22920,N_15029,N_16876);
nand U22921 (N_22921,N_15841,N_18753);
or U22922 (N_22922,N_19427,N_19543);
and U22923 (N_22923,N_16449,N_15974);
nor U22924 (N_22924,N_18122,N_16557);
or U22925 (N_22925,N_16541,N_15184);
xor U22926 (N_22926,N_15316,N_15174);
xor U22927 (N_22927,N_17263,N_16446);
or U22928 (N_22928,N_19288,N_18039);
or U22929 (N_22929,N_19465,N_17900);
or U22930 (N_22930,N_18914,N_16952);
nor U22931 (N_22931,N_16246,N_15349);
nor U22932 (N_22932,N_16798,N_17731);
xor U22933 (N_22933,N_19709,N_17693);
xor U22934 (N_22934,N_17354,N_17784);
nand U22935 (N_22935,N_15759,N_18082);
xnor U22936 (N_22936,N_18645,N_19310);
and U22937 (N_22937,N_17885,N_19830);
nand U22938 (N_22938,N_16281,N_15822);
nand U22939 (N_22939,N_17050,N_19602);
nand U22940 (N_22940,N_16128,N_16918);
and U22941 (N_22941,N_17971,N_16158);
nand U22942 (N_22942,N_16318,N_17646);
xnor U22943 (N_22943,N_19973,N_19472);
or U22944 (N_22944,N_17699,N_15778);
nand U22945 (N_22945,N_19849,N_16265);
xor U22946 (N_22946,N_19139,N_17051);
xor U22947 (N_22947,N_16996,N_19266);
nand U22948 (N_22948,N_15659,N_15019);
and U22949 (N_22949,N_17076,N_16123);
xnor U22950 (N_22950,N_18388,N_19413);
nor U22951 (N_22951,N_18320,N_15710);
xnor U22952 (N_22952,N_16499,N_18917);
or U22953 (N_22953,N_17750,N_18480);
and U22954 (N_22954,N_18938,N_17004);
or U22955 (N_22955,N_15311,N_16985);
nand U22956 (N_22956,N_15411,N_19097);
nand U22957 (N_22957,N_15884,N_19356);
and U22958 (N_22958,N_17633,N_19428);
nor U22959 (N_22959,N_15025,N_17755);
nor U22960 (N_22960,N_18765,N_16100);
xnor U22961 (N_22961,N_17018,N_16929);
or U22962 (N_22962,N_17728,N_16515);
and U22963 (N_22963,N_18400,N_19022);
xor U22964 (N_22964,N_16487,N_18879);
and U22965 (N_22965,N_19358,N_17841);
nand U22966 (N_22966,N_18222,N_17730);
nor U22967 (N_22967,N_18059,N_15290);
and U22968 (N_22968,N_15097,N_19474);
xnor U22969 (N_22969,N_15224,N_19344);
and U22970 (N_22970,N_18187,N_19298);
nand U22971 (N_22971,N_19827,N_15127);
nand U22972 (N_22972,N_17391,N_18515);
nor U22973 (N_22973,N_18250,N_17141);
or U22974 (N_22974,N_16088,N_19580);
nor U22975 (N_22975,N_17685,N_19379);
or U22976 (N_22976,N_19168,N_16436);
and U22977 (N_22977,N_16370,N_17369);
or U22978 (N_22978,N_19409,N_15018);
nand U22979 (N_22979,N_15806,N_17567);
and U22980 (N_22980,N_18799,N_17300);
or U22981 (N_22981,N_15763,N_19561);
or U22982 (N_22982,N_19494,N_18011);
xor U22983 (N_22983,N_18016,N_19070);
nand U22984 (N_22984,N_16308,N_18383);
and U22985 (N_22985,N_16581,N_17049);
or U22986 (N_22986,N_19340,N_19263);
or U22987 (N_22987,N_17999,N_16518);
nor U22988 (N_22988,N_16476,N_17901);
nand U22989 (N_22989,N_15485,N_16593);
or U22990 (N_22990,N_19493,N_19057);
xnor U22991 (N_22991,N_15881,N_18696);
and U22992 (N_22992,N_17165,N_19504);
xnor U22993 (N_22993,N_16328,N_16433);
nor U22994 (N_22994,N_16896,N_19682);
or U22995 (N_22995,N_18472,N_18678);
or U22996 (N_22996,N_15079,N_17181);
or U22997 (N_22997,N_15317,N_16645);
xnor U22998 (N_22998,N_19043,N_18984);
or U22999 (N_22999,N_17000,N_15382);
and U23000 (N_23000,N_18016,N_16591);
and U23001 (N_23001,N_17839,N_15843);
and U23002 (N_23002,N_18838,N_16210);
or U23003 (N_23003,N_19818,N_16742);
xnor U23004 (N_23004,N_16588,N_18042);
and U23005 (N_23005,N_15067,N_18487);
or U23006 (N_23006,N_19361,N_16782);
and U23007 (N_23007,N_17421,N_19436);
nand U23008 (N_23008,N_15447,N_19359);
and U23009 (N_23009,N_17920,N_18509);
and U23010 (N_23010,N_16056,N_16608);
nand U23011 (N_23011,N_18610,N_17966);
nor U23012 (N_23012,N_17667,N_17308);
nor U23013 (N_23013,N_17163,N_16000);
nor U23014 (N_23014,N_19103,N_18453);
nand U23015 (N_23015,N_17271,N_18852);
or U23016 (N_23016,N_16038,N_18848);
nor U23017 (N_23017,N_15641,N_18895);
or U23018 (N_23018,N_16454,N_17779);
xnor U23019 (N_23019,N_15181,N_17695);
nor U23020 (N_23020,N_17088,N_19187);
nor U23021 (N_23021,N_19491,N_15424);
nand U23022 (N_23022,N_17812,N_15427);
nor U23023 (N_23023,N_18270,N_16995);
and U23024 (N_23024,N_16723,N_19891);
or U23025 (N_23025,N_15124,N_18538);
nor U23026 (N_23026,N_18164,N_19811);
xnor U23027 (N_23027,N_15023,N_18462);
and U23028 (N_23028,N_19251,N_18344);
and U23029 (N_23029,N_17161,N_18427);
or U23030 (N_23030,N_16602,N_18504);
xor U23031 (N_23031,N_15420,N_17620);
nor U23032 (N_23032,N_15038,N_17812);
nand U23033 (N_23033,N_16445,N_17471);
and U23034 (N_23034,N_15527,N_19736);
or U23035 (N_23035,N_18369,N_15237);
xnor U23036 (N_23036,N_16908,N_18877);
and U23037 (N_23037,N_19563,N_16214);
xor U23038 (N_23038,N_16191,N_18135);
and U23039 (N_23039,N_17046,N_16159);
xnor U23040 (N_23040,N_16598,N_18889);
and U23041 (N_23041,N_15703,N_16047);
and U23042 (N_23042,N_19498,N_15910);
nor U23043 (N_23043,N_19415,N_15482);
nor U23044 (N_23044,N_17229,N_18547);
xnor U23045 (N_23045,N_17616,N_18704);
nand U23046 (N_23046,N_19785,N_18450);
xnor U23047 (N_23047,N_18648,N_17907);
or U23048 (N_23048,N_18463,N_15127);
or U23049 (N_23049,N_19283,N_17071);
and U23050 (N_23050,N_18139,N_17464);
xnor U23051 (N_23051,N_18358,N_19384);
and U23052 (N_23052,N_15865,N_17884);
and U23053 (N_23053,N_15013,N_19315);
or U23054 (N_23054,N_18614,N_18958);
nor U23055 (N_23055,N_17072,N_16245);
nor U23056 (N_23056,N_18590,N_15603);
nand U23057 (N_23057,N_19796,N_18121);
and U23058 (N_23058,N_18401,N_15610);
nor U23059 (N_23059,N_17605,N_17855);
and U23060 (N_23060,N_15515,N_16872);
xor U23061 (N_23061,N_15936,N_18423);
or U23062 (N_23062,N_18563,N_15533);
nor U23063 (N_23063,N_16969,N_19786);
nand U23064 (N_23064,N_15887,N_15896);
and U23065 (N_23065,N_16889,N_16052);
or U23066 (N_23066,N_19635,N_15067);
and U23067 (N_23067,N_17387,N_16222);
xor U23068 (N_23068,N_19730,N_15296);
xnor U23069 (N_23069,N_19770,N_16155);
xnor U23070 (N_23070,N_18209,N_19694);
and U23071 (N_23071,N_15381,N_17808);
nor U23072 (N_23072,N_15759,N_15233);
or U23073 (N_23073,N_17050,N_15636);
and U23074 (N_23074,N_17776,N_15687);
or U23075 (N_23075,N_17583,N_19667);
and U23076 (N_23076,N_17372,N_18409);
nor U23077 (N_23077,N_18454,N_19419);
or U23078 (N_23078,N_15595,N_16671);
nor U23079 (N_23079,N_17011,N_16501);
nor U23080 (N_23080,N_18224,N_19228);
nor U23081 (N_23081,N_17045,N_19372);
or U23082 (N_23082,N_16934,N_19755);
nand U23083 (N_23083,N_15798,N_16587);
and U23084 (N_23084,N_15280,N_18855);
or U23085 (N_23085,N_15335,N_19853);
or U23086 (N_23086,N_19774,N_18071);
or U23087 (N_23087,N_16611,N_16448);
nor U23088 (N_23088,N_15133,N_17498);
nand U23089 (N_23089,N_17672,N_17997);
nand U23090 (N_23090,N_15606,N_17606);
xnor U23091 (N_23091,N_19178,N_16704);
or U23092 (N_23092,N_18947,N_19421);
xnor U23093 (N_23093,N_18215,N_15129);
nand U23094 (N_23094,N_18860,N_17127);
or U23095 (N_23095,N_18872,N_17658);
and U23096 (N_23096,N_19366,N_18490);
nand U23097 (N_23097,N_18160,N_19358);
or U23098 (N_23098,N_16659,N_19114);
or U23099 (N_23099,N_18155,N_17140);
nand U23100 (N_23100,N_17869,N_16773);
or U23101 (N_23101,N_18991,N_18720);
or U23102 (N_23102,N_16538,N_15478);
or U23103 (N_23103,N_19426,N_15139);
or U23104 (N_23104,N_15840,N_18723);
or U23105 (N_23105,N_17651,N_16688);
and U23106 (N_23106,N_15725,N_18650);
or U23107 (N_23107,N_16797,N_19674);
nor U23108 (N_23108,N_19248,N_16088);
and U23109 (N_23109,N_17340,N_19629);
nor U23110 (N_23110,N_15767,N_19064);
nand U23111 (N_23111,N_19678,N_17462);
nor U23112 (N_23112,N_16260,N_15427);
or U23113 (N_23113,N_16785,N_17826);
or U23114 (N_23114,N_16308,N_15613);
xnor U23115 (N_23115,N_18628,N_16994);
and U23116 (N_23116,N_18702,N_17119);
nor U23117 (N_23117,N_19178,N_19512);
xnor U23118 (N_23118,N_15503,N_15499);
nor U23119 (N_23119,N_15632,N_15462);
or U23120 (N_23120,N_16236,N_17022);
nand U23121 (N_23121,N_19605,N_18140);
or U23122 (N_23122,N_15208,N_16468);
or U23123 (N_23123,N_16099,N_17836);
nand U23124 (N_23124,N_17846,N_16257);
xnor U23125 (N_23125,N_17220,N_18909);
nor U23126 (N_23126,N_16650,N_17312);
or U23127 (N_23127,N_18451,N_16497);
and U23128 (N_23128,N_18230,N_18746);
or U23129 (N_23129,N_15491,N_15276);
nand U23130 (N_23130,N_16923,N_17087);
nor U23131 (N_23131,N_15114,N_18188);
xnor U23132 (N_23132,N_15998,N_17843);
nand U23133 (N_23133,N_17863,N_16676);
nor U23134 (N_23134,N_17485,N_17786);
xor U23135 (N_23135,N_16132,N_15877);
nand U23136 (N_23136,N_19276,N_18106);
or U23137 (N_23137,N_15653,N_19110);
nor U23138 (N_23138,N_17919,N_18785);
or U23139 (N_23139,N_17059,N_18748);
xor U23140 (N_23140,N_18520,N_17054);
nor U23141 (N_23141,N_16962,N_18849);
xnor U23142 (N_23142,N_17152,N_16233);
and U23143 (N_23143,N_16579,N_16326);
xnor U23144 (N_23144,N_15031,N_17049);
nor U23145 (N_23145,N_18761,N_15443);
xor U23146 (N_23146,N_15321,N_15129);
and U23147 (N_23147,N_17571,N_18828);
nand U23148 (N_23148,N_18631,N_15540);
nand U23149 (N_23149,N_16614,N_17450);
or U23150 (N_23150,N_15337,N_19410);
nand U23151 (N_23151,N_15662,N_18042);
nand U23152 (N_23152,N_15613,N_17278);
nor U23153 (N_23153,N_16961,N_19130);
nor U23154 (N_23154,N_15857,N_19859);
xor U23155 (N_23155,N_16990,N_16382);
nor U23156 (N_23156,N_17834,N_15818);
and U23157 (N_23157,N_17935,N_19202);
or U23158 (N_23158,N_16531,N_19222);
xor U23159 (N_23159,N_19792,N_16140);
or U23160 (N_23160,N_19302,N_16431);
or U23161 (N_23161,N_18355,N_18575);
and U23162 (N_23162,N_16960,N_19494);
or U23163 (N_23163,N_17779,N_15040);
and U23164 (N_23164,N_15988,N_19049);
nor U23165 (N_23165,N_19504,N_17963);
and U23166 (N_23166,N_17228,N_19941);
xnor U23167 (N_23167,N_17714,N_15178);
or U23168 (N_23168,N_17442,N_16490);
xor U23169 (N_23169,N_16877,N_19858);
and U23170 (N_23170,N_19078,N_18983);
nand U23171 (N_23171,N_19753,N_15100);
nand U23172 (N_23172,N_19737,N_18369);
and U23173 (N_23173,N_15619,N_15514);
or U23174 (N_23174,N_16280,N_19965);
nor U23175 (N_23175,N_18527,N_15088);
nor U23176 (N_23176,N_15063,N_15262);
nor U23177 (N_23177,N_19262,N_16123);
or U23178 (N_23178,N_18045,N_16956);
xnor U23179 (N_23179,N_15223,N_15550);
xnor U23180 (N_23180,N_15016,N_19786);
xnor U23181 (N_23181,N_15507,N_16362);
and U23182 (N_23182,N_17481,N_18019);
nand U23183 (N_23183,N_16878,N_18275);
nand U23184 (N_23184,N_17125,N_16042);
and U23185 (N_23185,N_17903,N_18943);
or U23186 (N_23186,N_15089,N_18040);
nand U23187 (N_23187,N_15423,N_16314);
nor U23188 (N_23188,N_19340,N_19728);
nand U23189 (N_23189,N_17975,N_18016);
nor U23190 (N_23190,N_18971,N_19314);
nor U23191 (N_23191,N_15502,N_18004);
or U23192 (N_23192,N_18586,N_15983);
nor U23193 (N_23193,N_15507,N_16658);
nand U23194 (N_23194,N_19225,N_16627);
and U23195 (N_23195,N_19740,N_17541);
xor U23196 (N_23196,N_19214,N_17157);
xor U23197 (N_23197,N_17695,N_16516);
or U23198 (N_23198,N_19557,N_16642);
nand U23199 (N_23199,N_15262,N_17457);
nand U23200 (N_23200,N_17447,N_16524);
nor U23201 (N_23201,N_16143,N_17613);
and U23202 (N_23202,N_16647,N_18534);
nor U23203 (N_23203,N_16414,N_16684);
and U23204 (N_23204,N_19298,N_19462);
nor U23205 (N_23205,N_18113,N_18173);
nand U23206 (N_23206,N_16277,N_15968);
nand U23207 (N_23207,N_17018,N_15354);
nor U23208 (N_23208,N_15507,N_16983);
nor U23209 (N_23209,N_19664,N_19240);
nand U23210 (N_23210,N_15205,N_16071);
nand U23211 (N_23211,N_16504,N_19197);
or U23212 (N_23212,N_19688,N_17983);
and U23213 (N_23213,N_17353,N_17829);
nand U23214 (N_23214,N_16236,N_16944);
xnor U23215 (N_23215,N_18094,N_19010);
nand U23216 (N_23216,N_19497,N_19548);
nand U23217 (N_23217,N_19404,N_16515);
or U23218 (N_23218,N_17147,N_17178);
nand U23219 (N_23219,N_16407,N_18292);
nand U23220 (N_23220,N_18465,N_19759);
nor U23221 (N_23221,N_19119,N_19449);
and U23222 (N_23222,N_17553,N_18724);
and U23223 (N_23223,N_16359,N_15090);
nand U23224 (N_23224,N_19861,N_15366);
and U23225 (N_23225,N_19920,N_17795);
and U23226 (N_23226,N_16460,N_15193);
xor U23227 (N_23227,N_16860,N_18124);
or U23228 (N_23228,N_18055,N_18540);
nor U23229 (N_23229,N_18158,N_16326);
nor U23230 (N_23230,N_18639,N_18262);
nand U23231 (N_23231,N_19666,N_17658);
and U23232 (N_23232,N_19447,N_19630);
or U23233 (N_23233,N_18397,N_18275);
xnor U23234 (N_23234,N_19706,N_16654);
nor U23235 (N_23235,N_18724,N_18807);
nand U23236 (N_23236,N_17909,N_16860);
and U23237 (N_23237,N_17409,N_15147);
nand U23238 (N_23238,N_16462,N_16837);
xnor U23239 (N_23239,N_17872,N_15394);
nor U23240 (N_23240,N_18671,N_17990);
and U23241 (N_23241,N_18124,N_16732);
or U23242 (N_23242,N_18031,N_18206);
nor U23243 (N_23243,N_19941,N_18495);
and U23244 (N_23244,N_16419,N_18750);
nand U23245 (N_23245,N_16609,N_17139);
or U23246 (N_23246,N_17779,N_19579);
nor U23247 (N_23247,N_15770,N_19303);
nand U23248 (N_23248,N_15128,N_18585);
nor U23249 (N_23249,N_16455,N_15831);
nand U23250 (N_23250,N_19776,N_19345);
and U23251 (N_23251,N_18155,N_18883);
or U23252 (N_23252,N_15993,N_17797);
xor U23253 (N_23253,N_18932,N_19128);
or U23254 (N_23254,N_17115,N_15447);
nor U23255 (N_23255,N_15982,N_15091);
nand U23256 (N_23256,N_19301,N_16879);
nand U23257 (N_23257,N_19729,N_18987);
and U23258 (N_23258,N_16584,N_15907);
nor U23259 (N_23259,N_17230,N_17898);
nor U23260 (N_23260,N_16909,N_16838);
and U23261 (N_23261,N_16223,N_17204);
nor U23262 (N_23262,N_19400,N_18017);
or U23263 (N_23263,N_16202,N_19647);
nand U23264 (N_23264,N_19681,N_18872);
nand U23265 (N_23265,N_17733,N_17703);
nand U23266 (N_23266,N_15227,N_19383);
and U23267 (N_23267,N_18859,N_15505);
nand U23268 (N_23268,N_15005,N_15901);
nor U23269 (N_23269,N_18121,N_16396);
and U23270 (N_23270,N_15255,N_19669);
nor U23271 (N_23271,N_15539,N_16078);
and U23272 (N_23272,N_16253,N_16694);
and U23273 (N_23273,N_19564,N_18713);
nor U23274 (N_23274,N_16042,N_18226);
and U23275 (N_23275,N_18509,N_15721);
or U23276 (N_23276,N_16084,N_19548);
nor U23277 (N_23277,N_19156,N_15318);
nor U23278 (N_23278,N_19481,N_19303);
nand U23279 (N_23279,N_16414,N_18448);
nand U23280 (N_23280,N_16149,N_15423);
xor U23281 (N_23281,N_16774,N_17494);
xor U23282 (N_23282,N_15842,N_18847);
or U23283 (N_23283,N_16001,N_18824);
nand U23284 (N_23284,N_19813,N_19089);
xor U23285 (N_23285,N_15775,N_15935);
and U23286 (N_23286,N_15375,N_18338);
or U23287 (N_23287,N_17739,N_15541);
nand U23288 (N_23288,N_17665,N_19789);
and U23289 (N_23289,N_16226,N_19623);
and U23290 (N_23290,N_17928,N_19118);
nand U23291 (N_23291,N_17299,N_15559);
or U23292 (N_23292,N_19837,N_15891);
and U23293 (N_23293,N_16692,N_18252);
or U23294 (N_23294,N_19815,N_17210);
nand U23295 (N_23295,N_18234,N_19597);
and U23296 (N_23296,N_16853,N_19254);
and U23297 (N_23297,N_18597,N_18116);
or U23298 (N_23298,N_18265,N_18134);
xor U23299 (N_23299,N_16381,N_16120);
xnor U23300 (N_23300,N_18247,N_18642);
or U23301 (N_23301,N_16240,N_15780);
nand U23302 (N_23302,N_19931,N_16947);
and U23303 (N_23303,N_19115,N_17456);
nand U23304 (N_23304,N_18334,N_16704);
xnor U23305 (N_23305,N_15150,N_15031);
xor U23306 (N_23306,N_18913,N_15299);
and U23307 (N_23307,N_15891,N_19865);
and U23308 (N_23308,N_15159,N_18759);
nand U23309 (N_23309,N_19529,N_19881);
and U23310 (N_23310,N_17956,N_18941);
xor U23311 (N_23311,N_17180,N_16169);
or U23312 (N_23312,N_16341,N_16382);
and U23313 (N_23313,N_18714,N_19312);
nor U23314 (N_23314,N_18216,N_15322);
and U23315 (N_23315,N_16251,N_18396);
nand U23316 (N_23316,N_17514,N_19954);
or U23317 (N_23317,N_16576,N_16513);
nor U23318 (N_23318,N_15715,N_17222);
nor U23319 (N_23319,N_15472,N_15945);
or U23320 (N_23320,N_15606,N_17773);
and U23321 (N_23321,N_19968,N_18790);
xor U23322 (N_23322,N_15228,N_18541);
nand U23323 (N_23323,N_17174,N_18611);
xor U23324 (N_23324,N_19582,N_19022);
and U23325 (N_23325,N_19961,N_18877);
xnor U23326 (N_23326,N_15103,N_15901);
nand U23327 (N_23327,N_16030,N_16459);
or U23328 (N_23328,N_16783,N_19888);
nand U23329 (N_23329,N_18440,N_18317);
or U23330 (N_23330,N_17571,N_19552);
or U23331 (N_23331,N_18759,N_18405);
or U23332 (N_23332,N_16834,N_15294);
nor U23333 (N_23333,N_17504,N_19438);
nor U23334 (N_23334,N_16668,N_19634);
nand U23335 (N_23335,N_17432,N_18141);
nor U23336 (N_23336,N_19563,N_17241);
xor U23337 (N_23337,N_17570,N_16701);
and U23338 (N_23338,N_16476,N_19450);
or U23339 (N_23339,N_19874,N_18648);
and U23340 (N_23340,N_18362,N_18431);
nand U23341 (N_23341,N_19467,N_19472);
nor U23342 (N_23342,N_16220,N_17837);
xor U23343 (N_23343,N_17261,N_16605);
nand U23344 (N_23344,N_18494,N_16337);
nand U23345 (N_23345,N_19985,N_19556);
xor U23346 (N_23346,N_18591,N_19211);
or U23347 (N_23347,N_18795,N_17620);
nand U23348 (N_23348,N_15206,N_16037);
or U23349 (N_23349,N_17271,N_19839);
nand U23350 (N_23350,N_18093,N_17544);
and U23351 (N_23351,N_16612,N_18969);
or U23352 (N_23352,N_17133,N_19531);
nand U23353 (N_23353,N_18377,N_16192);
nor U23354 (N_23354,N_15005,N_16020);
or U23355 (N_23355,N_19376,N_19354);
and U23356 (N_23356,N_17675,N_19008);
or U23357 (N_23357,N_18471,N_19891);
nor U23358 (N_23358,N_15426,N_15809);
and U23359 (N_23359,N_15304,N_19057);
or U23360 (N_23360,N_16578,N_16028);
and U23361 (N_23361,N_17738,N_15417);
or U23362 (N_23362,N_16639,N_15951);
nand U23363 (N_23363,N_15999,N_15772);
nand U23364 (N_23364,N_15977,N_17292);
xnor U23365 (N_23365,N_17767,N_18529);
nor U23366 (N_23366,N_18848,N_19116);
nand U23367 (N_23367,N_19257,N_17707);
xor U23368 (N_23368,N_18194,N_16855);
nor U23369 (N_23369,N_16818,N_16006);
nor U23370 (N_23370,N_17466,N_17432);
xnor U23371 (N_23371,N_17557,N_15920);
and U23372 (N_23372,N_17206,N_16371);
nand U23373 (N_23373,N_19376,N_15708);
nand U23374 (N_23374,N_19707,N_16453);
nor U23375 (N_23375,N_15592,N_18138);
xnor U23376 (N_23376,N_17218,N_15981);
nor U23377 (N_23377,N_18201,N_19255);
or U23378 (N_23378,N_17072,N_16112);
and U23379 (N_23379,N_15992,N_18569);
nand U23380 (N_23380,N_15297,N_19942);
and U23381 (N_23381,N_16122,N_15553);
nor U23382 (N_23382,N_17961,N_15058);
or U23383 (N_23383,N_19301,N_17283);
or U23384 (N_23384,N_15141,N_19360);
and U23385 (N_23385,N_19243,N_16107);
xnor U23386 (N_23386,N_16173,N_18037);
xor U23387 (N_23387,N_15704,N_15898);
xor U23388 (N_23388,N_18149,N_16586);
or U23389 (N_23389,N_15451,N_15459);
nand U23390 (N_23390,N_17055,N_17465);
xnor U23391 (N_23391,N_16125,N_16091);
nand U23392 (N_23392,N_15901,N_17821);
or U23393 (N_23393,N_18093,N_16918);
xor U23394 (N_23394,N_15400,N_15715);
and U23395 (N_23395,N_15214,N_18351);
nor U23396 (N_23396,N_16549,N_17236);
and U23397 (N_23397,N_18427,N_18108);
nor U23398 (N_23398,N_15011,N_19215);
nor U23399 (N_23399,N_15670,N_16119);
nand U23400 (N_23400,N_18457,N_18424);
or U23401 (N_23401,N_19624,N_16464);
nand U23402 (N_23402,N_19857,N_15289);
or U23403 (N_23403,N_16222,N_16098);
nand U23404 (N_23404,N_15606,N_16504);
nand U23405 (N_23405,N_19019,N_18383);
nand U23406 (N_23406,N_19749,N_17676);
nor U23407 (N_23407,N_19304,N_15063);
and U23408 (N_23408,N_19218,N_17296);
nor U23409 (N_23409,N_15032,N_16075);
or U23410 (N_23410,N_15661,N_17910);
and U23411 (N_23411,N_19184,N_16361);
nor U23412 (N_23412,N_18896,N_16001);
nand U23413 (N_23413,N_16784,N_16465);
or U23414 (N_23414,N_19762,N_18929);
nor U23415 (N_23415,N_19369,N_15053);
xor U23416 (N_23416,N_16981,N_15141);
nor U23417 (N_23417,N_19870,N_19902);
or U23418 (N_23418,N_18686,N_18371);
nor U23419 (N_23419,N_15771,N_17760);
nand U23420 (N_23420,N_19513,N_16503);
xnor U23421 (N_23421,N_18214,N_19492);
or U23422 (N_23422,N_19854,N_15203);
nor U23423 (N_23423,N_16404,N_17604);
xor U23424 (N_23424,N_17385,N_18219);
xor U23425 (N_23425,N_16673,N_15767);
or U23426 (N_23426,N_19528,N_16993);
and U23427 (N_23427,N_18404,N_16710);
nor U23428 (N_23428,N_16021,N_15008);
xnor U23429 (N_23429,N_17468,N_15253);
nor U23430 (N_23430,N_17408,N_17763);
and U23431 (N_23431,N_15192,N_15082);
nand U23432 (N_23432,N_16485,N_18035);
xor U23433 (N_23433,N_16460,N_16929);
and U23434 (N_23434,N_19752,N_18765);
nand U23435 (N_23435,N_19546,N_18682);
xor U23436 (N_23436,N_16053,N_15250);
or U23437 (N_23437,N_16264,N_18425);
xor U23438 (N_23438,N_15433,N_17465);
nor U23439 (N_23439,N_18305,N_15941);
or U23440 (N_23440,N_17802,N_16161);
nor U23441 (N_23441,N_15490,N_15350);
or U23442 (N_23442,N_19173,N_19639);
nand U23443 (N_23443,N_19960,N_15772);
nor U23444 (N_23444,N_18089,N_15632);
nor U23445 (N_23445,N_18810,N_16918);
nor U23446 (N_23446,N_18196,N_18705);
xor U23447 (N_23447,N_15225,N_16094);
xnor U23448 (N_23448,N_15999,N_19615);
and U23449 (N_23449,N_16812,N_15211);
nor U23450 (N_23450,N_17048,N_19799);
nor U23451 (N_23451,N_15376,N_15850);
nor U23452 (N_23452,N_15396,N_15655);
and U23453 (N_23453,N_18892,N_19612);
nor U23454 (N_23454,N_18450,N_18033);
nor U23455 (N_23455,N_17256,N_16308);
and U23456 (N_23456,N_19293,N_17261);
and U23457 (N_23457,N_18561,N_16507);
or U23458 (N_23458,N_18345,N_15994);
and U23459 (N_23459,N_18553,N_15041);
xnor U23460 (N_23460,N_16913,N_15444);
xnor U23461 (N_23461,N_15697,N_19356);
nand U23462 (N_23462,N_18312,N_18181);
xor U23463 (N_23463,N_18229,N_17817);
and U23464 (N_23464,N_19300,N_19532);
and U23465 (N_23465,N_15489,N_16661);
and U23466 (N_23466,N_15892,N_16435);
nand U23467 (N_23467,N_15834,N_17469);
nor U23468 (N_23468,N_16545,N_19120);
nand U23469 (N_23469,N_18171,N_17257);
and U23470 (N_23470,N_19648,N_19711);
and U23471 (N_23471,N_19009,N_18109);
or U23472 (N_23472,N_19241,N_17823);
nor U23473 (N_23473,N_19312,N_15060);
xor U23474 (N_23474,N_18336,N_15730);
nor U23475 (N_23475,N_16505,N_18188);
xnor U23476 (N_23476,N_17088,N_16453);
or U23477 (N_23477,N_19861,N_17922);
xnor U23478 (N_23478,N_19477,N_18721);
nand U23479 (N_23479,N_18414,N_16041);
or U23480 (N_23480,N_18492,N_19739);
or U23481 (N_23481,N_15613,N_17005);
nor U23482 (N_23482,N_15951,N_15641);
xor U23483 (N_23483,N_17235,N_18103);
or U23484 (N_23484,N_18399,N_17735);
nor U23485 (N_23485,N_18524,N_18719);
nor U23486 (N_23486,N_18507,N_16026);
nand U23487 (N_23487,N_16496,N_16916);
or U23488 (N_23488,N_18061,N_18501);
xnor U23489 (N_23489,N_15196,N_16393);
nor U23490 (N_23490,N_18317,N_16124);
nor U23491 (N_23491,N_16936,N_15092);
or U23492 (N_23492,N_17686,N_17799);
xor U23493 (N_23493,N_17711,N_19523);
or U23494 (N_23494,N_19199,N_18629);
xnor U23495 (N_23495,N_18143,N_19004);
xnor U23496 (N_23496,N_15360,N_19955);
and U23497 (N_23497,N_19153,N_19970);
xnor U23498 (N_23498,N_17719,N_15171);
and U23499 (N_23499,N_15313,N_17266);
xor U23500 (N_23500,N_18592,N_18270);
and U23501 (N_23501,N_17565,N_15292);
xor U23502 (N_23502,N_19214,N_16525);
and U23503 (N_23503,N_15901,N_17302);
nand U23504 (N_23504,N_18976,N_16413);
or U23505 (N_23505,N_18445,N_19906);
or U23506 (N_23506,N_17567,N_18759);
and U23507 (N_23507,N_19599,N_19672);
and U23508 (N_23508,N_17780,N_18605);
nand U23509 (N_23509,N_16828,N_19235);
nand U23510 (N_23510,N_15719,N_19212);
nor U23511 (N_23511,N_19641,N_15474);
and U23512 (N_23512,N_15903,N_15862);
or U23513 (N_23513,N_17266,N_18770);
or U23514 (N_23514,N_17588,N_18327);
and U23515 (N_23515,N_19603,N_15175);
nor U23516 (N_23516,N_17810,N_18736);
nand U23517 (N_23517,N_15082,N_15324);
and U23518 (N_23518,N_17023,N_19913);
and U23519 (N_23519,N_18103,N_16114);
or U23520 (N_23520,N_15904,N_19731);
and U23521 (N_23521,N_19299,N_17585);
nor U23522 (N_23522,N_16268,N_18153);
nor U23523 (N_23523,N_15128,N_16161);
or U23524 (N_23524,N_19510,N_15146);
nand U23525 (N_23525,N_15228,N_16813);
or U23526 (N_23526,N_16193,N_15246);
and U23527 (N_23527,N_15602,N_16660);
or U23528 (N_23528,N_16989,N_19816);
nand U23529 (N_23529,N_18884,N_19142);
xor U23530 (N_23530,N_19378,N_15902);
and U23531 (N_23531,N_18317,N_17819);
and U23532 (N_23532,N_15426,N_18471);
xnor U23533 (N_23533,N_15383,N_18263);
xnor U23534 (N_23534,N_18549,N_15762);
nor U23535 (N_23535,N_15953,N_15802);
xnor U23536 (N_23536,N_18661,N_16578);
xnor U23537 (N_23537,N_19004,N_18402);
and U23538 (N_23538,N_17941,N_17547);
or U23539 (N_23539,N_18396,N_16740);
and U23540 (N_23540,N_17907,N_19225);
nand U23541 (N_23541,N_19636,N_16439);
or U23542 (N_23542,N_17808,N_17334);
nor U23543 (N_23543,N_15139,N_16935);
xnor U23544 (N_23544,N_15086,N_16299);
or U23545 (N_23545,N_17102,N_18579);
or U23546 (N_23546,N_19659,N_17119);
nor U23547 (N_23547,N_15834,N_19230);
and U23548 (N_23548,N_15602,N_19505);
or U23549 (N_23549,N_17183,N_15560);
nor U23550 (N_23550,N_17364,N_16182);
nand U23551 (N_23551,N_16769,N_17780);
or U23552 (N_23552,N_18414,N_16048);
nor U23553 (N_23553,N_17728,N_15591);
xnor U23554 (N_23554,N_15496,N_16921);
or U23555 (N_23555,N_15957,N_18761);
nor U23556 (N_23556,N_16878,N_18821);
xor U23557 (N_23557,N_19401,N_16469);
nor U23558 (N_23558,N_19361,N_15876);
or U23559 (N_23559,N_17706,N_16755);
and U23560 (N_23560,N_16753,N_15555);
nand U23561 (N_23561,N_18303,N_19502);
nand U23562 (N_23562,N_19888,N_15063);
xnor U23563 (N_23563,N_18826,N_16078);
xor U23564 (N_23564,N_15910,N_19142);
nand U23565 (N_23565,N_17356,N_15797);
nand U23566 (N_23566,N_18571,N_16532);
nor U23567 (N_23567,N_17007,N_18825);
and U23568 (N_23568,N_19016,N_16190);
and U23569 (N_23569,N_16974,N_18313);
nor U23570 (N_23570,N_16146,N_15783);
xor U23571 (N_23571,N_17784,N_15827);
nor U23572 (N_23572,N_17331,N_19407);
nand U23573 (N_23573,N_17403,N_15032);
and U23574 (N_23574,N_18184,N_18626);
xnor U23575 (N_23575,N_18473,N_18986);
nand U23576 (N_23576,N_18917,N_16632);
nand U23577 (N_23577,N_17918,N_19994);
and U23578 (N_23578,N_16513,N_15973);
nand U23579 (N_23579,N_16129,N_15478);
nor U23580 (N_23580,N_18470,N_16599);
nand U23581 (N_23581,N_17330,N_18219);
nand U23582 (N_23582,N_18626,N_17705);
and U23583 (N_23583,N_17853,N_19936);
xor U23584 (N_23584,N_17802,N_19295);
or U23585 (N_23585,N_18108,N_15449);
nand U23586 (N_23586,N_19901,N_18318);
or U23587 (N_23587,N_18625,N_17002);
and U23588 (N_23588,N_17474,N_18576);
nor U23589 (N_23589,N_16396,N_17122);
nor U23590 (N_23590,N_15619,N_16781);
xor U23591 (N_23591,N_16095,N_19851);
nor U23592 (N_23592,N_18543,N_17436);
nand U23593 (N_23593,N_17666,N_18179);
xor U23594 (N_23594,N_18576,N_16584);
nor U23595 (N_23595,N_15532,N_15344);
xor U23596 (N_23596,N_19235,N_17470);
or U23597 (N_23597,N_18252,N_19710);
and U23598 (N_23598,N_19987,N_17461);
or U23599 (N_23599,N_16579,N_16560);
or U23600 (N_23600,N_17854,N_17797);
nor U23601 (N_23601,N_15821,N_18517);
or U23602 (N_23602,N_15202,N_15280);
and U23603 (N_23603,N_16638,N_18572);
or U23604 (N_23604,N_16842,N_15138);
nand U23605 (N_23605,N_16071,N_19019);
xnor U23606 (N_23606,N_17134,N_15098);
nor U23607 (N_23607,N_15486,N_19239);
and U23608 (N_23608,N_16966,N_15349);
and U23609 (N_23609,N_17050,N_15653);
and U23610 (N_23610,N_18844,N_19752);
nand U23611 (N_23611,N_19343,N_18537);
nor U23612 (N_23612,N_17615,N_15323);
nand U23613 (N_23613,N_15479,N_19791);
and U23614 (N_23614,N_19082,N_15311);
nor U23615 (N_23615,N_18218,N_15585);
nand U23616 (N_23616,N_17091,N_16069);
and U23617 (N_23617,N_15366,N_16800);
nor U23618 (N_23618,N_18929,N_18434);
xnor U23619 (N_23619,N_17702,N_18046);
xor U23620 (N_23620,N_18920,N_18896);
or U23621 (N_23621,N_18134,N_18785);
nand U23622 (N_23622,N_18635,N_19018);
xor U23623 (N_23623,N_15772,N_16965);
nor U23624 (N_23624,N_19323,N_15708);
nand U23625 (N_23625,N_18122,N_18886);
and U23626 (N_23626,N_15654,N_19722);
xnor U23627 (N_23627,N_15112,N_15204);
nand U23628 (N_23628,N_18621,N_16371);
and U23629 (N_23629,N_17941,N_16657);
nor U23630 (N_23630,N_19871,N_15314);
xnor U23631 (N_23631,N_16762,N_18919);
nor U23632 (N_23632,N_19986,N_17085);
xnor U23633 (N_23633,N_17702,N_16264);
xnor U23634 (N_23634,N_16634,N_18155);
and U23635 (N_23635,N_18268,N_17997);
xnor U23636 (N_23636,N_16494,N_19633);
and U23637 (N_23637,N_17840,N_18049);
nand U23638 (N_23638,N_19843,N_16302);
or U23639 (N_23639,N_19118,N_15914);
nor U23640 (N_23640,N_17040,N_15623);
nand U23641 (N_23641,N_17909,N_17258);
or U23642 (N_23642,N_16511,N_17799);
nor U23643 (N_23643,N_18960,N_16429);
or U23644 (N_23644,N_16319,N_16978);
xnor U23645 (N_23645,N_17913,N_17087);
nand U23646 (N_23646,N_16694,N_16249);
and U23647 (N_23647,N_15514,N_16078);
nand U23648 (N_23648,N_17725,N_15715);
nor U23649 (N_23649,N_17974,N_15482);
xnor U23650 (N_23650,N_16061,N_18902);
xor U23651 (N_23651,N_18635,N_18092);
nor U23652 (N_23652,N_16213,N_18149);
nand U23653 (N_23653,N_18886,N_18053);
or U23654 (N_23654,N_17477,N_15379);
xnor U23655 (N_23655,N_18178,N_19133);
nand U23656 (N_23656,N_17474,N_19674);
nor U23657 (N_23657,N_15088,N_15379);
and U23658 (N_23658,N_16769,N_16428);
or U23659 (N_23659,N_16436,N_17097);
or U23660 (N_23660,N_16629,N_17143);
nor U23661 (N_23661,N_15271,N_18985);
xor U23662 (N_23662,N_15760,N_17717);
or U23663 (N_23663,N_15486,N_17633);
xnor U23664 (N_23664,N_19974,N_19312);
and U23665 (N_23665,N_19876,N_18543);
and U23666 (N_23666,N_18686,N_15400);
or U23667 (N_23667,N_15993,N_17063);
nor U23668 (N_23668,N_16026,N_17023);
xnor U23669 (N_23669,N_17751,N_15647);
and U23670 (N_23670,N_17555,N_15521);
and U23671 (N_23671,N_15866,N_16641);
nand U23672 (N_23672,N_17014,N_18228);
and U23673 (N_23673,N_18882,N_16142);
nor U23674 (N_23674,N_16499,N_15745);
nor U23675 (N_23675,N_18308,N_18270);
nor U23676 (N_23676,N_17996,N_19836);
nor U23677 (N_23677,N_19686,N_16732);
or U23678 (N_23678,N_15065,N_19758);
and U23679 (N_23679,N_17977,N_17135);
or U23680 (N_23680,N_19540,N_16360);
xor U23681 (N_23681,N_18097,N_15479);
nor U23682 (N_23682,N_17751,N_15290);
nor U23683 (N_23683,N_16399,N_16627);
or U23684 (N_23684,N_17396,N_16133);
xnor U23685 (N_23685,N_18453,N_19421);
nand U23686 (N_23686,N_18065,N_18597);
and U23687 (N_23687,N_15036,N_15690);
or U23688 (N_23688,N_16739,N_19276);
xnor U23689 (N_23689,N_16844,N_19702);
or U23690 (N_23690,N_16142,N_15600);
and U23691 (N_23691,N_17117,N_16878);
nand U23692 (N_23692,N_15386,N_18062);
nor U23693 (N_23693,N_17608,N_15719);
or U23694 (N_23694,N_18138,N_15557);
xor U23695 (N_23695,N_15255,N_19308);
and U23696 (N_23696,N_17657,N_17388);
nor U23697 (N_23697,N_16932,N_18325);
nor U23698 (N_23698,N_17499,N_17985);
or U23699 (N_23699,N_16762,N_18969);
nand U23700 (N_23700,N_16545,N_16132);
xor U23701 (N_23701,N_17045,N_18224);
nand U23702 (N_23702,N_19650,N_16373);
nand U23703 (N_23703,N_18228,N_15029);
or U23704 (N_23704,N_16648,N_15501);
or U23705 (N_23705,N_15366,N_15607);
nand U23706 (N_23706,N_16536,N_15569);
and U23707 (N_23707,N_19100,N_19601);
nand U23708 (N_23708,N_19516,N_19974);
nand U23709 (N_23709,N_18080,N_15722);
xnor U23710 (N_23710,N_16674,N_19988);
or U23711 (N_23711,N_18327,N_19359);
nor U23712 (N_23712,N_18739,N_15722);
nand U23713 (N_23713,N_18085,N_15394);
nand U23714 (N_23714,N_15567,N_18912);
and U23715 (N_23715,N_17812,N_17842);
xnor U23716 (N_23716,N_19461,N_17062);
or U23717 (N_23717,N_17336,N_19254);
and U23718 (N_23718,N_18679,N_19836);
nand U23719 (N_23719,N_19491,N_19803);
xor U23720 (N_23720,N_15881,N_19083);
or U23721 (N_23721,N_18597,N_19785);
or U23722 (N_23722,N_15253,N_18450);
nor U23723 (N_23723,N_15380,N_16160);
nand U23724 (N_23724,N_17029,N_19181);
xor U23725 (N_23725,N_15229,N_19127);
or U23726 (N_23726,N_15315,N_19263);
nor U23727 (N_23727,N_16063,N_16743);
xor U23728 (N_23728,N_15814,N_16283);
and U23729 (N_23729,N_15348,N_19122);
xor U23730 (N_23730,N_19077,N_17109);
or U23731 (N_23731,N_18594,N_17502);
or U23732 (N_23732,N_16003,N_16861);
and U23733 (N_23733,N_15107,N_19270);
or U23734 (N_23734,N_18419,N_15420);
xor U23735 (N_23735,N_17919,N_18309);
nand U23736 (N_23736,N_16816,N_16865);
and U23737 (N_23737,N_19450,N_16062);
and U23738 (N_23738,N_17648,N_19956);
and U23739 (N_23739,N_16996,N_15246);
nand U23740 (N_23740,N_16987,N_15839);
and U23741 (N_23741,N_15936,N_19505);
or U23742 (N_23742,N_15489,N_19575);
nor U23743 (N_23743,N_15399,N_16807);
nor U23744 (N_23744,N_18122,N_15522);
and U23745 (N_23745,N_19890,N_19284);
nand U23746 (N_23746,N_18842,N_17112);
nor U23747 (N_23747,N_19492,N_17934);
xnor U23748 (N_23748,N_15120,N_16553);
or U23749 (N_23749,N_16501,N_15803);
nand U23750 (N_23750,N_15299,N_15827);
nand U23751 (N_23751,N_15025,N_18192);
and U23752 (N_23752,N_15159,N_16717);
nor U23753 (N_23753,N_16475,N_15943);
nand U23754 (N_23754,N_17080,N_17719);
nor U23755 (N_23755,N_15692,N_19022);
or U23756 (N_23756,N_16650,N_16591);
xnor U23757 (N_23757,N_17548,N_17560);
nand U23758 (N_23758,N_19914,N_15047);
xor U23759 (N_23759,N_16765,N_15057);
or U23760 (N_23760,N_18626,N_16546);
nand U23761 (N_23761,N_18069,N_15718);
or U23762 (N_23762,N_19681,N_17908);
nor U23763 (N_23763,N_18431,N_15409);
or U23764 (N_23764,N_15296,N_18015);
nor U23765 (N_23765,N_17669,N_15440);
and U23766 (N_23766,N_19942,N_18460);
nand U23767 (N_23767,N_16175,N_17534);
and U23768 (N_23768,N_19351,N_19967);
or U23769 (N_23769,N_15787,N_16000);
xor U23770 (N_23770,N_18052,N_17255);
and U23771 (N_23771,N_19537,N_15262);
xor U23772 (N_23772,N_18430,N_17621);
and U23773 (N_23773,N_18042,N_18165);
or U23774 (N_23774,N_17532,N_18167);
nor U23775 (N_23775,N_15553,N_17275);
xor U23776 (N_23776,N_16604,N_19403);
or U23777 (N_23777,N_15653,N_15179);
and U23778 (N_23778,N_17098,N_17321);
xnor U23779 (N_23779,N_19594,N_17168);
or U23780 (N_23780,N_18172,N_17849);
and U23781 (N_23781,N_19768,N_19694);
xnor U23782 (N_23782,N_18218,N_17918);
nand U23783 (N_23783,N_17930,N_19071);
and U23784 (N_23784,N_15104,N_17765);
or U23785 (N_23785,N_19867,N_18957);
or U23786 (N_23786,N_18155,N_17508);
and U23787 (N_23787,N_17782,N_18334);
nand U23788 (N_23788,N_19562,N_18247);
and U23789 (N_23789,N_19957,N_17600);
and U23790 (N_23790,N_18197,N_19898);
nand U23791 (N_23791,N_17661,N_18841);
nand U23792 (N_23792,N_16744,N_16385);
xnor U23793 (N_23793,N_16423,N_15971);
or U23794 (N_23794,N_16858,N_19191);
xor U23795 (N_23795,N_18685,N_15502);
and U23796 (N_23796,N_18613,N_18578);
nor U23797 (N_23797,N_15962,N_15100);
nand U23798 (N_23798,N_18915,N_19483);
nor U23799 (N_23799,N_17211,N_15256);
xnor U23800 (N_23800,N_19695,N_16969);
nand U23801 (N_23801,N_15844,N_15895);
and U23802 (N_23802,N_18636,N_18692);
xnor U23803 (N_23803,N_18401,N_19783);
nand U23804 (N_23804,N_19522,N_19426);
and U23805 (N_23805,N_18963,N_19374);
nand U23806 (N_23806,N_17088,N_16132);
or U23807 (N_23807,N_17597,N_15313);
nor U23808 (N_23808,N_17215,N_18674);
nor U23809 (N_23809,N_16044,N_16882);
or U23810 (N_23810,N_17159,N_15303);
or U23811 (N_23811,N_18235,N_15454);
nor U23812 (N_23812,N_18938,N_17584);
xor U23813 (N_23813,N_16501,N_16822);
or U23814 (N_23814,N_16917,N_19693);
and U23815 (N_23815,N_16456,N_15170);
or U23816 (N_23816,N_18956,N_17279);
and U23817 (N_23817,N_17369,N_15320);
nor U23818 (N_23818,N_16139,N_17340);
nor U23819 (N_23819,N_19678,N_15751);
nor U23820 (N_23820,N_18331,N_15075);
xnor U23821 (N_23821,N_15495,N_16065);
xor U23822 (N_23822,N_15421,N_19748);
nand U23823 (N_23823,N_18749,N_17714);
and U23824 (N_23824,N_15541,N_17915);
xnor U23825 (N_23825,N_16909,N_17532);
or U23826 (N_23826,N_15254,N_18834);
or U23827 (N_23827,N_18914,N_17823);
xor U23828 (N_23828,N_19537,N_16946);
and U23829 (N_23829,N_19274,N_19127);
nand U23830 (N_23830,N_15677,N_16053);
xor U23831 (N_23831,N_16167,N_18310);
nor U23832 (N_23832,N_18494,N_16986);
nand U23833 (N_23833,N_18992,N_17929);
and U23834 (N_23834,N_17559,N_17385);
nand U23835 (N_23835,N_17344,N_19796);
and U23836 (N_23836,N_16843,N_16528);
nor U23837 (N_23837,N_17613,N_16679);
nand U23838 (N_23838,N_18030,N_19111);
nand U23839 (N_23839,N_15338,N_19636);
nor U23840 (N_23840,N_18075,N_16785);
nor U23841 (N_23841,N_19668,N_15284);
or U23842 (N_23842,N_17554,N_17556);
nor U23843 (N_23843,N_19152,N_19625);
xor U23844 (N_23844,N_19778,N_19537);
and U23845 (N_23845,N_17110,N_19241);
nand U23846 (N_23846,N_16052,N_16086);
nand U23847 (N_23847,N_17428,N_17638);
nor U23848 (N_23848,N_19085,N_18856);
nand U23849 (N_23849,N_18997,N_16898);
xnor U23850 (N_23850,N_15023,N_18856);
and U23851 (N_23851,N_18092,N_16579);
or U23852 (N_23852,N_15998,N_15307);
nor U23853 (N_23853,N_15914,N_19695);
nand U23854 (N_23854,N_15773,N_16006);
and U23855 (N_23855,N_16964,N_17026);
nor U23856 (N_23856,N_19809,N_16646);
nor U23857 (N_23857,N_18104,N_17548);
or U23858 (N_23858,N_17659,N_15587);
nor U23859 (N_23859,N_18797,N_18470);
nand U23860 (N_23860,N_19947,N_18976);
nor U23861 (N_23861,N_17439,N_17595);
nand U23862 (N_23862,N_17797,N_16371);
nor U23863 (N_23863,N_15077,N_19215);
xnor U23864 (N_23864,N_16317,N_15570);
or U23865 (N_23865,N_19758,N_19592);
nand U23866 (N_23866,N_15512,N_19409);
nor U23867 (N_23867,N_18149,N_15683);
nand U23868 (N_23868,N_18392,N_18233);
xnor U23869 (N_23869,N_18309,N_18260);
or U23870 (N_23870,N_17608,N_16058);
and U23871 (N_23871,N_16042,N_16848);
nor U23872 (N_23872,N_16195,N_17264);
and U23873 (N_23873,N_16392,N_17867);
nor U23874 (N_23874,N_16394,N_15234);
nand U23875 (N_23875,N_19516,N_19355);
xnor U23876 (N_23876,N_17052,N_16515);
and U23877 (N_23877,N_15315,N_17541);
nand U23878 (N_23878,N_19053,N_19778);
xnor U23879 (N_23879,N_15207,N_18610);
nor U23880 (N_23880,N_18880,N_17105);
and U23881 (N_23881,N_15357,N_19750);
or U23882 (N_23882,N_15601,N_19659);
and U23883 (N_23883,N_18240,N_16152);
nor U23884 (N_23884,N_19119,N_19825);
xor U23885 (N_23885,N_19765,N_19738);
and U23886 (N_23886,N_16235,N_18322);
nor U23887 (N_23887,N_17432,N_17391);
and U23888 (N_23888,N_16045,N_17812);
xor U23889 (N_23889,N_16449,N_17600);
xor U23890 (N_23890,N_19515,N_16103);
nand U23891 (N_23891,N_18915,N_19857);
or U23892 (N_23892,N_18710,N_16570);
nor U23893 (N_23893,N_17774,N_19788);
nand U23894 (N_23894,N_16582,N_16737);
or U23895 (N_23895,N_17064,N_17340);
or U23896 (N_23896,N_17273,N_19456);
xnor U23897 (N_23897,N_18766,N_19197);
xnor U23898 (N_23898,N_15171,N_19256);
nand U23899 (N_23899,N_17155,N_18562);
or U23900 (N_23900,N_15210,N_16938);
nand U23901 (N_23901,N_17865,N_19163);
nor U23902 (N_23902,N_17635,N_17447);
nor U23903 (N_23903,N_16376,N_17492);
nor U23904 (N_23904,N_16399,N_19383);
or U23905 (N_23905,N_19476,N_17297);
or U23906 (N_23906,N_17672,N_16908);
nand U23907 (N_23907,N_18507,N_16005);
xor U23908 (N_23908,N_15743,N_19400);
or U23909 (N_23909,N_17565,N_15674);
or U23910 (N_23910,N_16372,N_19323);
and U23911 (N_23911,N_15185,N_16759);
nor U23912 (N_23912,N_18427,N_15137);
nor U23913 (N_23913,N_16457,N_17140);
nor U23914 (N_23914,N_17351,N_15043);
and U23915 (N_23915,N_15215,N_16286);
nand U23916 (N_23916,N_16421,N_16732);
or U23917 (N_23917,N_16404,N_19021);
nand U23918 (N_23918,N_17513,N_17721);
xor U23919 (N_23919,N_18501,N_17670);
or U23920 (N_23920,N_18848,N_15863);
or U23921 (N_23921,N_19457,N_18713);
xnor U23922 (N_23922,N_15055,N_17551);
and U23923 (N_23923,N_15418,N_18449);
nor U23924 (N_23924,N_15600,N_17205);
and U23925 (N_23925,N_17590,N_17968);
nand U23926 (N_23926,N_19852,N_19116);
or U23927 (N_23927,N_19526,N_15117);
nor U23928 (N_23928,N_18767,N_19199);
nand U23929 (N_23929,N_16041,N_15072);
nor U23930 (N_23930,N_17055,N_15776);
and U23931 (N_23931,N_15764,N_17190);
and U23932 (N_23932,N_16401,N_19692);
nand U23933 (N_23933,N_16593,N_19853);
nor U23934 (N_23934,N_15483,N_18905);
xnor U23935 (N_23935,N_15418,N_18133);
or U23936 (N_23936,N_16092,N_15994);
nor U23937 (N_23937,N_18179,N_19481);
nor U23938 (N_23938,N_18892,N_18662);
nand U23939 (N_23939,N_19431,N_16668);
and U23940 (N_23940,N_19780,N_16841);
nor U23941 (N_23941,N_16793,N_17260);
xor U23942 (N_23942,N_19308,N_18730);
nand U23943 (N_23943,N_19871,N_15631);
nor U23944 (N_23944,N_19240,N_17259);
and U23945 (N_23945,N_15301,N_16165);
and U23946 (N_23946,N_19805,N_18707);
or U23947 (N_23947,N_17192,N_16321);
nor U23948 (N_23948,N_19091,N_18842);
nand U23949 (N_23949,N_18496,N_16663);
xnor U23950 (N_23950,N_18650,N_17031);
xnor U23951 (N_23951,N_16936,N_16690);
nor U23952 (N_23952,N_16809,N_15729);
nor U23953 (N_23953,N_18574,N_15607);
and U23954 (N_23954,N_19787,N_18947);
nand U23955 (N_23955,N_18558,N_19212);
nand U23956 (N_23956,N_16571,N_16361);
xor U23957 (N_23957,N_17303,N_18773);
nand U23958 (N_23958,N_19522,N_17374);
nand U23959 (N_23959,N_17332,N_19200);
nand U23960 (N_23960,N_19794,N_17645);
and U23961 (N_23961,N_17417,N_16610);
xnor U23962 (N_23962,N_19388,N_19968);
nand U23963 (N_23963,N_16993,N_18568);
nor U23964 (N_23964,N_15599,N_19283);
xnor U23965 (N_23965,N_15914,N_17477);
xnor U23966 (N_23966,N_18395,N_16505);
and U23967 (N_23967,N_15381,N_15797);
nor U23968 (N_23968,N_18328,N_18793);
or U23969 (N_23969,N_19685,N_15786);
nor U23970 (N_23970,N_15571,N_15932);
xor U23971 (N_23971,N_18233,N_16957);
and U23972 (N_23972,N_16630,N_19001);
nand U23973 (N_23973,N_17652,N_18500);
nor U23974 (N_23974,N_16562,N_17988);
nor U23975 (N_23975,N_15721,N_16755);
nand U23976 (N_23976,N_15842,N_17275);
xor U23977 (N_23977,N_19632,N_19940);
nor U23978 (N_23978,N_18220,N_17384);
nand U23979 (N_23979,N_17075,N_19927);
nand U23980 (N_23980,N_15065,N_19122);
and U23981 (N_23981,N_18618,N_19778);
or U23982 (N_23982,N_18295,N_17508);
nor U23983 (N_23983,N_19499,N_19947);
nor U23984 (N_23984,N_15255,N_19198);
xor U23985 (N_23985,N_17308,N_19342);
nand U23986 (N_23986,N_19335,N_16768);
and U23987 (N_23987,N_18977,N_19979);
and U23988 (N_23988,N_19204,N_19337);
xnor U23989 (N_23989,N_16288,N_16745);
nand U23990 (N_23990,N_17978,N_18484);
nand U23991 (N_23991,N_15739,N_19044);
nor U23992 (N_23992,N_15815,N_17518);
xnor U23993 (N_23993,N_16095,N_15399);
nor U23994 (N_23994,N_16699,N_16789);
nand U23995 (N_23995,N_16981,N_19707);
and U23996 (N_23996,N_15852,N_16519);
nor U23997 (N_23997,N_16543,N_19128);
xnor U23998 (N_23998,N_15080,N_17778);
nand U23999 (N_23999,N_19644,N_16114);
nand U24000 (N_24000,N_16554,N_17693);
nand U24001 (N_24001,N_19009,N_19610);
or U24002 (N_24002,N_15877,N_18237);
nor U24003 (N_24003,N_17778,N_15066);
and U24004 (N_24004,N_17257,N_17435);
nand U24005 (N_24005,N_19565,N_17452);
nor U24006 (N_24006,N_16837,N_16604);
nand U24007 (N_24007,N_15900,N_15627);
nand U24008 (N_24008,N_15658,N_18366);
or U24009 (N_24009,N_16713,N_19219);
xor U24010 (N_24010,N_18044,N_17776);
or U24011 (N_24011,N_19242,N_18311);
nor U24012 (N_24012,N_16892,N_16679);
nand U24013 (N_24013,N_17713,N_16297);
nand U24014 (N_24014,N_19751,N_17987);
nand U24015 (N_24015,N_15676,N_17878);
nor U24016 (N_24016,N_16581,N_19095);
nor U24017 (N_24017,N_16595,N_19080);
and U24018 (N_24018,N_17437,N_16158);
nor U24019 (N_24019,N_15272,N_16152);
nand U24020 (N_24020,N_19533,N_17713);
nand U24021 (N_24021,N_17682,N_17977);
nand U24022 (N_24022,N_16250,N_17209);
and U24023 (N_24023,N_15644,N_15581);
nor U24024 (N_24024,N_16831,N_19435);
nor U24025 (N_24025,N_15854,N_15092);
nand U24026 (N_24026,N_18017,N_16855);
or U24027 (N_24027,N_18240,N_19880);
and U24028 (N_24028,N_18002,N_15974);
nor U24029 (N_24029,N_15641,N_16427);
xor U24030 (N_24030,N_17880,N_15133);
xor U24031 (N_24031,N_15192,N_18700);
nand U24032 (N_24032,N_18279,N_15217);
nand U24033 (N_24033,N_17881,N_16272);
nor U24034 (N_24034,N_15925,N_15952);
or U24035 (N_24035,N_19368,N_17445);
and U24036 (N_24036,N_17606,N_15395);
or U24037 (N_24037,N_16679,N_15640);
or U24038 (N_24038,N_19645,N_17688);
xor U24039 (N_24039,N_19128,N_19948);
and U24040 (N_24040,N_19860,N_17524);
nand U24041 (N_24041,N_19745,N_16037);
nand U24042 (N_24042,N_17351,N_18227);
nand U24043 (N_24043,N_16280,N_18798);
nor U24044 (N_24044,N_16404,N_15437);
nor U24045 (N_24045,N_18196,N_18368);
or U24046 (N_24046,N_19070,N_17543);
nor U24047 (N_24047,N_15888,N_17129);
xnor U24048 (N_24048,N_19026,N_17879);
nor U24049 (N_24049,N_19500,N_18331);
nand U24050 (N_24050,N_15134,N_17930);
or U24051 (N_24051,N_18076,N_18811);
xor U24052 (N_24052,N_17093,N_15038);
nor U24053 (N_24053,N_19146,N_17139);
nor U24054 (N_24054,N_17672,N_16102);
or U24055 (N_24055,N_16436,N_17479);
or U24056 (N_24056,N_15149,N_15538);
nand U24057 (N_24057,N_15494,N_15107);
or U24058 (N_24058,N_15226,N_18406);
xnor U24059 (N_24059,N_16515,N_18639);
xor U24060 (N_24060,N_18365,N_17678);
nand U24061 (N_24061,N_15208,N_15716);
xnor U24062 (N_24062,N_18533,N_15978);
nor U24063 (N_24063,N_15386,N_19248);
nand U24064 (N_24064,N_17474,N_16301);
nor U24065 (N_24065,N_15703,N_15804);
or U24066 (N_24066,N_15348,N_16620);
and U24067 (N_24067,N_16380,N_16706);
and U24068 (N_24068,N_17831,N_19505);
xnor U24069 (N_24069,N_15115,N_19643);
or U24070 (N_24070,N_19440,N_15436);
and U24071 (N_24071,N_15289,N_15200);
or U24072 (N_24072,N_19518,N_16527);
nor U24073 (N_24073,N_19378,N_18262);
nand U24074 (N_24074,N_19979,N_17716);
xnor U24075 (N_24075,N_15920,N_17835);
nand U24076 (N_24076,N_15318,N_16851);
xor U24077 (N_24077,N_18315,N_17479);
nor U24078 (N_24078,N_17437,N_15991);
nand U24079 (N_24079,N_15407,N_18729);
nor U24080 (N_24080,N_18487,N_19895);
xnor U24081 (N_24081,N_16984,N_18570);
xnor U24082 (N_24082,N_18767,N_18239);
and U24083 (N_24083,N_18771,N_19632);
and U24084 (N_24084,N_17450,N_17422);
or U24085 (N_24085,N_16653,N_15150);
nor U24086 (N_24086,N_15411,N_19348);
nor U24087 (N_24087,N_16621,N_19653);
nand U24088 (N_24088,N_15255,N_17518);
and U24089 (N_24089,N_15331,N_17595);
xnor U24090 (N_24090,N_18731,N_15130);
xnor U24091 (N_24091,N_17423,N_18911);
nand U24092 (N_24092,N_19766,N_19740);
nand U24093 (N_24093,N_19316,N_19755);
and U24094 (N_24094,N_17588,N_15973);
nand U24095 (N_24095,N_18024,N_16820);
or U24096 (N_24096,N_15073,N_19842);
or U24097 (N_24097,N_16373,N_19548);
nor U24098 (N_24098,N_16434,N_19010);
xor U24099 (N_24099,N_16453,N_19508);
or U24100 (N_24100,N_18364,N_19144);
nor U24101 (N_24101,N_17047,N_17956);
and U24102 (N_24102,N_18473,N_16383);
nand U24103 (N_24103,N_16849,N_18839);
xor U24104 (N_24104,N_15497,N_19226);
xor U24105 (N_24105,N_16203,N_16582);
nand U24106 (N_24106,N_16035,N_16051);
nor U24107 (N_24107,N_18158,N_17634);
and U24108 (N_24108,N_19212,N_15803);
and U24109 (N_24109,N_17355,N_17344);
nor U24110 (N_24110,N_18678,N_19965);
and U24111 (N_24111,N_16670,N_17379);
and U24112 (N_24112,N_17241,N_16801);
xnor U24113 (N_24113,N_18079,N_16959);
xor U24114 (N_24114,N_19372,N_18000);
and U24115 (N_24115,N_18172,N_15162);
or U24116 (N_24116,N_18243,N_19875);
nor U24117 (N_24117,N_17194,N_16708);
xor U24118 (N_24118,N_16009,N_15326);
or U24119 (N_24119,N_16630,N_17274);
nand U24120 (N_24120,N_19509,N_16065);
nand U24121 (N_24121,N_16748,N_18382);
or U24122 (N_24122,N_16043,N_15873);
xnor U24123 (N_24123,N_15882,N_18521);
and U24124 (N_24124,N_19479,N_18119);
nand U24125 (N_24125,N_18284,N_17631);
nand U24126 (N_24126,N_19085,N_16041);
and U24127 (N_24127,N_15638,N_16902);
nand U24128 (N_24128,N_19016,N_15628);
xor U24129 (N_24129,N_16222,N_16240);
xnor U24130 (N_24130,N_15962,N_18148);
xnor U24131 (N_24131,N_15598,N_17003);
xnor U24132 (N_24132,N_17398,N_16126);
and U24133 (N_24133,N_19620,N_18764);
nor U24134 (N_24134,N_19885,N_15026);
nand U24135 (N_24135,N_19121,N_17903);
and U24136 (N_24136,N_16929,N_17906);
nand U24137 (N_24137,N_17926,N_16368);
nand U24138 (N_24138,N_18972,N_16478);
xnor U24139 (N_24139,N_19912,N_15211);
nand U24140 (N_24140,N_17679,N_15032);
nor U24141 (N_24141,N_19126,N_16450);
nor U24142 (N_24142,N_15203,N_17115);
and U24143 (N_24143,N_18702,N_18767);
xnor U24144 (N_24144,N_16242,N_18540);
nand U24145 (N_24145,N_17329,N_17411);
nor U24146 (N_24146,N_16064,N_15338);
and U24147 (N_24147,N_16232,N_15951);
xor U24148 (N_24148,N_16637,N_17853);
nor U24149 (N_24149,N_16289,N_15108);
or U24150 (N_24150,N_18305,N_18906);
and U24151 (N_24151,N_15711,N_18238);
xor U24152 (N_24152,N_15173,N_19746);
and U24153 (N_24153,N_17942,N_15379);
or U24154 (N_24154,N_18633,N_17628);
and U24155 (N_24155,N_17333,N_15812);
and U24156 (N_24156,N_17937,N_18360);
xnor U24157 (N_24157,N_16248,N_16356);
and U24158 (N_24158,N_19945,N_15892);
and U24159 (N_24159,N_18429,N_18458);
xor U24160 (N_24160,N_18532,N_15900);
nor U24161 (N_24161,N_15607,N_15961);
nor U24162 (N_24162,N_18431,N_19401);
nor U24163 (N_24163,N_18410,N_18260);
nor U24164 (N_24164,N_15230,N_18233);
nand U24165 (N_24165,N_17459,N_18516);
and U24166 (N_24166,N_16860,N_17345);
xnor U24167 (N_24167,N_16125,N_15048);
nand U24168 (N_24168,N_17922,N_15143);
nor U24169 (N_24169,N_19478,N_19288);
and U24170 (N_24170,N_15592,N_19921);
nor U24171 (N_24171,N_18716,N_18458);
and U24172 (N_24172,N_15269,N_18347);
xor U24173 (N_24173,N_17392,N_19428);
nand U24174 (N_24174,N_17064,N_15623);
and U24175 (N_24175,N_16642,N_17847);
nand U24176 (N_24176,N_19590,N_15448);
and U24177 (N_24177,N_19975,N_16207);
xnor U24178 (N_24178,N_16240,N_15822);
and U24179 (N_24179,N_18496,N_15025);
nor U24180 (N_24180,N_16232,N_19978);
nand U24181 (N_24181,N_16585,N_17003);
xor U24182 (N_24182,N_16621,N_16251);
nand U24183 (N_24183,N_17254,N_15531);
nand U24184 (N_24184,N_18680,N_17854);
nor U24185 (N_24185,N_16356,N_16686);
or U24186 (N_24186,N_16225,N_19107);
nor U24187 (N_24187,N_18150,N_15634);
or U24188 (N_24188,N_15299,N_17560);
xor U24189 (N_24189,N_16283,N_17069);
nor U24190 (N_24190,N_19210,N_16293);
nor U24191 (N_24191,N_19932,N_16775);
nand U24192 (N_24192,N_16745,N_19401);
nand U24193 (N_24193,N_16143,N_17843);
xor U24194 (N_24194,N_17137,N_18481);
xor U24195 (N_24195,N_17278,N_15158);
and U24196 (N_24196,N_16401,N_15628);
nand U24197 (N_24197,N_17746,N_18435);
and U24198 (N_24198,N_17352,N_17966);
xnor U24199 (N_24199,N_18070,N_17887);
nand U24200 (N_24200,N_15271,N_19194);
nand U24201 (N_24201,N_18208,N_16015);
nand U24202 (N_24202,N_16411,N_17329);
xor U24203 (N_24203,N_17562,N_16110);
or U24204 (N_24204,N_19358,N_16387);
nand U24205 (N_24205,N_15241,N_17499);
and U24206 (N_24206,N_16419,N_15771);
or U24207 (N_24207,N_17863,N_17955);
xnor U24208 (N_24208,N_16557,N_18276);
and U24209 (N_24209,N_16432,N_16962);
nor U24210 (N_24210,N_18349,N_17295);
nor U24211 (N_24211,N_15624,N_16910);
xor U24212 (N_24212,N_19297,N_17742);
nor U24213 (N_24213,N_17119,N_16009);
xor U24214 (N_24214,N_18123,N_17165);
or U24215 (N_24215,N_17155,N_15316);
nand U24216 (N_24216,N_15832,N_15840);
xnor U24217 (N_24217,N_18292,N_16489);
and U24218 (N_24218,N_18095,N_18620);
nor U24219 (N_24219,N_18541,N_18719);
nor U24220 (N_24220,N_17337,N_16150);
nand U24221 (N_24221,N_16042,N_18049);
and U24222 (N_24222,N_17713,N_18125);
and U24223 (N_24223,N_19588,N_15547);
or U24224 (N_24224,N_18077,N_17597);
nor U24225 (N_24225,N_19466,N_18675);
nor U24226 (N_24226,N_17837,N_15207);
nor U24227 (N_24227,N_16455,N_19310);
nand U24228 (N_24228,N_18602,N_19481);
nor U24229 (N_24229,N_18786,N_15482);
xnor U24230 (N_24230,N_15758,N_16569);
nand U24231 (N_24231,N_15179,N_17591);
nor U24232 (N_24232,N_18496,N_19902);
and U24233 (N_24233,N_19557,N_17717);
nand U24234 (N_24234,N_15598,N_18866);
nor U24235 (N_24235,N_15150,N_16057);
nand U24236 (N_24236,N_19737,N_17869);
xor U24237 (N_24237,N_19187,N_15822);
or U24238 (N_24238,N_15858,N_17446);
or U24239 (N_24239,N_17144,N_19132);
nor U24240 (N_24240,N_18699,N_16308);
nor U24241 (N_24241,N_17875,N_18511);
xor U24242 (N_24242,N_18523,N_16465);
or U24243 (N_24243,N_15850,N_17101);
nand U24244 (N_24244,N_15312,N_17862);
or U24245 (N_24245,N_19368,N_19311);
or U24246 (N_24246,N_18831,N_19018);
nor U24247 (N_24247,N_16456,N_18527);
and U24248 (N_24248,N_18260,N_17335);
nand U24249 (N_24249,N_19481,N_17508);
xnor U24250 (N_24250,N_15877,N_16442);
nand U24251 (N_24251,N_18928,N_19375);
nor U24252 (N_24252,N_18781,N_18349);
nor U24253 (N_24253,N_19301,N_15705);
xor U24254 (N_24254,N_17763,N_18665);
nor U24255 (N_24255,N_19582,N_19747);
xnor U24256 (N_24256,N_18718,N_16894);
and U24257 (N_24257,N_19895,N_19088);
nand U24258 (N_24258,N_19368,N_15780);
and U24259 (N_24259,N_18545,N_19130);
xor U24260 (N_24260,N_18284,N_19025);
xor U24261 (N_24261,N_18436,N_19279);
nand U24262 (N_24262,N_16124,N_15678);
and U24263 (N_24263,N_18263,N_15411);
nand U24264 (N_24264,N_16321,N_19117);
nand U24265 (N_24265,N_16813,N_17249);
nand U24266 (N_24266,N_19322,N_15375);
xor U24267 (N_24267,N_15672,N_17702);
or U24268 (N_24268,N_18800,N_15954);
nor U24269 (N_24269,N_19999,N_16364);
nand U24270 (N_24270,N_17991,N_16572);
nand U24271 (N_24271,N_17397,N_16149);
nand U24272 (N_24272,N_16405,N_17271);
nor U24273 (N_24273,N_18636,N_17532);
nand U24274 (N_24274,N_19672,N_17669);
nor U24275 (N_24275,N_18457,N_17724);
xor U24276 (N_24276,N_17882,N_16858);
xnor U24277 (N_24277,N_17141,N_18757);
nor U24278 (N_24278,N_15592,N_19270);
xor U24279 (N_24279,N_18772,N_19179);
or U24280 (N_24280,N_19611,N_15185);
nor U24281 (N_24281,N_15541,N_19205);
nor U24282 (N_24282,N_18985,N_15033);
xnor U24283 (N_24283,N_15915,N_18865);
xnor U24284 (N_24284,N_19576,N_15449);
and U24285 (N_24285,N_19211,N_16659);
or U24286 (N_24286,N_18439,N_18653);
xor U24287 (N_24287,N_17952,N_15686);
or U24288 (N_24288,N_18189,N_17195);
xnor U24289 (N_24289,N_16135,N_15250);
and U24290 (N_24290,N_16994,N_16959);
xor U24291 (N_24291,N_16624,N_16807);
nor U24292 (N_24292,N_19320,N_16553);
and U24293 (N_24293,N_18261,N_17656);
nor U24294 (N_24294,N_15440,N_18367);
xor U24295 (N_24295,N_15362,N_19975);
xor U24296 (N_24296,N_15615,N_17868);
or U24297 (N_24297,N_15445,N_19952);
and U24298 (N_24298,N_15221,N_18999);
nor U24299 (N_24299,N_19493,N_16557);
or U24300 (N_24300,N_15950,N_16658);
or U24301 (N_24301,N_18411,N_19870);
or U24302 (N_24302,N_15408,N_19797);
or U24303 (N_24303,N_17300,N_19260);
or U24304 (N_24304,N_16974,N_17809);
and U24305 (N_24305,N_17695,N_15486);
nor U24306 (N_24306,N_15917,N_15878);
xnor U24307 (N_24307,N_15494,N_18083);
nand U24308 (N_24308,N_18259,N_15831);
nand U24309 (N_24309,N_17293,N_16681);
nand U24310 (N_24310,N_17615,N_19573);
or U24311 (N_24311,N_15313,N_19212);
xor U24312 (N_24312,N_17805,N_16893);
or U24313 (N_24313,N_19170,N_17612);
nor U24314 (N_24314,N_19918,N_18036);
or U24315 (N_24315,N_17638,N_19498);
xor U24316 (N_24316,N_18047,N_18337);
nand U24317 (N_24317,N_15242,N_15276);
nor U24318 (N_24318,N_15861,N_18755);
or U24319 (N_24319,N_18662,N_16368);
nand U24320 (N_24320,N_19038,N_15843);
and U24321 (N_24321,N_16367,N_17667);
nor U24322 (N_24322,N_16346,N_15833);
and U24323 (N_24323,N_17131,N_15447);
xor U24324 (N_24324,N_18892,N_15600);
nand U24325 (N_24325,N_17596,N_16360);
and U24326 (N_24326,N_19030,N_16564);
nor U24327 (N_24327,N_18409,N_15679);
xor U24328 (N_24328,N_17929,N_16133);
and U24329 (N_24329,N_19653,N_18167);
and U24330 (N_24330,N_19956,N_17121);
nand U24331 (N_24331,N_15197,N_17798);
or U24332 (N_24332,N_18409,N_16668);
nor U24333 (N_24333,N_17217,N_16267);
nor U24334 (N_24334,N_19180,N_17761);
nor U24335 (N_24335,N_19721,N_17499);
xnor U24336 (N_24336,N_15004,N_16725);
nand U24337 (N_24337,N_16422,N_19636);
nand U24338 (N_24338,N_19722,N_15656);
and U24339 (N_24339,N_17251,N_17052);
xor U24340 (N_24340,N_17226,N_17792);
nand U24341 (N_24341,N_18480,N_17333);
nand U24342 (N_24342,N_18633,N_18688);
nand U24343 (N_24343,N_19130,N_15613);
nand U24344 (N_24344,N_19673,N_17270);
and U24345 (N_24345,N_15389,N_17190);
nand U24346 (N_24346,N_16105,N_19661);
and U24347 (N_24347,N_15205,N_18514);
nand U24348 (N_24348,N_19249,N_16038);
xnor U24349 (N_24349,N_19752,N_19891);
nor U24350 (N_24350,N_16305,N_18856);
nand U24351 (N_24351,N_15672,N_18840);
and U24352 (N_24352,N_18984,N_15490);
or U24353 (N_24353,N_19097,N_16569);
nand U24354 (N_24354,N_16458,N_18038);
nand U24355 (N_24355,N_15240,N_17908);
nor U24356 (N_24356,N_15892,N_15061);
nand U24357 (N_24357,N_15855,N_17871);
or U24358 (N_24358,N_17248,N_16626);
nand U24359 (N_24359,N_16818,N_16852);
nor U24360 (N_24360,N_15115,N_16692);
xnor U24361 (N_24361,N_15217,N_18977);
or U24362 (N_24362,N_18324,N_18885);
and U24363 (N_24363,N_19350,N_16337);
nand U24364 (N_24364,N_15889,N_16420);
nand U24365 (N_24365,N_16395,N_19095);
or U24366 (N_24366,N_19995,N_15961);
xnor U24367 (N_24367,N_19144,N_16215);
nor U24368 (N_24368,N_19201,N_17885);
xnor U24369 (N_24369,N_15779,N_19046);
nor U24370 (N_24370,N_16774,N_19940);
nor U24371 (N_24371,N_18263,N_15866);
xor U24372 (N_24372,N_15409,N_15981);
xor U24373 (N_24373,N_16184,N_16225);
and U24374 (N_24374,N_17310,N_17766);
and U24375 (N_24375,N_15724,N_19969);
nor U24376 (N_24376,N_17938,N_18041);
xnor U24377 (N_24377,N_19241,N_15516);
nor U24378 (N_24378,N_15578,N_15015);
nand U24379 (N_24379,N_19489,N_18112);
nor U24380 (N_24380,N_15943,N_16866);
nand U24381 (N_24381,N_19615,N_18211);
nor U24382 (N_24382,N_15589,N_19498);
and U24383 (N_24383,N_17947,N_18078);
or U24384 (N_24384,N_15407,N_17043);
nand U24385 (N_24385,N_17661,N_18669);
and U24386 (N_24386,N_17326,N_16928);
nand U24387 (N_24387,N_17824,N_15050);
nand U24388 (N_24388,N_19484,N_19630);
or U24389 (N_24389,N_19397,N_19096);
or U24390 (N_24390,N_16005,N_18355);
or U24391 (N_24391,N_15179,N_17284);
nor U24392 (N_24392,N_17037,N_18736);
or U24393 (N_24393,N_18351,N_19732);
xor U24394 (N_24394,N_18847,N_15015);
nand U24395 (N_24395,N_19376,N_17124);
nand U24396 (N_24396,N_18934,N_19123);
nand U24397 (N_24397,N_15222,N_17230);
xnor U24398 (N_24398,N_17271,N_17189);
nand U24399 (N_24399,N_16480,N_17502);
nor U24400 (N_24400,N_15969,N_16369);
or U24401 (N_24401,N_18230,N_16934);
nor U24402 (N_24402,N_15965,N_19556);
nor U24403 (N_24403,N_15512,N_18525);
nor U24404 (N_24404,N_18014,N_18167);
nand U24405 (N_24405,N_18370,N_16824);
nand U24406 (N_24406,N_16899,N_18151);
and U24407 (N_24407,N_16178,N_17945);
nor U24408 (N_24408,N_17075,N_15200);
nand U24409 (N_24409,N_18957,N_18715);
or U24410 (N_24410,N_19174,N_18851);
nand U24411 (N_24411,N_16669,N_19944);
nor U24412 (N_24412,N_16995,N_15549);
or U24413 (N_24413,N_15364,N_18748);
xor U24414 (N_24414,N_15450,N_16203);
and U24415 (N_24415,N_15320,N_19772);
xnor U24416 (N_24416,N_15081,N_18610);
and U24417 (N_24417,N_19428,N_17299);
nand U24418 (N_24418,N_16015,N_16712);
nand U24419 (N_24419,N_15741,N_16986);
and U24420 (N_24420,N_17434,N_19715);
nand U24421 (N_24421,N_17856,N_16001);
or U24422 (N_24422,N_15684,N_18764);
nand U24423 (N_24423,N_19100,N_19374);
or U24424 (N_24424,N_18525,N_15390);
nand U24425 (N_24425,N_17927,N_15375);
xor U24426 (N_24426,N_19712,N_19872);
or U24427 (N_24427,N_16543,N_16911);
nor U24428 (N_24428,N_18591,N_16923);
or U24429 (N_24429,N_19929,N_15554);
and U24430 (N_24430,N_17651,N_16527);
or U24431 (N_24431,N_15027,N_19866);
xnor U24432 (N_24432,N_19081,N_16109);
or U24433 (N_24433,N_17600,N_19627);
or U24434 (N_24434,N_17650,N_16851);
nand U24435 (N_24435,N_16727,N_16530);
nor U24436 (N_24436,N_15399,N_19019);
nor U24437 (N_24437,N_19985,N_18993);
or U24438 (N_24438,N_16925,N_15463);
or U24439 (N_24439,N_18849,N_15028);
nand U24440 (N_24440,N_18324,N_18714);
and U24441 (N_24441,N_17461,N_18861);
and U24442 (N_24442,N_15940,N_19014);
nor U24443 (N_24443,N_18571,N_15991);
or U24444 (N_24444,N_18177,N_19142);
or U24445 (N_24445,N_15675,N_17892);
or U24446 (N_24446,N_18668,N_15385);
nor U24447 (N_24447,N_18016,N_15330);
nand U24448 (N_24448,N_16515,N_17476);
and U24449 (N_24449,N_16585,N_19540);
xnor U24450 (N_24450,N_15248,N_18184);
xor U24451 (N_24451,N_15329,N_19488);
nand U24452 (N_24452,N_19697,N_16004);
xnor U24453 (N_24453,N_18906,N_19781);
xor U24454 (N_24454,N_15466,N_18265);
and U24455 (N_24455,N_17802,N_17879);
and U24456 (N_24456,N_18529,N_15185);
xor U24457 (N_24457,N_19450,N_16793);
xor U24458 (N_24458,N_16158,N_17778);
and U24459 (N_24459,N_15320,N_19417);
nand U24460 (N_24460,N_19127,N_19638);
or U24461 (N_24461,N_19336,N_16935);
or U24462 (N_24462,N_17734,N_19981);
and U24463 (N_24463,N_19634,N_17988);
nand U24464 (N_24464,N_16433,N_16334);
or U24465 (N_24465,N_16345,N_16699);
xnor U24466 (N_24466,N_17914,N_16663);
or U24467 (N_24467,N_17398,N_16534);
nor U24468 (N_24468,N_15980,N_16618);
or U24469 (N_24469,N_15453,N_18369);
xor U24470 (N_24470,N_16059,N_16704);
or U24471 (N_24471,N_19849,N_19870);
and U24472 (N_24472,N_16140,N_16133);
nand U24473 (N_24473,N_19359,N_15285);
xnor U24474 (N_24474,N_19816,N_17459);
and U24475 (N_24475,N_16988,N_16238);
xor U24476 (N_24476,N_17751,N_15856);
nand U24477 (N_24477,N_15313,N_19720);
or U24478 (N_24478,N_19783,N_19277);
xor U24479 (N_24479,N_17660,N_17522);
xnor U24480 (N_24480,N_15771,N_18339);
nand U24481 (N_24481,N_19273,N_19928);
nand U24482 (N_24482,N_19903,N_18242);
xor U24483 (N_24483,N_18348,N_15438);
and U24484 (N_24484,N_15806,N_15989);
nand U24485 (N_24485,N_18018,N_15230);
or U24486 (N_24486,N_17617,N_16079);
or U24487 (N_24487,N_19159,N_17767);
nand U24488 (N_24488,N_17903,N_19005);
nor U24489 (N_24489,N_19653,N_16265);
or U24490 (N_24490,N_18595,N_19261);
nand U24491 (N_24491,N_15793,N_18865);
and U24492 (N_24492,N_17793,N_16180);
nor U24493 (N_24493,N_17580,N_17889);
nor U24494 (N_24494,N_19470,N_16839);
and U24495 (N_24495,N_19326,N_16075);
and U24496 (N_24496,N_18904,N_19747);
or U24497 (N_24497,N_17280,N_19963);
and U24498 (N_24498,N_18000,N_17463);
xor U24499 (N_24499,N_17463,N_17780);
nand U24500 (N_24500,N_17999,N_16409);
and U24501 (N_24501,N_18286,N_17384);
xnor U24502 (N_24502,N_15957,N_15415);
xor U24503 (N_24503,N_16746,N_17620);
nand U24504 (N_24504,N_16969,N_19689);
nand U24505 (N_24505,N_19475,N_16138);
and U24506 (N_24506,N_18635,N_16072);
xnor U24507 (N_24507,N_19290,N_16494);
nor U24508 (N_24508,N_17014,N_17375);
xnor U24509 (N_24509,N_18275,N_18801);
xor U24510 (N_24510,N_18858,N_15780);
xnor U24511 (N_24511,N_16234,N_17085);
nor U24512 (N_24512,N_16127,N_18401);
and U24513 (N_24513,N_17008,N_16469);
xor U24514 (N_24514,N_16803,N_16517);
or U24515 (N_24515,N_19262,N_15258);
and U24516 (N_24516,N_19477,N_16623);
nand U24517 (N_24517,N_19228,N_17510);
nor U24518 (N_24518,N_15267,N_19729);
nor U24519 (N_24519,N_18215,N_18716);
and U24520 (N_24520,N_15020,N_18709);
nand U24521 (N_24521,N_19074,N_19171);
xor U24522 (N_24522,N_15898,N_18308);
xnor U24523 (N_24523,N_18204,N_17576);
or U24524 (N_24524,N_15679,N_15498);
or U24525 (N_24525,N_17187,N_18841);
nor U24526 (N_24526,N_16591,N_17287);
or U24527 (N_24527,N_18371,N_15810);
or U24528 (N_24528,N_17813,N_17578);
or U24529 (N_24529,N_17062,N_18282);
or U24530 (N_24530,N_15024,N_15214);
and U24531 (N_24531,N_17668,N_17939);
xor U24532 (N_24532,N_17319,N_18340);
or U24533 (N_24533,N_16710,N_18524);
nand U24534 (N_24534,N_17783,N_16278);
and U24535 (N_24535,N_15265,N_18379);
nand U24536 (N_24536,N_19566,N_16477);
nand U24537 (N_24537,N_17246,N_19961);
nand U24538 (N_24538,N_19854,N_18546);
nor U24539 (N_24539,N_19423,N_18908);
xnor U24540 (N_24540,N_18649,N_15888);
and U24541 (N_24541,N_19596,N_16619);
or U24542 (N_24542,N_18591,N_15218);
xor U24543 (N_24543,N_16382,N_15195);
and U24544 (N_24544,N_18102,N_16294);
nand U24545 (N_24545,N_19675,N_19370);
nor U24546 (N_24546,N_18334,N_16332);
or U24547 (N_24547,N_17437,N_17314);
nor U24548 (N_24548,N_15585,N_15874);
and U24549 (N_24549,N_16704,N_15965);
xnor U24550 (N_24550,N_19348,N_17630);
or U24551 (N_24551,N_18314,N_19694);
or U24552 (N_24552,N_18139,N_19837);
nor U24553 (N_24553,N_16620,N_17018);
nand U24554 (N_24554,N_19994,N_17147);
nor U24555 (N_24555,N_18747,N_16707);
xnor U24556 (N_24556,N_19895,N_17429);
or U24557 (N_24557,N_17804,N_19521);
or U24558 (N_24558,N_15599,N_17905);
nand U24559 (N_24559,N_17568,N_16189);
nor U24560 (N_24560,N_17059,N_15283);
nand U24561 (N_24561,N_19281,N_16788);
or U24562 (N_24562,N_19756,N_19044);
xor U24563 (N_24563,N_19997,N_17473);
xor U24564 (N_24564,N_17535,N_16838);
or U24565 (N_24565,N_18421,N_17147);
xnor U24566 (N_24566,N_19792,N_18846);
and U24567 (N_24567,N_19732,N_18913);
or U24568 (N_24568,N_18652,N_18729);
and U24569 (N_24569,N_16235,N_18472);
or U24570 (N_24570,N_16578,N_15425);
and U24571 (N_24571,N_19652,N_18443);
xnor U24572 (N_24572,N_19881,N_16317);
xor U24573 (N_24573,N_18184,N_19165);
nand U24574 (N_24574,N_16648,N_18442);
nand U24575 (N_24575,N_19218,N_19236);
or U24576 (N_24576,N_17837,N_18761);
and U24577 (N_24577,N_15285,N_15992);
nand U24578 (N_24578,N_15754,N_17305);
or U24579 (N_24579,N_17060,N_17861);
xor U24580 (N_24580,N_16540,N_15428);
nand U24581 (N_24581,N_15615,N_17998);
nand U24582 (N_24582,N_17269,N_15697);
and U24583 (N_24583,N_16041,N_15180);
nand U24584 (N_24584,N_16185,N_16621);
or U24585 (N_24585,N_15243,N_19897);
nor U24586 (N_24586,N_16368,N_16435);
xnor U24587 (N_24587,N_17281,N_15000);
nor U24588 (N_24588,N_15968,N_17942);
xor U24589 (N_24589,N_17417,N_18956);
nand U24590 (N_24590,N_18386,N_15874);
and U24591 (N_24591,N_15577,N_19857);
and U24592 (N_24592,N_19178,N_18221);
nand U24593 (N_24593,N_18027,N_16565);
nor U24594 (N_24594,N_16617,N_17978);
nor U24595 (N_24595,N_18579,N_18555);
xor U24596 (N_24596,N_19773,N_16369);
and U24597 (N_24597,N_17927,N_17439);
or U24598 (N_24598,N_18293,N_18178);
nand U24599 (N_24599,N_18417,N_15489);
or U24600 (N_24600,N_18164,N_15170);
nor U24601 (N_24601,N_17920,N_19436);
and U24602 (N_24602,N_19829,N_17562);
nor U24603 (N_24603,N_16847,N_15688);
and U24604 (N_24604,N_15727,N_15267);
xnor U24605 (N_24605,N_15605,N_18318);
xor U24606 (N_24606,N_16723,N_18279);
or U24607 (N_24607,N_15479,N_16824);
or U24608 (N_24608,N_17011,N_19679);
nor U24609 (N_24609,N_15203,N_16263);
or U24610 (N_24610,N_16772,N_16923);
nor U24611 (N_24611,N_17985,N_17896);
or U24612 (N_24612,N_18712,N_18999);
or U24613 (N_24613,N_19508,N_16393);
or U24614 (N_24614,N_19043,N_17939);
xnor U24615 (N_24615,N_16411,N_15876);
and U24616 (N_24616,N_18436,N_16179);
xnor U24617 (N_24617,N_15092,N_15486);
xor U24618 (N_24618,N_19246,N_15499);
nand U24619 (N_24619,N_18690,N_19045);
nand U24620 (N_24620,N_16023,N_19700);
nor U24621 (N_24621,N_16742,N_17995);
and U24622 (N_24622,N_16895,N_17608);
or U24623 (N_24623,N_17313,N_18245);
xnor U24624 (N_24624,N_19546,N_19483);
and U24625 (N_24625,N_18224,N_18903);
or U24626 (N_24626,N_17667,N_15134);
nor U24627 (N_24627,N_16849,N_15979);
nand U24628 (N_24628,N_18906,N_17205);
nand U24629 (N_24629,N_19082,N_17766);
nand U24630 (N_24630,N_18422,N_15312);
or U24631 (N_24631,N_15652,N_15307);
nand U24632 (N_24632,N_16448,N_16641);
nor U24633 (N_24633,N_17776,N_19106);
and U24634 (N_24634,N_16864,N_16234);
and U24635 (N_24635,N_17072,N_18302);
and U24636 (N_24636,N_17587,N_19575);
xnor U24637 (N_24637,N_19281,N_16020);
or U24638 (N_24638,N_19229,N_16313);
nand U24639 (N_24639,N_16006,N_17916);
nor U24640 (N_24640,N_15464,N_19728);
or U24641 (N_24641,N_18327,N_18559);
nor U24642 (N_24642,N_15296,N_16214);
and U24643 (N_24643,N_17345,N_19063);
xor U24644 (N_24644,N_19684,N_18734);
or U24645 (N_24645,N_17595,N_18740);
xnor U24646 (N_24646,N_17974,N_15438);
xnor U24647 (N_24647,N_15113,N_17016);
nand U24648 (N_24648,N_15850,N_15710);
and U24649 (N_24649,N_16360,N_18593);
nand U24650 (N_24650,N_19380,N_18960);
or U24651 (N_24651,N_16941,N_15263);
nor U24652 (N_24652,N_18495,N_16398);
or U24653 (N_24653,N_15037,N_17163);
nand U24654 (N_24654,N_19255,N_18097);
nor U24655 (N_24655,N_18985,N_19320);
nand U24656 (N_24656,N_17679,N_15269);
and U24657 (N_24657,N_17147,N_15239);
nor U24658 (N_24658,N_15465,N_19715);
or U24659 (N_24659,N_17256,N_18910);
nor U24660 (N_24660,N_18774,N_16861);
nor U24661 (N_24661,N_19330,N_18792);
nor U24662 (N_24662,N_17939,N_17193);
xor U24663 (N_24663,N_18533,N_15916);
nor U24664 (N_24664,N_18289,N_15158);
xor U24665 (N_24665,N_15806,N_16579);
or U24666 (N_24666,N_18102,N_17006);
or U24667 (N_24667,N_17284,N_17444);
or U24668 (N_24668,N_15130,N_16898);
nor U24669 (N_24669,N_16417,N_17469);
and U24670 (N_24670,N_16030,N_17086);
or U24671 (N_24671,N_18783,N_17883);
nor U24672 (N_24672,N_18826,N_19727);
nand U24673 (N_24673,N_18490,N_17795);
nand U24674 (N_24674,N_17182,N_17527);
nor U24675 (N_24675,N_18392,N_17051);
xor U24676 (N_24676,N_17007,N_15620);
xnor U24677 (N_24677,N_15037,N_19473);
nand U24678 (N_24678,N_18887,N_19233);
or U24679 (N_24679,N_19342,N_18108);
xnor U24680 (N_24680,N_16818,N_19124);
nand U24681 (N_24681,N_19758,N_17313);
and U24682 (N_24682,N_16654,N_16788);
nand U24683 (N_24683,N_17359,N_15974);
nor U24684 (N_24684,N_19138,N_15675);
nor U24685 (N_24685,N_16255,N_18393);
or U24686 (N_24686,N_17083,N_18823);
or U24687 (N_24687,N_17698,N_17922);
or U24688 (N_24688,N_17254,N_16940);
or U24689 (N_24689,N_18695,N_17825);
and U24690 (N_24690,N_16398,N_17423);
xor U24691 (N_24691,N_19067,N_18637);
nor U24692 (N_24692,N_16411,N_16505);
nand U24693 (N_24693,N_17218,N_18530);
nand U24694 (N_24694,N_16353,N_17597);
and U24695 (N_24695,N_18155,N_18212);
nand U24696 (N_24696,N_18056,N_15203);
nor U24697 (N_24697,N_19673,N_18011);
nor U24698 (N_24698,N_17449,N_15876);
nand U24699 (N_24699,N_17928,N_17324);
nand U24700 (N_24700,N_16297,N_19770);
or U24701 (N_24701,N_16030,N_17190);
or U24702 (N_24702,N_15893,N_16606);
and U24703 (N_24703,N_19814,N_17725);
nor U24704 (N_24704,N_19237,N_16499);
or U24705 (N_24705,N_18173,N_15529);
xnor U24706 (N_24706,N_17702,N_15254);
nor U24707 (N_24707,N_19752,N_19724);
nor U24708 (N_24708,N_16158,N_18592);
nor U24709 (N_24709,N_18664,N_19057);
nand U24710 (N_24710,N_16469,N_18210);
and U24711 (N_24711,N_16368,N_17106);
xnor U24712 (N_24712,N_17720,N_17666);
xnor U24713 (N_24713,N_19788,N_17986);
nor U24714 (N_24714,N_19863,N_18833);
xor U24715 (N_24715,N_15663,N_19569);
nand U24716 (N_24716,N_19246,N_19990);
or U24717 (N_24717,N_19888,N_16899);
and U24718 (N_24718,N_16815,N_18734);
nor U24719 (N_24719,N_18706,N_15509);
xor U24720 (N_24720,N_17266,N_15033);
or U24721 (N_24721,N_18505,N_18021);
xor U24722 (N_24722,N_17285,N_18962);
nor U24723 (N_24723,N_15782,N_15207);
nor U24724 (N_24724,N_15670,N_16772);
nor U24725 (N_24725,N_16261,N_16277);
and U24726 (N_24726,N_15583,N_18028);
and U24727 (N_24727,N_18640,N_17602);
nor U24728 (N_24728,N_18237,N_18888);
and U24729 (N_24729,N_16979,N_17333);
or U24730 (N_24730,N_17979,N_18383);
and U24731 (N_24731,N_18341,N_18250);
nor U24732 (N_24732,N_18378,N_18071);
nor U24733 (N_24733,N_16539,N_19376);
or U24734 (N_24734,N_17960,N_15882);
nand U24735 (N_24735,N_16358,N_17015);
or U24736 (N_24736,N_19227,N_19993);
or U24737 (N_24737,N_18334,N_17384);
xor U24738 (N_24738,N_16614,N_18131);
xor U24739 (N_24739,N_19280,N_19155);
nor U24740 (N_24740,N_15536,N_18686);
or U24741 (N_24741,N_15882,N_18588);
or U24742 (N_24742,N_18092,N_18860);
or U24743 (N_24743,N_16934,N_15186);
and U24744 (N_24744,N_15603,N_16294);
or U24745 (N_24745,N_17097,N_19006);
nand U24746 (N_24746,N_16760,N_17594);
or U24747 (N_24747,N_15127,N_18327);
and U24748 (N_24748,N_15713,N_17852);
or U24749 (N_24749,N_19090,N_15609);
or U24750 (N_24750,N_17620,N_17457);
or U24751 (N_24751,N_16665,N_18462);
nand U24752 (N_24752,N_17585,N_19633);
or U24753 (N_24753,N_18239,N_16873);
nor U24754 (N_24754,N_18603,N_18674);
and U24755 (N_24755,N_16424,N_18083);
nor U24756 (N_24756,N_17630,N_17093);
and U24757 (N_24757,N_18598,N_15323);
nand U24758 (N_24758,N_16006,N_19632);
or U24759 (N_24759,N_19143,N_15665);
nand U24760 (N_24760,N_16968,N_16213);
nand U24761 (N_24761,N_17367,N_18166);
xnor U24762 (N_24762,N_17543,N_16243);
nor U24763 (N_24763,N_15895,N_16635);
nand U24764 (N_24764,N_19187,N_15316);
or U24765 (N_24765,N_15340,N_15610);
nand U24766 (N_24766,N_15957,N_15870);
nor U24767 (N_24767,N_15385,N_15241);
nand U24768 (N_24768,N_18150,N_16428);
nor U24769 (N_24769,N_16103,N_19063);
nor U24770 (N_24770,N_17428,N_16439);
or U24771 (N_24771,N_16953,N_16548);
and U24772 (N_24772,N_17010,N_15349);
or U24773 (N_24773,N_16957,N_18853);
xnor U24774 (N_24774,N_17329,N_16898);
and U24775 (N_24775,N_19262,N_18401);
and U24776 (N_24776,N_16613,N_15216);
xor U24777 (N_24777,N_18316,N_18737);
nor U24778 (N_24778,N_18945,N_18768);
xnor U24779 (N_24779,N_16082,N_15189);
or U24780 (N_24780,N_16846,N_16753);
and U24781 (N_24781,N_19863,N_17401);
nor U24782 (N_24782,N_18850,N_15791);
nand U24783 (N_24783,N_19777,N_18949);
nor U24784 (N_24784,N_17572,N_17764);
xor U24785 (N_24785,N_18904,N_16056);
xnor U24786 (N_24786,N_15050,N_17350);
or U24787 (N_24787,N_16928,N_16543);
nand U24788 (N_24788,N_16942,N_17109);
or U24789 (N_24789,N_18659,N_15830);
or U24790 (N_24790,N_15262,N_19655);
nor U24791 (N_24791,N_19032,N_17225);
nand U24792 (N_24792,N_19402,N_16156);
and U24793 (N_24793,N_18562,N_18286);
nand U24794 (N_24794,N_15782,N_18248);
and U24795 (N_24795,N_17512,N_18189);
nor U24796 (N_24796,N_18520,N_17659);
xnor U24797 (N_24797,N_18099,N_18281);
or U24798 (N_24798,N_15340,N_16434);
and U24799 (N_24799,N_18993,N_15643);
nor U24800 (N_24800,N_19250,N_15302);
nor U24801 (N_24801,N_19303,N_18732);
nand U24802 (N_24802,N_17836,N_17259);
or U24803 (N_24803,N_19345,N_15012);
nor U24804 (N_24804,N_19967,N_19087);
nand U24805 (N_24805,N_16224,N_17572);
and U24806 (N_24806,N_18240,N_17503);
nor U24807 (N_24807,N_15816,N_19618);
xnor U24808 (N_24808,N_16385,N_17615);
and U24809 (N_24809,N_19502,N_18925);
nor U24810 (N_24810,N_17757,N_18477);
nor U24811 (N_24811,N_17429,N_16466);
xor U24812 (N_24812,N_16685,N_17808);
xnor U24813 (N_24813,N_19467,N_19332);
nor U24814 (N_24814,N_16975,N_19899);
or U24815 (N_24815,N_15952,N_18661);
xnor U24816 (N_24816,N_18917,N_18355);
nand U24817 (N_24817,N_18727,N_17759);
nand U24818 (N_24818,N_19822,N_18106);
and U24819 (N_24819,N_15488,N_19053);
or U24820 (N_24820,N_18187,N_19434);
xnor U24821 (N_24821,N_17180,N_16471);
nand U24822 (N_24822,N_16972,N_15284);
nor U24823 (N_24823,N_18639,N_16420);
and U24824 (N_24824,N_16746,N_17426);
nand U24825 (N_24825,N_16264,N_15133);
nand U24826 (N_24826,N_19727,N_17465);
xor U24827 (N_24827,N_18812,N_18196);
or U24828 (N_24828,N_17462,N_19828);
or U24829 (N_24829,N_17175,N_18351);
or U24830 (N_24830,N_16227,N_18658);
nor U24831 (N_24831,N_17222,N_17499);
or U24832 (N_24832,N_15576,N_19393);
or U24833 (N_24833,N_15132,N_18893);
nand U24834 (N_24834,N_16013,N_18496);
xor U24835 (N_24835,N_16287,N_17061);
xor U24836 (N_24836,N_18881,N_15859);
and U24837 (N_24837,N_18808,N_18200);
and U24838 (N_24838,N_19060,N_16381);
xnor U24839 (N_24839,N_16933,N_18267);
xor U24840 (N_24840,N_18815,N_15070);
nor U24841 (N_24841,N_15511,N_16383);
and U24842 (N_24842,N_16824,N_17828);
or U24843 (N_24843,N_17023,N_19834);
or U24844 (N_24844,N_15220,N_18795);
nor U24845 (N_24845,N_16772,N_16346);
nor U24846 (N_24846,N_19217,N_18152);
nor U24847 (N_24847,N_15165,N_17677);
or U24848 (N_24848,N_18959,N_17413);
and U24849 (N_24849,N_18752,N_15836);
nand U24850 (N_24850,N_19783,N_15707);
and U24851 (N_24851,N_17002,N_18347);
xnor U24852 (N_24852,N_16938,N_19269);
or U24853 (N_24853,N_19583,N_16286);
nor U24854 (N_24854,N_18382,N_19955);
or U24855 (N_24855,N_16684,N_16577);
and U24856 (N_24856,N_15701,N_18103);
nor U24857 (N_24857,N_17809,N_18840);
and U24858 (N_24858,N_17782,N_16668);
xnor U24859 (N_24859,N_18135,N_15258);
and U24860 (N_24860,N_15435,N_19114);
or U24861 (N_24861,N_17752,N_15113);
and U24862 (N_24862,N_17564,N_15598);
or U24863 (N_24863,N_18691,N_18321);
xnor U24864 (N_24864,N_17771,N_17552);
nand U24865 (N_24865,N_17538,N_17461);
or U24866 (N_24866,N_17809,N_16616);
nand U24867 (N_24867,N_16731,N_19581);
nand U24868 (N_24868,N_17226,N_16495);
xnor U24869 (N_24869,N_17525,N_19610);
nand U24870 (N_24870,N_17861,N_15270);
nand U24871 (N_24871,N_18285,N_17628);
or U24872 (N_24872,N_16410,N_17881);
and U24873 (N_24873,N_19100,N_18451);
xor U24874 (N_24874,N_19047,N_17033);
nor U24875 (N_24875,N_18698,N_18158);
and U24876 (N_24876,N_17957,N_15186);
xnor U24877 (N_24877,N_16490,N_15439);
xnor U24878 (N_24878,N_19850,N_18680);
nand U24879 (N_24879,N_17700,N_19598);
nor U24880 (N_24880,N_17280,N_17522);
nand U24881 (N_24881,N_15021,N_18940);
or U24882 (N_24882,N_18886,N_16669);
nand U24883 (N_24883,N_19313,N_15697);
or U24884 (N_24884,N_16907,N_18568);
and U24885 (N_24885,N_17420,N_15214);
or U24886 (N_24886,N_18098,N_17371);
or U24887 (N_24887,N_18812,N_19758);
xor U24888 (N_24888,N_15225,N_16897);
nor U24889 (N_24889,N_18581,N_15566);
or U24890 (N_24890,N_18113,N_19772);
nand U24891 (N_24891,N_15344,N_19768);
nand U24892 (N_24892,N_15677,N_19761);
xor U24893 (N_24893,N_17624,N_16781);
nor U24894 (N_24894,N_19654,N_17785);
and U24895 (N_24895,N_18697,N_17382);
and U24896 (N_24896,N_18463,N_18311);
or U24897 (N_24897,N_19528,N_17183);
and U24898 (N_24898,N_16479,N_18734);
xnor U24899 (N_24899,N_17171,N_16089);
xor U24900 (N_24900,N_17036,N_15442);
xor U24901 (N_24901,N_17524,N_19499);
or U24902 (N_24902,N_15825,N_18571);
and U24903 (N_24903,N_15447,N_17090);
nor U24904 (N_24904,N_16677,N_19463);
xor U24905 (N_24905,N_15746,N_17435);
nand U24906 (N_24906,N_17447,N_18397);
xor U24907 (N_24907,N_16735,N_16238);
nor U24908 (N_24908,N_19077,N_15399);
and U24909 (N_24909,N_17104,N_19099);
xor U24910 (N_24910,N_16491,N_15726);
and U24911 (N_24911,N_17857,N_16225);
or U24912 (N_24912,N_15258,N_17300);
nand U24913 (N_24913,N_17019,N_15848);
nor U24914 (N_24914,N_19571,N_15734);
nand U24915 (N_24915,N_19461,N_15863);
and U24916 (N_24916,N_16387,N_16220);
and U24917 (N_24917,N_17753,N_17786);
nand U24918 (N_24918,N_15372,N_15480);
xor U24919 (N_24919,N_18824,N_16733);
nand U24920 (N_24920,N_15483,N_15634);
nor U24921 (N_24921,N_19272,N_19697);
and U24922 (N_24922,N_16063,N_16837);
and U24923 (N_24923,N_17495,N_19521);
nor U24924 (N_24924,N_18516,N_15770);
xor U24925 (N_24925,N_18443,N_18102);
nor U24926 (N_24926,N_17333,N_18895);
and U24927 (N_24927,N_15057,N_18672);
and U24928 (N_24928,N_17316,N_19502);
or U24929 (N_24929,N_18971,N_15873);
and U24930 (N_24930,N_15996,N_16368);
nor U24931 (N_24931,N_17745,N_15707);
and U24932 (N_24932,N_16289,N_18117);
xor U24933 (N_24933,N_17855,N_16700);
or U24934 (N_24934,N_16187,N_19362);
or U24935 (N_24935,N_19239,N_15190);
xor U24936 (N_24936,N_19516,N_19447);
nor U24937 (N_24937,N_19221,N_19448);
or U24938 (N_24938,N_15374,N_17780);
or U24939 (N_24939,N_15230,N_16182);
nor U24940 (N_24940,N_15481,N_19769);
xor U24941 (N_24941,N_16523,N_16521);
xnor U24942 (N_24942,N_18227,N_18136);
nand U24943 (N_24943,N_19299,N_15063);
nor U24944 (N_24944,N_18467,N_17802);
or U24945 (N_24945,N_17856,N_17402);
and U24946 (N_24946,N_17854,N_17880);
nand U24947 (N_24947,N_15147,N_18668);
and U24948 (N_24948,N_18296,N_17195);
and U24949 (N_24949,N_19582,N_19866);
and U24950 (N_24950,N_15530,N_17623);
nor U24951 (N_24951,N_18728,N_15210);
nand U24952 (N_24952,N_15512,N_15488);
nand U24953 (N_24953,N_18529,N_19083);
xor U24954 (N_24954,N_16978,N_18738);
nand U24955 (N_24955,N_18544,N_19261);
and U24956 (N_24956,N_17923,N_16848);
nand U24957 (N_24957,N_16905,N_17277);
or U24958 (N_24958,N_15671,N_17080);
or U24959 (N_24959,N_15631,N_18421);
xnor U24960 (N_24960,N_18742,N_19952);
nor U24961 (N_24961,N_15052,N_17582);
nand U24962 (N_24962,N_15915,N_19047);
nand U24963 (N_24963,N_17256,N_17533);
nor U24964 (N_24964,N_19400,N_15518);
or U24965 (N_24965,N_18681,N_19717);
nand U24966 (N_24966,N_15824,N_19079);
xnor U24967 (N_24967,N_18442,N_18946);
and U24968 (N_24968,N_15555,N_17374);
nand U24969 (N_24969,N_19741,N_18927);
nor U24970 (N_24970,N_19586,N_15303);
and U24971 (N_24971,N_15248,N_17428);
nor U24972 (N_24972,N_16535,N_17475);
or U24973 (N_24973,N_16875,N_18932);
nand U24974 (N_24974,N_17353,N_19056);
or U24975 (N_24975,N_17671,N_17863);
nor U24976 (N_24976,N_17400,N_16166);
nand U24977 (N_24977,N_18430,N_18466);
or U24978 (N_24978,N_19825,N_17496);
xor U24979 (N_24979,N_15046,N_19269);
xnor U24980 (N_24980,N_17361,N_16683);
or U24981 (N_24981,N_18952,N_17856);
or U24982 (N_24982,N_15772,N_16558);
xor U24983 (N_24983,N_15030,N_19292);
and U24984 (N_24984,N_15335,N_18699);
nor U24985 (N_24985,N_16054,N_18273);
xnor U24986 (N_24986,N_18757,N_19092);
nor U24987 (N_24987,N_19217,N_17775);
xnor U24988 (N_24988,N_16790,N_16968);
xor U24989 (N_24989,N_19212,N_15585);
or U24990 (N_24990,N_17151,N_15097);
xnor U24991 (N_24991,N_16010,N_19068);
and U24992 (N_24992,N_19694,N_16970);
nand U24993 (N_24993,N_18222,N_17270);
and U24994 (N_24994,N_17070,N_19795);
nand U24995 (N_24995,N_15525,N_17274);
or U24996 (N_24996,N_17982,N_18600);
xnor U24997 (N_24997,N_17598,N_15220);
nand U24998 (N_24998,N_16111,N_19045);
xnor U24999 (N_24999,N_15304,N_17729);
nand U25000 (N_25000,N_23079,N_24811);
or U25001 (N_25001,N_20707,N_22706);
and U25002 (N_25002,N_20579,N_20733);
nand U25003 (N_25003,N_24870,N_20340);
and U25004 (N_25004,N_21739,N_20725);
nand U25005 (N_25005,N_21789,N_23077);
nand U25006 (N_25006,N_22131,N_24031);
nand U25007 (N_25007,N_21147,N_20095);
and U25008 (N_25008,N_20378,N_21812);
xor U25009 (N_25009,N_20213,N_23496);
nand U25010 (N_25010,N_20215,N_24421);
nor U25011 (N_25011,N_20559,N_21023);
or U25012 (N_25012,N_23540,N_21935);
xnor U25013 (N_25013,N_24224,N_24473);
xnor U25014 (N_25014,N_20483,N_21199);
xor U25015 (N_25015,N_23579,N_21528);
nor U25016 (N_25016,N_22342,N_24877);
and U25017 (N_25017,N_20909,N_21165);
nor U25018 (N_25018,N_23239,N_22176);
nand U25019 (N_25019,N_24586,N_23379);
nand U25020 (N_25020,N_22705,N_22430);
or U25021 (N_25021,N_24374,N_21437);
or U25022 (N_25022,N_24447,N_22134);
and U25023 (N_25023,N_22228,N_24982);
and U25024 (N_25024,N_23783,N_23662);
or U25025 (N_25025,N_23700,N_23698);
or U25026 (N_25026,N_20060,N_23293);
and U25027 (N_25027,N_24449,N_20938);
nand U25028 (N_25028,N_23021,N_22344);
or U25029 (N_25029,N_21021,N_24973);
nor U25030 (N_25030,N_24034,N_24007);
xnor U25031 (N_25031,N_23915,N_24839);
nand U25032 (N_25032,N_20085,N_22335);
xnor U25033 (N_25033,N_21954,N_22460);
or U25034 (N_25034,N_20253,N_22000);
xor U25035 (N_25035,N_20871,N_21681);
nor U25036 (N_25036,N_20341,N_24550);
or U25037 (N_25037,N_21409,N_20965);
xnor U25038 (N_25038,N_21003,N_21560);
or U25039 (N_25039,N_23005,N_24732);
or U25040 (N_25040,N_22455,N_20638);
or U25041 (N_25041,N_24604,N_23420);
nand U25042 (N_25042,N_21218,N_24438);
or U25043 (N_25043,N_20678,N_23311);
or U25044 (N_25044,N_22038,N_21322);
nor U25045 (N_25045,N_23345,N_21007);
xnor U25046 (N_25046,N_23686,N_23096);
nand U25047 (N_25047,N_23946,N_24532);
nor U25048 (N_25048,N_24615,N_20175);
nor U25049 (N_25049,N_22899,N_23369);
nor U25050 (N_25050,N_21672,N_23826);
nand U25051 (N_25051,N_22163,N_24859);
nand U25052 (N_25052,N_21770,N_22249);
and U25053 (N_25053,N_23512,N_20408);
and U25054 (N_25054,N_20220,N_20100);
or U25055 (N_25055,N_23377,N_22402);
nor U25056 (N_25056,N_20715,N_22754);
and U25057 (N_25057,N_24320,N_20154);
and U25058 (N_25058,N_20192,N_20371);
or U25059 (N_25059,N_22803,N_21067);
xor U25060 (N_25060,N_23484,N_20151);
or U25061 (N_25061,N_24233,N_22942);
xnor U25062 (N_25062,N_24630,N_24898);
and U25063 (N_25063,N_24836,N_20551);
nand U25064 (N_25064,N_21821,N_20696);
nand U25065 (N_25065,N_24886,N_21638);
nor U25066 (N_25066,N_21291,N_21829);
nand U25067 (N_25067,N_20432,N_21644);
or U25068 (N_25068,N_23214,N_22216);
xnor U25069 (N_25069,N_23551,N_23749);
and U25070 (N_25070,N_23865,N_24976);
and U25071 (N_25071,N_22900,N_20475);
and U25072 (N_25072,N_21267,N_23268);
or U25073 (N_25073,N_21004,N_24940);
or U25074 (N_25074,N_21828,N_20501);
nand U25075 (N_25075,N_20621,N_20488);
and U25076 (N_25076,N_22734,N_24009);
and U25077 (N_25077,N_20236,N_21832);
nor U25078 (N_25078,N_20446,N_24652);
nand U25079 (N_25079,N_22516,N_22094);
or U25080 (N_25080,N_21036,N_23258);
nor U25081 (N_25081,N_20655,N_20173);
nor U25082 (N_25082,N_22322,N_20476);
or U25083 (N_25083,N_21738,N_23889);
xnor U25084 (N_25084,N_20402,N_20109);
and U25085 (N_25085,N_24749,N_20147);
nand U25086 (N_25086,N_24085,N_21584);
nor U25087 (N_25087,N_20206,N_23559);
nor U25088 (N_25088,N_22640,N_20700);
and U25089 (N_25089,N_20503,N_21498);
xnor U25090 (N_25090,N_23591,N_24515);
nand U25091 (N_25091,N_22477,N_21262);
xor U25092 (N_25092,N_24977,N_22487);
nand U25093 (N_25093,N_23733,N_21532);
or U25094 (N_25094,N_22639,N_23296);
nand U25095 (N_25095,N_22667,N_22977);
nand U25096 (N_25096,N_21453,N_24408);
nand U25097 (N_25097,N_22982,N_23404);
or U25098 (N_25098,N_21966,N_20900);
xor U25099 (N_25099,N_24376,N_22817);
or U25100 (N_25100,N_24847,N_23548);
nand U25101 (N_25101,N_20401,N_23186);
and U25102 (N_25102,N_21546,N_21176);
nand U25103 (N_25103,N_21677,N_20334);
nand U25104 (N_25104,N_22510,N_21772);
xnor U25105 (N_25105,N_20803,N_24993);
and U25106 (N_25106,N_22921,N_24777);
nand U25107 (N_25107,N_24162,N_20308);
nor U25108 (N_25108,N_24778,N_23613);
or U25109 (N_25109,N_23805,N_24834);
or U25110 (N_25110,N_21970,N_23951);
or U25111 (N_25111,N_20016,N_21509);
nor U25112 (N_25112,N_24319,N_23665);
and U25113 (N_25113,N_22913,N_20400);
and U25114 (N_25114,N_20079,N_24776);
and U25115 (N_25115,N_22010,N_24808);
xnor U25116 (N_25116,N_24584,N_24311);
and U25117 (N_25117,N_21104,N_21731);
nand U25118 (N_25118,N_23978,N_23285);
or U25119 (N_25119,N_20982,N_23328);
xnor U25120 (N_25120,N_23460,N_23273);
nor U25121 (N_25121,N_23067,N_22148);
nand U25122 (N_25122,N_20366,N_23059);
and U25123 (N_25123,N_21850,N_22215);
nor U25124 (N_25124,N_22703,N_24582);
nand U25125 (N_25125,N_22443,N_24930);
xor U25126 (N_25126,N_23489,N_21319);
or U25127 (N_25127,N_21796,N_24842);
nand U25128 (N_25128,N_22239,N_23706);
xnor U25129 (N_25129,N_23996,N_21467);
and U25130 (N_25130,N_20823,N_21892);
nor U25131 (N_25131,N_20801,N_22542);
or U25132 (N_25132,N_21006,N_24139);
nand U25133 (N_25133,N_24618,N_20327);
or U25134 (N_25134,N_24503,N_22585);
xnor U25135 (N_25135,N_24869,N_20697);
nor U25136 (N_25136,N_21541,N_24444);
nor U25137 (N_25137,N_23305,N_24362);
xnor U25138 (N_25138,N_24213,N_23942);
or U25139 (N_25139,N_22794,N_20421);
nand U25140 (N_25140,N_23469,N_24094);
nand U25141 (N_25141,N_24664,N_22425);
nor U25142 (N_25142,N_20228,N_24648);
or U25143 (N_25143,N_24414,N_23202);
or U25144 (N_25144,N_22623,N_20728);
and U25145 (N_25145,N_22728,N_21281);
nand U25146 (N_25146,N_24453,N_24632);
or U25147 (N_25147,N_20156,N_22145);
and U25148 (N_25148,N_22528,N_24791);
or U25149 (N_25149,N_21429,N_23923);
nor U25150 (N_25150,N_23012,N_22405);
nor U25151 (N_25151,N_22688,N_23794);
nor U25152 (N_25152,N_24691,N_24764);
or U25153 (N_25153,N_20836,N_24783);
nor U25154 (N_25154,N_20122,N_20407);
xor U25155 (N_25155,N_23791,N_22770);
nand U25156 (N_25156,N_24557,N_24167);
and U25157 (N_25157,N_24159,N_23854);
nand U25158 (N_25158,N_24310,N_21028);
and U25159 (N_25159,N_20758,N_22690);
or U25160 (N_25160,N_22541,N_23103);
xnor U25161 (N_25161,N_24678,N_22065);
and U25162 (N_25162,N_20952,N_24639);
nor U25163 (N_25163,N_21612,N_20703);
or U25164 (N_25164,N_20591,N_24774);
and U25165 (N_25165,N_22363,N_23054);
nor U25166 (N_25166,N_22588,N_24125);
nand U25167 (N_25167,N_21562,N_22272);
nand U25168 (N_25168,N_20118,N_20325);
and U25169 (N_25169,N_21286,N_23307);
nor U25170 (N_25170,N_22472,N_23860);
and U25171 (N_25171,N_22298,N_20108);
xor U25172 (N_25172,N_22896,N_22151);
nand U25173 (N_25173,N_20333,N_20873);
nor U25174 (N_25174,N_20044,N_21486);
or U25175 (N_25175,N_21714,N_22593);
nand U25176 (N_25176,N_21160,N_21988);
xnor U25177 (N_25177,N_22241,N_23809);
xnor U25178 (N_25178,N_21666,N_22212);
nor U25179 (N_25179,N_22649,N_21412);
nor U25180 (N_25180,N_20693,N_24270);
nand U25181 (N_25181,N_20264,N_24357);
nor U25182 (N_25182,N_24535,N_21786);
xor U25183 (N_25183,N_22491,N_20338);
nor U25184 (N_25184,N_23112,N_24264);
nor U25185 (N_25185,N_21591,N_21623);
and U25186 (N_25186,N_21872,N_24546);
or U25187 (N_25187,N_21060,N_24028);
or U25188 (N_25188,N_21436,N_24580);
xor U25189 (N_25189,N_22143,N_24258);
xnor U25190 (N_25190,N_23542,N_23395);
nor U25191 (N_25191,N_20549,N_22079);
nor U25192 (N_25192,N_20106,N_21462);
and U25193 (N_25193,N_21057,N_20732);
nand U25194 (N_25194,N_20928,N_20411);
nor U25195 (N_25195,N_24479,N_20025);
nor U25196 (N_25196,N_24069,N_23736);
xnor U25197 (N_25197,N_24267,N_20508);
and U25198 (N_25198,N_20119,N_24140);
xnor U25199 (N_25199,N_24927,N_23324);
or U25200 (N_25200,N_20478,N_21233);
or U25201 (N_25201,N_21902,N_21080);
or U25202 (N_25202,N_20813,N_21611);
nand U25203 (N_25203,N_21269,N_21408);
or U25204 (N_25204,N_20820,N_21953);
xnor U25205 (N_25205,N_23141,N_22988);
nor U25206 (N_25206,N_23819,N_22799);
and U25207 (N_25207,N_20981,N_24370);
or U25208 (N_25208,N_20645,N_20116);
and U25209 (N_25209,N_21815,N_20365);
or U25210 (N_25210,N_20137,N_21209);
or U25211 (N_25211,N_20917,N_24385);
nor U25212 (N_25212,N_20767,N_20959);
nor U25213 (N_25213,N_24731,N_20642);
and U25214 (N_25214,N_22650,N_21143);
nor U25215 (N_25215,N_22167,N_20690);
and U25216 (N_25216,N_20738,N_20633);
or U25217 (N_25217,N_22610,N_23456);
xor U25218 (N_25218,N_23066,N_22328);
nor U25219 (N_25219,N_20515,N_21764);
or U25220 (N_25220,N_22409,N_23892);
and U25221 (N_25221,N_20632,N_21665);
nor U25222 (N_25222,N_22692,N_24323);
and U25223 (N_25223,N_21097,N_21774);
or U25224 (N_25224,N_22677,N_21840);
nor U25225 (N_25225,N_21676,N_22397);
or U25226 (N_25226,N_21943,N_22012);
xor U25227 (N_25227,N_23343,N_20331);
nor U25228 (N_25228,N_23424,N_22671);
and U25229 (N_25229,N_24480,N_22424);
or U25230 (N_25230,N_20737,N_24809);
and U25231 (N_25231,N_22445,N_20679);
nor U25232 (N_25232,N_21159,N_21008);
nand U25233 (N_25233,N_22313,N_20187);
nand U25234 (N_25234,N_24396,N_20208);
or U25235 (N_25235,N_22822,N_22108);
or U25236 (N_25236,N_20948,N_21752);
and U25237 (N_25237,N_20027,N_21535);
nor U25238 (N_25238,N_23333,N_21607);
nor U25239 (N_25239,N_21108,N_24205);
nand U25240 (N_25240,N_22380,N_21765);
nor U25241 (N_25241,N_22932,N_20272);
xnor U25242 (N_25242,N_21551,N_23695);
nor U25243 (N_25243,N_21873,N_23020);
nand U25244 (N_25244,N_22251,N_23742);
and U25245 (N_25245,N_21507,N_23175);
nand U25246 (N_25246,N_24921,N_21635);
and U25247 (N_25247,N_20763,N_23385);
xor U25248 (N_25248,N_20218,N_24063);
xnor U25249 (N_25249,N_21382,N_20362);
or U25250 (N_25250,N_24722,N_20103);
nor U25251 (N_25251,N_20356,N_21581);
xnor U25252 (N_25252,N_24670,N_22598);
xor U25253 (N_25253,N_21245,N_20266);
and U25254 (N_25254,N_20500,N_24888);
and U25255 (N_25255,N_20162,N_20915);
or U25256 (N_25256,N_23786,N_22435);
or U25257 (N_25257,N_23832,N_20851);
or U25258 (N_25258,N_20453,N_24945);
xnor U25259 (N_25259,N_22992,N_22165);
or U25260 (N_25260,N_22985,N_21307);
or U25261 (N_25261,N_24173,N_20854);
xor U25262 (N_25262,N_20399,N_24278);
and U25263 (N_25263,N_22261,N_24908);
or U25264 (N_25264,N_21805,N_24342);
nand U25265 (N_25265,N_22871,N_20412);
and U25266 (N_25266,N_20934,N_20513);
and U25267 (N_25267,N_24341,N_20904);
nor U25268 (N_25268,N_22604,N_20870);
xor U25269 (N_25269,N_21250,N_23200);
nor U25270 (N_25270,N_21346,N_23183);
xor U25271 (N_25271,N_20950,N_21554);
nand U25272 (N_25272,N_22776,N_22501);
nor U25273 (N_25273,N_23022,N_23035);
xnor U25274 (N_25274,N_24938,N_20604);
or U25275 (N_25275,N_22087,N_23234);
nand U25276 (N_25276,N_20166,N_22037);
or U25277 (N_25277,N_23666,N_20350);
or U25278 (N_25278,N_24553,N_20744);
xnor U25279 (N_25279,N_22950,N_23121);
xnor U25280 (N_25280,N_24710,N_20564);
xnor U25281 (N_25281,N_23499,N_22696);
and U25282 (N_25282,N_21087,N_23939);
nand U25283 (N_25283,N_20382,N_24784);
xnor U25284 (N_25284,N_20742,N_24292);
nand U25285 (N_25285,N_21602,N_23004);
nand U25286 (N_25286,N_22007,N_23509);
nand U25287 (N_25287,N_21019,N_20720);
and U25288 (N_25288,N_22918,N_24299);
or U25289 (N_25289,N_20473,N_23914);
nand U25290 (N_25290,N_24241,N_24057);
xor U25291 (N_25291,N_21625,N_21440);
nand U25292 (N_25292,N_24084,N_20302);
nor U25293 (N_25293,N_24529,N_24860);
nand U25294 (N_25294,N_21733,N_24166);
and U25295 (N_25295,N_24617,N_21134);
xnor U25296 (N_25296,N_21481,N_23431);
xnor U25297 (N_25297,N_21180,N_21646);
xor U25298 (N_25298,N_20837,N_24038);
and U25299 (N_25299,N_21972,N_24683);
and U25300 (N_25300,N_21010,N_21070);
xor U25301 (N_25301,N_24955,N_20385);
nand U25302 (N_25302,N_23006,N_23956);
or U25303 (N_25303,N_23415,N_23494);
or U25304 (N_25304,N_21787,N_21356);
nor U25305 (N_25305,N_21015,N_23884);
xnor U25306 (N_25306,N_20469,N_20342);
or U25307 (N_25307,N_21634,N_20189);
xor U25308 (N_25308,N_21388,N_23954);
nand U25309 (N_25309,N_24464,N_23435);
or U25310 (N_25310,N_24690,N_24829);
nand U25311 (N_25311,N_21597,N_21277);
nor U25312 (N_25312,N_22157,N_21013);
and U25313 (N_25313,N_21848,N_20439);
or U25314 (N_25314,N_23359,N_22778);
nor U25315 (N_25315,N_20739,N_24493);
and U25316 (N_25316,N_20148,N_21982);
nor U25317 (N_25317,N_22810,N_23891);
xor U25318 (N_25318,N_24720,N_24100);
and U25319 (N_25319,N_20277,N_22872);
xnor U25320 (N_25320,N_23936,N_21038);
or U25321 (N_25321,N_24407,N_24637);
nor U25322 (N_25322,N_21565,N_20096);
nand U25323 (N_25323,N_20883,N_21707);
and U25324 (N_25324,N_21193,N_23229);
nand U25325 (N_25325,N_23085,N_24257);
or U25326 (N_25326,N_20072,N_21167);
nor U25327 (N_25327,N_21282,N_22707);
xor U25328 (N_25328,N_23432,N_24855);
xor U25329 (N_25329,N_23668,N_24935);
and U25330 (N_25330,N_23215,N_20456);
xor U25331 (N_25331,N_21803,N_24857);
and U25332 (N_25332,N_20171,N_20988);
xnor U25333 (N_25333,N_23885,N_23075);
or U25334 (N_25334,N_20177,N_20230);
or U25335 (N_25335,N_21398,N_23701);
xor U25336 (N_25336,N_23152,N_22139);
nor U25337 (N_25337,N_20750,N_20319);
and U25338 (N_25338,N_20927,N_22193);
or U25339 (N_25339,N_22168,N_21136);
and U25340 (N_25340,N_24765,N_24390);
or U25341 (N_25341,N_24075,N_23194);
nor U25342 (N_25342,N_21480,N_21129);
or U25343 (N_25343,N_23032,N_21457);
xor U25344 (N_25344,N_23501,N_20993);
nor U25345 (N_25345,N_23381,N_21867);
or U25346 (N_25346,N_20355,N_22359);
nand U25347 (N_25347,N_20903,N_24246);
and U25348 (N_25348,N_24519,N_23949);
xnor U25349 (N_25349,N_23840,N_24215);
nand U25350 (N_25350,N_20433,N_20512);
or U25351 (N_25351,N_23441,N_24295);
nor U25352 (N_25352,N_20262,N_20451);
and U25353 (N_25353,N_20799,N_21368);
nand U25354 (N_25354,N_23882,N_23127);
nor U25355 (N_25355,N_20202,N_23161);
nand U25356 (N_25356,N_23257,N_21247);
nand U25357 (N_25357,N_24450,N_20083);
nand U25358 (N_25358,N_22791,N_21278);
or U25359 (N_25359,N_20797,N_21582);
nand U25360 (N_25360,N_22779,N_22732);
and U25361 (N_25361,N_24244,N_23045);
nand U25362 (N_25362,N_21074,N_24271);
nor U25363 (N_25363,N_24329,N_20076);
and U25364 (N_25364,N_24203,N_24207);
nor U25365 (N_25365,N_20448,N_23836);
nand U25366 (N_25366,N_22373,N_20358);
and U25367 (N_25367,N_23696,N_23741);
and U25368 (N_25368,N_22971,N_23052);
or U25369 (N_25369,N_23301,N_22551);
xnor U25370 (N_25370,N_24497,N_24810);
nor U25371 (N_25371,N_21678,N_21637);
and U25372 (N_25372,N_22571,N_22508);
nor U25373 (N_25373,N_20425,N_23259);
nand U25374 (N_25374,N_22194,N_22751);
and U25375 (N_25375,N_20650,N_24466);
or U25376 (N_25376,N_23216,N_22225);
and U25377 (N_25377,N_20858,N_20905);
and U25378 (N_25378,N_22310,N_22600);
xnor U25379 (N_25379,N_24923,N_22815);
or U25380 (N_25380,N_21654,N_24850);
or U25381 (N_25381,N_21066,N_21161);
xnor U25382 (N_25382,N_22539,N_21920);
nor U25383 (N_25383,N_23189,N_24204);
nor U25384 (N_25384,N_24538,N_20681);
and U25385 (N_25385,N_23750,N_24440);
xor U25386 (N_25386,N_21339,N_23875);
nand U25387 (N_25387,N_22597,N_24255);
nor U25388 (N_25388,N_22916,N_22956);
or U25389 (N_25389,N_24906,N_23777);
nand U25390 (N_25390,N_22886,N_20388);
nand U25391 (N_25391,N_20997,N_21993);
and U25392 (N_25392,N_23876,N_21253);
or U25393 (N_25393,N_20946,N_22333);
or U25394 (N_25394,N_22155,N_21775);
nor U25395 (N_25395,N_22426,N_22820);
or U25396 (N_25396,N_22323,N_21293);
xnor U25397 (N_25397,N_24049,N_20683);
and U25398 (N_25398,N_21076,N_24136);
and U25399 (N_25399,N_23410,N_23461);
xnor U25400 (N_25400,N_23523,N_22868);
xnor U25401 (N_25401,N_22753,N_20040);
xor U25402 (N_25402,N_24435,N_21170);
and U25403 (N_25403,N_24891,N_20879);
nand U25404 (N_25404,N_24965,N_22264);
or U25405 (N_25405,N_22968,N_22917);
xor U25406 (N_25406,N_23960,N_21360);
or U25407 (N_25407,N_24781,N_20393);
and U25408 (N_25408,N_20901,N_21397);
or U25409 (N_25409,N_24415,N_21987);
nor U25410 (N_25410,N_24876,N_20567);
nand U25411 (N_25411,N_22031,N_21925);
xor U25412 (N_25412,N_20051,N_21751);
and U25413 (N_25413,N_22800,N_23557);
nand U25414 (N_25414,N_21410,N_23010);
xnor U25415 (N_25415,N_21425,N_20863);
or U25416 (N_25416,N_22898,N_21556);
nand U25417 (N_25417,N_20450,N_22574);
or U25418 (N_25418,N_20140,N_21434);
xor U25419 (N_25419,N_23237,N_24812);
nor U25420 (N_25420,N_24423,N_23147);
or U25421 (N_25421,N_22944,N_21794);
or U25422 (N_25422,N_21373,N_22417);
and U25423 (N_25423,N_24117,N_23877);
xor U25424 (N_25424,N_21862,N_22920);
nor U25425 (N_25425,N_20753,N_21355);
and U25426 (N_25426,N_23294,N_20465);
nand U25427 (N_25427,N_20844,N_20182);
and U25428 (N_25428,N_22523,N_21609);
or U25429 (N_25429,N_21913,N_20541);
nand U25430 (N_25430,N_21485,N_21506);
xnor U25431 (N_25431,N_23197,N_22080);
nor U25432 (N_25432,N_21626,N_23247);
nand U25433 (N_25433,N_22580,N_21690);
xor U25434 (N_25434,N_23961,N_20613);
and U25435 (N_25435,N_24872,N_22881);
nand U25436 (N_25436,N_22697,N_22869);
or U25437 (N_25437,N_23680,N_21261);
and U25438 (N_25438,N_23473,N_24608);
xnor U25439 (N_25439,N_20894,N_24095);
xnor U25440 (N_25440,N_21085,N_24609);
nor U25441 (N_25441,N_22495,N_21403);
and U25442 (N_25442,N_23262,N_22897);
or U25443 (N_25443,N_21141,N_22568);
or U25444 (N_25444,N_20379,N_20620);
xnor U25445 (N_25445,N_24429,N_20916);
xnor U25446 (N_25446,N_22774,N_22535);
nor U25447 (N_25447,N_24642,N_22275);
nor U25448 (N_25448,N_23195,N_23344);
nand U25449 (N_25449,N_23793,N_24250);
or U25450 (N_25450,N_22329,N_21118);
or U25451 (N_25451,N_23718,N_24455);
xor U25452 (N_25452,N_20110,N_20849);
nor U25453 (N_25453,N_22129,N_23399);
or U25454 (N_25454,N_21287,N_20881);
xor U25455 (N_25455,N_21592,N_23988);
nand U25456 (N_25456,N_24564,N_23539);
and U25457 (N_25457,N_21710,N_21657);
and U25458 (N_25458,N_23129,N_22556);
xor U25459 (N_25459,N_21510,N_23353);
or U25460 (N_25460,N_24992,N_22098);
or U25461 (N_25461,N_23198,N_22724);
and U25462 (N_25462,N_21912,N_20794);
or U25463 (N_25463,N_20969,N_24787);
xor U25464 (N_25464,N_23228,N_21761);
nand U25465 (N_25465,N_22747,N_24296);
and U25466 (N_25466,N_24266,N_22638);
nand U25467 (N_25467,N_20691,N_23170);
nand U25468 (N_25468,N_20018,N_21686);
and U25469 (N_25469,N_23064,N_22399);
nor U25470 (N_25470,N_20472,N_21220);
xnor U25471 (N_25471,N_22708,N_24950);
xnor U25472 (N_25472,N_22721,N_21310);
nand U25473 (N_25473,N_23472,N_23057);
or U25474 (N_25474,N_22104,N_20880);
nor U25475 (N_25475,N_22970,N_23537);
nand U25476 (N_25476,N_20217,N_23100);
nand U25477 (N_25477,N_24828,N_20831);
or U25478 (N_25478,N_20482,N_21120);
nor U25479 (N_25479,N_20158,N_23336);
xnor U25480 (N_25480,N_21195,N_21194);
xor U25481 (N_25481,N_21239,N_21938);
nor U25482 (N_25482,N_24767,N_24635);
nor U25483 (N_25483,N_22736,N_20674);
and U25484 (N_25484,N_20194,N_23974);
xor U25485 (N_25485,N_23737,N_24897);
and U25486 (N_25486,N_21914,N_22940);
nand U25487 (N_25487,N_21022,N_24107);
nand U25488 (N_25488,N_21596,N_21991);
nand U25489 (N_25489,N_23113,N_20507);
and U25490 (N_25490,N_20431,N_20525);
nand U25491 (N_25491,N_21026,N_23502);
nand U25492 (N_25492,N_22825,N_20770);
nand U25493 (N_25493,N_24996,N_24513);
and U25494 (N_25494,N_23271,N_21564);
and U25495 (N_25495,N_23992,N_21213);
and U25496 (N_25496,N_21309,N_21313);
nand U25497 (N_25497,N_22097,N_20689);
nand U25498 (N_25498,N_22518,N_24730);
nand U25499 (N_25499,N_20430,N_20145);
or U25500 (N_25500,N_20301,N_21709);
and U25501 (N_25501,N_20682,N_20375);
or U25502 (N_25502,N_23372,N_23585);
and U25503 (N_25503,N_20816,N_22759);
nand U25504 (N_25504,N_20022,N_21699);
xnor U25505 (N_25505,N_21936,N_23150);
nand U25506 (N_25506,N_22208,N_22713);
or U25507 (N_25507,N_20712,N_22880);
nand U25508 (N_25508,N_21948,N_24947);
or U25509 (N_25509,N_20281,N_24381);
and U25510 (N_25510,N_20526,N_20590);
or U25511 (N_25511,N_23890,N_24879);
nand U25512 (N_25512,N_21240,N_23589);
nand U25513 (N_25513,N_21303,N_22735);
nand U25514 (N_25514,N_21056,N_21332);
or U25515 (N_25515,N_20639,N_21754);
and U25516 (N_25516,N_21593,N_21522);
and U25517 (N_25517,N_22545,N_22538);
nor U25518 (N_25518,N_22878,N_22339);
xor U25519 (N_25519,N_21910,N_24733);
nand U25520 (N_25520,N_21660,N_23581);
nor U25521 (N_25521,N_22998,N_21869);
or U25522 (N_25522,N_21769,N_24330);
nor U25523 (N_25523,N_24451,N_23528);
and U25524 (N_25524,N_24017,N_22188);
nand U25525 (N_25525,N_20454,N_24280);
xor U25526 (N_25526,N_22726,N_22805);
nor U25527 (N_25527,N_21915,N_23620);
or U25528 (N_25528,N_20467,N_24309);
or U25529 (N_25529,N_22265,N_20010);
nand U25530 (N_25530,N_23221,N_22927);
and U25531 (N_25531,N_20941,N_20536);
nor U25532 (N_25532,N_20254,N_21380);
or U25533 (N_25533,N_20289,N_21427);
and U25534 (N_25534,N_23265,N_24082);
or U25535 (N_25535,N_23756,N_23564);
xor U25536 (N_25536,N_22376,N_21523);
nand U25537 (N_25537,N_21971,N_24956);
nand U25538 (N_25538,N_23011,N_21241);
or U25539 (N_25539,N_23872,N_21883);
nand U25540 (N_25540,N_22461,N_23526);
xnor U25541 (N_25541,N_21571,N_20933);
nand U25542 (N_25542,N_23157,N_23144);
nand U25543 (N_25543,N_23864,N_24236);
nand U25544 (N_25544,N_24928,N_24137);
xnor U25545 (N_25545,N_20389,N_20374);
xnor U25546 (N_25546,N_22566,N_23790);
or U25547 (N_25547,N_20517,N_21338);
or U25548 (N_25548,N_20443,N_23430);
xor U25549 (N_25549,N_20872,N_24624);
and U25550 (N_25550,N_21858,N_23060);
nor U25551 (N_25551,N_24641,N_24384);
and U25552 (N_25552,N_21330,N_24995);
nand U25553 (N_25553,N_21391,N_23203);
nand U25554 (N_25554,N_21092,N_20945);
and U25555 (N_25555,N_24556,N_23488);
nor U25556 (N_25556,N_21078,N_24001);
or U25557 (N_25557,N_21471,N_24378);
and U25558 (N_25558,N_24225,N_21148);
nand U25559 (N_25559,N_22925,N_20918);
nor U25560 (N_25560,N_20726,N_24799);
nor U25561 (N_25561,N_20838,N_22857);
nand U25562 (N_25562,N_24397,N_24587);
nand U25563 (N_25563,N_24030,N_20986);
or U25564 (N_25564,N_21779,N_23277);
nand U25565 (N_25565,N_22773,N_23684);
nand U25566 (N_25566,N_23310,N_20314);
and U25567 (N_25567,N_20554,N_21909);
nor U25568 (N_25568,N_22798,N_20684);
nand U25569 (N_25569,N_20692,N_22159);
nor U25570 (N_25570,N_23361,N_22107);
and U25571 (N_25571,N_21455,N_22242);
nand U25572 (N_25572,N_20504,N_21392);
xor U25573 (N_25573,N_23637,N_20477);
nand U25574 (N_25574,N_22358,N_24875);
and U25575 (N_25575,N_21830,N_23894);
nand U25576 (N_25576,N_21511,N_22449);
or U25577 (N_25577,N_20013,N_21301);
or U25578 (N_25578,N_22002,N_23339);
xnor U25579 (N_25579,N_22276,N_22230);
xor U25580 (N_25580,N_20706,N_22498);
and U25581 (N_25581,N_24042,N_21918);
and U25582 (N_25582,N_23766,N_22214);
nand U25583 (N_25583,N_23248,N_23058);
nor U25584 (N_25584,N_22255,N_23402);
or U25585 (N_25585,N_20131,N_24704);
nand U25586 (N_25586,N_23474,N_22750);
and U25587 (N_25587,N_22146,N_24734);
or U25588 (N_25588,N_22806,N_20398);
or U25589 (N_25589,N_23480,N_20603);
and U25590 (N_25590,N_23137,N_24316);
and U25591 (N_25591,N_22961,N_20973);
and U25592 (N_25592,N_20368,N_21572);
and U25593 (N_25593,N_21773,N_22256);
or U25594 (N_25594,N_23508,N_21713);
nor U25595 (N_25595,N_21210,N_20573);
xor U25596 (N_25596,N_21073,N_21876);
or U25597 (N_25597,N_20466,N_20074);
nand U25598 (N_25598,N_22245,N_23846);
nor U25599 (N_25599,N_21265,N_20181);
nand U25600 (N_25600,N_24018,N_20976);
nor U25601 (N_25601,N_22457,N_24638);
xnor U25602 (N_25602,N_24975,N_23541);
nor U25603 (N_25603,N_21358,N_21696);
nand U25604 (N_25604,N_24610,N_24116);
and U25605 (N_25605,N_20003,N_24958);
xnor U25606 (N_25606,N_21745,N_24782);
or U25607 (N_25607,N_20357,N_23967);
xnor U25608 (N_25608,N_24050,N_23321);
nand U25609 (N_25609,N_23835,N_21688);
nor U25610 (N_25610,N_24000,N_20832);
or U25611 (N_25611,N_24178,N_23495);
and U25612 (N_25612,N_21870,N_20210);
or U25613 (N_25613,N_21144,N_23807);
or U25614 (N_25614,N_22672,N_20954);
or U25615 (N_25615,N_22285,N_23828);
or U25616 (N_25616,N_23730,N_21335);
and U25617 (N_25617,N_23483,N_22848);
xor U25618 (N_25618,N_21156,N_20207);
nor U25619 (N_25619,N_24668,N_20347);
or U25620 (N_25620,N_24495,N_22199);
nand U25621 (N_25621,N_20174,N_24467);
nor U25622 (N_25622,N_22679,N_22466);
and U25623 (N_25623,N_22111,N_20830);
xor U25624 (N_25624,N_24919,N_21549);
and U25625 (N_25625,N_22994,N_22123);
and U25626 (N_25626,N_21737,N_24441);
nor U25627 (N_25627,N_23993,N_23796);
nor U25628 (N_25628,N_21311,N_22605);
or U25629 (N_25629,N_20967,N_21272);
and U25630 (N_25630,N_24092,N_22808);
nand U25631 (N_25631,N_21759,N_22049);
xnor U25632 (N_25632,N_21960,N_20034);
nor U25633 (N_25633,N_20394,N_24790);
xor U25634 (N_25634,N_22365,N_22475);
or U25635 (N_25635,N_23146,N_23212);
and U25636 (N_25636,N_20699,N_21370);
nor U25637 (N_25637,N_22234,N_24263);
or U25638 (N_25638,N_22309,N_23405);
nand U25639 (N_25639,N_20136,N_22206);
nor U25640 (N_25640,N_22785,N_23610);
xnor U25641 (N_25641,N_21259,N_20353);
or U25642 (N_25642,N_21051,N_22709);
and U25643 (N_25643,N_20211,N_24416);
nand U25644 (N_25644,N_20267,N_22056);
xnor U25645 (N_25645,N_20716,N_22938);
or U25646 (N_25646,N_24830,N_20305);
and U25647 (N_25647,N_22356,N_20867);
and U25648 (N_25648,N_22468,N_23887);
nand U25649 (N_25649,N_22957,N_23753);
nand U25650 (N_25650,N_23675,N_22448);
and U25651 (N_25651,N_20345,N_20814);
and U25652 (N_25652,N_22887,N_21314);
xnor U25653 (N_25653,N_23302,N_21415);
or U25654 (N_25654,N_22928,N_24366);
xor U25655 (N_25655,N_24628,N_23869);
nor U25656 (N_25656,N_22619,N_20313);
and U25657 (N_25657,N_21633,N_23636);
and U25658 (N_25658,N_20736,N_20862);
nor U25659 (N_25659,N_21285,N_20577);
xnor U25660 (N_25660,N_23329,N_23180);
and U25661 (N_25661,N_23487,N_21705);
or U25662 (N_25662,N_20542,N_21069);
xor U25663 (N_25663,N_22042,N_24091);
nor U25664 (N_25664,N_21306,N_22385);
or U25665 (N_25665,N_24090,N_22819);
nor U25666 (N_25666,N_20120,N_21297);
nand U25667 (N_25667,N_22020,N_23109);
and U25668 (N_25668,N_22976,N_21041);
or U25669 (N_25669,N_22217,N_20745);
or U25670 (N_25670,N_22626,N_23644);
or U25671 (N_25671,N_22832,N_20602);
and U25672 (N_25672,N_23352,N_23387);
nand U25673 (N_25673,N_21542,N_22364);
nor U25674 (N_25674,N_24098,N_24738);
xor U25675 (N_25675,N_23176,N_23759);
nor U25676 (N_25676,N_21656,N_24819);
nand U25677 (N_25677,N_21939,N_21887);
nor U25678 (N_25678,N_20659,N_24118);
xor U25679 (N_25679,N_24102,N_22220);
or U25680 (N_25680,N_21885,N_21817);
and U25681 (N_25681,N_21226,N_24592);
nor U25682 (N_25682,N_23422,N_23110);
or U25683 (N_25683,N_23457,N_23827);
nor U25684 (N_25684,N_24399,N_20318);
nor U25685 (N_25685,N_20943,N_22043);
nor U25686 (N_25686,N_24806,N_20168);
nor U25687 (N_25687,N_20575,N_21615);
nor U25688 (N_25688,N_24939,N_24824);
or U25689 (N_25689,N_20200,N_21559);
or U25690 (N_25690,N_24112,N_24155);
nand U25691 (N_25691,N_22951,N_24045);
or U25692 (N_25692,N_22771,N_21047);
nand U25693 (N_25693,N_23728,N_24413);
nand U25694 (N_25694,N_22067,N_21050);
and U25695 (N_25695,N_24032,N_21255);
nand U25696 (N_25696,N_23621,N_24978);
and U25697 (N_25697,N_23845,N_23207);
nand U25698 (N_25698,N_24521,N_23181);
and U25699 (N_25699,N_20902,N_21124);
nor U25700 (N_25700,N_24644,N_20533);
and U25701 (N_25701,N_20505,N_24967);
and U25702 (N_25702,N_24729,N_21898);
xnor U25703 (N_25703,N_23151,N_21394);
and U25704 (N_25704,N_23446,N_23019);
nand U25705 (N_25705,N_20817,N_21406);
or U25706 (N_25706,N_21652,N_23230);
and U25707 (N_25707,N_20821,N_22090);
nor U25708 (N_25708,N_24991,N_20989);
nand U25709 (N_25709,N_22250,N_22743);
and U25710 (N_25710,N_20607,N_22209);
nand U25711 (N_25711,N_24147,N_20747);
xor U25712 (N_25712,N_21955,N_20782);
xnor U25713 (N_25713,N_21231,N_23652);
xor U25714 (N_25714,N_20808,N_22702);
and U25715 (N_25715,N_20086,N_24674);
nor U25716 (N_25716,N_22792,N_24141);
nand U25717 (N_25717,N_22772,N_22218);
or U25718 (N_25718,N_21469,N_24540);
nor U25719 (N_25719,N_23513,N_20532);
and U25720 (N_25720,N_23752,N_23855);
nor U25721 (N_25721,N_22033,N_20983);
or U25722 (N_25722,N_24542,N_23511);
nor U25723 (N_25723,N_24578,N_21729);
and U25724 (N_25724,N_22787,N_20658);
xnor U25725 (N_25725,N_20764,N_24386);
and U25726 (N_25726,N_23921,N_22698);
nor U25727 (N_25727,N_23363,N_23356);
or U25728 (N_25728,N_24103,N_21037);
or U25729 (N_25729,N_23870,N_24013);
and U25730 (N_25730,N_21616,N_22586);
xor U25731 (N_25731,N_22577,N_23055);
nand U25732 (N_25732,N_23406,N_23319);
xor U25733 (N_25733,N_24008,N_22205);
nor U25734 (N_25734,N_22689,N_23569);
nor U25735 (N_25735,N_22133,N_23450);
xor U25736 (N_25736,N_24383,N_24951);
nand U25737 (N_25737,N_20069,N_20608);
and U25738 (N_25738,N_23808,N_24350);
or U25739 (N_25739,N_21519,N_23284);
nor U25740 (N_25740,N_21990,N_23428);
xor U25741 (N_25741,N_23593,N_22001);
or U25742 (N_25742,N_22764,N_22026);
xor U25743 (N_25743,N_24531,N_24331);
nand U25744 (N_25744,N_24518,N_22219);
nor U25745 (N_25745,N_22327,N_23619);
and U25746 (N_25746,N_22095,N_22073);
and U25747 (N_25747,N_21323,N_24322);
nor U25748 (N_25748,N_23280,N_20186);
xnor U25749 (N_25749,N_23546,N_20247);
nand U25750 (N_25750,N_20078,N_21734);
nand U25751 (N_25751,N_22048,N_23602);
nand U25752 (N_25752,N_22818,N_20265);
and U25753 (N_25753,N_24465,N_22838);
xnor U25754 (N_25754,N_21651,N_20866);
and U25755 (N_25755,N_23182,N_23713);
or U25756 (N_25756,N_20735,N_23475);
xnor U25757 (N_25757,N_20000,N_21300);
nand U25758 (N_25758,N_24229,N_24700);
nand U25759 (N_25759,N_22740,N_20641);
or U25760 (N_25760,N_21009,N_24483);
or U25761 (N_25761,N_21171,N_20793);
nor U25762 (N_25762,N_21780,N_24702);
and U25763 (N_25763,N_24798,N_24336);
and U25764 (N_25764,N_22281,N_23088);
nand U25765 (N_25765,N_20321,N_20686);
nand U25766 (N_25766,N_21075,N_23745);
or U25767 (N_25767,N_22652,N_24354);
xnor U25768 (N_25768,N_22846,N_20778);
nand U25769 (N_25769,N_20364,N_24217);
and U25770 (N_25770,N_24281,N_23097);
xor U25771 (N_25771,N_20440,N_21177);
nor U25772 (N_25772,N_22919,N_22704);
nand U25773 (N_25773,N_24590,N_22653);
and U25774 (N_25774,N_21655,N_23639);
nor U25775 (N_25775,N_21550,N_23140);
xnor U25776 (N_25776,N_22204,N_22473);
and U25777 (N_25777,N_22336,N_24152);
or U25778 (N_25778,N_23671,N_20059);
or U25779 (N_25779,N_21100,N_24677);
nand U25780 (N_25780,N_22029,N_21538);
or U25781 (N_25781,N_22074,N_23649);
nor U25782 (N_25782,N_22646,N_21956);
nand U25783 (N_25783,N_23640,N_22297);
xor U25784 (N_25784,N_20675,N_24932);
xnor U25785 (N_25785,N_21389,N_22851);
nor U25786 (N_25786,N_23798,N_24054);
nor U25787 (N_25787,N_20204,N_22714);
nor U25788 (N_25788,N_20640,N_23434);
or U25789 (N_25789,N_22070,N_20285);
xor U25790 (N_25790,N_23560,N_24815);
nand U25791 (N_25791,N_20130,N_21816);
or U25792 (N_25792,N_22354,N_21130);
nor U25793 (N_25793,N_21378,N_24524);
xnor U25794 (N_25794,N_20636,N_23238);
and U25795 (N_25795,N_24901,N_21351);
xnor U25796 (N_25796,N_23895,N_21768);
nand U25797 (N_25797,N_21501,N_24698);
and U25798 (N_25798,N_24805,N_24883);
xnor U25799 (N_25799,N_22563,N_22307);
nor U25800 (N_25800,N_20576,N_24933);
nor U25801 (N_25801,N_23519,N_23655);
or U25802 (N_25802,N_21223,N_24252);
nand U25803 (N_25803,N_21736,N_23455);
nor U25804 (N_25804,N_23851,N_22332);
and U25805 (N_25805,N_23952,N_23580);
nand U25806 (N_25806,N_20534,N_24245);
xnor U25807 (N_25807,N_22233,N_23252);
nor U25808 (N_25808,N_21715,N_21859);
nor U25809 (N_25809,N_22554,N_21430);
and U25810 (N_25810,N_24941,N_23091);
or U25811 (N_25811,N_23968,N_21361);
nor U25812 (N_25812,N_23831,N_23241);
and U25813 (N_25813,N_20561,N_21106);
nand U25814 (N_25814,N_22306,N_24621);
and U25815 (N_25815,N_24368,N_20953);
or U25816 (N_25816,N_24345,N_21476);
nand U25817 (N_25817,N_24555,N_20391);
and U25818 (N_25818,N_20198,N_20176);
nor U25819 (N_25819,N_21543,N_21601);
xnor U25820 (N_25820,N_22122,N_21173);
nor U25821 (N_25821,N_22513,N_20627);
or U25822 (N_25822,N_23710,N_23735);
nor U25823 (N_25823,N_22185,N_20610);
or U25824 (N_25824,N_22174,N_20543);
or U25825 (N_25825,N_21483,N_24827);
or U25826 (N_25826,N_20768,N_21107);
xor U25827 (N_25827,N_21151,N_22540);
and U25828 (N_25828,N_21861,N_23168);
nand U25829 (N_25829,N_20584,N_24496);
xor U25830 (N_25830,N_23048,N_23747);
nand U25831 (N_25831,N_22189,N_22236);
nor U25832 (N_25832,N_24138,N_22173);
nor U25833 (N_25833,N_23858,N_20295);
nand U25834 (N_25834,N_21639,N_20926);
nor U25835 (N_25835,N_22062,N_21679);
xor U25836 (N_25836,N_23179,N_20857);
or U25837 (N_25837,N_21603,N_22369);
and U25838 (N_25838,N_21632,N_22161);
xor U25839 (N_25839,N_23545,N_23108);
nor U25840 (N_25840,N_22213,N_23950);
or U25841 (N_25841,N_23467,N_24291);
or U25842 (N_25842,N_23153,N_21536);
nor U25843 (N_25843,N_21533,N_24104);
nor U25844 (N_25844,N_22483,N_20212);
and U25845 (N_25845,N_20141,N_22393);
nor U25846 (N_25846,N_22407,N_21963);
xor U25847 (N_25847,N_20773,N_22969);
or U25848 (N_25848,N_20968,N_20307);
or U25849 (N_25849,N_22064,N_21622);
xnor U25850 (N_25850,N_24153,N_22720);
nor U25851 (N_25851,N_23647,N_24984);
and U25852 (N_25852,N_22153,N_24835);
and U25853 (N_25853,N_20805,N_21524);
and U25854 (N_25854,N_22400,N_24474);
nor U25855 (N_25855,N_22178,N_20417);
or U25856 (N_25856,N_20878,N_20282);
or U25857 (N_25857,N_22334,N_23925);
nand U25858 (N_25858,N_24253,N_23787);
xnor U25859 (N_25859,N_21619,N_21329);
nand U25860 (N_25860,N_23267,N_22660);
xnor U25861 (N_25861,N_24742,N_21468);
and U25862 (N_25862,N_21874,N_24667);
nand U25863 (N_25863,N_21900,N_23712);
nor U25864 (N_25864,N_24887,N_22057);
or U25865 (N_25865,N_24074,N_22530);
nor U25866 (N_25866,N_22482,N_24616);
nor U25867 (N_25867,N_20518,N_22659);
nor U25868 (N_25868,N_24127,N_24896);
nor U25869 (N_25869,N_21094,N_23232);
nor U25870 (N_25870,N_24706,N_21513);
nor U25871 (N_25871,N_21324,N_23847);
or U25872 (N_25872,N_23881,N_21600);
and U25873 (N_25873,N_24846,N_24488);
and U25874 (N_25874,N_24954,N_23236);
xnor U25875 (N_25875,N_21112,N_21701);
xnor U25876 (N_25876,N_23780,N_23063);
xnor U25877 (N_25877,N_23883,N_21880);
nor U25878 (N_25878,N_23122,N_24994);
nor U25879 (N_25879,N_24696,N_22282);
and U25880 (N_25880,N_20092,N_22582);
or U25881 (N_25881,N_22685,N_22303);
xnor U25882 (N_25882,N_22931,N_22386);
nand U25883 (N_25883,N_23989,N_24347);
and U25884 (N_25884,N_23863,N_24223);
xor U25885 (N_25885,N_20581,N_22040);
nand U25886 (N_25886,N_23130,N_24307);
nand U25887 (N_25887,N_23003,N_22439);
xor U25888 (N_25888,N_21585,N_23761);
or U25889 (N_25889,N_21196,N_21450);
and U25890 (N_25890,N_24403,N_20259);
and U25891 (N_25891,N_24997,N_22305);
xor U25892 (N_25892,N_20239,N_21103);
xor U25893 (N_25893,N_22288,N_21640);
or U25894 (N_25894,N_23068,N_21237);
xnor U25895 (N_25895,N_24420,N_22532);
or U25896 (N_25896,N_23527,N_23837);
or U25897 (N_25897,N_23588,N_24235);
nor U25898 (N_25898,N_24333,N_23346);
nor U25899 (N_25899,N_21068,N_20644);
or U25900 (N_25900,N_20435,N_24425);
nor U25901 (N_25901,N_23812,N_24633);
nor U25902 (N_25902,N_24816,N_20947);
nand U25903 (N_25903,N_23553,N_22525);
nor U25904 (N_25904,N_22030,N_20359);
nand U25905 (N_25905,N_20628,N_23378);
xor U25906 (N_25906,N_20184,N_21234);
or U25907 (N_25907,N_20114,N_23282);
xor U25908 (N_25908,N_21014,N_24158);
or U25909 (N_25909,N_20656,N_20828);
nand U25910 (N_25910,N_22569,N_22999);
or U25911 (N_25911,N_23490,N_20936);
and U25912 (N_25912,N_23746,N_22118);
nor U25913 (N_25913,N_22441,N_20511);
or U25914 (N_25914,N_20719,N_20646);
and U25915 (N_25915,N_24431,N_21539);
nor U25916 (N_25916,N_20702,N_24579);
and U25917 (N_25917,N_24003,N_24334);
nand U25918 (N_25918,N_20344,N_21445);
xnor U25919 (N_25919,N_24763,N_24755);
or U25920 (N_25920,N_22960,N_20492);
nand U25921 (N_25921,N_21553,N_21172);
xor U25922 (N_25922,N_23552,N_21350);
and U25923 (N_25923,N_24963,N_24968);
nand U25924 (N_25924,N_21674,N_23053);
nor U25925 (N_25925,N_21814,N_23478);
or U25926 (N_25926,N_22962,N_22267);
nand U25927 (N_25927,N_24914,N_24097);
nor U25928 (N_25928,N_22515,N_24597);
and U25929 (N_25929,N_24209,N_23497);
xnor U25930 (N_25930,N_24769,N_23204);
nand U25931 (N_25931,N_24684,N_21820);
or U25932 (N_25932,N_24766,N_23682);
and U25933 (N_25933,N_21478,N_21851);
nand U25934 (N_25934,N_24789,N_20071);
nor U25935 (N_25935,N_20491,N_22078);
xor U25936 (N_25936,N_23681,N_24522);
nor U25937 (N_25937,N_24016,N_24142);
or U25938 (N_25938,N_23806,N_21807);
xnor U25939 (N_25939,N_20367,N_22427);
or U25940 (N_25940,N_21257,N_22259);
xnor U25941 (N_25941,N_23222,N_21363);
xnor U25942 (N_25942,N_23932,N_21061);
nor U25943 (N_25943,N_22058,N_24364);
xor U25944 (N_25944,N_24663,N_20677);
nand U25945 (N_25945,N_24129,N_24389);
and U25946 (N_25946,N_24300,N_20931);
and U25947 (N_25947,N_20932,N_22112);
and U25948 (N_25948,N_21294,N_23685);
nor U25949 (N_25949,N_20405,N_24156);
nor U25950 (N_25950,N_21276,N_20538);
or U25951 (N_25951,N_22366,N_23479);
xnor U25952 (N_25952,N_24983,N_24115);
nor U25953 (N_25953,N_21547,N_24574);
or U25954 (N_25954,N_20452,N_24754);
nor U25955 (N_25955,N_22936,N_21647);
nor U25956 (N_25956,N_23940,N_24206);
nor U25957 (N_25957,N_23768,N_22934);
nand U25958 (N_25958,N_20792,N_22280);
nor U25959 (N_25959,N_21965,N_23465);
or U25960 (N_25960,N_20991,N_24528);
nor U25961 (N_25961,N_23772,N_22845);
and U25962 (N_25962,N_23722,N_21251);
nand U25963 (N_25963,N_20426,N_22745);
nor U25964 (N_25964,N_21146,N_22587);
nand U25965 (N_25965,N_23187,N_22401);
nand U25966 (N_25966,N_21781,N_22826);
nor U25967 (N_25967,N_24033,N_20695);
nand U25968 (N_25968,N_21669,N_20833);
and U25969 (N_25969,N_22763,N_21182);
or U25970 (N_25970,N_24779,N_21446);
nand U25971 (N_25971,N_22738,N_22420);
xor U25972 (N_25972,N_21033,N_20229);
nand U25973 (N_25973,N_20605,N_20528);
xor U25974 (N_25974,N_22695,N_24514);
nor U25975 (N_25975,N_21030,N_24286);
or U25976 (N_25976,N_22370,N_21904);
nand U25977 (N_25977,N_24643,N_21853);
and U25978 (N_25978,N_22050,N_21292);
or U25979 (N_25979,N_24881,N_20756);
and U25980 (N_25980,N_21521,N_22912);
and U25981 (N_25981,N_22717,N_23565);
nor U25982 (N_25982,N_24076,N_21166);
xor U25983 (N_25983,N_23013,N_20807);
and U25984 (N_25984,N_20540,N_24989);
or U25985 (N_25985,N_20979,N_23522);
or U25986 (N_25986,N_23316,N_23471);
and U25987 (N_25987,N_22347,N_20252);
and U25988 (N_25988,N_23566,N_21032);
nand U25989 (N_25989,N_24964,N_20335);
nor U25990 (N_25990,N_20037,N_23124);
nand U25991 (N_25991,N_22109,N_22854);
nor U25992 (N_25992,N_22180,N_24259);
and U25993 (N_25993,N_24227,N_24070);
nand U25994 (N_25994,N_23853,N_21157);
or U25995 (N_25995,N_22235,N_20806);
nor U25996 (N_25996,N_22948,N_20755);
or U25997 (N_25997,N_20354,N_24577);
xnor U25998 (N_25998,N_20809,N_22802);
nor U25999 (N_25999,N_23231,N_20222);
xor U26000 (N_26000,N_22082,N_24462);
nor U26001 (N_26001,N_24187,N_21207);
or U26002 (N_26002,N_20387,N_22183);
nor U26003 (N_26003,N_23111,N_20648);
nand U26004 (N_26004,N_22890,N_20622);
or U26005 (N_26005,N_21767,N_22723);
nor U26006 (N_26006,N_24231,N_23957);
nand U26007 (N_26007,N_23622,N_22655);
and U26008 (N_26008,N_20133,N_20462);
or U26009 (N_26009,N_23934,N_20552);
and U26010 (N_26010,N_22419,N_24520);
or U26011 (N_26011,N_21500,N_22666);
or U26012 (N_26012,N_22436,N_20005);
xor U26013 (N_26013,N_23817,N_24325);
nor U26014 (N_26014,N_22645,N_22694);
nor U26015 (N_26015,N_22664,N_23507);
or U26016 (N_26016,N_21340,N_21331);
xnor U26017 (N_26017,N_21505,N_21941);
nand U26018 (N_26018,N_21793,N_22179);
nand U26019 (N_26019,N_22611,N_22680);
nor U26020 (N_26020,N_22733,N_21002);
xnor U26021 (N_26021,N_22589,N_20153);
nor U26022 (N_26022,N_20170,N_24840);
nand U26023 (N_26023,N_23947,N_20293);
xnor U26024 (N_26024,N_24471,N_23370);
nor U26025 (N_26025,N_21992,N_23983);
xnor U26026 (N_26026,N_22231,N_21479);
or U26027 (N_26027,N_22777,N_21178);
and U26028 (N_26028,N_21362,N_24602);
and U26029 (N_26029,N_20751,N_24867);
xor U26030 (N_26030,N_20713,N_22175);
nor U26031 (N_26031,N_24672,N_22422);
xor U26032 (N_26032,N_24024,N_23648);
nand U26033 (N_26033,N_23444,N_24547);
or U26034 (N_26034,N_20068,N_23654);
and U26035 (N_26035,N_24511,N_23504);
xnor U26036 (N_26036,N_22681,N_20061);
nor U26037 (N_26037,N_21235,N_22828);
nand U26038 (N_26038,N_24534,N_23089);
or U26039 (N_26039,N_22989,N_20775);
and U26040 (N_26040,N_22670,N_21886);
and U26041 (N_26041,N_21833,N_23083);
and U26042 (N_26042,N_21720,N_24725);
or U26043 (N_26043,N_21268,N_23171);
xor U26044 (N_26044,N_20080,N_23158);
xor U26045 (N_26045,N_20336,N_22340);
xnor U26046 (N_26046,N_20922,N_21753);
or U26047 (N_26047,N_21215,N_23717);
nor U26048 (N_26048,N_24899,N_22795);
xor U26049 (N_26049,N_20586,N_24459);
and U26050 (N_26050,N_20132,N_21045);
nor U26051 (N_26051,N_23813,N_22463);
and U26052 (N_26052,N_24796,N_23635);
xor U26053 (N_26053,N_24803,N_24620);
xnor U26054 (N_26054,N_22360,N_23861);
or U26055 (N_26055,N_22338,N_23789);
and U26056 (N_26056,N_20972,N_22924);
xnor U26057 (N_26057,N_24558,N_23505);
or U26058 (N_26058,N_22493,N_20616);
or U26059 (N_26059,N_24948,N_20913);
and U26060 (N_26060,N_24093,N_20685);
nor U26061 (N_26061,N_21881,N_23799);
and U26062 (N_26062,N_23364,N_21933);
and U26063 (N_26063,N_20601,N_21353);
or U26064 (N_26064,N_23672,N_21648);
and U26065 (N_26065,N_24172,N_20062);
nand U26066 (N_26066,N_24837,N_23571);
and U26067 (N_26067,N_22617,N_24802);
or U26068 (N_26068,N_24353,N_21438);
nor U26069 (N_26069,N_21662,N_21922);
xor U26070 (N_26070,N_24360,N_24053);
or U26071 (N_26071,N_21290,N_20580);
and U26072 (N_26072,N_21049,N_21762);
nor U26073 (N_26073,N_24393,N_24843);
nor U26074 (N_26074,N_22371,N_20626);
nor U26075 (N_26075,N_22907,N_20493);
and U26076 (N_26076,N_24043,N_21179);
xor U26077 (N_26077,N_20718,N_23210);
or U26078 (N_26078,N_24569,N_24131);
nor U26079 (N_26079,N_21947,N_23139);
and U26080 (N_26080,N_22531,N_22149);
and U26081 (N_26081,N_22317,N_24671);
nor U26082 (N_26082,N_22575,N_24044);
xnor U26083 (N_26083,N_23002,N_20306);
nand U26084 (N_26084,N_24629,N_20785);
and U26085 (N_26085,N_20288,N_22156);
nand U26086 (N_26086,N_20942,N_21490);
and U26087 (N_26087,N_21724,N_24746);
nor U26088 (N_26088,N_23317,N_24405);
or U26089 (N_26089,N_23556,N_24771);
xor U26090 (N_26090,N_21186,N_23081);
and U26091 (N_26091,N_21969,N_20964);
xnor U26092 (N_26092,N_22434,N_20144);
nor U26093 (N_26093,N_23114,N_23763);
or U26094 (N_26094,N_22612,N_20935);
xnor U26095 (N_26095,N_24505,N_22859);
nand U26096 (N_26096,N_23309,N_20788);
xnor U26097 (N_26097,N_24148,N_24713);
and U26098 (N_26098,N_20091,N_21620);
and U26099 (N_26099,N_20595,N_22641);
nor U26100 (N_26100,N_23645,N_23598);
or U26101 (N_26101,N_21187,N_23774);
or U26102 (N_26102,N_22181,N_21631);
nor U26103 (N_26103,N_20152,N_24352);
xor U26104 (N_26104,N_23116,N_23517);
nand U26105 (N_26105,N_23320,N_22858);
nand U26106 (N_26106,N_23673,N_21102);
or U26107 (N_26107,N_24196,N_21221);
xor U26108 (N_26108,N_22421,N_21852);
nor U26109 (N_26109,N_20565,N_23998);
and U26110 (N_26110,N_21386,N_21424);
or U26111 (N_26111,N_23899,N_20142);
or U26112 (N_26112,N_22063,N_21957);
xnor U26113 (N_26113,N_20654,N_24500);
or U26114 (N_26114,N_24492,N_20052);
nor U26115 (N_26115,N_23366,N_20496);
or U26116 (N_26116,N_21798,N_21072);
and U26117 (N_26117,N_21692,N_23715);
nand U26118 (N_26118,N_24631,N_24962);
nand U26119 (N_26119,N_20839,N_21275);
nor U26120 (N_26120,N_22278,N_22138);
or U26121 (N_26121,N_24719,N_24707);
or U26122 (N_26122,N_23033,N_22849);
or U26123 (N_26123,N_21735,N_20117);
xor U26124 (N_26124,N_23943,N_22416);
nor U26125 (N_26125,N_23442,N_22381);
nand U26126 (N_26126,N_22974,N_20524);
and U26127 (N_26127,N_24676,N_23407);
nand U26128 (N_26128,N_24369,N_24998);
and U26129 (N_26129,N_20629,N_23920);
nand U26130 (N_26130,N_24669,N_21364);
xnor U26131 (N_26131,N_23126,N_24080);
nand U26132 (N_26132,N_20637,N_23397);
or U26133 (N_26133,N_24611,N_20088);
nand U26134 (N_26134,N_21308,N_21096);
and U26135 (N_26135,N_20081,N_24915);
nor U26136 (N_26136,N_22768,N_24351);
nor U26137 (N_26137,N_24181,N_24373);
or U26138 (N_26138,N_20138,N_23191);
nor U26139 (N_26139,N_22384,N_23985);
and U26140 (N_26140,N_22479,N_22905);
nand U26141 (N_26141,N_23930,N_23958);
xor U26142 (N_26142,N_21926,N_20036);
or U26143 (N_26143,N_24909,N_21018);
or U26144 (N_26144,N_21723,N_21518);
xor U26145 (N_26145,N_23263,N_21273);
nand U26146 (N_26146,N_21402,N_24890);
and U26147 (N_26147,N_21153,N_23627);
nor U26148 (N_26148,N_24662,N_22410);
nor U26149 (N_26149,N_23547,N_22302);
nand U26150 (N_26150,N_23842,N_21945);
or U26151 (N_26151,N_23823,N_23871);
or U26152 (N_26152,N_23286,N_24411);
or U26153 (N_26153,N_24687,N_20634);
nor U26154 (N_26154,N_20271,N_24468);
or U26155 (N_26155,N_22454,N_22377);
xnor U26156 (N_26156,N_24189,N_23976);
and U26157 (N_26157,N_20415,N_24367);
nand U26158 (N_26158,N_21448,N_23699);
nand U26159 (N_26159,N_20774,N_24338);
xnor U26160 (N_26160,N_22867,N_23340);
nor U26161 (N_26161,N_22790,N_22154);
and U26162 (N_26162,N_22471,N_20047);
or U26163 (N_26163,N_20652,N_23638);
and U26164 (N_26164,N_20510,N_21375);
nor U26165 (N_26165,N_20164,N_22987);
or U26166 (N_26166,N_22841,N_21274);
or U26167 (N_26167,N_24133,N_22068);
or U26168 (N_26168,N_24601,N_20330);
xnor U26169 (N_26169,N_21289,N_23612);
and U26170 (N_26170,N_21325,N_24566);
and U26171 (N_26171,N_22207,N_22260);
or U26172 (N_26172,N_23966,N_22367);
xor U26173 (N_26173,N_22521,N_21650);
xnor U26174 (N_26174,N_24482,N_20811);
nand U26175 (N_26175,N_20363,N_20847);
and U26176 (N_26176,N_24646,N_20598);
nand U26177 (N_26177,N_20101,N_23041);
and U26178 (N_26178,N_23288,N_24885);
nand U26179 (N_26179,N_23334,N_21029);
and U26180 (N_26180,N_24826,N_21877);
xor U26181 (N_26181,N_21627,N_21411);
and U26182 (N_26182,N_21458,N_24015);
or U26183 (N_26183,N_23901,N_23325);
or U26184 (N_26184,N_20669,N_23607);
and U26185 (N_26185,N_20582,N_22911);
nor U26186 (N_26186,N_24073,N_22766);
and U26187 (N_26187,N_20907,N_24606);
nor U26188 (N_26188,N_21354,N_24660);
and U26189 (N_26189,N_21579,N_21569);
nor U26190 (N_26190,N_22490,N_20214);
nor U26191 (N_26191,N_24201,N_21164);
nand U26192 (N_26192,N_20531,N_24078);
and U26193 (N_26193,N_20882,N_23029);
nand U26194 (N_26194,N_22548,N_24910);
xnor U26195 (N_26195,N_22474,N_22990);
and U26196 (N_26196,N_21663,N_24953);
or U26197 (N_26197,N_21968,N_21843);
xor U26198 (N_26198,N_24174,N_21271);
xnor U26199 (N_26199,N_21895,N_23624);
nor U26200 (N_26200,N_22458,N_20134);
and U26201 (N_26201,N_23447,N_20842);
xor U26202 (N_26202,N_21695,N_23658);
nand U26203 (N_26203,N_22438,N_23412);
nor U26204 (N_26204,N_21063,N_22923);
nor U26205 (N_26205,N_24959,N_22570);
nand U26206 (N_26206,N_24079,N_23670);
and U26207 (N_26207,N_20861,N_23184);
nor U26208 (N_26208,N_21341,N_20273);
and U26209 (N_26209,N_22864,N_22683);
or U26210 (N_26210,N_23464,N_22480);
and U26211 (N_26211,N_23650,N_21981);
or U26212 (N_26212,N_20899,N_20975);
nand U26213 (N_26213,N_23778,N_20250);
nor U26214 (N_26214,N_21034,N_21185);
and U26215 (N_26215,N_23955,N_20843);
nand U26216 (N_26216,N_20328,N_22749);
nand U26217 (N_26217,N_22596,N_20672);
xor U26218 (N_26218,N_23136,N_21426);
nand U26219 (N_26219,N_23605,N_22533);
nand U26220 (N_26220,N_24753,N_24113);
nand U26221 (N_26221,N_20209,N_20812);
xor U26222 (N_26222,N_21989,N_23491);
nand U26223 (N_26223,N_20395,N_20315);
nand U26224 (N_26224,N_21983,N_23278);
xor U26225 (N_26225,N_20868,N_20045);
and U26226 (N_26226,N_24006,N_23575);
xor U26227 (N_26227,N_23466,N_24305);
nor U26228 (N_26228,N_21689,N_22914);
nor U26229 (N_26229,N_20082,N_23323);
and U26230 (N_26230,N_20098,N_23015);
and U26231 (N_26231,N_21381,N_23896);
or U26232 (N_26232,N_20287,N_23072);
and U26233 (N_26233,N_23452,N_23143);
nand U26234 (N_26234,N_24198,N_21799);
and U26235 (N_26235,N_21320,N_24058);
and U26236 (N_26236,N_20249,N_20617);
xnor U26237 (N_26237,N_23331,N_20694);
nand U26238 (N_26238,N_24348,N_24472);
nand U26239 (N_26239,N_23574,N_22391);
or U26240 (N_26240,N_22850,N_22955);
and U26241 (N_26241,N_23938,N_24712);
nand U26242 (N_26242,N_21344,N_24344);
nor U26243 (N_26243,N_20104,N_23970);
or U26244 (N_26244,N_21263,N_23811);
or U26245 (N_26245,N_21979,N_24406);
xor U26246 (N_26246,N_24589,N_22537);
xnor U26247 (N_26247,N_21610,N_24499);
xnor U26248 (N_26248,N_21043,N_24294);
nor U26249 (N_26249,N_20850,N_24243);
nand U26250 (N_26250,N_23414,N_21150);
or U26251 (N_26251,N_24813,N_23614);
and U26252 (N_26252,N_22973,N_21826);
nor U26253 (N_26253,N_20017,N_24168);
nor U26254 (N_26254,N_23390,N_22357);
nor U26255 (N_26255,N_20701,N_21819);
xor U26256 (N_26256,N_21126,N_20925);
nand U26257 (N_26257,N_20244,N_24952);
nand U26258 (N_26258,N_20373,N_22202);
nor U26259 (N_26259,N_21661,N_21693);
or U26260 (N_26260,N_22876,N_21191);
nor U26261 (N_26261,N_23568,N_22440);
xnor U26262 (N_26262,N_24056,N_22609);
or U26263 (N_26263,N_23810,N_24326);
nand U26264 (N_26264,N_23944,N_22700);
nor U26265 (N_26265,N_20384,N_21973);
nand U26266 (N_26266,N_21443,N_20449);
or U26267 (N_26267,N_20460,N_23708);
nand U26268 (N_26268,N_24750,N_24265);
or U26269 (N_26269,N_21071,N_23716);
or U26270 (N_26270,N_24949,N_22866);
nand U26271 (N_26271,N_24448,N_23242);
nand U26272 (N_26272,N_21813,N_22254);
nand U26273 (N_26273,N_21048,N_23185);
nor U26274 (N_26274,N_20420,N_22895);
and U26275 (N_26275,N_22464,N_21342);
and U26276 (N_26276,N_24599,N_22716);
xnor U26277 (N_26277,N_23246,N_21934);
nor U26278 (N_26278,N_23829,N_21742);
xnor U26279 (N_26279,N_20390,N_20660);
or U26280 (N_26280,N_20066,N_21192);
nor U26281 (N_26281,N_23919,N_21746);
nor U26282 (N_26282,N_22137,N_23094);
xor U26283 (N_26283,N_20804,N_20073);
or U26284 (N_26284,N_23500,N_22823);
or U26285 (N_26285,N_21090,N_24856);
or U26286 (N_26286,N_22089,N_20741);
nand U26287 (N_26287,N_22404,N_21621);
xor U26288 (N_26288,N_21025,N_24613);
nor U26289 (N_26289,N_20437,N_23731);
and U26290 (N_26290,N_23689,N_24709);
nor U26291 (N_26291,N_20920,N_22748);
nor U26292 (N_26292,N_23727,N_24445);
nor U26293 (N_26293,N_24697,N_22836);
nor U26294 (N_26294,N_23857,N_22238);
or U26295 (N_26295,N_23255,N_20961);
and U26296 (N_26296,N_21227,N_21667);
nand U26297 (N_26297,N_20724,N_22782);
or U26298 (N_26298,N_21517,N_21552);
nand U26299 (N_26299,N_21256,N_20490);
nand U26300 (N_26300,N_24363,N_20578);
or U26301 (N_26301,N_21125,N_20759);
or U26302 (N_26302,N_24804,N_22066);
xnor U26303 (N_26303,N_21834,N_20343);
and U26304 (N_26304,N_24356,N_20530);
nand U26305 (N_26305,N_24293,N_23964);
xnor U26306 (N_26306,N_23720,N_24339);
nand U26307 (N_26307,N_24288,N_22978);
nand U26308 (N_26308,N_21664,N_20455);
nor U26309 (N_26309,N_24491,N_20562);
nor U26310 (N_26310,N_23037,N_20055);
nand U26311 (N_26311,N_20860,N_21577);
nor U26312 (N_26312,N_22092,N_20463);
and U26313 (N_26313,N_23028,N_23367);
nand U26314 (N_26314,N_24986,N_24186);
nand U26315 (N_26315,N_20203,N_22232);
or U26316 (N_26316,N_24068,N_22616);
and U26317 (N_26317,N_23977,N_20921);
nand U26318 (N_26318,N_24422,N_24903);
nor U26319 (N_26319,N_21238,N_23779);
xnor U26320 (N_26320,N_21818,N_22620);
nand U26321 (N_26321,N_20107,N_22873);
nand U26322 (N_26322,N_20834,N_21919);
and U26323 (N_26323,N_20480,N_21225);
or U26324 (N_26324,N_22351,N_22901);
and U26325 (N_26325,N_23167,N_23873);
xnor U26326 (N_26326,N_24688,N_20255);
nor U26327 (N_26327,N_24844,N_24027);
and U26328 (N_26328,N_23449,N_22469);
nand U26329 (N_26329,N_22447,N_24210);
nor U26330 (N_26330,N_21645,N_20196);
xor U26331 (N_26331,N_22579,N_21557);
nor U26332 (N_26332,N_23485,N_24969);
and U26333 (N_26333,N_20951,N_21184);
nand U26334 (N_26334,N_22283,N_23850);
and U26335 (N_26335,N_20332,N_23418);
xor U26336 (N_26336,N_21529,N_23243);
and U26337 (N_26337,N_20784,N_21137);
xor U26338 (N_26338,N_24041,N_24848);
or U26339 (N_26339,N_24002,N_22741);
nand U26340 (N_26340,N_23740,N_20160);
and U26341 (N_26341,N_24694,N_22879);
nor U26342 (N_26342,N_21822,N_24934);
nor U26343 (N_26343,N_23618,N_24841);
or U26344 (N_26344,N_20201,N_23532);
nor U26345 (N_26345,N_21749,N_23192);
xor U26346 (N_26346,N_24313,N_20275);
and U26347 (N_26347,N_20270,N_23905);
nand U26348 (N_26348,N_23578,N_21433);
nand U26349 (N_26349,N_23213,N_20007);
nand U26350 (N_26350,N_20392,N_20777);
xnor U26351 (N_26351,N_23082,N_24751);
nand U26352 (N_26352,N_20569,N_22744);
nand U26353 (N_26353,N_22059,N_24111);
xnor U26354 (N_26354,N_22286,N_23911);
or U26355 (N_26355,N_24715,N_24987);
nor U26356 (N_26356,N_24838,N_20372);
nand U26357 (N_26357,N_23383,N_23330);
nor U26358 (N_26358,N_22804,N_20396);
xor U26359 (N_26359,N_24931,N_21316);
and U26360 (N_26360,N_23767,N_20795);
xnor U26361 (N_26361,N_24026,N_22158);
nand U26362 (N_26362,N_23038,N_21797);
and U26363 (N_26363,N_20429,N_22893);
xor U26364 (N_26364,N_24797,N_24463);
and U26365 (N_26365,N_21888,N_23909);
nor U26366 (N_26366,N_24487,N_23634);
or U26367 (N_26367,N_24651,N_20070);
nor U26368 (N_26368,N_22953,N_24974);
and U26369 (N_26369,N_22674,N_23771);
and U26370 (N_26370,N_24485,N_24605);
nand U26371 (N_26371,N_24035,N_22355);
or U26372 (N_26372,N_23426,N_22476);
xor U26373 (N_26373,N_22997,N_22197);
nor U26374 (N_26374,N_22840,N_20593);
xor U26375 (N_26375,N_22018,N_24536);
nor U26376 (N_26376,N_23279,N_20419);
xnor U26377 (N_26377,N_24327,N_22352);
and U26378 (N_26378,N_21604,N_20663);
and U26379 (N_26379,N_22451,N_22045);
xor U26380 (N_26380,N_22258,N_22277);
xor U26381 (N_26381,N_22196,N_20416);
nor U26382 (N_26382,N_24716,N_23567);
nand U26383 (N_26383,N_22550,N_23524);
and U26384 (N_26384,N_22144,N_23090);
xnor U26385 (N_26385,N_23849,N_22187);
or U26386 (N_26386,N_22829,N_24565);
xor U26387 (N_26387,N_23935,N_21181);
nand U26388 (N_26388,N_23086,N_23726);
or U26389 (N_26389,N_22894,N_24567);
nand U26390 (N_26390,N_21857,N_21980);
and U26391 (N_26391,N_21222,N_23928);
nor U26392 (N_26392,N_22226,N_20923);
nand U26393 (N_26393,N_21064,N_20781);
xnor U26394 (N_26394,N_22929,N_21419);
or U26395 (N_26395,N_22330,N_23355);
or U26396 (N_26396,N_22014,N_20115);
nand U26397 (N_26397,N_23036,N_22628);
and U26398 (N_26398,N_20688,N_20428);
or U26399 (N_26399,N_22016,N_21154);
nor U26400 (N_26400,N_21675,N_24072);
or U26401 (N_26401,N_22293,N_21447);
and U26402 (N_26402,N_24377,N_21691);
or U26403 (N_26403,N_20422,N_24498);
and U26404 (N_26404,N_21844,N_23351);
nor U26405 (N_26405,N_21174,N_21790);
and U26406 (N_26406,N_24088,N_22411);
or U26407 (N_26407,N_20874,N_22203);
or U26408 (N_26408,N_20631,N_22909);
or U26409 (N_26409,N_23225,N_22634);
and U26410 (N_26410,N_20471,N_22348);
nand U26411 (N_26411,N_20643,N_24501);
nand U26412 (N_26412,N_22517,N_24337);
and U26413 (N_26413,N_21784,N_23049);
or U26414 (N_26414,N_22135,N_20566);
nand U26415 (N_26415,N_22294,N_22247);
nand U26416 (N_26416,N_22651,N_20351);
xor U26417 (N_26417,N_23824,N_21413);
xor U26418 (N_26418,N_22676,N_20161);
nand U26419 (N_26419,N_24430,N_23440);
xor U26420 (N_26420,N_20754,N_23535);
and U26421 (N_26421,N_24457,N_24864);
nor U26422 (N_26422,N_23481,N_21168);
nor U26423 (N_26423,N_21404,N_24904);
nand U26424 (N_26424,N_24060,N_24193);
and U26425 (N_26425,N_22047,N_22722);
nand U26426 (N_26426,N_22289,N_23609);
and U26427 (N_26427,N_21374,N_21390);
nor U26428 (N_26428,N_24443,N_24570);
nor U26429 (N_26429,N_23795,N_22546);
nor U26430 (N_26430,N_20057,N_22937);
and U26431 (N_26431,N_24283,N_22943);
xor U26432 (N_26432,N_21280,N_24849);
xor U26433 (N_26433,N_20502,N_22908);
nor U26434 (N_26434,N_22874,N_24285);
or U26435 (N_26435,N_21974,N_23781);
or U26436 (N_26436,N_22011,N_24149);
and U26437 (N_26437,N_20855,N_21418);
nor U26438 (N_26438,N_21421,N_20232);
xor U26439 (N_26439,N_23972,N_21489);
or U26440 (N_26440,N_23738,N_23218);
or U26441 (N_26441,N_21131,N_24436);
or U26442 (N_26442,N_23590,N_22211);
nor U26443 (N_26443,N_20279,N_24272);
and U26444 (N_26444,N_23101,N_21704);
or U26445 (N_26445,N_24685,N_23001);
nand U26446 (N_26446,N_21499,N_21393);
nand U26447 (N_26447,N_20056,N_22319);
nand U26448 (N_26448,N_21937,N_22291);
xor U26449 (N_26449,N_23838,N_23291);
nand U26450 (N_26450,N_22615,N_24105);
or U26451 (N_26451,N_21928,N_20568);
and U26452 (N_26452,N_22627,N_24768);
nor U26453 (N_26453,N_23815,N_22966);
and U26454 (N_26454,N_21254,N_23596);
xnor U26455 (N_26455,N_21855,N_24188);
and U26456 (N_26456,N_21951,N_21312);
xor U26457 (N_26457,N_24526,N_22023);
and U26458 (N_26458,N_23503,N_23549);
and U26459 (N_26459,N_20303,N_24625);
nor U26460 (N_26460,N_22979,N_21587);
xor U26461 (N_26461,N_22986,N_20225);
nand U26462 (N_26462,N_20829,N_20980);
nand U26463 (N_26463,N_24647,N_23667);
nand U26464 (N_26464,N_24736,N_24199);
xor U26465 (N_26465,N_24021,N_22603);
xor U26466 (N_26466,N_24394,N_20102);
or U26467 (N_26467,N_20840,N_20852);
xnor U26468 (N_26468,N_22833,N_20635);
nand U26469 (N_26469,N_20030,N_21464);
xnor U26470 (N_26470,N_22847,N_24432);
or U26471 (N_26471,N_21279,N_22553);
and U26472 (N_26472,N_23980,N_20971);
or U26473 (N_26473,N_20892,N_21079);
nor U26474 (N_26474,N_23142,N_21994);
nand U26475 (N_26475,N_24833,N_24701);
or U26476 (N_26476,N_23573,N_21923);
and U26477 (N_26477,N_20783,N_21740);
and U26478 (N_26478,N_21871,N_21809);
xnor U26479 (N_26479,N_21202,N_23270);
or U26480 (N_26480,N_24854,N_20323);
xnor U26481 (N_26481,N_21778,N_21806);
nor U26482 (N_26482,N_22028,N_21482);
or U26483 (N_26483,N_24912,N_24332);
nor U26484 (N_26484,N_21224,N_22520);
nand U26485 (N_26485,N_22719,N_24108);
and U26486 (N_26486,N_23084,N_21264);
nor U26487 (N_26487,N_24575,N_23651);
nor U26488 (N_26488,N_21246,N_20423);
and U26489 (N_26489,N_20729,N_24135);
xnor U26490 (N_26490,N_20529,N_20790);
nor U26491 (N_26491,N_21906,N_20410);
and U26492 (N_26492,N_20216,N_22362);
nand U26493 (N_26493,N_23597,N_23516);
xor U26494 (N_26494,N_20064,N_22171);
xor U26495 (N_26495,N_23250,N_21258);
xor U26496 (N_26496,N_21698,N_21946);
or U26497 (N_26497,N_23209,N_21525);
nor U26498 (N_26498,N_22564,N_21152);
nor U26499 (N_26499,N_22633,N_23862);
and U26500 (N_26500,N_21785,N_22906);
xor U26501 (N_26501,N_21530,N_22076);
nand U26502 (N_26502,N_22017,N_22561);
or U26503 (N_26503,N_21252,N_22299);
nor U26504 (N_26504,N_24490,N_20054);
xnor U26505 (N_26505,N_23416,N_22958);
or U26506 (N_26506,N_20238,N_20522);
or U26507 (N_26507,N_20864,N_20826);
xor U26508 (N_26508,N_21758,N_20441);
xnor U26509 (N_26509,N_22534,N_20383);
xor U26510 (N_26510,N_23040,N_20031);
nor U26511 (N_26511,N_22842,N_22164);
nor U26512 (N_26512,N_22126,N_23867);
or U26513 (N_26513,N_23859,N_20029);
or U26514 (N_26514,N_24165,N_21685);
or U26515 (N_26515,N_20309,N_22132);
xnor U26516 (N_26516,N_24568,N_22665);
xor U26517 (N_26517,N_22599,N_21942);
nor U26518 (N_26518,N_20486,N_24679);
nor U26519 (N_26519,N_20944,N_20299);
or U26520 (N_26520,N_24936,N_24728);
nand U26521 (N_26521,N_21123,N_21114);
nand U26522 (N_26522,N_22786,N_24051);
xnor U26523 (N_26523,N_22888,N_23802);
xnor U26524 (N_26524,N_23897,N_21149);
xor U26525 (N_26525,N_22114,N_20960);
and U26526 (N_26526,N_20558,N_20042);
xnor U26527 (N_26527,N_21422,N_24052);
xnor U26528 (N_26528,N_24892,N_20962);
nand U26529 (N_26529,N_23299,N_20169);
or U26530 (N_26530,N_23386,N_22142);
nand U26531 (N_26531,N_23690,N_22983);
nand U26532 (N_26532,N_24929,N_22263);
nor U26533 (N_26533,N_22343,N_20197);
nand U26534 (N_26534,N_21158,N_24184);
nor U26535 (N_26535,N_23034,N_21189);
nor U26536 (N_26536,N_22446,N_24748);
or U26537 (N_26537,N_20269,N_20865);
nand U26538 (N_26538,N_23269,N_23893);
and U26539 (N_26539,N_20487,N_23244);
nand U26540 (N_26540,N_20779,N_22052);
or U26541 (N_26541,N_22514,N_24419);
or U26542 (N_26542,N_21343,N_20606);
nand U26543 (N_26543,N_22390,N_22136);
or U26544 (N_26544,N_23533,N_23419);
xor U26545 (N_26545,N_20470,N_23758);
nand U26546 (N_26546,N_21317,N_21984);
nand U26547 (N_26547,N_21243,N_20300);
nand U26548 (N_26548,N_20722,N_22903);
nor U26549 (N_26549,N_24190,N_23971);
xor U26550 (N_26550,N_24218,N_20278);
nand U26551 (N_26551,N_23403,N_22731);
nor U26552 (N_26552,N_21387,N_20545);
and U26553 (N_26553,N_21206,N_24543);
nand U26554 (N_26554,N_21288,N_24595);
nor U26555 (N_26555,N_20159,N_20673);
or U26556 (N_26556,N_20268,N_21295);
or U26557 (N_26557,N_24623,N_21260);
xor U26558 (N_26558,N_22054,N_20930);
and U26559 (N_26559,N_20623,N_22526);
or U26560 (N_26560,N_21544,N_22875);
nand U26561 (N_26561,N_20179,N_20583);
xnor U26562 (N_26562,N_21296,N_21944);
nand U26563 (N_26563,N_22963,N_22304);
xnor U26564 (N_26564,N_22607,N_24757);
xnor U26565 (N_26565,N_23801,N_21999);
or U26566 (N_26566,N_20283,N_22403);
nand U26567 (N_26567,N_22450,N_21649);
nor U26568 (N_26568,N_22429,N_24260);
nor U26569 (N_26569,N_23117,N_21907);
and U26570 (N_26570,N_22223,N_24433);
and U26571 (N_26571,N_22926,N_21420);
xor U26572 (N_26572,N_23453,N_21566);
nand U26573 (N_26573,N_20329,N_24279);
nand U26574 (N_26574,N_23913,N_24412);
nand U26575 (N_26575,N_22039,N_24773);
xor U26576 (N_26576,N_23154,N_22522);
xor U26577 (N_26577,N_20924,N_21095);
xor U26578 (N_26578,N_22993,N_22105);
nand U26579 (N_26579,N_23679,N_24180);
xnor U26580 (N_26580,N_21741,N_22300);
nor U26581 (N_26581,N_21460,N_22024);
xor U26582 (N_26582,N_23373,N_20819);
nor U26583 (N_26583,N_22271,N_22324);
and U26584 (N_26584,N_21864,N_24122);
nand U26585 (N_26585,N_21537,N_21217);
nand U26586 (N_26586,N_23922,N_23775);
nor U26587 (N_26587,N_21384,N_23626);
or U26588 (N_26588,N_22486,N_21595);
xnor U26589 (N_26589,N_22863,N_22933);
or U26590 (N_26590,N_23274,N_23314);
xnor U26591 (N_26591,N_24525,N_23705);
nor U26592 (N_26592,N_22492,N_20067);
or U26593 (N_26593,N_21128,N_23135);
and U26594 (N_26594,N_24047,N_23400);
nand U26595 (N_26595,N_24151,N_22341);
nand U26596 (N_26596,N_22497,N_21456);
nor U26597 (N_26597,N_21766,N_24456);
xor U26598 (N_26598,N_20084,N_23459);
or U26599 (N_26599,N_20651,N_24308);
and U26600 (N_26600,N_23337,N_20058);
and U26601 (N_26601,N_23601,N_22524);
xor U26602 (N_26602,N_21035,N_21896);
nor U26603 (N_26603,N_23694,N_24735);
nand U26604 (N_26604,N_24268,N_21232);
nand U26605 (N_26605,N_22041,N_20094);
or U26606 (N_26606,N_23674,N_21976);
and U26607 (N_26607,N_23965,N_21801);
nor U26608 (N_26608,N_24645,N_24686);
nor U26609 (N_26609,N_21495,N_24290);
nor U26610 (N_26610,N_24121,N_24596);
nand U26611 (N_26611,N_22718,N_22954);
and U26612 (N_26612,N_23723,N_24287);
nand U26613 (N_26613,N_22106,N_20662);
xor U26614 (N_26614,N_24083,N_21614);
nand U26615 (N_26615,N_21318,N_23572);
xnor U26616 (N_26616,N_22172,N_22488);
or U26617 (N_26617,N_24424,N_23792);
xor U26618 (N_26618,N_24801,N_21924);
nand U26619 (N_26619,N_23095,N_21841);
xor U26620 (N_26620,N_20772,N_24905);
nand U26621 (N_26621,N_22883,N_20520);
nor U26622 (N_26622,N_20661,N_21836);
and U26623 (N_26623,N_20403,N_24379);
nand U26624 (N_26624,N_22691,N_20887);
nor U26625 (N_26625,N_22635,N_20205);
xnor U26626 (N_26626,N_24066,N_20705);
xor U26627 (N_26627,N_22947,N_20885);
or U26628 (N_26628,N_20614,N_20185);
xnor U26629 (N_26629,N_23256,N_20035);
nor U26630 (N_26630,N_20296,N_23903);
xnor U26631 (N_26631,N_21728,N_22656);
nand U26632 (N_26632,N_24355,N_20006);
or U26633 (N_26633,N_22432,N_21771);
and U26634 (N_26634,N_22318,N_23520);
and U26635 (N_26635,N_23550,N_24530);
nand U26636 (N_26636,N_23959,N_22102);
xnor U26637 (N_26637,N_20574,N_21122);
and U26638 (N_26638,N_22368,N_20041);
or U26639 (N_26639,N_23931,N_24681);
nor U26640 (N_26640,N_23916,N_23145);
and U26641 (N_26641,N_20226,N_22746);
nand U26642 (N_26642,N_24614,N_23555);
and U26643 (N_26643,N_21917,N_20065);
xnor U26644 (N_26644,N_20859,N_20908);
nor U26645 (N_26645,N_23785,N_20889);
and U26646 (N_26646,N_23118,N_23009);
or U26647 (N_26647,N_23046,N_23839);
and U26648 (N_26648,N_21905,N_23784);
and U26649 (N_26649,N_23997,N_21366);
xor U26650 (N_26650,N_20897,N_24036);
xnor U26651 (N_26651,N_20957,N_22086);
and U26652 (N_26652,N_21516,N_24242);
xnor U26653 (N_26653,N_20996,N_21835);
xor U26654 (N_26654,N_21016,N_22637);
xnor U26655 (N_26655,N_21491,N_20521);
xor U26656 (N_26656,N_20178,N_20995);
or U26657 (N_26657,N_20316,N_22252);
nand U26658 (N_26658,N_23615,N_22711);
or U26659 (N_26659,N_24957,N_22005);
or U26660 (N_26660,N_21400,N_20223);
nand U26661 (N_26661,N_20949,N_23703);
nor U26662 (N_26662,N_21395,N_23616);
xor U26663 (N_26663,N_20317,N_23398);
or U26664 (N_26664,N_20188,N_23413);
nand U26665 (N_26665,N_20630,N_21399);
xnor U26666 (N_26666,N_23227,N_24023);
or U26667 (N_26667,N_20157,N_23226);
and U26668 (N_26668,N_23987,N_24699);
and U26669 (N_26669,N_21594,N_24752);
xor U26670 (N_26670,N_21012,N_22184);
nor U26671 (N_26671,N_21908,N_24780);
and U26672 (N_26672,N_22110,N_22321);
nor U26673 (N_26673,N_20676,N_22812);
or U26674 (N_26674,N_22124,N_24972);
nor U26675 (N_26675,N_22113,N_22834);
nor U26676 (N_26676,N_23663,N_21893);
nor U26677 (N_26677,N_23592,N_22262);
or U26678 (N_26678,N_22345,N_21683);
nor U26679 (N_26679,N_22595,N_23423);
and U26680 (N_26680,N_24062,N_24409);
nor U26681 (N_26681,N_23629,N_24689);
nand U26682 (N_26682,N_23751,N_23563);
and U26683 (N_26683,N_20183,N_22100);
xnor U26684 (N_26684,N_24554,N_23584);
nand U26685 (N_26685,N_23660,N_20555);
nand U26686 (N_26686,N_21712,N_22021);
nor U26687 (N_26687,N_24970,N_24942);
nand U26688 (N_26688,N_23743,N_24533);
and U26689 (N_26689,N_20386,N_21496);
xor U26690 (N_26690,N_21748,N_24818);
xnor U26691 (N_26691,N_23595,N_22843);
or U26692 (N_26692,N_24317,N_20193);
and U26693 (N_26693,N_22959,N_21121);
nand U26694 (N_26694,N_21091,N_22789);
and U26695 (N_26695,N_24395,N_23169);
nand U26696 (N_26696,N_24303,N_20625);
nand U26697 (N_26697,N_20053,N_23276);
or U26698 (N_26698,N_20746,N_23577);
nand U26699 (N_26699,N_20557,N_21684);
or U26700 (N_26700,N_23289,N_20668);
nor U26701 (N_26701,N_21526,N_24230);
or U26702 (N_26702,N_24545,N_23178);
xnor U26703 (N_26703,N_20825,N_22821);
nor U26704 (N_26704,N_21270,N_22147);
nand U26705 (N_26705,N_20539,N_22022);
and U26706 (N_26706,N_23482,N_22852);
nand U26707 (N_26707,N_21839,N_24274);
or U26708 (N_26708,N_23734,N_21930);
and U26709 (N_26709,N_22101,N_21618);
or U26710 (N_26710,N_21792,N_22658);
nor U26711 (N_26711,N_24852,N_22519);
xor U26712 (N_26712,N_24216,N_21459);
xor U26713 (N_26713,N_20043,N_22761);
nand U26714 (N_26714,N_20704,N_21949);
xnor U26715 (N_26715,N_21249,N_23797);
nand U26716 (N_26716,N_21040,N_24943);
nor U26717 (N_26717,N_23119,N_20009);
nand U26718 (N_26718,N_20761,N_24551);
and U26719 (N_26719,N_22549,N_22775);
nand U26720 (N_26720,N_21304,N_23776);
nand U26721 (N_26721,N_21613,N_22855);
xnor U26722 (N_26722,N_22006,N_20619);
xnor U26723 (N_26723,N_24398,N_22573);
nand U26724 (N_26724,N_21315,N_21856);
and U26725 (N_26725,N_24055,N_20165);
nor U26726 (N_26726,N_24324,N_23754);
nor U26727 (N_26727,N_20413,N_21212);
nand U26728 (N_26728,N_22504,N_22077);
xor U26729 (N_26729,N_24387,N_24183);
or U26730 (N_26730,N_24985,N_20910);
and U26731 (N_26731,N_21711,N_24832);
and U26732 (N_26732,N_21299,N_22547);
or U26733 (N_26733,N_23166,N_22229);
xnor U26734 (N_26734,N_22642,N_20324);
xor U26735 (N_26735,N_22915,N_23249);
nor U26736 (N_26736,N_22682,N_23027);
nor U26737 (N_26737,N_24759,N_22125);
xor U26738 (N_26738,N_24510,N_23253);
or U26739 (N_26739,N_20798,N_20242);
xnor U26740 (N_26740,N_20709,N_24907);
nand U26741 (N_26741,N_20664,N_20670);
or U26742 (N_26742,N_22127,N_24745);
nor U26743 (N_26743,N_22946,N_22769);
and U26744 (N_26744,N_23087,N_24077);
xnor U26745 (N_26745,N_23312,N_20352);
nor U26746 (N_26746,N_21997,N_21098);
nand U26747 (N_26747,N_23969,N_20464);
or U26748 (N_26748,N_22618,N_21493);
nand U26749 (N_26749,N_22312,N_20815);
nor U26750 (N_26750,N_23525,N_22654);
or U26751 (N_26751,N_21011,N_20099);
xor U26752 (N_26752,N_21027,N_24607);
and U26753 (N_26753,N_23042,N_23755);
xnor U26754 (N_26754,N_23092,N_24226);
and U26755 (N_26755,N_22572,N_21555);
nor U26756 (N_26756,N_21589,N_20093);
or U26757 (N_26757,N_21345,N_21414);
and U26758 (N_26758,N_22140,N_21727);
xnor U26759 (N_26759,N_22816,N_20727);
and U26760 (N_26760,N_22922,N_21244);
and U26761 (N_26761,N_23617,N_21719);
and U26762 (N_26762,N_24814,N_23693);
or U26763 (N_26763,N_23880,N_20611);
xor U26764 (N_26764,N_20653,N_21721);
or U26765 (N_26765,N_24314,N_21573);
or U26766 (N_26766,N_22835,N_21717);
or U26767 (N_26767,N_24046,N_23900);
nand U26768 (N_26768,N_21487,N_23788);
nand U26769 (N_26769,N_21996,N_23260);
nor U26770 (N_26770,N_23739,N_22072);
or U26771 (N_26771,N_20749,N_22201);
xor U26772 (N_26772,N_20886,N_21747);
and U26773 (N_26773,N_20290,N_21901);
xnor U26774 (N_26774,N_23632,N_23454);
and U26775 (N_26775,N_21545,N_23396);
and U26776 (N_26776,N_22831,N_22500);
and U26777 (N_26777,N_22884,N_21110);
nand U26778 (N_26778,N_24737,N_23678);
or U26779 (N_26779,N_22965,N_21561);
and U26780 (N_26780,N_21065,N_23721);
nand U26781 (N_26781,N_24273,N_24382);
xnor U26782 (N_26782,N_23886,N_20123);
nand U26783 (N_26783,N_24858,N_23725);
or U26784 (N_26784,N_21298,N_20298);
xor U26785 (N_26785,N_20731,N_20026);
nor U26786 (N_26786,N_23155,N_21643);
or U26787 (N_26787,N_20097,N_24191);
or U26788 (N_26788,N_24894,N_21682);
xor U26789 (N_26789,N_20893,N_20698);
nand U26790 (N_26790,N_21838,N_22536);
xnor U26791 (N_26791,N_22512,N_21636);
and U26792 (N_26792,N_21725,N_22388);
xor U26793 (N_26793,N_24560,N_20721);
nor U26794 (N_26794,N_21583,N_21204);
or U26795 (N_26795,N_24619,N_23350);
xor U26796 (N_26796,N_21921,N_20089);
nand U26797 (N_26797,N_23342,N_20771);
nand U26798 (N_26798,N_24656,N_23360);
or U26799 (N_26799,N_24476,N_23697);
or U26800 (N_26800,N_23719,N_20665);
or U26801 (N_26801,N_21197,N_21052);
and U26802 (N_26802,N_24442,N_22387);
or U26803 (N_26803,N_20748,N_20050);
nand U26804 (N_26804,N_24185,N_24552);
nor U26805 (N_26805,N_21336,N_23105);
or U26806 (N_26806,N_22811,N_21242);
or U26807 (N_26807,N_20129,N_22372);
nand U26808 (N_26808,N_21929,N_22071);
nor U26809 (N_26809,N_23962,N_20760);
or U26810 (N_26810,N_20424,N_22311);
xor U26811 (N_26811,N_22581,N_20113);
or U26812 (N_26812,N_20418,N_23659);
and U26813 (N_26813,N_21219,N_20550);
nand U26814 (N_26814,N_22141,N_21891);
or U26815 (N_26815,N_20112,N_21140);
or U26816 (N_26816,N_22428,N_24261);
xnor U26817 (N_26817,N_22560,N_22578);
xor U26818 (N_26818,N_23492,N_24461);
or U26819 (N_26819,N_24823,N_24920);
or U26820 (N_26820,N_21630,N_22198);
and U26821 (N_26821,N_24591,N_24913);
xnor U26822 (N_26822,N_23866,N_24695);
and U26823 (N_26823,N_24371,N_23531);
or U26824 (N_26824,N_20376,N_22499);
xor U26825 (N_26825,N_21824,N_20848);
xnor U26826 (N_26826,N_21062,N_22891);
nand U26827 (N_26827,N_21372,N_21333);
xnor U26828 (N_26828,N_21039,N_22622);
or U26829 (N_26829,N_20438,N_23973);
nand U26830 (N_26830,N_23814,N_24865);
nor U26831 (N_26831,N_22781,N_21376);
and U26832 (N_26832,N_20019,N_23910);
nand U26833 (N_26833,N_22543,N_21932);
nand U26834 (N_26834,N_21442,N_23576);
and U26835 (N_26835,N_21115,N_23587);
nand U26836 (N_26836,N_24653,N_21540);
or U26837 (N_26837,N_23165,N_23080);
and U26838 (N_26838,N_22083,N_24177);
xnor U26839 (N_26839,N_23543,N_22496);
nand U26840 (N_26840,N_22758,N_24600);
or U26841 (N_26841,N_21046,N_23570);
and U26842 (N_26842,N_21810,N_21962);
nor U26843 (N_26843,N_21105,N_20481);
nand U26844 (N_26844,N_22583,N_22200);
nand U26845 (N_26845,N_23357,N_21465);
nand U26846 (N_26846,N_23281,N_20257);
and U26847 (N_26847,N_20624,N_21431);
xnor U26848 (N_26848,N_22120,N_24219);
nand U26849 (N_26849,N_22902,N_24658);
nor U26850 (N_26850,N_22755,N_20978);
nand U26851 (N_26851,N_24175,N_23732);
nand U26852 (N_26852,N_20835,N_24889);
or U26853 (N_26853,N_22621,N_24794);
or U26854 (N_26854,N_21842,N_21371);
or U26855 (N_26855,N_21653,N_24603);
and U26856 (N_26856,N_20404,N_24220);
nand U26857 (N_26857,N_21673,N_23999);
and U26858 (N_26858,N_21031,N_22710);
or U26859 (N_26859,N_23704,N_21205);
nand U26860 (N_26860,N_21477,N_22503);
nor U26861 (N_26861,N_20227,N_24343);
or U26862 (N_26862,N_22801,N_21534);
nor U26863 (N_26863,N_22555,N_22494);
nor U26864 (N_26864,N_22459,N_24132);
xnor U26865 (N_26865,N_22796,N_24902);
and U26866 (N_26866,N_24494,N_20241);
nor U26867 (N_26867,N_23159,N_20126);
and U26868 (N_26868,N_22559,N_22856);
or U26869 (N_26869,N_24900,N_24675);
and U26870 (N_26870,N_24302,N_22035);
and U26871 (N_26871,N_20090,N_21132);
xor U26872 (N_26872,N_24349,N_23656);
or U26873 (N_26873,N_20523,N_20360);
nor U26874 (N_26874,N_23062,N_20261);
and U26875 (N_26875,N_24071,N_22941);
nor U26876 (N_26876,N_24211,N_21017);
or U26877 (N_26877,N_21624,N_24758);
or U26878 (N_26878,N_20020,N_20172);
and U26879 (N_26879,N_22287,N_23188);
xnor U26880 (N_26880,N_20105,N_23631);
and U26881 (N_26881,N_23371,N_21054);
xnor U26882 (N_26882,N_21347,N_23298);
xor U26883 (N_26883,N_20039,N_22044);
and U26884 (N_26884,N_22756,N_20752);
nand U26885 (N_26885,N_23018,N_22861);
nor U26886 (N_26886,N_22984,N_23308);
nor U26887 (N_26887,N_24726,N_22632);
nand U26888 (N_26888,N_23844,N_24741);
nor U26889 (N_26889,N_20038,N_21995);
and U26890 (N_26890,N_21417,N_21198);
nand U26891 (N_26891,N_23874,N_23937);
or U26892 (N_26892,N_22025,N_20322);
xnor U26893 (N_26893,N_24365,N_22019);
and U26894 (N_26894,N_23290,N_24061);
and U26895 (N_26895,N_23235,N_23498);
nor U26896 (N_26896,N_24195,N_24401);
or U26897 (N_26897,N_24666,N_20012);
nor U26898 (N_26898,N_21760,N_24484);
nor U26899 (N_26899,N_21680,N_22279);
nand U26900 (N_26900,N_23643,N_21086);
xnor U26901 (N_26901,N_22824,N_21508);
nor U26902 (N_26902,N_21162,N_22830);
xnor U26903 (N_26903,N_20890,N_24040);
xnor U26904 (N_26904,N_23199,N_24144);
and U26905 (N_26905,N_23272,N_20444);
nand U26906 (N_26906,N_21133,N_22415);
nor U26907 (N_26907,N_20955,N_23427);
or U26908 (N_26908,N_21494,N_24988);
or U26909 (N_26909,N_20377,N_20723);
nor U26910 (N_26910,N_20427,N_21229);
nand U26911 (N_26911,N_22844,N_20409);
nor U26912 (N_26912,N_20436,N_20856);
xor U26913 (N_26913,N_23327,N_23128);
xor U26914 (N_26914,N_23536,N_22413);
nand U26915 (N_26915,N_22590,N_22191);
nand U26916 (N_26916,N_23506,N_21763);
nand U26917 (N_26917,N_24306,N_24315);
nor U26918 (N_26918,N_20612,N_24598);
or U26919 (N_26919,N_20553,N_22442);
xor U26920 (N_26920,N_24086,N_24893);
and U26921 (N_26921,N_22669,N_24256);
nor U26922 (N_26922,N_24380,N_21423);
nor U26923 (N_26923,N_20380,N_22003);
xor U26924 (N_26924,N_21116,N_23888);
nand U26925 (N_26925,N_23990,N_21461);
or U26926 (N_26926,N_20008,N_21884);
and U26927 (N_26927,N_20286,N_22160);
and U26928 (N_26928,N_21978,N_22630);
nor U26929 (N_26929,N_23391,N_22061);
xnor U26930 (N_26930,N_20547,N_21284);
nor U26931 (N_26931,N_22121,N_24202);
or U26932 (N_26932,N_22662,N_22712);
nand U26933 (N_26933,N_22009,N_20014);
nand U26934 (N_26934,N_22663,N_23493);
or U26935 (N_26935,N_24110,N_20349);
nand U26936 (N_26936,N_21083,N_21642);
nand U26937 (N_26937,N_22552,N_24563);
nor U26938 (N_26938,N_24426,N_24817);
nor U26939 (N_26939,N_20339,N_20570);
xor U26940 (N_26940,N_24404,N_24627);
nand U26941 (N_26941,N_24249,N_24822);
or U26942 (N_26942,N_21791,N_22296);
and U26943 (N_26943,N_21823,N_24960);
nor U26944 (N_26944,N_20337,N_22797);
or U26945 (N_26945,N_24163,N_21163);
nand U26946 (N_26946,N_24561,N_20966);
nand U26947 (N_26947,N_21208,N_21687);
xor U26948 (N_26948,N_24853,N_23205);
nor U26949 (N_26949,N_22270,N_24239);
nor U26950 (N_26950,N_22389,N_23927);
and U26951 (N_26951,N_20001,N_24114);
xnor U26952 (N_26952,N_23374,N_22361);
or U26953 (N_26953,N_21708,N_22567);
xnor U26954 (N_26954,N_24212,N_23429);
or U26955 (N_26955,N_23401,N_20326);
and U26956 (N_26956,N_21590,N_20891);
and U26957 (N_26957,N_22119,N_24756);
and U26958 (N_26958,N_20292,N_24649);
xnor U26959 (N_26959,N_22995,N_24693);
and U26960 (N_26960,N_21668,N_22594);
nand U26961 (N_26961,N_20710,N_22008);
and U26962 (N_26962,N_22051,N_23657);
xnor U26963 (N_26963,N_24269,N_22657);
or U26964 (N_26964,N_20827,N_21608);
or U26965 (N_26965,N_21800,N_24507);
nand U26966 (N_26966,N_23313,N_21228);
and U26967 (N_26967,N_20786,N_23393);
or U26968 (N_26968,N_22485,N_23115);
nor U26969 (N_26969,N_24301,N_22608);
xnor U26970 (N_26970,N_24439,N_22509);
nand U26971 (N_26971,N_22715,N_22169);
xnor U26972 (N_26972,N_24937,N_21750);
and U26973 (N_26973,N_22115,N_23661);
nor U26974 (N_26974,N_21169,N_23600);
nand U26975 (N_26975,N_21574,N_23608);
nand U26976 (N_26976,N_23688,N_21811);
xor U26977 (N_26977,N_24106,N_23031);
xor U26978 (N_26978,N_20657,N_23051);
or U26979 (N_26979,N_21337,N_22675);
xor U26980 (N_26980,N_20769,N_22182);
xnor U26981 (N_26981,N_23201,N_24145);
and U26982 (N_26982,N_20548,N_21428);
xor U26983 (N_26983,N_23132,N_22290);
or U26984 (N_26984,N_24262,N_23816);
nand U26985 (N_26985,N_23133,N_23702);
xor U26986 (N_26986,N_22673,N_23843);
xor U26987 (N_26987,N_22565,N_21958);
or U26988 (N_26988,N_21959,N_24372);
nand U26989 (N_26989,N_20021,N_22877);
and U26990 (N_26990,N_21605,N_23160);
xor U26991 (N_26991,N_21396,N_22631);
nor U26992 (N_26992,N_24868,N_21706);
nor U26993 (N_26993,N_21576,N_24160);
or U26994 (N_26994,N_22053,N_21058);
nand U26995 (N_26995,N_23341,N_20876);
nand U26996 (N_26996,N_24714,N_20434);
nor U26997 (N_26997,N_23818,N_22452);
xnor U26998 (N_26998,N_24548,N_23211);
nand U26999 (N_26999,N_23770,N_22584);
and U27000 (N_27000,N_23208,N_23856);
nand U27001 (N_27001,N_21203,N_20199);
and U27002 (N_27002,N_24304,N_22346);
nand U27003 (N_27003,N_24717,N_24489);
or U27004 (N_27004,N_23233,N_23762);
or U27005 (N_27005,N_20246,N_22325);
and U27006 (N_27006,N_22784,N_24099);
and U27007 (N_27007,N_23220,N_23261);
xor U27008 (N_27008,N_20139,N_21401);
xor U27009 (N_27009,N_24795,N_20877);
nor U27010 (N_27010,N_24727,N_21575);
nand U27011 (N_27011,N_23583,N_23437);
and U27012 (N_27012,N_22793,N_22378);
xnor U27013 (N_27013,N_24634,N_24926);
or U27014 (N_27014,N_23375,N_21084);
nand U27015 (N_27015,N_23918,N_21441);
and U27016 (N_27016,N_23303,N_20730);
or U27017 (N_27017,N_20596,N_23295);
nor U27018 (N_27018,N_21726,N_20791);
and U27019 (N_27019,N_21214,N_23833);
xnor U27020 (N_27020,N_23093,N_22967);
xnor U27021 (N_27021,N_23104,N_21617);
and U27022 (N_27022,N_22027,N_20708);
nand U27023 (N_27023,N_22648,N_22248);
nor U27024 (N_27024,N_24014,N_24544);
nand U27025 (N_27025,N_22467,N_20381);
xnor U27026 (N_27026,N_21449,N_24862);
xnor U27027 (N_27027,N_23653,N_20149);
xor U27028 (N_27028,N_20977,N_23963);
or U27029 (N_27029,N_21474,N_24037);
or U27030 (N_27030,N_24194,N_23240);
nor U27031 (N_27031,N_20914,N_21383);
nand U27032 (N_27032,N_23365,N_20898);
or U27033 (N_27033,N_20221,N_21998);
xor U27034 (N_27034,N_23926,N_23007);
nand U27035 (N_27035,N_20714,N_20489);
nor U27036 (N_27036,N_23254,N_23008);
nor U27037 (N_27037,N_23677,N_21847);
nor U27038 (N_27038,N_23376,N_20818);
or U27039 (N_27039,N_24506,N_20457);
or U27040 (N_27040,N_22807,N_21897);
xor U27041 (N_27041,N_22431,N_20312);
nor U27042 (N_27042,N_24793,N_20459);
xor U27043 (N_27043,N_21903,N_20075);
nand U27044 (N_27044,N_23026,N_20011);
or U27045 (N_27045,N_23558,N_24682);
xor U27046 (N_27046,N_22687,N_22964);
or U27047 (N_27047,N_23421,N_20397);
or U27048 (N_27048,N_23024,N_20810);
or U27049 (N_27049,N_20762,N_21964);
and U27050 (N_27050,N_21042,N_21138);
and U27051 (N_27051,N_20587,N_24549);
xnor U27052 (N_27052,N_21327,N_20940);
nand U27053 (N_27053,N_24182,N_23451);
and U27054 (N_27054,N_23848,N_23148);
xor U27055 (N_27055,N_20589,N_20875);
nand U27056 (N_27056,N_22392,N_23724);
and U27057 (N_27057,N_21109,N_22507);
xor U27058 (N_27058,N_21531,N_20592);
nand U27059 (N_27059,N_23070,N_22444);
or U27060 (N_27060,N_20556,N_23692);
nor U27061 (N_27061,N_24775,N_24460);
and U27062 (N_27062,N_23417,N_21878);
nand U27063 (N_27063,N_24762,N_21359);
or U27064 (N_27064,N_21407,N_20260);
and U27065 (N_27065,N_24861,N_24109);
or U27066 (N_27066,N_22505,N_20544);
nor U27067 (N_27067,N_23448,N_24845);
and U27068 (N_27068,N_24340,N_24388);
nor U27069 (N_27069,N_21302,N_22991);
nand U27070 (N_27070,N_22668,N_20369);
nor U27071 (N_27071,N_22601,N_21504);
nor U27072 (N_27072,N_23830,N_23744);
nor U27073 (N_27073,N_22788,N_21348);
or U27074 (N_27074,N_21860,N_22046);
and U27075 (N_27075,N_24477,N_21081);
nand U27076 (N_27076,N_20585,N_21755);
nand U27077 (N_27077,N_24831,N_21369);
nor U27078 (N_27078,N_21385,N_22981);
or U27079 (N_27079,N_21879,N_24475);
xor U27080 (N_27080,N_21940,N_23073);
or U27081 (N_27081,N_21188,N_24208);
xnor U27082 (N_27082,N_23292,N_20671);
xor U27083 (N_27083,N_23438,N_22130);
nor U27084 (N_27084,N_22862,N_24251);
or U27085 (N_27085,N_24458,N_20615);
or U27086 (N_27086,N_22320,N_20237);
xor U27087 (N_27087,N_21567,N_22224);
or U27088 (N_27088,N_20046,N_20468);
xnor U27089 (N_27089,N_23975,N_21671);
and U27090 (N_27090,N_23676,N_21777);
nor U27091 (N_27091,N_21694,N_21452);
nor U27092 (N_27092,N_22326,N_23050);
or U27093 (N_27093,N_20912,N_23245);
or U27094 (N_27094,N_23908,N_23515);
xor U27095 (N_27095,N_23991,N_20146);
xnor U27096 (N_27096,N_23409,N_22374);
and U27097 (N_27097,N_24922,N_24297);
nor U27098 (N_27098,N_21470,N_20240);
xnor U27099 (N_27099,N_22085,N_21155);
nor U27100 (N_27100,N_21175,N_20999);
xor U27101 (N_27101,N_23603,N_24571);
or U27102 (N_27102,N_20888,N_24358);
nand U27103 (N_27103,N_20499,N_21444);
and U27104 (N_27104,N_22562,N_22190);
or U27105 (N_27105,N_21024,N_21889);
nor U27106 (N_27106,N_24661,N_20757);
nor U27107 (N_27107,N_23362,N_23518);
nand U27108 (N_27108,N_23757,N_22614);
xor U27109 (N_27109,N_24640,N_21216);
nor U27110 (N_27110,N_20600,N_24228);
or U27111 (N_27111,N_21201,N_23223);
nand U27112 (N_27112,N_23623,N_24665);
or U27113 (N_27113,N_24400,N_23979);
or U27114 (N_27114,N_22186,N_23206);
xnor U27115 (N_27115,N_22470,N_20015);
nor U27116 (N_27116,N_21890,N_22699);
or U27117 (N_27117,N_22150,N_21899);
or U27118 (N_27118,N_24593,N_24282);
nor U27119 (N_27119,N_21451,N_20667);
nand U27120 (N_27120,N_23388,N_24486);
or U27121 (N_27121,N_24744,N_20535);
and U27122 (N_27122,N_22103,N_21416);
xnor U27123 (N_27123,N_22910,N_22210);
and U27124 (N_27124,N_23098,N_24469);
or U27125 (N_27125,N_22643,N_24359);
nor U27126 (N_27126,N_22701,N_20447);
and U27127 (N_27127,N_20150,N_23348);
nor U27128 (N_27128,N_21334,N_23530);
or U27129 (N_27129,N_20509,N_21088);
and U27130 (N_27130,N_23907,N_24583);
xnor U27131 (N_27131,N_22418,N_20800);
nor U27132 (N_27132,N_22752,N_24537);
nor U27133 (N_27133,N_22170,N_23642);
xor U27134 (N_27134,N_24924,N_21520);
nor U27135 (N_27135,N_22809,N_22602);
nor U27136 (N_27136,N_22678,N_24004);
nand U27137 (N_27137,N_23687,N_24276);
xor U27138 (N_27138,N_22481,N_24101);
nor U27139 (N_27139,N_21099,N_20234);
xor U27140 (N_27140,N_21599,N_24392);
nor U27141 (N_27141,N_23868,N_24626);
nor U27142 (N_27142,N_24081,N_22693);
and U27143 (N_27143,N_24786,N_21783);
nor U27144 (N_27144,N_23102,N_20195);
xor U27145 (N_27145,N_24277,N_24990);
xnor U27146 (N_27146,N_24871,N_20484);
xor U27147 (N_27147,N_24119,N_24541);
or U27148 (N_27148,N_20002,N_24065);
nand U27149 (N_27149,N_21000,N_21641);
nor U27150 (N_27150,N_21512,N_22730);
and U27151 (N_27151,N_20958,N_22382);
or U27152 (N_27152,N_24884,N_24248);
and U27153 (N_27153,N_21001,N_20494);
nor U27154 (N_27154,N_24418,N_24820);
or U27155 (N_27155,N_23384,N_24705);
and U27156 (N_27156,N_22865,N_22870);
nor U27157 (N_27157,N_23630,N_24572);
and U27158 (N_27158,N_21349,N_24417);
xnor U27159 (N_27159,N_24232,N_23707);
xor U27160 (N_27160,N_20263,N_23392);
and U27161 (N_27161,N_24895,N_21405);
and U27162 (N_27162,N_22116,N_21986);
or U27163 (N_27163,N_23349,N_20276);
xor U27164 (N_27164,N_20024,N_21586);
and U27165 (N_27165,N_24179,N_21985);
or U27166 (N_27166,N_20571,N_21111);
xor U27167 (N_27167,N_20994,N_20845);
and U27168 (N_27168,N_20789,N_20311);
nand U27169 (N_27169,N_21514,N_20802);
nor U27170 (N_27170,N_22952,N_23538);
xnor U27171 (N_27171,N_22462,N_21788);
nor U27172 (N_27172,N_21454,N_24402);
and U27173 (N_27173,N_23380,N_22814);
or U27174 (N_27174,N_24275,N_21473);
and U27175 (N_27175,N_22813,N_23411);
and U27176 (N_27176,N_24120,N_22350);
nand U27177 (N_27177,N_24925,N_23711);
and U27178 (N_27178,N_21142,N_24361);
xor U27179 (N_27179,N_20896,N_24788);
nand U27180 (N_27180,N_21703,N_21804);
or U27181 (N_27181,N_21352,N_21379);
or U27182 (N_27182,N_22613,N_22949);
xor U27183 (N_27183,N_24284,N_21367);
and U27184 (N_27184,N_23394,N_21077);
xor U27185 (N_27185,N_24200,N_22529);
xnor U27186 (N_27186,N_22257,N_21808);
or U27187 (N_27187,N_20143,N_21101);
nor U27188 (N_27188,N_20572,N_21950);
or U27189 (N_27189,N_24761,N_20111);
and U27190 (N_27190,N_20618,N_20514);
xnor U27191 (N_27191,N_24502,N_22274);
nand U27192 (N_27192,N_21977,N_22221);
nand U27193 (N_27193,N_21568,N_24089);
nand U27194 (N_27194,N_20743,N_21606);
xor U27195 (N_27195,N_23912,N_21463);
nor U27196 (N_27196,N_20361,N_23904);
nand U27197 (N_27197,N_23074,N_21795);
xor U27198 (N_27198,N_23929,N_22783);
xnor U27199 (N_27199,N_23138,N_23347);
and U27200 (N_27200,N_23099,N_21055);
xor U27201 (N_27201,N_23436,N_20248);
nor U27202 (N_27202,N_22576,N_22013);
nor U27203 (N_27203,N_24123,N_23714);
nand U27204 (N_27204,N_24792,N_24918);
or U27205 (N_27205,N_21802,N_20445);
xnor U27206 (N_27206,N_23898,N_22839);
nor U27207 (N_27207,N_23134,N_20127);
and U27208 (N_27208,N_20167,N_24770);
and U27209 (N_27209,N_20597,N_20497);
or U27210 (N_27210,N_21776,N_21875);
xnor U27211 (N_27211,N_20740,N_20990);
or U27212 (N_27212,N_23953,N_24654);
or U27213 (N_27213,N_20906,N_23106);
xnor U27214 (N_27214,N_22882,N_23264);
nand U27215 (N_27215,N_21365,N_24067);
nand U27216 (N_27216,N_23304,N_22243);
and U27217 (N_27217,N_22727,N_23368);
and U27218 (N_27218,N_21722,N_24739);
and U27219 (N_27219,N_23544,N_24010);
xor U27220 (N_27220,N_21044,N_23691);
and U27221 (N_27221,N_23906,N_21927);
xnor U27222 (N_27222,N_24039,N_24254);
or U27223 (N_27223,N_22506,N_22930);
xor U27224 (N_27224,N_24134,N_20516);
nor U27225 (N_27225,N_23933,N_21503);
nand U27226 (N_27226,N_24427,N_23462);
and U27227 (N_27227,N_21718,N_23120);
nand U27228 (N_27228,N_23358,N_21894);
nor U27229 (N_27229,N_21782,N_23825);
xnor U27230 (N_27230,N_23948,N_22379);
and U27231 (N_27231,N_23382,N_23510);
or U27232 (N_27232,N_23039,N_20235);
nand U27233 (N_27233,N_20919,N_22557);
or U27234 (N_27234,N_22780,N_24800);
or U27235 (N_27235,N_23163,N_22395);
or U27236 (N_27236,N_23425,N_24005);
xnor U27237 (N_27237,N_21578,N_23834);
or U27238 (N_27238,N_24979,N_20929);
nand U27239 (N_27239,N_20077,N_21283);
nor U27240 (N_27240,N_24760,N_22316);
or U27241 (N_27241,N_22084,N_20780);
nor U27242 (N_27242,N_23641,N_22268);
xnor U27243 (N_27243,N_24512,N_23902);
and U27244 (N_27244,N_22273,N_24747);
xnor U27245 (N_27245,N_22237,N_21093);
or U27246 (N_27246,N_22266,N_24999);
xor U27247 (N_27247,N_20233,N_20320);
nor U27248 (N_27248,N_22661,N_21082);
nand U27249 (N_27249,N_21846,N_22453);
or U27250 (N_27250,N_21628,N_23149);
nor U27251 (N_27251,N_21916,N_22315);
and U27252 (N_27252,N_22406,N_20028);
or U27253 (N_27253,N_23275,N_21466);
nor U27254 (N_27254,N_22889,N_24946);
xor U27255 (N_27255,N_24238,N_23941);
nor U27256 (N_27256,N_23445,N_20765);
or U27257 (N_27257,N_23529,N_23287);
xnor U27258 (N_27258,N_24328,N_23016);
nand U27259 (N_27259,N_22088,N_20992);
and U27260 (N_27260,N_23251,N_24025);
and U27261 (N_27261,N_20734,N_24214);
nor U27262 (N_27262,N_23917,N_20853);
nand U27263 (N_27263,N_23071,N_23852);
nand U27264 (N_27264,N_21975,N_24410);
nor U27265 (N_27265,N_23354,N_22408);
or U27266 (N_27266,N_22757,N_21845);
nand U27267 (N_27267,N_20310,N_22244);
nand U27268 (N_27268,N_21580,N_23030);
or U27269 (N_27269,N_23468,N_20304);
or U27270 (N_27270,N_24723,N_24523);
nor U27271 (N_27271,N_24011,N_22117);
nand U27272 (N_27272,N_20414,N_21730);
nor U27273 (N_27273,N_22337,N_23599);
or U27274 (N_27274,N_22177,N_24878);
nor U27275 (N_27275,N_21059,N_23782);
xnor U27276 (N_27276,N_24612,N_21911);
and U27277 (N_27277,N_21119,N_23562);
nand U27278 (N_27278,N_20822,N_24318);
and U27279 (N_27279,N_22767,N_21882);
or U27280 (N_27280,N_23628,N_23172);
and U27281 (N_27281,N_24539,N_22240);
and U27282 (N_27282,N_22892,N_22349);
and U27283 (N_27283,N_23764,N_20869);
nor U27284 (N_27284,N_21702,N_24012);
and U27285 (N_27285,N_22093,N_23804);
nand U27286 (N_27286,N_24150,N_22394);
nand U27287 (N_27287,N_22591,N_20163);
xnor U27288 (N_27288,N_23076,N_24585);
or U27289 (N_27289,N_23683,N_23190);
nand U27290 (N_27290,N_23047,N_20297);
xnor U27291 (N_27291,N_20687,N_21230);
and U27292 (N_27292,N_23625,N_23554);
nand U27293 (N_27293,N_22295,N_24622);
or U27294 (N_27294,N_24096,N_20498);
nor U27295 (N_27295,N_20032,N_21053);
nand U27296 (N_27296,N_23306,N_24825);
nand U27297 (N_27297,N_22152,N_22099);
or U27298 (N_27298,N_21488,N_20063);
nand U27299 (N_27299,N_22624,N_23604);
and U27300 (N_27300,N_22527,N_20256);
nand U27301 (N_27301,N_21497,N_24454);
xnor U27302 (N_27302,N_24298,N_23709);
or U27303 (N_27303,N_24470,N_22765);
nand U27304 (N_27304,N_21659,N_20125);
nand U27305 (N_27305,N_24192,N_20599);
xor U27306 (N_27306,N_21831,N_23196);
xnor U27307 (N_27307,N_24130,N_24944);
or U27308 (N_27308,N_20442,N_23056);
or U27309 (N_27309,N_23219,N_21145);
xnor U27310 (N_27310,N_23017,N_22644);
and U27311 (N_27311,N_20970,N_20609);
or U27312 (N_27312,N_22827,N_21598);
and U27313 (N_27313,N_21825,N_21475);
or U27314 (N_27314,N_23338,N_24161);
or U27315 (N_27315,N_23514,N_23994);
nand U27316 (N_27316,N_24064,N_24863);
nand U27317 (N_27317,N_20939,N_23283);
nor U27318 (N_27318,N_22980,N_23773);
nor U27319 (N_27319,N_20563,N_23300);
nand U27320 (N_27320,N_24234,N_24873);
or U27321 (N_27321,N_20458,N_24321);
nor U27322 (N_27322,N_24019,N_24171);
and U27323 (N_27323,N_21266,N_23521);
or U27324 (N_27324,N_22060,N_22939);
and U27325 (N_27325,N_21756,N_20911);
nor U27326 (N_27326,N_21548,N_21200);
and U27327 (N_27327,N_22433,N_22331);
or U27328 (N_27328,N_22398,N_21432);
xor U27329 (N_27329,N_21952,N_24721);
nor U27330 (N_27330,N_22606,N_21863);
and U27331 (N_27331,N_24966,N_23879);
or U27332 (N_27332,N_21716,N_21484);
or U27333 (N_27333,N_24504,N_24516);
xnor U27334 (N_27334,N_23173,N_24022);
nand U27335 (N_27335,N_22742,N_24882);
and U27336 (N_27336,N_24673,N_24517);
xor U27337 (N_27337,N_20506,N_23984);
nand U27338 (N_27338,N_24146,N_22739);
and U27339 (N_27339,N_23748,N_22729);
nor U27340 (N_27340,N_21868,N_20841);
xor U27341 (N_27341,N_24222,N_24708);
nor U27342 (N_27342,N_23611,N_24020);
and U27343 (N_27343,N_23945,N_22478);
xor U27344 (N_27344,N_23318,N_22860);
xnor U27345 (N_27345,N_20274,N_23561);
xor U27346 (N_27346,N_23326,N_20461);
nand U27347 (N_27347,N_22081,N_21127);
nand U27348 (N_27348,N_24785,N_24391);
xnor U27349 (N_27349,N_22308,N_24312);
nand U27350 (N_27350,N_23023,N_21757);
or U27351 (N_27351,N_24170,N_24240);
and U27352 (N_27352,N_22412,N_20846);
or U27353 (N_27353,N_23821,N_23841);
nor U27354 (N_27354,N_24588,N_23800);
or U27355 (N_27355,N_20588,N_20087);
and U27356 (N_27356,N_24509,N_21139);
and U27357 (N_27357,N_24143,N_20987);
nor U27358 (N_27358,N_21744,N_20348);
and U27359 (N_27359,N_20895,N_20251);
nand U27360 (N_27360,N_24124,N_21854);
nand U27361 (N_27361,N_22375,N_22069);
and U27362 (N_27362,N_24650,N_21658);
and U27363 (N_27363,N_21472,N_24655);
nor U27364 (N_27364,N_21439,N_23646);
and U27365 (N_27365,N_20666,N_20711);
nand U27366 (N_27366,N_24154,N_22091);
and U27367 (N_27367,N_21570,N_24169);
xor U27368 (N_27368,N_24821,N_21183);
nor U27369 (N_27369,N_23217,N_23025);
nand U27370 (N_27370,N_20049,N_24157);
and U27371 (N_27371,N_22246,N_22972);
nor U27372 (N_27372,N_20963,N_22853);
nor U27373 (N_27373,N_22502,N_24851);
nand U27374 (N_27374,N_20243,N_22544);
nor U27375 (N_27375,N_21515,N_24659);
xnor U27376 (N_27376,N_20787,N_20023);
nand U27377 (N_27377,N_20937,N_23664);
nand U27378 (N_27378,N_21866,N_20495);
nand U27379 (N_27379,N_24221,N_24452);
and U27380 (N_27380,N_21967,N_22456);
or U27381 (N_27381,N_20594,N_23477);
and U27382 (N_27382,N_23606,N_21931);
nand U27383 (N_27383,N_20224,N_23297);
nand U27384 (N_27384,N_23582,N_20370);
nand U27385 (N_27385,N_22253,N_21326);
xnor U27386 (N_27386,N_23443,N_22192);
nand U27387 (N_27387,N_23131,N_24434);
and U27388 (N_27388,N_23463,N_22383);
xnor U27389 (N_27389,N_24711,N_24375);
xor U27390 (N_27390,N_21236,N_24743);
and U27391 (N_27391,N_20766,N_21732);
and U27392 (N_27392,N_21865,N_24247);
xnor U27393 (N_27393,N_24581,N_24911);
xor U27394 (N_27394,N_23586,N_24807);
xor U27395 (N_27395,N_23924,N_22292);
xnor U27396 (N_27396,N_20560,N_20121);
or U27397 (N_27397,N_20474,N_23069);
nand U27398 (N_27398,N_21113,N_24740);
nand U27399 (N_27399,N_20219,N_24636);
xnor U27400 (N_27400,N_22396,N_22314);
and U27401 (N_27401,N_23065,N_20155);
nor U27402 (N_27402,N_23389,N_20884);
nand U27403 (N_27403,N_23332,N_23803);
and U27404 (N_27404,N_22636,N_24087);
nor U27405 (N_27405,N_24562,N_23014);
nand U27406 (N_27406,N_21435,N_24335);
or U27407 (N_27407,N_23822,N_23878);
nand U27408 (N_27408,N_21563,N_24980);
nor U27409 (N_27409,N_20984,N_20231);
nor U27410 (N_27410,N_20546,N_24916);
and U27411 (N_27411,N_21328,N_21135);
nor U27412 (N_27412,N_22166,N_22686);
nand U27413 (N_27413,N_22284,N_20647);
xor U27414 (N_27414,N_22511,N_22885);
nand U27415 (N_27415,N_21117,N_23107);
xor U27416 (N_27416,N_23125,N_24059);
xnor U27417 (N_27417,N_20974,N_24126);
and U27418 (N_27418,N_24428,N_22647);
or U27419 (N_27419,N_23986,N_20180);
nor U27420 (N_27420,N_24508,N_20124);
and U27421 (N_27421,N_20033,N_22414);
xnor U27422 (N_27422,N_22935,N_24527);
or U27423 (N_27423,N_20191,N_22465);
and U27424 (N_27424,N_24724,N_21211);
xnor U27425 (N_27425,N_20479,N_23044);
nor U27426 (N_27426,N_20245,N_23224);
and U27427 (N_27427,N_21089,N_21743);
or U27428 (N_27428,N_22629,N_22034);
and U27429 (N_27429,N_20537,N_20284);
nand U27430 (N_27430,N_24981,N_23193);
or U27431 (N_27431,N_20527,N_23156);
or U27432 (N_27432,N_20519,N_21248);
nor U27433 (N_27433,N_22075,N_24128);
nand U27434 (N_27434,N_23164,N_21321);
xor U27435 (N_27435,N_24164,N_23043);
nand U27436 (N_27436,N_24657,N_22015);
or U27437 (N_27437,N_23322,N_21588);
nand U27438 (N_27438,N_24692,N_24917);
or U27439 (N_27439,N_23078,N_22128);
nor U27440 (N_27440,N_24289,N_20406);
nand U27441 (N_27441,N_22301,N_23486);
and U27442 (N_27442,N_23995,N_22996);
nand U27443 (N_27443,N_20280,N_21849);
nand U27444 (N_27444,N_21827,N_23594);
nor U27445 (N_27445,N_24048,N_23433);
nor U27446 (N_27446,N_20004,N_20485);
and U27447 (N_27447,N_22558,N_21700);
nand U27448 (N_27448,N_22945,N_22684);
and U27449 (N_27449,N_20998,N_23669);
xor U27450 (N_27450,N_22032,N_24961);
or U27451 (N_27451,N_23820,N_20346);
xor U27452 (N_27452,N_22489,N_21961);
xor U27453 (N_27453,N_22625,N_22096);
xnor U27454 (N_27454,N_23123,N_24718);
and U27455 (N_27455,N_21837,N_22353);
xnor U27456 (N_27456,N_24874,N_20776);
and U27457 (N_27457,N_23174,N_21492);
nand U27458 (N_27458,N_24481,N_22269);
and U27459 (N_27459,N_20128,N_21305);
and U27460 (N_27460,N_24772,N_22592);
xor U27461 (N_27461,N_24576,N_24197);
xor U27462 (N_27462,N_24446,N_20985);
and U27463 (N_27463,N_23981,N_23439);
or U27464 (N_27464,N_24029,N_22004);
or U27465 (N_27465,N_23476,N_23000);
and U27466 (N_27466,N_20680,N_23534);
nand U27467 (N_27467,N_24680,N_24437);
or U27468 (N_27468,N_20956,N_23061);
and U27469 (N_27469,N_23408,N_22055);
or U27470 (N_27470,N_24866,N_23177);
xnor U27471 (N_27471,N_23470,N_24573);
and U27472 (N_27472,N_22837,N_23633);
or U27473 (N_27473,N_23982,N_23458);
nor U27474 (N_27474,N_21558,N_20258);
or U27475 (N_27475,N_21357,N_22036);
nand U27476 (N_27476,N_22437,N_23266);
and U27477 (N_27477,N_21377,N_23315);
nor U27478 (N_27478,N_21527,N_21005);
nor U27479 (N_27479,N_24971,N_23765);
xnor U27480 (N_27480,N_23729,N_20135);
nor U27481 (N_27481,N_24346,N_22725);
nor U27482 (N_27482,N_21020,N_24880);
nor U27483 (N_27483,N_23760,N_22484);
or U27484 (N_27484,N_24703,N_23335);
nand U27485 (N_27485,N_24594,N_22195);
nor U27486 (N_27486,N_23162,N_22904);
and U27487 (N_27487,N_21502,N_22227);
nor U27488 (N_27488,N_22162,N_22423);
nor U27489 (N_27489,N_20796,N_20649);
nor U27490 (N_27490,N_20294,N_22975);
nand U27491 (N_27491,N_20048,N_20824);
nor U27492 (N_27492,N_22760,N_20717);
and U27493 (N_27493,N_23769,N_20291);
nand U27494 (N_27494,N_20190,N_21670);
xor U27495 (N_27495,N_24559,N_21190);
and U27496 (N_27496,N_22222,N_22737);
or U27497 (N_27497,N_24237,N_21697);
xor U27498 (N_27498,N_24176,N_21629);
xor U27499 (N_27499,N_24478,N_22762);
and U27500 (N_27500,N_21975,N_21267);
xnor U27501 (N_27501,N_21964,N_20056);
and U27502 (N_27502,N_23516,N_21419);
nand U27503 (N_27503,N_22726,N_22612);
xor U27504 (N_27504,N_22282,N_23979);
and U27505 (N_27505,N_23969,N_23444);
and U27506 (N_27506,N_21443,N_24836);
or U27507 (N_27507,N_21998,N_22405);
nand U27508 (N_27508,N_23058,N_24476);
nor U27509 (N_27509,N_20375,N_21265);
nor U27510 (N_27510,N_23661,N_22618);
or U27511 (N_27511,N_23556,N_21578);
nor U27512 (N_27512,N_21462,N_21472);
nand U27513 (N_27513,N_23710,N_22622);
and U27514 (N_27514,N_24919,N_21523);
or U27515 (N_27515,N_20206,N_21555);
nor U27516 (N_27516,N_23070,N_23565);
xor U27517 (N_27517,N_24540,N_24622);
nand U27518 (N_27518,N_20365,N_21797);
xor U27519 (N_27519,N_24772,N_20192);
and U27520 (N_27520,N_22322,N_21602);
nand U27521 (N_27521,N_24796,N_23429);
and U27522 (N_27522,N_23747,N_23461);
and U27523 (N_27523,N_23131,N_23242);
nor U27524 (N_27524,N_20670,N_21805);
and U27525 (N_27525,N_21439,N_23957);
and U27526 (N_27526,N_22863,N_20762);
nor U27527 (N_27527,N_22129,N_23538);
or U27528 (N_27528,N_22721,N_21792);
or U27529 (N_27529,N_24084,N_21298);
and U27530 (N_27530,N_21105,N_24983);
nand U27531 (N_27531,N_22312,N_22375);
xnor U27532 (N_27532,N_24724,N_23582);
or U27533 (N_27533,N_21261,N_21626);
nor U27534 (N_27534,N_23147,N_24417);
or U27535 (N_27535,N_21687,N_23145);
nand U27536 (N_27536,N_21285,N_23707);
nor U27537 (N_27537,N_23981,N_21077);
xnor U27538 (N_27538,N_21947,N_24724);
nand U27539 (N_27539,N_20211,N_24635);
xnor U27540 (N_27540,N_22159,N_23241);
and U27541 (N_27541,N_23478,N_20668);
or U27542 (N_27542,N_20774,N_23395);
nand U27543 (N_27543,N_20388,N_22012);
xor U27544 (N_27544,N_23607,N_20448);
xor U27545 (N_27545,N_20184,N_24403);
xnor U27546 (N_27546,N_21515,N_23598);
or U27547 (N_27547,N_21642,N_21673);
or U27548 (N_27548,N_22595,N_21696);
and U27549 (N_27549,N_20860,N_20674);
or U27550 (N_27550,N_24894,N_24792);
nand U27551 (N_27551,N_23705,N_21434);
nor U27552 (N_27552,N_24185,N_24334);
xnor U27553 (N_27553,N_24558,N_22972);
nand U27554 (N_27554,N_24814,N_22002);
nor U27555 (N_27555,N_23990,N_22844);
and U27556 (N_27556,N_20911,N_20255);
nand U27557 (N_27557,N_24312,N_22796);
xnor U27558 (N_27558,N_23284,N_24983);
or U27559 (N_27559,N_23894,N_23258);
nor U27560 (N_27560,N_24775,N_23925);
and U27561 (N_27561,N_24627,N_24784);
or U27562 (N_27562,N_21413,N_20438);
nand U27563 (N_27563,N_23199,N_22954);
xnor U27564 (N_27564,N_20226,N_20029);
nand U27565 (N_27565,N_20352,N_24429);
and U27566 (N_27566,N_21915,N_20006);
and U27567 (N_27567,N_24732,N_22293);
xnor U27568 (N_27568,N_22942,N_24749);
nor U27569 (N_27569,N_21155,N_23377);
or U27570 (N_27570,N_21202,N_20904);
nor U27571 (N_27571,N_22371,N_23268);
and U27572 (N_27572,N_23876,N_22382);
xor U27573 (N_27573,N_24565,N_23074);
or U27574 (N_27574,N_22536,N_22010);
nand U27575 (N_27575,N_24743,N_23629);
nor U27576 (N_27576,N_20380,N_23397);
and U27577 (N_27577,N_21762,N_21459);
nand U27578 (N_27578,N_22969,N_24226);
and U27579 (N_27579,N_23235,N_20548);
xor U27580 (N_27580,N_22378,N_20272);
nor U27581 (N_27581,N_21338,N_20983);
or U27582 (N_27582,N_21117,N_24752);
xor U27583 (N_27583,N_21651,N_23583);
and U27584 (N_27584,N_21584,N_20572);
and U27585 (N_27585,N_24022,N_24839);
xor U27586 (N_27586,N_20731,N_20433);
nand U27587 (N_27587,N_22256,N_22862);
nand U27588 (N_27588,N_23401,N_20452);
xnor U27589 (N_27589,N_22636,N_23647);
nor U27590 (N_27590,N_22499,N_23145);
and U27591 (N_27591,N_24856,N_21997);
nor U27592 (N_27592,N_22651,N_21882);
nor U27593 (N_27593,N_24434,N_21913);
xnor U27594 (N_27594,N_21212,N_22047);
nor U27595 (N_27595,N_21703,N_23621);
nor U27596 (N_27596,N_21588,N_22091);
nor U27597 (N_27597,N_24146,N_23002);
nand U27598 (N_27598,N_24926,N_24638);
or U27599 (N_27599,N_20902,N_20111);
or U27600 (N_27600,N_24023,N_20506);
nor U27601 (N_27601,N_20685,N_20462);
xnor U27602 (N_27602,N_24407,N_23891);
nor U27603 (N_27603,N_24164,N_21472);
and U27604 (N_27604,N_24197,N_20781);
xor U27605 (N_27605,N_24595,N_21944);
nand U27606 (N_27606,N_23028,N_21488);
nor U27607 (N_27607,N_24558,N_24608);
and U27608 (N_27608,N_22505,N_22154);
nor U27609 (N_27609,N_24834,N_21442);
nand U27610 (N_27610,N_24857,N_24417);
xnor U27611 (N_27611,N_21570,N_24558);
or U27612 (N_27612,N_22234,N_20051);
nand U27613 (N_27613,N_20372,N_22764);
xnor U27614 (N_27614,N_23636,N_21261);
xnor U27615 (N_27615,N_22047,N_21448);
nand U27616 (N_27616,N_21563,N_22744);
nor U27617 (N_27617,N_22779,N_21994);
nor U27618 (N_27618,N_22468,N_23077);
nand U27619 (N_27619,N_23027,N_22313);
nand U27620 (N_27620,N_23810,N_24562);
nand U27621 (N_27621,N_22089,N_23209);
or U27622 (N_27622,N_20629,N_20146);
and U27623 (N_27623,N_24558,N_21128);
or U27624 (N_27624,N_22503,N_20058);
and U27625 (N_27625,N_24314,N_24829);
or U27626 (N_27626,N_20067,N_20488);
xnor U27627 (N_27627,N_24073,N_23910);
and U27628 (N_27628,N_23423,N_20836);
nor U27629 (N_27629,N_22288,N_22665);
nand U27630 (N_27630,N_23842,N_24662);
xor U27631 (N_27631,N_23100,N_22738);
and U27632 (N_27632,N_22291,N_24485);
and U27633 (N_27633,N_21994,N_23099);
nor U27634 (N_27634,N_22659,N_22336);
xnor U27635 (N_27635,N_21936,N_22170);
xnor U27636 (N_27636,N_23665,N_24311);
nand U27637 (N_27637,N_24571,N_23101);
or U27638 (N_27638,N_24931,N_23559);
and U27639 (N_27639,N_22542,N_22479);
nand U27640 (N_27640,N_22514,N_21503);
nand U27641 (N_27641,N_23215,N_20105);
and U27642 (N_27642,N_23305,N_21656);
and U27643 (N_27643,N_20018,N_21110);
nand U27644 (N_27644,N_23391,N_23617);
xor U27645 (N_27645,N_20167,N_22528);
nand U27646 (N_27646,N_21891,N_22918);
nor U27647 (N_27647,N_20094,N_20082);
xor U27648 (N_27648,N_20367,N_21330);
xnor U27649 (N_27649,N_20366,N_24507);
and U27650 (N_27650,N_24152,N_20578);
xnor U27651 (N_27651,N_23364,N_21316);
nor U27652 (N_27652,N_21887,N_24255);
nand U27653 (N_27653,N_21911,N_22906);
xnor U27654 (N_27654,N_22940,N_24837);
or U27655 (N_27655,N_23586,N_23054);
nor U27656 (N_27656,N_22094,N_21942);
or U27657 (N_27657,N_20277,N_21351);
nand U27658 (N_27658,N_23387,N_21476);
xnor U27659 (N_27659,N_22158,N_24346);
or U27660 (N_27660,N_21571,N_20082);
nor U27661 (N_27661,N_24544,N_23897);
nand U27662 (N_27662,N_20046,N_20514);
or U27663 (N_27663,N_24847,N_20436);
and U27664 (N_27664,N_24306,N_23618);
xor U27665 (N_27665,N_22638,N_24913);
nand U27666 (N_27666,N_20915,N_24440);
nand U27667 (N_27667,N_21458,N_20588);
nor U27668 (N_27668,N_24190,N_23212);
nand U27669 (N_27669,N_23178,N_24756);
or U27670 (N_27670,N_24745,N_20126);
nand U27671 (N_27671,N_22672,N_20024);
and U27672 (N_27672,N_20904,N_24162);
nand U27673 (N_27673,N_22809,N_24911);
nor U27674 (N_27674,N_21812,N_23715);
xor U27675 (N_27675,N_21388,N_23990);
xor U27676 (N_27676,N_21092,N_21217);
and U27677 (N_27677,N_20350,N_23529);
xor U27678 (N_27678,N_20247,N_21494);
or U27679 (N_27679,N_22333,N_24025);
or U27680 (N_27680,N_22929,N_23600);
xor U27681 (N_27681,N_23645,N_21598);
nand U27682 (N_27682,N_20470,N_24376);
xor U27683 (N_27683,N_22226,N_24110);
and U27684 (N_27684,N_24479,N_20695);
or U27685 (N_27685,N_21414,N_21889);
nand U27686 (N_27686,N_22237,N_24031);
nor U27687 (N_27687,N_23522,N_20301);
nor U27688 (N_27688,N_20383,N_22069);
nand U27689 (N_27689,N_22740,N_20577);
nand U27690 (N_27690,N_22076,N_23126);
xor U27691 (N_27691,N_22257,N_21277);
and U27692 (N_27692,N_21401,N_22936);
xnor U27693 (N_27693,N_21109,N_23737);
nor U27694 (N_27694,N_23840,N_22503);
nor U27695 (N_27695,N_23849,N_22239);
xnor U27696 (N_27696,N_23040,N_22888);
xor U27697 (N_27697,N_23191,N_22599);
nand U27698 (N_27698,N_23559,N_20817);
nor U27699 (N_27699,N_22258,N_22749);
nand U27700 (N_27700,N_23232,N_24567);
and U27701 (N_27701,N_20565,N_22088);
or U27702 (N_27702,N_24478,N_22703);
nor U27703 (N_27703,N_22299,N_22808);
nand U27704 (N_27704,N_22196,N_24648);
xor U27705 (N_27705,N_21651,N_24450);
and U27706 (N_27706,N_20193,N_24564);
or U27707 (N_27707,N_22960,N_22291);
xor U27708 (N_27708,N_24613,N_21411);
nor U27709 (N_27709,N_22557,N_21376);
xor U27710 (N_27710,N_22758,N_21343);
xor U27711 (N_27711,N_23303,N_20131);
nand U27712 (N_27712,N_20193,N_23707);
xor U27713 (N_27713,N_24682,N_21277);
nand U27714 (N_27714,N_22883,N_23147);
nor U27715 (N_27715,N_21409,N_22349);
xor U27716 (N_27716,N_20169,N_24247);
nor U27717 (N_27717,N_24290,N_23317);
or U27718 (N_27718,N_21350,N_21481);
xor U27719 (N_27719,N_20074,N_22420);
xor U27720 (N_27720,N_22088,N_21426);
xnor U27721 (N_27721,N_22879,N_23083);
xor U27722 (N_27722,N_21478,N_23268);
xor U27723 (N_27723,N_22961,N_20188);
or U27724 (N_27724,N_20121,N_21109);
or U27725 (N_27725,N_21782,N_23412);
xor U27726 (N_27726,N_22396,N_21011);
and U27727 (N_27727,N_24895,N_21228);
xnor U27728 (N_27728,N_23752,N_22590);
or U27729 (N_27729,N_22927,N_22783);
and U27730 (N_27730,N_20103,N_20267);
and U27731 (N_27731,N_22131,N_22900);
xnor U27732 (N_27732,N_22654,N_22034);
xnor U27733 (N_27733,N_24434,N_24401);
nor U27734 (N_27734,N_23710,N_21848);
or U27735 (N_27735,N_22123,N_24153);
or U27736 (N_27736,N_22990,N_24789);
nand U27737 (N_27737,N_20582,N_23882);
xnor U27738 (N_27738,N_21181,N_24168);
xnor U27739 (N_27739,N_21476,N_24905);
nand U27740 (N_27740,N_23227,N_20058);
or U27741 (N_27741,N_21393,N_23344);
nor U27742 (N_27742,N_23417,N_21096);
and U27743 (N_27743,N_24437,N_20313);
nor U27744 (N_27744,N_20939,N_23048);
xnor U27745 (N_27745,N_23641,N_20584);
nor U27746 (N_27746,N_23569,N_23093);
nand U27747 (N_27747,N_22873,N_20568);
nor U27748 (N_27748,N_24459,N_24343);
nand U27749 (N_27749,N_24134,N_20800);
xnor U27750 (N_27750,N_23923,N_21951);
xor U27751 (N_27751,N_24034,N_24932);
nand U27752 (N_27752,N_21230,N_22968);
nand U27753 (N_27753,N_24190,N_23835);
or U27754 (N_27754,N_23840,N_23940);
or U27755 (N_27755,N_24877,N_22268);
nand U27756 (N_27756,N_21122,N_24092);
or U27757 (N_27757,N_24737,N_23310);
xnor U27758 (N_27758,N_24493,N_20767);
or U27759 (N_27759,N_24916,N_24010);
nor U27760 (N_27760,N_24910,N_22281);
nand U27761 (N_27761,N_22149,N_22933);
nor U27762 (N_27762,N_20036,N_22167);
xor U27763 (N_27763,N_20182,N_22523);
nand U27764 (N_27764,N_24665,N_23189);
and U27765 (N_27765,N_24112,N_21294);
nor U27766 (N_27766,N_24946,N_22571);
or U27767 (N_27767,N_20445,N_22854);
and U27768 (N_27768,N_20725,N_22934);
and U27769 (N_27769,N_21307,N_21048);
nor U27770 (N_27770,N_22217,N_23994);
xnor U27771 (N_27771,N_20028,N_22503);
or U27772 (N_27772,N_24477,N_20680);
xor U27773 (N_27773,N_22724,N_20078);
or U27774 (N_27774,N_23751,N_21047);
nor U27775 (N_27775,N_23351,N_24015);
and U27776 (N_27776,N_24928,N_22647);
nand U27777 (N_27777,N_21873,N_21910);
or U27778 (N_27778,N_24178,N_24032);
xnor U27779 (N_27779,N_23478,N_24254);
nand U27780 (N_27780,N_20035,N_21201);
xor U27781 (N_27781,N_24042,N_21958);
nand U27782 (N_27782,N_20691,N_21595);
or U27783 (N_27783,N_20144,N_20167);
and U27784 (N_27784,N_20693,N_21051);
and U27785 (N_27785,N_20565,N_24539);
nor U27786 (N_27786,N_20977,N_21378);
and U27787 (N_27787,N_23712,N_24027);
nand U27788 (N_27788,N_21558,N_20154);
and U27789 (N_27789,N_23523,N_23163);
and U27790 (N_27790,N_22701,N_23191);
nor U27791 (N_27791,N_21203,N_21688);
or U27792 (N_27792,N_21693,N_21077);
xor U27793 (N_27793,N_24545,N_23235);
nand U27794 (N_27794,N_23196,N_24549);
nand U27795 (N_27795,N_20107,N_20405);
nor U27796 (N_27796,N_21550,N_24742);
nor U27797 (N_27797,N_21686,N_21337);
nand U27798 (N_27798,N_22049,N_24934);
or U27799 (N_27799,N_21030,N_24444);
or U27800 (N_27800,N_21555,N_22632);
nand U27801 (N_27801,N_20555,N_20282);
and U27802 (N_27802,N_24530,N_20660);
nand U27803 (N_27803,N_23704,N_21536);
nor U27804 (N_27804,N_22556,N_23060);
nand U27805 (N_27805,N_20273,N_22388);
or U27806 (N_27806,N_22840,N_21862);
xnor U27807 (N_27807,N_22849,N_22990);
and U27808 (N_27808,N_21044,N_23085);
or U27809 (N_27809,N_24143,N_23196);
nand U27810 (N_27810,N_24152,N_20105);
nand U27811 (N_27811,N_23674,N_23912);
and U27812 (N_27812,N_21831,N_24701);
nand U27813 (N_27813,N_20211,N_20711);
xor U27814 (N_27814,N_20026,N_22806);
nor U27815 (N_27815,N_22724,N_20928);
nor U27816 (N_27816,N_21749,N_22493);
xor U27817 (N_27817,N_24048,N_20348);
nor U27818 (N_27818,N_22357,N_24639);
nand U27819 (N_27819,N_20397,N_24981);
or U27820 (N_27820,N_20377,N_20102);
and U27821 (N_27821,N_23037,N_23136);
and U27822 (N_27822,N_21276,N_23443);
and U27823 (N_27823,N_24220,N_22079);
or U27824 (N_27824,N_21209,N_20797);
xnor U27825 (N_27825,N_20241,N_22971);
and U27826 (N_27826,N_24948,N_20413);
nand U27827 (N_27827,N_21256,N_24001);
and U27828 (N_27828,N_21098,N_20011);
xnor U27829 (N_27829,N_22632,N_20340);
and U27830 (N_27830,N_21575,N_20195);
nor U27831 (N_27831,N_21856,N_24631);
or U27832 (N_27832,N_22356,N_23254);
or U27833 (N_27833,N_23102,N_22886);
and U27834 (N_27834,N_20683,N_21711);
nor U27835 (N_27835,N_20651,N_21016);
nor U27836 (N_27836,N_22548,N_24091);
and U27837 (N_27837,N_24592,N_21222);
and U27838 (N_27838,N_24995,N_20231);
and U27839 (N_27839,N_24525,N_20278);
and U27840 (N_27840,N_20224,N_21748);
xnor U27841 (N_27841,N_22235,N_21510);
xnor U27842 (N_27842,N_22893,N_23845);
and U27843 (N_27843,N_22974,N_20274);
nand U27844 (N_27844,N_23130,N_23844);
or U27845 (N_27845,N_23834,N_23572);
nor U27846 (N_27846,N_24277,N_23555);
xnor U27847 (N_27847,N_22099,N_21208);
and U27848 (N_27848,N_23192,N_24397);
or U27849 (N_27849,N_21808,N_22002);
nand U27850 (N_27850,N_24379,N_22555);
nor U27851 (N_27851,N_23798,N_22973);
or U27852 (N_27852,N_23048,N_24091);
xnor U27853 (N_27853,N_23963,N_20138);
or U27854 (N_27854,N_20745,N_21731);
nand U27855 (N_27855,N_22813,N_20505);
or U27856 (N_27856,N_20214,N_24479);
nor U27857 (N_27857,N_21014,N_24616);
nor U27858 (N_27858,N_20461,N_24894);
nand U27859 (N_27859,N_23325,N_23860);
nand U27860 (N_27860,N_24698,N_23496);
xnor U27861 (N_27861,N_21940,N_21953);
xnor U27862 (N_27862,N_24583,N_22566);
nand U27863 (N_27863,N_20561,N_20973);
xor U27864 (N_27864,N_24305,N_23526);
and U27865 (N_27865,N_20036,N_24586);
and U27866 (N_27866,N_22825,N_21312);
nor U27867 (N_27867,N_20997,N_21137);
nand U27868 (N_27868,N_21336,N_21615);
nor U27869 (N_27869,N_23525,N_21426);
or U27870 (N_27870,N_23530,N_23221);
xnor U27871 (N_27871,N_23048,N_23783);
and U27872 (N_27872,N_22555,N_22707);
and U27873 (N_27873,N_22633,N_24420);
and U27874 (N_27874,N_22129,N_22309);
nor U27875 (N_27875,N_23182,N_21800);
nand U27876 (N_27876,N_20583,N_21856);
nand U27877 (N_27877,N_20671,N_20714);
or U27878 (N_27878,N_20789,N_20005);
nor U27879 (N_27879,N_23578,N_24033);
and U27880 (N_27880,N_22211,N_23810);
nand U27881 (N_27881,N_20012,N_21471);
xor U27882 (N_27882,N_23725,N_24364);
nand U27883 (N_27883,N_20300,N_23785);
nand U27884 (N_27884,N_24593,N_22465);
and U27885 (N_27885,N_22022,N_22274);
nand U27886 (N_27886,N_20995,N_24415);
and U27887 (N_27887,N_24791,N_23031);
or U27888 (N_27888,N_22551,N_23239);
nand U27889 (N_27889,N_21257,N_23019);
nand U27890 (N_27890,N_21821,N_22413);
nor U27891 (N_27891,N_21774,N_21666);
nand U27892 (N_27892,N_24135,N_23548);
or U27893 (N_27893,N_20538,N_24264);
nor U27894 (N_27894,N_22976,N_24688);
xor U27895 (N_27895,N_23288,N_21038);
and U27896 (N_27896,N_23750,N_21543);
xor U27897 (N_27897,N_22311,N_23123);
and U27898 (N_27898,N_24944,N_22858);
or U27899 (N_27899,N_24861,N_22686);
nor U27900 (N_27900,N_21434,N_24510);
or U27901 (N_27901,N_22941,N_20237);
and U27902 (N_27902,N_20828,N_24474);
or U27903 (N_27903,N_22550,N_24224);
xnor U27904 (N_27904,N_23978,N_23496);
nor U27905 (N_27905,N_22195,N_23810);
or U27906 (N_27906,N_23857,N_24267);
xnor U27907 (N_27907,N_21750,N_23223);
nor U27908 (N_27908,N_20362,N_20580);
or U27909 (N_27909,N_20252,N_22107);
or U27910 (N_27910,N_24613,N_22757);
or U27911 (N_27911,N_21310,N_20437);
xnor U27912 (N_27912,N_24639,N_24918);
nor U27913 (N_27913,N_20863,N_20077);
nand U27914 (N_27914,N_21038,N_21845);
and U27915 (N_27915,N_23987,N_22519);
and U27916 (N_27916,N_21169,N_23861);
and U27917 (N_27917,N_24708,N_23676);
and U27918 (N_27918,N_24480,N_22115);
nor U27919 (N_27919,N_23964,N_21018);
or U27920 (N_27920,N_23973,N_21947);
nor U27921 (N_27921,N_24267,N_23696);
nand U27922 (N_27922,N_21686,N_20382);
nor U27923 (N_27923,N_21876,N_20840);
xnor U27924 (N_27924,N_24827,N_24489);
and U27925 (N_27925,N_20568,N_21265);
nor U27926 (N_27926,N_22444,N_22750);
and U27927 (N_27927,N_22674,N_22469);
or U27928 (N_27928,N_24662,N_20300);
xor U27929 (N_27929,N_21688,N_21633);
nand U27930 (N_27930,N_20149,N_22043);
nand U27931 (N_27931,N_22930,N_20217);
or U27932 (N_27932,N_21554,N_20199);
or U27933 (N_27933,N_22476,N_24114);
or U27934 (N_27934,N_24958,N_20080);
xor U27935 (N_27935,N_23268,N_21076);
nand U27936 (N_27936,N_24139,N_23673);
nor U27937 (N_27937,N_20575,N_22533);
or U27938 (N_27938,N_20066,N_22134);
or U27939 (N_27939,N_23127,N_22025);
and U27940 (N_27940,N_24361,N_23168);
xor U27941 (N_27941,N_21933,N_22355);
xnor U27942 (N_27942,N_20082,N_20939);
xor U27943 (N_27943,N_23076,N_21037);
nor U27944 (N_27944,N_21647,N_24543);
nor U27945 (N_27945,N_24152,N_21236);
xnor U27946 (N_27946,N_21719,N_24856);
or U27947 (N_27947,N_20408,N_24956);
or U27948 (N_27948,N_21806,N_24687);
and U27949 (N_27949,N_22054,N_24041);
nand U27950 (N_27950,N_24155,N_20976);
nor U27951 (N_27951,N_21878,N_23448);
or U27952 (N_27952,N_20880,N_24494);
nor U27953 (N_27953,N_22941,N_22754);
xor U27954 (N_27954,N_20045,N_22440);
or U27955 (N_27955,N_24277,N_24495);
xnor U27956 (N_27956,N_24721,N_23602);
nand U27957 (N_27957,N_24403,N_21716);
and U27958 (N_27958,N_21585,N_20417);
xnor U27959 (N_27959,N_24571,N_20103);
nand U27960 (N_27960,N_24196,N_21283);
nand U27961 (N_27961,N_20630,N_21869);
nand U27962 (N_27962,N_24763,N_22698);
and U27963 (N_27963,N_20957,N_24773);
nor U27964 (N_27964,N_24052,N_24084);
nor U27965 (N_27965,N_23043,N_23088);
xor U27966 (N_27966,N_22565,N_22355);
and U27967 (N_27967,N_22883,N_23707);
or U27968 (N_27968,N_20543,N_22533);
nor U27969 (N_27969,N_21678,N_23968);
nor U27970 (N_27970,N_21264,N_24843);
nand U27971 (N_27971,N_23099,N_22731);
and U27972 (N_27972,N_23930,N_24837);
or U27973 (N_27973,N_20092,N_21149);
nand U27974 (N_27974,N_21570,N_22409);
nand U27975 (N_27975,N_24491,N_20590);
and U27976 (N_27976,N_23008,N_22565);
xor U27977 (N_27977,N_22217,N_22948);
nand U27978 (N_27978,N_20228,N_24220);
and U27979 (N_27979,N_24731,N_23790);
or U27980 (N_27980,N_21833,N_24620);
nand U27981 (N_27981,N_21122,N_22983);
or U27982 (N_27982,N_20908,N_23124);
and U27983 (N_27983,N_24103,N_20937);
xnor U27984 (N_27984,N_20097,N_23170);
and U27985 (N_27985,N_24855,N_20976);
nor U27986 (N_27986,N_21588,N_21444);
or U27987 (N_27987,N_24534,N_21726);
xor U27988 (N_27988,N_21313,N_21941);
nor U27989 (N_27989,N_20509,N_24944);
nand U27990 (N_27990,N_20813,N_23515);
nand U27991 (N_27991,N_24675,N_21435);
and U27992 (N_27992,N_20389,N_20404);
xnor U27993 (N_27993,N_21728,N_21246);
nor U27994 (N_27994,N_22320,N_24941);
or U27995 (N_27995,N_24355,N_22753);
nand U27996 (N_27996,N_24043,N_21715);
or U27997 (N_27997,N_24904,N_21030);
nor U27998 (N_27998,N_24254,N_20764);
or U27999 (N_27999,N_20674,N_22255);
xnor U28000 (N_28000,N_21733,N_24634);
or U28001 (N_28001,N_23418,N_21957);
nand U28002 (N_28002,N_24013,N_21072);
xnor U28003 (N_28003,N_22661,N_24626);
nor U28004 (N_28004,N_22747,N_22760);
nand U28005 (N_28005,N_22584,N_21591);
nor U28006 (N_28006,N_22237,N_21589);
or U28007 (N_28007,N_23873,N_21095);
nand U28008 (N_28008,N_24982,N_20639);
and U28009 (N_28009,N_23014,N_23481);
or U28010 (N_28010,N_20949,N_21776);
nor U28011 (N_28011,N_21611,N_24934);
nor U28012 (N_28012,N_20311,N_21399);
xnor U28013 (N_28013,N_22716,N_20097);
xnor U28014 (N_28014,N_22942,N_21246);
or U28015 (N_28015,N_24023,N_23922);
nand U28016 (N_28016,N_23140,N_22666);
xor U28017 (N_28017,N_24541,N_22169);
nor U28018 (N_28018,N_23878,N_23514);
or U28019 (N_28019,N_23638,N_23273);
or U28020 (N_28020,N_22324,N_24302);
nand U28021 (N_28021,N_24817,N_22992);
and U28022 (N_28022,N_20837,N_23549);
xor U28023 (N_28023,N_20514,N_23180);
nand U28024 (N_28024,N_20605,N_22680);
nand U28025 (N_28025,N_21047,N_21910);
xnor U28026 (N_28026,N_22555,N_24092);
and U28027 (N_28027,N_20414,N_22089);
or U28028 (N_28028,N_20690,N_20988);
nand U28029 (N_28029,N_24206,N_23491);
or U28030 (N_28030,N_23737,N_23429);
or U28031 (N_28031,N_21748,N_20958);
nand U28032 (N_28032,N_23490,N_20194);
nor U28033 (N_28033,N_22031,N_23486);
and U28034 (N_28034,N_20181,N_20663);
nor U28035 (N_28035,N_22602,N_23890);
or U28036 (N_28036,N_21653,N_23224);
and U28037 (N_28037,N_24065,N_21271);
and U28038 (N_28038,N_20584,N_23090);
xor U28039 (N_28039,N_22622,N_23576);
xnor U28040 (N_28040,N_22704,N_23452);
and U28041 (N_28041,N_20838,N_24929);
or U28042 (N_28042,N_23161,N_23857);
nor U28043 (N_28043,N_21755,N_23475);
nor U28044 (N_28044,N_21098,N_22839);
and U28045 (N_28045,N_20933,N_22020);
nor U28046 (N_28046,N_24586,N_21637);
and U28047 (N_28047,N_22023,N_21043);
xnor U28048 (N_28048,N_24758,N_20681);
nand U28049 (N_28049,N_21330,N_21349);
xor U28050 (N_28050,N_22537,N_23918);
nor U28051 (N_28051,N_21824,N_22286);
xnor U28052 (N_28052,N_21459,N_22928);
xnor U28053 (N_28053,N_20665,N_21336);
nand U28054 (N_28054,N_22425,N_24421);
or U28055 (N_28055,N_20117,N_23474);
nor U28056 (N_28056,N_22092,N_24062);
nor U28057 (N_28057,N_24203,N_24408);
nand U28058 (N_28058,N_22615,N_20473);
nor U28059 (N_28059,N_21047,N_21213);
and U28060 (N_28060,N_21197,N_20994);
or U28061 (N_28061,N_24609,N_20883);
and U28062 (N_28062,N_22306,N_22912);
nor U28063 (N_28063,N_20939,N_22910);
nand U28064 (N_28064,N_24182,N_24049);
nor U28065 (N_28065,N_23124,N_21313);
nand U28066 (N_28066,N_20762,N_24773);
nand U28067 (N_28067,N_21543,N_20668);
nand U28068 (N_28068,N_20429,N_23601);
or U28069 (N_28069,N_20399,N_23192);
nor U28070 (N_28070,N_21024,N_24118);
nand U28071 (N_28071,N_22073,N_22871);
nor U28072 (N_28072,N_21485,N_22208);
nor U28073 (N_28073,N_22121,N_23521);
nand U28074 (N_28074,N_23859,N_22026);
or U28075 (N_28075,N_21775,N_22731);
xnor U28076 (N_28076,N_22845,N_24086);
and U28077 (N_28077,N_21181,N_20966);
nand U28078 (N_28078,N_24013,N_21336);
xor U28079 (N_28079,N_23551,N_22655);
nor U28080 (N_28080,N_20700,N_22849);
nand U28081 (N_28081,N_21693,N_23229);
or U28082 (N_28082,N_22318,N_20704);
xor U28083 (N_28083,N_22137,N_20613);
and U28084 (N_28084,N_24986,N_22949);
xor U28085 (N_28085,N_24736,N_21385);
or U28086 (N_28086,N_23848,N_23064);
and U28087 (N_28087,N_20621,N_23368);
and U28088 (N_28088,N_23374,N_22985);
xnor U28089 (N_28089,N_22293,N_22682);
xor U28090 (N_28090,N_22523,N_20260);
nand U28091 (N_28091,N_24192,N_23603);
or U28092 (N_28092,N_22483,N_20088);
or U28093 (N_28093,N_22330,N_22263);
nand U28094 (N_28094,N_20654,N_23382);
xor U28095 (N_28095,N_23345,N_23662);
xnor U28096 (N_28096,N_22163,N_23200);
and U28097 (N_28097,N_22614,N_20440);
nor U28098 (N_28098,N_20642,N_23789);
nor U28099 (N_28099,N_22142,N_24407);
nor U28100 (N_28100,N_21710,N_20286);
nand U28101 (N_28101,N_24542,N_22044);
nor U28102 (N_28102,N_23766,N_22379);
nor U28103 (N_28103,N_24215,N_21717);
or U28104 (N_28104,N_21831,N_21273);
nand U28105 (N_28105,N_22056,N_20099);
and U28106 (N_28106,N_20602,N_24101);
nor U28107 (N_28107,N_21880,N_20006);
nor U28108 (N_28108,N_21040,N_20870);
nand U28109 (N_28109,N_24858,N_22222);
and U28110 (N_28110,N_22103,N_20542);
xnor U28111 (N_28111,N_22013,N_20669);
or U28112 (N_28112,N_24222,N_20154);
nand U28113 (N_28113,N_22761,N_24739);
or U28114 (N_28114,N_22167,N_20415);
nor U28115 (N_28115,N_23023,N_21717);
nor U28116 (N_28116,N_21436,N_20625);
and U28117 (N_28117,N_23473,N_24138);
or U28118 (N_28118,N_24092,N_24748);
nor U28119 (N_28119,N_22784,N_24218);
or U28120 (N_28120,N_24586,N_21023);
nand U28121 (N_28121,N_24616,N_23830);
xnor U28122 (N_28122,N_24190,N_23268);
or U28123 (N_28123,N_23805,N_20483);
xnor U28124 (N_28124,N_21799,N_21704);
or U28125 (N_28125,N_21263,N_22187);
nand U28126 (N_28126,N_24502,N_24109);
or U28127 (N_28127,N_24493,N_24037);
or U28128 (N_28128,N_22562,N_22420);
nor U28129 (N_28129,N_20263,N_21989);
nand U28130 (N_28130,N_24233,N_20026);
xnor U28131 (N_28131,N_20766,N_20990);
nand U28132 (N_28132,N_22638,N_22666);
and U28133 (N_28133,N_23199,N_20344);
xor U28134 (N_28134,N_23189,N_23887);
and U28135 (N_28135,N_20156,N_24770);
nand U28136 (N_28136,N_22448,N_23838);
and U28137 (N_28137,N_24767,N_24073);
nor U28138 (N_28138,N_20727,N_20744);
xor U28139 (N_28139,N_21378,N_23836);
xor U28140 (N_28140,N_23882,N_21199);
and U28141 (N_28141,N_20103,N_24341);
or U28142 (N_28142,N_24284,N_24369);
nand U28143 (N_28143,N_20224,N_23278);
nand U28144 (N_28144,N_23930,N_22643);
nand U28145 (N_28145,N_23023,N_21237);
nor U28146 (N_28146,N_21795,N_24195);
xnor U28147 (N_28147,N_24523,N_21201);
and U28148 (N_28148,N_22175,N_21959);
xor U28149 (N_28149,N_22152,N_21199);
xnor U28150 (N_28150,N_20441,N_23658);
xnor U28151 (N_28151,N_20971,N_22667);
xnor U28152 (N_28152,N_24235,N_24210);
xor U28153 (N_28153,N_23187,N_20893);
nand U28154 (N_28154,N_23420,N_21317);
and U28155 (N_28155,N_20203,N_21248);
and U28156 (N_28156,N_21851,N_22398);
nand U28157 (N_28157,N_21559,N_21348);
xor U28158 (N_28158,N_24195,N_21646);
nand U28159 (N_28159,N_23462,N_20522);
nand U28160 (N_28160,N_23813,N_23383);
xnor U28161 (N_28161,N_24599,N_21592);
or U28162 (N_28162,N_22753,N_24576);
and U28163 (N_28163,N_23783,N_20481);
or U28164 (N_28164,N_23592,N_24115);
or U28165 (N_28165,N_21709,N_20281);
or U28166 (N_28166,N_21391,N_22520);
or U28167 (N_28167,N_20220,N_20542);
or U28168 (N_28168,N_22006,N_22882);
and U28169 (N_28169,N_23757,N_24108);
or U28170 (N_28170,N_23621,N_20340);
nor U28171 (N_28171,N_24171,N_20156);
or U28172 (N_28172,N_21753,N_24058);
xnor U28173 (N_28173,N_21171,N_20445);
and U28174 (N_28174,N_20335,N_24741);
xnor U28175 (N_28175,N_22757,N_21187);
nor U28176 (N_28176,N_22466,N_21530);
xnor U28177 (N_28177,N_21240,N_21802);
xor U28178 (N_28178,N_21943,N_23810);
or U28179 (N_28179,N_24799,N_23954);
nand U28180 (N_28180,N_21367,N_24175);
nor U28181 (N_28181,N_20566,N_23247);
nor U28182 (N_28182,N_20493,N_24043);
and U28183 (N_28183,N_24108,N_23093);
or U28184 (N_28184,N_20003,N_21320);
nor U28185 (N_28185,N_22706,N_20904);
xnor U28186 (N_28186,N_23247,N_24609);
nor U28187 (N_28187,N_23991,N_21717);
and U28188 (N_28188,N_23641,N_21799);
xor U28189 (N_28189,N_22653,N_23801);
nand U28190 (N_28190,N_24854,N_24708);
and U28191 (N_28191,N_20460,N_24928);
nand U28192 (N_28192,N_21027,N_24488);
or U28193 (N_28193,N_20193,N_20204);
nand U28194 (N_28194,N_22698,N_20675);
and U28195 (N_28195,N_22204,N_20391);
xor U28196 (N_28196,N_24821,N_20725);
nand U28197 (N_28197,N_22593,N_24070);
nand U28198 (N_28198,N_20857,N_21153);
nand U28199 (N_28199,N_23587,N_20641);
xnor U28200 (N_28200,N_21549,N_21941);
nand U28201 (N_28201,N_23685,N_24854);
or U28202 (N_28202,N_22109,N_22452);
nand U28203 (N_28203,N_20701,N_24696);
and U28204 (N_28204,N_23005,N_21173);
or U28205 (N_28205,N_23429,N_24838);
nor U28206 (N_28206,N_24794,N_22851);
nand U28207 (N_28207,N_21865,N_21589);
nand U28208 (N_28208,N_21111,N_23862);
or U28209 (N_28209,N_22073,N_20437);
and U28210 (N_28210,N_21070,N_22151);
and U28211 (N_28211,N_22167,N_20984);
nand U28212 (N_28212,N_21371,N_21521);
nor U28213 (N_28213,N_21867,N_23228);
nand U28214 (N_28214,N_22997,N_22433);
nor U28215 (N_28215,N_21817,N_22286);
nand U28216 (N_28216,N_21028,N_24790);
or U28217 (N_28217,N_24201,N_22373);
or U28218 (N_28218,N_23481,N_24843);
xnor U28219 (N_28219,N_20167,N_20890);
xnor U28220 (N_28220,N_24094,N_20151);
nand U28221 (N_28221,N_21700,N_24661);
nand U28222 (N_28222,N_21150,N_21183);
and U28223 (N_28223,N_22665,N_20030);
nor U28224 (N_28224,N_21270,N_20738);
or U28225 (N_28225,N_21880,N_24398);
and U28226 (N_28226,N_24155,N_24322);
nand U28227 (N_28227,N_20782,N_21828);
nor U28228 (N_28228,N_23848,N_24286);
nor U28229 (N_28229,N_24483,N_24024);
xor U28230 (N_28230,N_20311,N_23376);
xnor U28231 (N_28231,N_22475,N_23635);
xnor U28232 (N_28232,N_21878,N_23280);
nor U28233 (N_28233,N_24355,N_20672);
and U28234 (N_28234,N_20089,N_21282);
nor U28235 (N_28235,N_20118,N_22969);
and U28236 (N_28236,N_20834,N_23531);
and U28237 (N_28237,N_24053,N_24065);
nand U28238 (N_28238,N_24788,N_21704);
nor U28239 (N_28239,N_21169,N_20611);
nand U28240 (N_28240,N_23983,N_21642);
xnor U28241 (N_28241,N_22281,N_22417);
nand U28242 (N_28242,N_20055,N_22667);
xor U28243 (N_28243,N_21793,N_21795);
nor U28244 (N_28244,N_20394,N_22142);
nand U28245 (N_28245,N_22014,N_20643);
and U28246 (N_28246,N_20422,N_22633);
and U28247 (N_28247,N_23570,N_24865);
and U28248 (N_28248,N_23923,N_23249);
or U28249 (N_28249,N_21564,N_24695);
or U28250 (N_28250,N_20407,N_21299);
and U28251 (N_28251,N_22720,N_24777);
or U28252 (N_28252,N_20583,N_20378);
or U28253 (N_28253,N_23278,N_20812);
nand U28254 (N_28254,N_21704,N_23664);
xnor U28255 (N_28255,N_20533,N_21765);
and U28256 (N_28256,N_24280,N_23831);
xor U28257 (N_28257,N_24244,N_24466);
nand U28258 (N_28258,N_22579,N_24037);
and U28259 (N_28259,N_22441,N_22988);
nand U28260 (N_28260,N_24542,N_24277);
nor U28261 (N_28261,N_22742,N_23249);
or U28262 (N_28262,N_24613,N_21402);
or U28263 (N_28263,N_21173,N_24424);
nor U28264 (N_28264,N_23722,N_24663);
and U28265 (N_28265,N_21401,N_20149);
nand U28266 (N_28266,N_23501,N_20749);
or U28267 (N_28267,N_20862,N_21412);
nand U28268 (N_28268,N_24519,N_22940);
and U28269 (N_28269,N_21949,N_23062);
xnor U28270 (N_28270,N_24254,N_22725);
xor U28271 (N_28271,N_22859,N_21367);
or U28272 (N_28272,N_21195,N_20256);
xor U28273 (N_28273,N_23408,N_20038);
nor U28274 (N_28274,N_20176,N_21532);
xnor U28275 (N_28275,N_24765,N_21626);
nand U28276 (N_28276,N_21656,N_20830);
nor U28277 (N_28277,N_23786,N_22839);
or U28278 (N_28278,N_22522,N_24214);
nor U28279 (N_28279,N_23019,N_23023);
and U28280 (N_28280,N_24756,N_22412);
and U28281 (N_28281,N_22402,N_24368);
and U28282 (N_28282,N_21822,N_20126);
or U28283 (N_28283,N_24483,N_22272);
nor U28284 (N_28284,N_23190,N_24021);
nor U28285 (N_28285,N_21232,N_24056);
xor U28286 (N_28286,N_24202,N_23093);
nand U28287 (N_28287,N_20510,N_24303);
nor U28288 (N_28288,N_23014,N_20910);
nor U28289 (N_28289,N_24111,N_24969);
nand U28290 (N_28290,N_20561,N_22549);
nand U28291 (N_28291,N_24198,N_24327);
and U28292 (N_28292,N_20866,N_24145);
nand U28293 (N_28293,N_22615,N_20368);
or U28294 (N_28294,N_23009,N_20205);
nand U28295 (N_28295,N_22781,N_23837);
nor U28296 (N_28296,N_21202,N_23697);
or U28297 (N_28297,N_20849,N_20162);
nand U28298 (N_28298,N_23229,N_20979);
xor U28299 (N_28299,N_21972,N_23786);
xor U28300 (N_28300,N_24345,N_23234);
nand U28301 (N_28301,N_24536,N_21009);
or U28302 (N_28302,N_24996,N_24194);
nand U28303 (N_28303,N_21084,N_21495);
and U28304 (N_28304,N_22504,N_24743);
or U28305 (N_28305,N_23911,N_24727);
nand U28306 (N_28306,N_24904,N_21536);
nor U28307 (N_28307,N_22847,N_24193);
nor U28308 (N_28308,N_24026,N_21774);
nor U28309 (N_28309,N_24084,N_22686);
or U28310 (N_28310,N_22338,N_24703);
or U28311 (N_28311,N_23187,N_24840);
nand U28312 (N_28312,N_22991,N_22957);
nor U28313 (N_28313,N_23162,N_20578);
or U28314 (N_28314,N_20941,N_21180);
nand U28315 (N_28315,N_22235,N_20775);
or U28316 (N_28316,N_23892,N_20895);
or U28317 (N_28317,N_20801,N_20572);
nand U28318 (N_28318,N_20432,N_23294);
nand U28319 (N_28319,N_20584,N_23895);
nand U28320 (N_28320,N_24619,N_21042);
xor U28321 (N_28321,N_22068,N_21771);
xnor U28322 (N_28322,N_21904,N_22043);
nor U28323 (N_28323,N_20837,N_21692);
nor U28324 (N_28324,N_22628,N_23715);
nor U28325 (N_28325,N_24025,N_20542);
nor U28326 (N_28326,N_24665,N_24431);
and U28327 (N_28327,N_20137,N_24246);
and U28328 (N_28328,N_24894,N_20846);
or U28329 (N_28329,N_23627,N_21803);
xnor U28330 (N_28330,N_21758,N_23801);
or U28331 (N_28331,N_23796,N_22239);
nor U28332 (N_28332,N_24738,N_23010);
xor U28333 (N_28333,N_22718,N_24499);
and U28334 (N_28334,N_22456,N_23009);
nor U28335 (N_28335,N_23152,N_21034);
nand U28336 (N_28336,N_23638,N_20409);
or U28337 (N_28337,N_21335,N_21425);
xor U28338 (N_28338,N_22646,N_20622);
nor U28339 (N_28339,N_24294,N_24496);
xor U28340 (N_28340,N_23437,N_24375);
nor U28341 (N_28341,N_24444,N_21972);
or U28342 (N_28342,N_21940,N_21642);
xnor U28343 (N_28343,N_21320,N_22489);
nand U28344 (N_28344,N_23763,N_24774);
nor U28345 (N_28345,N_22611,N_23899);
nand U28346 (N_28346,N_24077,N_21328);
xor U28347 (N_28347,N_20892,N_22450);
nor U28348 (N_28348,N_21489,N_21637);
nand U28349 (N_28349,N_21616,N_23082);
or U28350 (N_28350,N_20589,N_23146);
xor U28351 (N_28351,N_20880,N_20550);
and U28352 (N_28352,N_21111,N_23176);
and U28353 (N_28353,N_20871,N_20062);
xor U28354 (N_28354,N_20305,N_20175);
nand U28355 (N_28355,N_24893,N_20792);
nor U28356 (N_28356,N_20557,N_22043);
or U28357 (N_28357,N_23343,N_21117);
xor U28358 (N_28358,N_22716,N_21514);
nand U28359 (N_28359,N_21649,N_24931);
nand U28360 (N_28360,N_24054,N_21843);
nand U28361 (N_28361,N_23729,N_21519);
nor U28362 (N_28362,N_24391,N_24198);
xor U28363 (N_28363,N_22492,N_22115);
and U28364 (N_28364,N_23279,N_22278);
nand U28365 (N_28365,N_24055,N_20746);
nor U28366 (N_28366,N_21884,N_20633);
xor U28367 (N_28367,N_24836,N_22233);
and U28368 (N_28368,N_20917,N_21619);
or U28369 (N_28369,N_22762,N_23103);
nor U28370 (N_28370,N_21867,N_24178);
nor U28371 (N_28371,N_23678,N_20208);
nand U28372 (N_28372,N_23195,N_24273);
xnor U28373 (N_28373,N_20923,N_22588);
xor U28374 (N_28374,N_20601,N_22243);
and U28375 (N_28375,N_21133,N_23984);
xnor U28376 (N_28376,N_20030,N_24422);
or U28377 (N_28377,N_22571,N_21289);
xnor U28378 (N_28378,N_24380,N_24889);
or U28379 (N_28379,N_21259,N_24805);
nand U28380 (N_28380,N_22130,N_21755);
and U28381 (N_28381,N_22334,N_21705);
nor U28382 (N_28382,N_24350,N_22234);
nand U28383 (N_28383,N_20332,N_23740);
xnor U28384 (N_28384,N_21685,N_22846);
or U28385 (N_28385,N_23995,N_21338);
nor U28386 (N_28386,N_21934,N_24920);
nor U28387 (N_28387,N_22422,N_21526);
nand U28388 (N_28388,N_23269,N_20787);
xor U28389 (N_28389,N_22509,N_21300);
nand U28390 (N_28390,N_24902,N_20849);
and U28391 (N_28391,N_21305,N_24195);
nor U28392 (N_28392,N_24564,N_23884);
nor U28393 (N_28393,N_23582,N_21305);
nand U28394 (N_28394,N_23725,N_23661);
and U28395 (N_28395,N_23649,N_23239);
nand U28396 (N_28396,N_24593,N_21397);
xnor U28397 (N_28397,N_22496,N_24152);
xnor U28398 (N_28398,N_20486,N_21842);
nor U28399 (N_28399,N_21227,N_22929);
or U28400 (N_28400,N_23488,N_20919);
or U28401 (N_28401,N_24914,N_20907);
or U28402 (N_28402,N_20817,N_24830);
nor U28403 (N_28403,N_23605,N_20328);
nor U28404 (N_28404,N_23725,N_22889);
and U28405 (N_28405,N_24299,N_22414);
or U28406 (N_28406,N_22561,N_24898);
or U28407 (N_28407,N_21680,N_20303);
and U28408 (N_28408,N_23324,N_22841);
xnor U28409 (N_28409,N_24789,N_21654);
xnor U28410 (N_28410,N_20971,N_22780);
nor U28411 (N_28411,N_24142,N_20402);
and U28412 (N_28412,N_21653,N_23119);
or U28413 (N_28413,N_24906,N_20751);
or U28414 (N_28414,N_22123,N_20430);
nor U28415 (N_28415,N_21230,N_23711);
nand U28416 (N_28416,N_24330,N_24285);
nand U28417 (N_28417,N_22608,N_20249);
nand U28418 (N_28418,N_20799,N_22338);
and U28419 (N_28419,N_21207,N_23330);
nor U28420 (N_28420,N_22617,N_20995);
and U28421 (N_28421,N_24387,N_20410);
nand U28422 (N_28422,N_20922,N_21183);
nand U28423 (N_28423,N_22632,N_21288);
nand U28424 (N_28424,N_22105,N_24503);
nand U28425 (N_28425,N_20632,N_24345);
xnor U28426 (N_28426,N_21544,N_22411);
xnor U28427 (N_28427,N_24906,N_23561);
nor U28428 (N_28428,N_24861,N_21551);
xnor U28429 (N_28429,N_20766,N_22602);
nor U28430 (N_28430,N_23178,N_22373);
xnor U28431 (N_28431,N_24943,N_20778);
and U28432 (N_28432,N_23480,N_21812);
or U28433 (N_28433,N_22249,N_22020);
nor U28434 (N_28434,N_24613,N_20963);
nand U28435 (N_28435,N_24078,N_20881);
nand U28436 (N_28436,N_23163,N_20550);
nor U28437 (N_28437,N_22565,N_20524);
nor U28438 (N_28438,N_20686,N_21583);
nor U28439 (N_28439,N_23253,N_24982);
nor U28440 (N_28440,N_24336,N_21596);
nor U28441 (N_28441,N_24943,N_20718);
and U28442 (N_28442,N_20005,N_20479);
and U28443 (N_28443,N_21071,N_22171);
xnor U28444 (N_28444,N_21737,N_23418);
and U28445 (N_28445,N_20921,N_23986);
nand U28446 (N_28446,N_20518,N_21812);
xnor U28447 (N_28447,N_24209,N_24439);
and U28448 (N_28448,N_22984,N_20263);
xnor U28449 (N_28449,N_20286,N_21120);
nor U28450 (N_28450,N_24839,N_22689);
nand U28451 (N_28451,N_21527,N_21953);
xnor U28452 (N_28452,N_22626,N_24330);
and U28453 (N_28453,N_24324,N_22792);
or U28454 (N_28454,N_22269,N_22891);
and U28455 (N_28455,N_21587,N_21967);
and U28456 (N_28456,N_23512,N_23075);
nand U28457 (N_28457,N_21262,N_24830);
nor U28458 (N_28458,N_24542,N_24085);
nand U28459 (N_28459,N_24828,N_24974);
xnor U28460 (N_28460,N_21374,N_21726);
xor U28461 (N_28461,N_24723,N_20574);
nor U28462 (N_28462,N_20201,N_21052);
nor U28463 (N_28463,N_21285,N_20935);
nor U28464 (N_28464,N_22330,N_24187);
nor U28465 (N_28465,N_23021,N_23545);
nor U28466 (N_28466,N_21725,N_22839);
xor U28467 (N_28467,N_23346,N_20079);
nand U28468 (N_28468,N_23292,N_24550);
and U28469 (N_28469,N_22532,N_21132);
nor U28470 (N_28470,N_20955,N_24744);
nand U28471 (N_28471,N_24935,N_20307);
nand U28472 (N_28472,N_21322,N_23748);
xnor U28473 (N_28473,N_22187,N_21890);
or U28474 (N_28474,N_24356,N_22760);
xnor U28475 (N_28475,N_20473,N_21001);
nor U28476 (N_28476,N_23878,N_20751);
nor U28477 (N_28477,N_20038,N_22624);
or U28478 (N_28478,N_23620,N_23337);
xor U28479 (N_28479,N_21477,N_21513);
xor U28480 (N_28480,N_24483,N_24528);
xnor U28481 (N_28481,N_20913,N_22821);
xnor U28482 (N_28482,N_23676,N_23471);
nand U28483 (N_28483,N_22498,N_23125);
nand U28484 (N_28484,N_21819,N_20545);
and U28485 (N_28485,N_24334,N_22831);
or U28486 (N_28486,N_21937,N_24520);
nand U28487 (N_28487,N_20843,N_23281);
nor U28488 (N_28488,N_22110,N_22683);
nor U28489 (N_28489,N_24810,N_23309);
and U28490 (N_28490,N_24015,N_22173);
nand U28491 (N_28491,N_20613,N_24065);
nor U28492 (N_28492,N_20117,N_22176);
xnor U28493 (N_28493,N_22203,N_20246);
xnor U28494 (N_28494,N_20928,N_23405);
nand U28495 (N_28495,N_20741,N_22184);
nand U28496 (N_28496,N_20890,N_22233);
nor U28497 (N_28497,N_21402,N_21979);
nand U28498 (N_28498,N_22396,N_24094);
nor U28499 (N_28499,N_24642,N_22666);
xnor U28500 (N_28500,N_22623,N_22048);
xnor U28501 (N_28501,N_22245,N_23039);
xnor U28502 (N_28502,N_20288,N_23588);
and U28503 (N_28503,N_20362,N_23186);
nand U28504 (N_28504,N_21918,N_23347);
xor U28505 (N_28505,N_22501,N_20063);
nand U28506 (N_28506,N_22531,N_22929);
or U28507 (N_28507,N_24769,N_23604);
xnor U28508 (N_28508,N_22930,N_23594);
xnor U28509 (N_28509,N_22577,N_23941);
xor U28510 (N_28510,N_23170,N_22297);
or U28511 (N_28511,N_20337,N_20748);
nor U28512 (N_28512,N_23780,N_20539);
nand U28513 (N_28513,N_24027,N_24250);
nand U28514 (N_28514,N_24166,N_23676);
nor U28515 (N_28515,N_22688,N_20285);
or U28516 (N_28516,N_23677,N_21529);
xor U28517 (N_28517,N_23355,N_22023);
nand U28518 (N_28518,N_21309,N_20714);
xor U28519 (N_28519,N_24573,N_24990);
or U28520 (N_28520,N_24568,N_20641);
and U28521 (N_28521,N_23436,N_21928);
xnor U28522 (N_28522,N_24433,N_23174);
or U28523 (N_28523,N_24205,N_24094);
and U28524 (N_28524,N_24513,N_20029);
nand U28525 (N_28525,N_23017,N_23833);
nand U28526 (N_28526,N_22606,N_21146);
or U28527 (N_28527,N_20081,N_21879);
or U28528 (N_28528,N_23706,N_23961);
nand U28529 (N_28529,N_20863,N_21322);
or U28530 (N_28530,N_22796,N_20014);
and U28531 (N_28531,N_21609,N_21618);
and U28532 (N_28532,N_24764,N_20942);
or U28533 (N_28533,N_24942,N_21484);
nor U28534 (N_28534,N_21633,N_23525);
nand U28535 (N_28535,N_22912,N_23538);
nand U28536 (N_28536,N_22968,N_20189);
or U28537 (N_28537,N_22804,N_22969);
nor U28538 (N_28538,N_20512,N_24732);
or U28539 (N_28539,N_22467,N_21902);
and U28540 (N_28540,N_24841,N_21327);
xor U28541 (N_28541,N_23973,N_23825);
nand U28542 (N_28542,N_20738,N_20665);
nand U28543 (N_28543,N_20004,N_22148);
nand U28544 (N_28544,N_24674,N_24749);
nand U28545 (N_28545,N_22357,N_23349);
nor U28546 (N_28546,N_24531,N_23203);
xor U28547 (N_28547,N_22645,N_22868);
xor U28548 (N_28548,N_23215,N_24872);
xnor U28549 (N_28549,N_24451,N_24097);
nor U28550 (N_28550,N_23604,N_21951);
nand U28551 (N_28551,N_23339,N_21975);
and U28552 (N_28552,N_21116,N_21076);
nor U28553 (N_28553,N_22538,N_24060);
nor U28554 (N_28554,N_24347,N_21699);
nand U28555 (N_28555,N_21355,N_22990);
nor U28556 (N_28556,N_21469,N_20582);
or U28557 (N_28557,N_22578,N_20806);
xnor U28558 (N_28558,N_23911,N_24851);
nand U28559 (N_28559,N_20965,N_22274);
nor U28560 (N_28560,N_23773,N_20538);
xnor U28561 (N_28561,N_22321,N_22007);
nor U28562 (N_28562,N_20925,N_24727);
and U28563 (N_28563,N_21623,N_23117);
nand U28564 (N_28564,N_23161,N_21429);
nor U28565 (N_28565,N_23258,N_24004);
or U28566 (N_28566,N_22977,N_20411);
or U28567 (N_28567,N_22086,N_24042);
nor U28568 (N_28568,N_23865,N_20408);
nand U28569 (N_28569,N_21550,N_23227);
nor U28570 (N_28570,N_21958,N_24244);
nor U28571 (N_28571,N_21521,N_21020);
and U28572 (N_28572,N_22423,N_23258);
or U28573 (N_28573,N_20972,N_24150);
and U28574 (N_28574,N_24581,N_22130);
and U28575 (N_28575,N_22418,N_24995);
xor U28576 (N_28576,N_21310,N_22622);
or U28577 (N_28577,N_21622,N_22654);
or U28578 (N_28578,N_23149,N_20236);
nand U28579 (N_28579,N_24382,N_24038);
xor U28580 (N_28580,N_21532,N_23519);
or U28581 (N_28581,N_21839,N_23367);
nand U28582 (N_28582,N_24628,N_23962);
or U28583 (N_28583,N_20307,N_24843);
nand U28584 (N_28584,N_20983,N_20903);
xor U28585 (N_28585,N_20439,N_24694);
or U28586 (N_28586,N_20162,N_21886);
xnor U28587 (N_28587,N_24761,N_20757);
nand U28588 (N_28588,N_23955,N_22950);
xnor U28589 (N_28589,N_22527,N_22865);
nor U28590 (N_28590,N_22368,N_20983);
nand U28591 (N_28591,N_22915,N_23565);
or U28592 (N_28592,N_20966,N_24559);
nand U28593 (N_28593,N_20782,N_20961);
nor U28594 (N_28594,N_22141,N_22702);
or U28595 (N_28595,N_20772,N_23306);
or U28596 (N_28596,N_23405,N_21329);
xor U28597 (N_28597,N_24288,N_20019);
and U28598 (N_28598,N_22427,N_24125);
or U28599 (N_28599,N_21741,N_20060);
and U28600 (N_28600,N_21754,N_23525);
nor U28601 (N_28601,N_24437,N_22920);
and U28602 (N_28602,N_20856,N_20474);
nor U28603 (N_28603,N_23164,N_24616);
nor U28604 (N_28604,N_21202,N_24326);
or U28605 (N_28605,N_20788,N_23094);
and U28606 (N_28606,N_20424,N_22486);
nor U28607 (N_28607,N_21171,N_20957);
nor U28608 (N_28608,N_20254,N_22138);
or U28609 (N_28609,N_21544,N_24668);
xnor U28610 (N_28610,N_22369,N_20690);
nor U28611 (N_28611,N_21822,N_20179);
or U28612 (N_28612,N_20590,N_24105);
and U28613 (N_28613,N_20240,N_23767);
and U28614 (N_28614,N_22803,N_21604);
nand U28615 (N_28615,N_22919,N_23968);
or U28616 (N_28616,N_22967,N_20212);
or U28617 (N_28617,N_22791,N_20022);
or U28618 (N_28618,N_22853,N_24995);
and U28619 (N_28619,N_23920,N_21066);
nor U28620 (N_28620,N_24588,N_21750);
nand U28621 (N_28621,N_20591,N_24529);
nor U28622 (N_28622,N_23779,N_24940);
or U28623 (N_28623,N_21590,N_24900);
xnor U28624 (N_28624,N_20787,N_23684);
and U28625 (N_28625,N_22226,N_23502);
nor U28626 (N_28626,N_23339,N_23229);
and U28627 (N_28627,N_24509,N_21416);
and U28628 (N_28628,N_21524,N_22355);
nand U28629 (N_28629,N_20616,N_22610);
or U28630 (N_28630,N_20044,N_24349);
xnor U28631 (N_28631,N_21834,N_22948);
xnor U28632 (N_28632,N_21275,N_24446);
xor U28633 (N_28633,N_22368,N_20662);
and U28634 (N_28634,N_20757,N_23244);
nor U28635 (N_28635,N_21555,N_24263);
and U28636 (N_28636,N_24179,N_24688);
and U28637 (N_28637,N_21493,N_23295);
or U28638 (N_28638,N_23919,N_21880);
or U28639 (N_28639,N_22452,N_23407);
or U28640 (N_28640,N_20933,N_22545);
or U28641 (N_28641,N_22518,N_24767);
and U28642 (N_28642,N_20926,N_20430);
and U28643 (N_28643,N_20502,N_24273);
and U28644 (N_28644,N_23645,N_24271);
nand U28645 (N_28645,N_22072,N_21368);
nand U28646 (N_28646,N_22325,N_22846);
xor U28647 (N_28647,N_23582,N_21545);
xnor U28648 (N_28648,N_22918,N_24361);
or U28649 (N_28649,N_22468,N_22331);
nor U28650 (N_28650,N_23089,N_24160);
and U28651 (N_28651,N_21744,N_20037);
nor U28652 (N_28652,N_21072,N_24733);
or U28653 (N_28653,N_24372,N_21388);
nand U28654 (N_28654,N_21423,N_22591);
nand U28655 (N_28655,N_22569,N_23720);
and U28656 (N_28656,N_22435,N_21726);
or U28657 (N_28657,N_24226,N_22179);
and U28658 (N_28658,N_21203,N_21245);
nand U28659 (N_28659,N_24383,N_20593);
nor U28660 (N_28660,N_23491,N_24241);
or U28661 (N_28661,N_20618,N_24890);
or U28662 (N_28662,N_22168,N_24626);
xor U28663 (N_28663,N_22672,N_20507);
and U28664 (N_28664,N_20620,N_21293);
nand U28665 (N_28665,N_21326,N_24464);
nand U28666 (N_28666,N_20103,N_24156);
or U28667 (N_28667,N_22620,N_23588);
nor U28668 (N_28668,N_20971,N_21557);
and U28669 (N_28669,N_21710,N_21645);
nand U28670 (N_28670,N_23080,N_23090);
or U28671 (N_28671,N_21451,N_23992);
nand U28672 (N_28672,N_24553,N_24303);
xor U28673 (N_28673,N_24310,N_23591);
and U28674 (N_28674,N_24229,N_23021);
nand U28675 (N_28675,N_24688,N_22627);
nand U28676 (N_28676,N_22492,N_20208);
nor U28677 (N_28677,N_20701,N_23202);
nand U28678 (N_28678,N_20521,N_22159);
and U28679 (N_28679,N_22874,N_23053);
nor U28680 (N_28680,N_21572,N_24057);
nor U28681 (N_28681,N_23504,N_24168);
or U28682 (N_28682,N_24938,N_20777);
xnor U28683 (N_28683,N_22451,N_22478);
and U28684 (N_28684,N_22755,N_24059);
nor U28685 (N_28685,N_21549,N_21636);
or U28686 (N_28686,N_23371,N_20611);
and U28687 (N_28687,N_20996,N_21982);
nand U28688 (N_28688,N_20244,N_23519);
xor U28689 (N_28689,N_20370,N_22489);
xnor U28690 (N_28690,N_20847,N_21729);
or U28691 (N_28691,N_22065,N_23225);
nand U28692 (N_28692,N_20371,N_21613);
nor U28693 (N_28693,N_24794,N_23651);
and U28694 (N_28694,N_23538,N_21199);
xnor U28695 (N_28695,N_22680,N_21004);
xor U28696 (N_28696,N_23890,N_21808);
and U28697 (N_28697,N_22606,N_23522);
and U28698 (N_28698,N_21815,N_24932);
and U28699 (N_28699,N_23430,N_22437);
and U28700 (N_28700,N_20445,N_21942);
nor U28701 (N_28701,N_21232,N_22202);
xnor U28702 (N_28702,N_22614,N_21997);
nand U28703 (N_28703,N_23389,N_23164);
nand U28704 (N_28704,N_24651,N_21994);
and U28705 (N_28705,N_21429,N_20788);
xor U28706 (N_28706,N_20220,N_24721);
nor U28707 (N_28707,N_23449,N_23545);
or U28708 (N_28708,N_20617,N_20651);
or U28709 (N_28709,N_22498,N_24659);
nand U28710 (N_28710,N_22723,N_24971);
or U28711 (N_28711,N_23452,N_23649);
nor U28712 (N_28712,N_21609,N_21594);
or U28713 (N_28713,N_22767,N_20503);
or U28714 (N_28714,N_21408,N_22580);
nand U28715 (N_28715,N_21345,N_21850);
xnor U28716 (N_28716,N_24410,N_24926);
nor U28717 (N_28717,N_21968,N_22238);
nor U28718 (N_28718,N_20357,N_24857);
and U28719 (N_28719,N_20848,N_21392);
nand U28720 (N_28720,N_22895,N_20316);
nor U28721 (N_28721,N_21773,N_23519);
nand U28722 (N_28722,N_21668,N_24304);
nand U28723 (N_28723,N_21787,N_24045);
and U28724 (N_28724,N_23275,N_24109);
nor U28725 (N_28725,N_20480,N_21390);
nor U28726 (N_28726,N_23115,N_21514);
or U28727 (N_28727,N_24742,N_21710);
xor U28728 (N_28728,N_23813,N_23721);
nand U28729 (N_28729,N_22974,N_20123);
and U28730 (N_28730,N_20291,N_21673);
nand U28731 (N_28731,N_20712,N_24297);
nand U28732 (N_28732,N_24335,N_23597);
or U28733 (N_28733,N_20948,N_20696);
nand U28734 (N_28734,N_22937,N_21017);
or U28735 (N_28735,N_24538,N_20501);
nor U28736 (N_28736,N_20324,N_20718);
nand U28737 (N_28737,N_24420,N_21562);
xnor U28738 (N_28738,N_23676,N_23901);
or U28739 (N_28739,N_22740,N_21268);
or U28740 (N_28740,N_20192,N_22106);
or U28741 (N_28741,N_23997,N_22516);
or U28742 (N_28742,N_20672,N_20574);
or U28743 (N_28743,N_24595,N_23098);
xor U28744 (N_28744,N_24491,N_20418);
and U28745 (N_28745,N_23903,N_21029);
nand U28746 (N_28746,N_23861,N_22889);
nor U28747 (N_28747,N_21470,N_22963);
xnor U28748 (N_28748,N_21921,N_24996);
xnor U28749 (N_28749,N_22479,N_20761);
nand U28750 (N_28750,N_24380,N_21070);
nor U28751 (N_28751,N_22490,N_22087);
and U28752 (N_28752,N_22684,N_23919);
xnor U28753 (N_28753,N_21546,N_22028);
nor U28754 (N_28754,N_20542,N_21818);
and U28755 (N_28755,N_22901,N_23139);
and U28756 (N_28756,N_21424,N_24546);
nor U28757 (N_28757,N_20123,N_21951);
and U28758 (N_28758,N_20548,N_24766);
or U28759 (N_28759,N_24538,N_21735);
xnor U28760 (N_28760,N_21228,N_24465);
xor U28761 (N_28761,N_22016,N_20021);
xnor U28762 (N_28762,N_21720,N_20616);
or U28763 (N_28763,N_21857,N_20166);
nand U28764 (N_28764,N_24722,N_22458);
nand U28765 (N_28765,N_24070,N_20252);
or U28766 (N_28766,N_21686,N_23369);
nor U28767 (N_28767,N_24699,N_20169);
or U28768 (N_28768,N_20777,N_20327);
and U28769 (N_28769,N_20212,N_21969);
or U28770 (N_28770,N_22364,N_21147);
nand U28771 (N_28771,N_21541,N_22322);
xnor U28772 (N_28772,N_22434,N_23537);
or U28773 (N_28773,N_22555,N_24448);
xnor U28774 (N_28774,N_21464,N_22606);
nand U28775 (N_28775,N_23393,N_22217);
and U28776 (N_28776,N_20452,N_20394);
or U28777 (N_28777,N_24566,N_24523);
and U28778 (N_28778,N_21263,N_23978);
nor U28779 (N_28779,N_20894,N_23386);
xnor U28780 (N_28780,N_22794,N_24022);
or U28781 (N_28781,N_23381,N_23533);
xor U28782 (N_28782,N_23077,N_21805);
nand U28783 (N_28783,N_23262,N_20578);
xnor U28784 (N_28784,N_23448,N_21784);
and U28785 (N_28785,N_21973,N_23759);
or U28786 (N_28786,N_22067,N_24395);
and U28787 (N_28787,N_21819,N_22175);
nor U28788 (N_28788,N_22376,N_24823);
xnor U28789 (N_28789,N_24654,N_21865);
and U28790 (N_28790,N_21881,N_20143);
nand U28791 (N_28791,N_24319,N_20477);
xnor U28792 (N_28792,N_23765,N_22943);
nand U28793 (N_28793,N_21961,N_24439);
and U28794 (N_28794,N_22243,N_20793);
and U28795 (N_28795,N_22030,N_20939);
or U28796 (N_28796,N_20084,N_23381);
nand U28797 (N_28797,N_23590,N_21530);
nand U28798 (N_28798,N_20483,N_21134);
nand U28799 (N_28799,N_24666,N_24742);
nand U28800 (N_28800,N_20726,N_24506);
xor U28801 (N_28801,N_21193,N_23121);
or U28802 (N_28802,N_20814,N_24198);
or U28803 (N_28803,N_21922,N_24534);
xor U28804 (N_28804,N_20787,N_21174);
and U28805 (N_28805,N_23295,N_22810);
and U28806 (N_28806,N_21983,N_21307);
and U28807 (N_28807,N_20143,N_24393);
and U28808 (N_28808,N_23845,N_20147);
nand U28809 (N_28809,N_23304,N_23923);
or U28810 (N_28810,N_22880,N_20730);
xor U28811 (N_28811,N_20992,N_21175);
nor U28812 (N_28812,N_21899,N_24410);
or U28813 (N_28813,N_24920,N_22118);
nand U28814 (N_28814,N_21834,N_20866);
or U28815 (N_28815,N_24939,N_22340);
nand U28816 (N_28816,N_20865,N_20949);
and U28817 (N_28817,N_22593,N_21059);
nand U28818 (N_28818,N_22752,N_24030);
or U28819 (N_28819,N_23753,N_22568);
nor U28820 (N_28820,N_21161,N_23744);
xor U28821 (N_28821,N_24574,N_20161);
nor U28822 (N_28822,N_20926,N_22313);
nor U28823 (N_28823,N_21031,N_23501);
or U28824 (N_28824,N_24489,N_24898);
and U28825 (N_28825,N_20934,N_24596);
and U28826 (N_28826,N_22541,N_23792);
nand U28827 (N_28827,N_20445,N_22247);
or U28828 (N_28828,N_22599,N_22611);
or U28829 (N_28829,N_23574,N_24209);
and U28830 (N_28830,N_23081,N_24959);
and U28831 (N_28831,N_23762,N_21046);
xor U28832 (N_28832,N_23396,N_21325);
or U28833 (N_28833,N_20793,N_24170);
or U28834 (N_28834,N_23054,N_23019);
or U28835 (N_28835,N_21306,N_22112);
or U28836 (N_28836,N_21675,N_23534);
xnor U28837 (N_28837,N_22544,N_22093);
or U28838 (N_28838,N_23738,N_20157);
nor U28839 (N_28839,N_22804,N_22137);
nand U28840 (N_28840,N_24904,N_24950);
nor U28841 (N_28841,N_22131,N_20137);
or U28842 (N_28842,N_20188,N_23101);
xnor U28843 (N_28843,N_22366,N_21320);
nor U28844 (N_28844,N_23011,N_21232);
nor U28845 (N_28845,N_23273,N_24462);
or U28846 (N_28846,N_20645,N_21674);
and U28847 (N_28847,N_23613,N_24259);
or U28848 (N_28848,N_22461,N_21033);
nand U28849 (N_28849,N_20385,N_21594);
and U28850 (N_28850,N_22051,N_21577);
nand U28851 (N_28851,N_20478,N_20530);
xnor U28852 (N_28852,N_20005,N_21199);
and U28853 (N_28853,N_20748,N_20723);
xor U28854 (N_28854,N_20603,N_22209);
nand U28855 (N_28855,N_23552,N_21483);
and U28856 (N_28856,N_21105,N_22113);
and U28857 (N_28857,N_23080,N_23732);
and U28858 (N_28858,N_20048,N_20558);
xor U28859 (N_28859,N_23197,N_23068);
and U28860 (N_28860,N_20362,N_22894);
nor U28861 (N_28861,N_24651,N_22398);
nor U28862 (N_28862,N_20900,N_20806);
or U28863 (N_28863,N_24469,N_21756);
xor U28864 (N_28864,N_24147,N_23013);
nand U28865 (N_28865,N_22542,N_24747);
nand U28866 (N_28866,N_24268,N_22764);
nand U28867 (N_28867,N_20502,N_21745);
and U28868 (N_28868,N_24790,N_20413);
or U28869 (N_28869,N_20057,N_22269);
or U28870 (N_28870,N_24958,N_21745);
nor U28871 (N_28871,N_24963,N_24941);
nor U28872 (N_28872,N_22428,N_23438);
nor U28873 (N_28873,N_24893,N_20919);
nor U28874 (N_28874,N_22361,N_21328);
nor U28875 (N_28875,N_20222,N_23439);
nand U28876 (N_28876,N_24387,N_24482);
nor U28877 (N_28877,N_20783,N_23710);
and U28878 (N_28878,N_23492,N_21956);
xnor U28879 (N_28879,N_23442,N_22729);
xor U28880 (N_28880,N_23192,N_23186);
nand U28881 (N_28881,N_20321,N_23308);
and U28882 (N_28882,N_20076,N_20898);
nor U28883 (N_28883,N_24710,N_20711);
or U28884 (N_28884,N_21404,N_24793);
and U28885 (N_28885,N_24990,N_21289);
and U28886 (N_28886,N_23937,N_20715);
and U28887 (N_28887,N_22023,N_20635);
or U28888 (N_28888,N_21097,N_24275);
or U28889 (N_28889,N_22285,N_21301);
xor U28890 (N_28890,N_23474,N_24414);
and U28891 (N_28891,N_21014,N_22287);
or U28892 (N_28892,N_24586,N_21436);
nand U28893 (N_28893,N_24000,N_24022);
nor U28894 (N_28894,N_22719,N_21622);
nand U28895 (N_28895,N_23262,N_23593);
xor U28896 (N_28896,N_23305,N_24615);
nor U28897 (N_28897,N_24152,N_23044);
or U28898 (N_28898,N_22235,N_23315);
and U28899 (N_28899,N_21604,N_23901);
and U28900 (N_28900,N_24750,N_23578);
and U28901 (N_28901,N_21318,N_22822);
and U28902 (N_28902,N_20249,N_24817);
nand U28903 (N_28903,N_24751,N_24155);
xor U28904 (N_28904,N_22300,N_22827);
and U28905 (N_28905,N_24310,N_22038);
and U28906 (N_28906,N_21509,N_22225);
nand U28907 (N_28907,N_24651,N_23407);
nor U28908 (N_28908,N_23590,N_20879);
nor U28909 (N_28909,N_24480,N_20577);
xnor U28910 (N_28910,N_22630,N_21112);
or U28911 (N_28911,N_24055,N_24620);
and U28912 (N_28912,N_20263,N_22059);
nor U28913 (N_28913,N_22536,N_21549);
nor U28914 (N_28914,N_22419,N_24456);
nor U28915 (N_28915,N_20504,N_24317);
and U28916 (N_28916,N_22321,N_24174);
xnor U28917 (N_28917,N_24350,N_23380);
xnor U28918 (N_28918,N_23745,N_23076);
and U28919 (N_28919,N_21154,N_20607);
nand U28920 (N_28920,N_22722,N_21706);
xnor U28921 (N_28921,N_22137,N_21310);
xor U28922 (N_28922,N_22370,N_23039);
and U28923 (N_28923,N_22841,N_24940);
xnor U28924 (N_28924,N_21059,N_24981);
nor U28925 (N_28925,N_22014,N_20728);
or U28926 (N_28926,N_24638,N_20268);
nor U28927 (N_28927,N_23174,N_24878);
xor U28928 (N_28928,N_20093,N_24954);
and U28929 (N_28929,N_22791,N_21075);
nor U28930 (N_28930,N_20376,N_20378);
nand U28931 (N_28931,N_21195,N_23550);
xnor U28932 (N_28932,N_21791,N_23399);
xor U28933 (N_28933,N_22229,N_24476);
nand U28934 (N_28934,N_21719,N_24744);
or U28935 (N_28935,N_21643,N_21811);
nand U28936 (N_28936,N_22435,N_23063);
xor U28937 (N_28937,N_20201,N_22336);
nor U28938 (N_28938,N_21922,N_23466);
nor U28939 (N_28939,N_24591,N_21846);
xor U28940 (N_28940,N_20116,N_21691);
nor U28941 (N_28941,N_24646,N_24912);
and U28942 (N_28942,N_23556,N_21188);
or U28943 (N_28943,N_24250,N_24908);
nand U28944 (N_28944,N_24112,N_23105);
nand U28945 (N_28945,N_22704,N_21294);
or U28946 (N_28946,N_21244,N_21843);
and U28947 (N_28947,N_24669,N_23159);
nor U28948 (N_28948,N_21155,N_23253);
nor U28949 (N_28949,N_20039,N_22674);
nor U28950 (N_28950,N_22708,N_23158);
nor U28951 (N_28951,N_24665,N_22940);
and U28952 (N_28952,N_23751,N_24409);
nand U28953 (N_28953,N_24740,N_21294);
nand U28954 (N_28954,N_21478,N_21954);
nor U28955 (N_28955,N_20590,N_20384);
and U28956 (N_28956,N_20606,N_24717);
xnor U28957 (N_28957,N_24133,N_21413);
or U28958 (N_28958,N_20624,N_20425);
xor U28959 (N_28959,N_22852,N_21740);
or U28960 (N_28960,N_21400,N_22542);
nor U28961 (N_28961,N_24605,N_24341);
and U28962 (N_28962,N_22222,N_20227);
and U28963 (N_28963,N_24534,N_20129);
xnor U28964 (N_28964,N_24932,N_24863);
nor U28965 (N_28965,N_22480,N_20594);
xnor U28966 (N_28966,N_23315,N_24430);
and U28967 (N_28967,N_20225,N_22702);
xor U28968 (N_28968,N_23659,N_24167);
xnor U28969 (N_28969,N_21433,N_21973);
or U28970 (N_28970,N_23342,N_23812);
and U28971 (N_28971,N_24564,N_24492);
and U28972 (N_28972,N_20480,N_21153);
nand U28973 (N_28973,N_23180,N_23277);
or U28974 (N_28974,N_22031,N_22552);
nor U28975 (N_28975,N_21384,N_24574);
xor U28976 (N_28976,N_24770,N_20380);
and U28977 (N_28977,N_24824,N_23622);
nor U28978 (N_28978,N_23546,N_22087);
xor U28979 (N_28979,N_21487,N_24869);
or U28980 (N_28980,N_21175,N_24236);
nor U28981 (N_28981,N_22218,N_22123);
nor U28982 (N_28982,N_23780,N_23156);
nand U28983 (N_28983,N_20151,N_23451);
and U28984 (N_28984,N_24707,N_20083);
nand U28985 (N_28985,N_20949,N_22817);
or U28986 (N_28986,N_22922,N_22310);
xnor U28987 (N_28987,N_23225,N_24078);
and U28988 (N_28988,N_23968,N_23769);
xor U28989 (N_28989,N_20147,N_23159);
xor U28990 (N_28990,N_23112,N_20067);
xor U28991 (N_28991,N_21493,N_22797);
xnor U28992 (N_28992,N_22509,N_24509);
nor U28993 (N_28993,N_22533,N_22901);
nor U28994 (N_28994,N_23120,N_23516);
or U28995 (N_28995,N_21853,N_21432);
nor U28996 (N_28996,N_21159,N_23579);
nand U28997 (N_28997,N_21982,N_23386);
nand U28998 (N_28998,N_24996,N_23229);
nor U28999 (N_28999,N_20759,N_22249);
nor U29000 (N_29000,N_20232,N_23391);
and U29001 (N_29001,N_21817,N_20245);
xor U29002 (N_29002,N_23099,N_22661);
xor U29003 (N_29003,N_24534,N_21089);
or U29004 (N_29004,N_23309,N_21739);
xnor U29005 (N_29005,N_23339,N_21896);
nor U29006 (N_29006,N_23011,N_20152);
nor U29007 (N_29007,N_20898,N_24698);
and U29008 (N_29008,N_21101,N_20171);
nor U29009 (N_29009,N_24436,N_20770);
or U29010 (N_29010,N_23420,N_24013);
nand U29011 (N_29011,N_20184,N_20430);
nor U29012 (N_29012,N_21893,N_24338);
nand U29013 (N_29013,N_20596,N_22487);
xor U29014 (N_29014,N_21975,N_22778);
and U29015 (N_29015,N_24614,N_23553);
or U29016 (N_29016,N_21610,N_20034);
nand U29017 (N_29017,N_21346,N_22186);
xor U29018 (N_29018,N_24233,N_24791);
nand U29019 (N_29019,N_20763,N_22511);
or U29020 (N_29020,N_23660,N_23760);
and U29021 (N_29021,N_20819,N_20498);
xor U29022 (N_29022,N_20403,N_24868);
and U29023 (N_29023,N_21765,N_23606);
and U29024 (N_29024,N_22075,N_24474);
and U29025 (N_29025,N_21923,N_21636);
xor U29026 (N_29026,N_22022,N_20884);
or U29027 (N_29027,N_20594,N_23238);
xnor U29028 (N_29028,N_21192,N_20311);
nor U29029 (N_29029,N_21397,N_24471);
nor U29030 (N_29030,N_21683,N_23422);
nor U29031 (N_29031,N_20424,N_24741);
nand U29032 (N_29032,N_21146,N_21966);
and U29033 (N_29033,N_24095,N_22894);
or U29034 (N_29034,N_21955,N_21577);
or U29035 (N_29035,N_24137,N_23514);
xor U29036 (N_29036,N_24128,N_20039);
xor U29037 (N_29037,N_22182,N_23981);
xor U29038 (N_29038,N_21886,N_24273);
nand U29039 (N_29039,N_23807,N_21658);
and U29040 (N_29040,N_21776,N_22198);
xor U29041 (N_29041,N_21645,N_21365);
xor U29042 (N_29042,N_22011,N_21528);
nor U29043 (N_29043,N_20663,N_24746);
nand U29044 (N_29044,N_22311,N_22243);
xnor U29045 (N_29045,N_22407,N_20350);
or U29046 (N_29046,N_24760,N_23898);
xor U29047 (N_29047,N_20716,N_24587);
xor U29048 (N_29048,N_21974,N_22614);
xor U29049 (N_29049,N_21211,N_23810);
and U29050 (N_29050,N_20578,N_23919);
xor U29051 (N_29051,N_20972,N_20606);
or U29052 (N_29052,N_24768,N_23792);
nand U29053 (N_29053,N_23416,N_20843);
nor U29054 (N_29054,N_22587,N_22121);
and U29055 (N_29055,N_20089,N_24141);
nor U29056 (N_29056,N_22266,N_23518);
and U29057 (N_29057,N_24643,N_22804);
nand U29058 (N_29058,N_20655,N_23145);
nor U29059 (N_29059,N_22704,N_24966);
or U29060 (N_29060,N_23424,N_20239);
xnor U29061 (N_29061,N_23689,N_20999);
nor U29062 (N_29062,N_22989,N_22796);
and U29063 (N_29063,N_23798,N_20226);
xor U29064 (N_29064,N_20004,N_21407);
or U29065 (N_29065,N_20748,N_23810);
or U29066 (N_29066,N_20858,N_21671);
or U29067 (N_29067,N_23260,N_22512);
nor U29068 (N_29068,N_22874,N_23337);
and U29069 (N_29069,N_24590,N_22894);
or U29070 (N_29070,N_24954,N_21423);
xor U29071 (N_29071,N_22362,N_21954);
and U29072 (N_29072,N_21026,N_21465);
xor U29073 (N_29073,N_24829,N_21395);
or U29074 (N_29074,N_20925,N_20620);
nand U29075 (N_29075,N_24093,N_20363);
nand U29076 (N_29076,N_23450,N_20768);
or U29077 (N_29077,N_22907,N_23028);
and U29078 (N_29078,N_23162,N_20445);
nor U29079 (N_29079,N_23290,N_21262);
and U29080 (N_29080,N_24268,N_24326);
xor U29081 (N_29081,N_20915,N_24786);
xnor U29082 (N_29082,N_20896,N_22461);
xnor U29083 (N_29083,N_22841,N_23271);
xnor U29084 (N_29084,N_21210,N_21757);
nand U29085 (N_29085,N_22160,N_22290);
or U29086 (N_29086,N_20048,N_22011);
and U29087 (N_29087,N_21762,N_21102);
nor U29088 (N_29088,N_20666,N_24092);
or U29089 (N_29089,N_20236,N_20850);
xnor U29090 (N_29090,N_23868,N_21706);
nand U29091 (N_29091,N_24874,N_23253);
xnor U29092 (N_29092,N_23722,N_20164);
xor U29093 (N_29093,N_21524,N_22114);
nand U29094 (N_29094,N_22725,N_22974);
xnor U29095 (N_29095,N_21257,N_20973);
nor U29096 (N_29096,N_21407,N_21239);
xnor U29097 (N_29097,N_20298,N_23246);
and U29098 (N_29098,N_20943,N_22368);
nor U29099 (N_29099,N_20357,N_22411);
or U29100 (N_29100,N_23451,N_20568);
xnor U29101 (N_29101,N_20827,N_20075);
and U29102 (N_29102,N_21176,N_24383);
or U29103 (N_29103,N_21023,N_20137);
xnor U29104 (N_29104,N_21096,N_22901);
nor U29105 (N_29105,N_24229,N_21147);
nor U29106 (N_29106,N_20731,N_24626);
nand U29107 (N_29107,N_20250,N_21104);
xor U29108 (N_29108,N_22579,N_23419);
and U29109 (N_29109,N_21842,N_23743);
nand U29110 (N_29110,N_22978,N_21194);
or U29111 (N_29111,N_22654,N_22504);
and U29112 (N_29112,N_24247,N_20597);
or U29113 (N_29113,N_24588,N_21154);
xor U29114 (N_29114,N_22719,N_23656);
or U29115 (N_29115,N_22611,N_23719);
and U29116 (N_29116,N_24266,N_23176);
nand U29117 (N_29117,N_24822,N_20707);
and U29118 (N_29118,N_23961,N_21425);
xnor U29119 (N_29119,N_22627,N_20219);
nand U29120 (N_29120,N_22455,N_22181);
nand U29121 (N_29121,N_21079,N_21049);
xnor U29122 (N_29122,N_23567,N_24806);
or U29123 (N_29123,N_23683,N_20585);
or U29124 (N_29124,N_20441,N_24307);
xnor U29125 (N_29125,N_24256,N_23079);
nor U29126 (N_29126,N_20175,N_22474);
nand U29127 (N_29127,N_20352,N_22434);
nand U29128 (N_29128,N_23720,N_23701);
or U29129 (N_29129,N_22556,N_23751);
or U29130 (N_29130,N_21839,N_22604);
and U29131 (N_29131,N_23899,N_24195);
and U29132 (N_29132,N_20742,N_22182);
or U29133 (N_29133,N_20554,N_23805);
or U29134 (N_29134,N_24086,N_22024);
or U29135 (N_29135,N_24839,N_20848);
and U29136 (N_29136,N_20079,N_23373);
and U29137 (N_29137,N_21209,N_21145);
or U29138 (N_29138,N_23781,N_24173);
nor U29139 (N_29139,N_24263,N_21052);
xnor U29140 (N_29140,N_23204,N_24685);
xnor U29141 (N_29141,N_23813,N_21304);
and U29142 (N_29142,N_23332,N_21979);
or U29143 (N_29143,N_21263,N_21228);
nand U29144 (N_29144,N_22539,N_20968);
xor U29145 (N_29145,N_20484,N_22984);
nor U29146 (N_29146,N_20984,N_23631);
and U29147 (N_29147,N_20916,N_22909);
and U29148 (N_29148,N_22141,N_24433);
and U29149 (N_29149,N_20205,N_23365);
nand U29150 (N_29150,N_22439,N_23702);
nand U29151 (N_29151,N_22028,N_21629);
xnor U29152 (N_29152,N_21909,N_23064);
nor U29153 (N_29153,N_20410,N_23612);
or U29154 (N_29154,N_24005,N_20268);
nand U29155 (N_29155,N_22910,N_21848);
xor U29156 (N_29156,N_23532,N_20644);
or U29157 (N_29157,N_23754,N_24507);
xnor U29158 (N_29158,N_20293,N_23506);
xnor U29159 (N_29159,N_21478,N_24371);
xnor U29160 (N_29160,N_23433,N_22430);
or U29161 (N_29161,N_24681,N_22939);
nand U29162 (N_29162,N_22516,N_21094);
xor U29163 (N_29163,N_20472,N_21568);
or U29164 (N_29164,N_24522,N_24968);
or U29165 (N_29165,N_21877,N_20494);
or U29166 (N_29166,N_22182,N_23915);
nand U29167 (N_29167,N_23225,N_24879);
xnor U29168 (N_29168,N_24644,N_21445);
or U29169 (N_29169,N_23173,N_23875);
xor U29170 (N_29170,N_23763,N_24358);
and U29171 (N_29171,N_21389,N_22073);
nor U29172 (N_29172,N_21680,N_23128);
or U29173 (N_29173,N_20115,N_22968);
and U29174 (N_29174,N_24642,N_21110);
and U29175 (N_29175,N_20841,N_20635);
or U29176 (N_29176,N_24742,N_22968);
xor U29177 (N_29177,N_20031,N_22137);
nand U29178 (N_29178,N_22768,N_23415);
or U29179 (N_29179,N_21599,N_20533);
nor U29180 (N_29180,N_22695,N_22988);
or U29181 (N_29181,N_23023,N_22117);
nand U29182 (N_29182,N_22111,N_22568);
nand U29183 (N_29183,N_21249,N_24454);
nor U29184 (N_29184,N_22878,N_22734);
nor U29185 (N_29185,N_24537,N_20073);
or U29186 (N_29186,N_24332,N_24726);
xnor U29187 (N_29187,N_24984,N_23040);
nand U29188 (N_29188,N_24687,N_21136);
nand U29189 (N_29189,N_24299,N_23306);
nand U29190 (N_29190,N_21643,N_21579);
nor U29191 (N_29191,N_22496,N_20520);
nand U29192 (N_29192,N_22556,N_23937);
nor U29193 (N_29193,N_22839,N_20482);
or U29194 (N_29194,N_23203,N_22906);
nand U29195 (N_29195,N_20390,N_23418);
nor U29196 (N_29196,N_23541,N_24100);
or U29197 (N_29197,N_20856,N_21277);
nand U29198 (N_29198,N_21450,N_22827);
xnor U29199 (N_29199,N_21959,N_24087);
nand U29200 (N_29200,N_23971,N_21312);
or U29201 (N_29201,N_22444,N_23797);
or U29202 (N_29202,N_23525,N_21575);
or U29203 (N_29203,N_21663,N_21103);
xor U29204 (N_29204,N_23195,N_23483);
nor U29205 (N_29205,N_22602,N_22288);
xor U29206 (N_29206,N_23341,N_24296);
nand U29207 (N_29207,N_23615,N_24667);
nand U29208 (N_29208,N_24691,N_23816);
nor U29209 (N_29209,N_24801,N_22515);
xnor U29210 (N_29210,N_24941,N_22757);
and U29211 (N_29211,N_21260,N_22359);
nor U29212 (N_29212,N_22842,N_21581);
xor U29213 (N_29213,N_24290,N_21681);
xor U29214 (N_29214,N_23250,N_24878);
nand U29215 (N_29215,N_20161,N_22781);
or U29216 (N_29216,N_21340,N_21970);
xor U29217 (N_29217,N_20744,N_22853);
nor U29218 (N_29218,N_22110,N_23641);
nand U29219 (N_29219,N_21512,N_21793);
nor U29220 (N_29220,N_22742,N_24173);
and U29221 (N_29221,N_23834,N_24453);
xnor U29222 (N_29222,N_20316,N_21596);
nor U29223 (N_29223,N_24121,N_22390);
nand U29224 (N_29224,N_21367,N_22827);
or U29225 (N_29225,N_21976,N_22163);
or U29226 (N_29226,N_22833,N_21926);
or U29227 (N_29227,N_21505,N_22331);
and U29228 (N_29228,N_21821,N_23763);
xnor U29229 (N_29229,N_20591,N_21553);
nand U29230 (N_29230,N_20313,N_24837);
xnor U29231 (N_29231,N_23599,N_20575);
and U29232 (N_29232,N_24468,N_21327);
or U29233 (N_29233,N_23107,N_21138);
nor U29234 (N_29234,N_20030,N_20216);
or U29235 (N_29235,N_23137,N_24118);
and U29236 (N_29236,N_22680,N_24169);
and U29237 (N_29237,N_23571,N_24429);
and U29238 (N_29238,N_22476,N_24130);
xor U29239 (N_29239,N_22032,N_20854);
xor U29240 (N_29240,N_21123,N_22138);
and U29241 (N_29241,N_21067,N_22118);
and U29242 (N_29242,N_21833,N_23869);
and U29243 (N_29243,N_22782,N_24919);
nor U29244 (N_29244,N_22697,N_21027);
and U29245 (N_29245,N_21000,N_23223);
or U29246 (N_29246,N_21400,N_24762);
nor U29247 (N_29247,N_24563,N_21898);
or U29248 (N_29248,N_23148,N_20691);
and U29249 (N_29249,N_24535,N_24656);
or U29250 (N_29250,N_24200,N_22311);
xor U29251 (N_29251,N_23076,N_23721);
nor U29252 (N_29252,N_22771,N_21498);
nand U29253 (N_29253,N_23590,N_23712);
nand U29254 (N_29254,N_22859,N_20945);
and U29255 (N_29255,N_24435,N_22613);
nand U29256 (N_29256,N_21229,N_23536);
nand U29257 (N_29257,N_20515,N_20513);
or U29258 (N_29258,N_22995,N_21378);
nor U29259 (N_29259,N_21080,N_22242);
or U29260 (N_29260,N_24700,N_23494);
nor U29261 (N_29261,N_20549,N_24103);
or U29262 (N_29262,N_24560,N_23402);
nor U29263 (N_29263,N_22058,N_22591);
xor U29264 (N_29264,N_22257,N_24087);
or U29265 (N_29265,N_24183,N_24875);
xnor U29266 (N_29266,N_22487,N_20423);
or U29267 (N_29267,N_21890,N_23084);
nor U29268 (N_29268,N_23309,N_20338);
nand U29269 (N_29269,N_22438,N_24968);
and U29270 (N_29270,N_20030,N_20281);
xnor U29271 (N_29271,N_21929,N_23798);
and U29272 (N_29272,N_22867,N_21096);
xor U29273 (N_29273,N_20459,N_24228);
nor U29274 (N_29274,N_24020,N_24647);
nor U29275 (N_29275,N_24657,N_23223);
nand U29276 (N_29276,N_21997,N_24717);
or U29277 (N_29277,N_23587,N_21849);
or U29278 (N_29278,N_22285,N_21494);
nand U29279 (N_29279,N_23949,N_21481);
nor U29280 (N_29280,N_21142,N_23658);
or U29281 (N_29281,N_21901,N_23016);
or U29282 (N_29282,N_24194,N_24012);
xnor U29283 (N_29283,N_21715,N_21725);
and U29284 (N_29284,N_23399,N_23498);
nor U29285 (N_29285,N_23547,N_21632);
nand U29286 (N_29286,N_24644,N_23283);
xnor U29287 (N_29287,N_23862,N_22366);
xnor U29288 (N_29288,N_22091,N_24880);
and U29289 (N_29289,N_23019,N_22557);
or U29290 (N_29290,N_20565,N_20823);
nand U29291 (N_29291,N_22741,N_24484);
xnor U29292 (N_29292,N_23502,N_20883);
xnor U29293 (N_29293,N_23127,N_22841);
nand U29294 (N_29294,N_20556,N_20649);
or U29295 (N_29295,N_22120,N_22252);
xnor U29296 (N_29296,N_21720,N_20796);
nand U29297 (N_29297,N_23799,N_21466);
nor U29298 (N_29298,N_20197,N_24068);
or U29299 (N_29299,N_22893,N_23416);
or U29300 (N_29300,N_22460,N_22007);
and U29301 (N_29301,N_20034,N_21737);
or U29302 (N_29302,N_20340,N_24722);
nor U29303 (N_29303,N_20379,N_21444);
nand U29304 (N_29304,N_20261,N_24137);
or U29305 (N_29305,N_23638,N_23459);
nand U29306 (N_29306,N_22989,N_22110);
xor U29307 (N_29307,N_20830,N_21644);
xnor U29308 (N_29308,N_21341,N_23791);
xnor U29309 (N_29309,N_20115,N_20849);
nand U29310 (N_29310,N_22359,N_21491);
nand U29311 (N_29311,N_24863,N_20229);
nor U29312 (N_29312,N_20707,N_20599);
nand U29313 (N_29313,N_22172,N_23949);
nand U29314 (N_29314,N_23023,N_24800);
nand U29315 (N_29315,N_24788,N_23622);
and U29316 (N_29316,N_20478,N_22112);
nand U29317 (N_29317,N_20117,N_20481);
xnor U29318 (N_29318,N_20874,N_24822);
and U29319 (N_29319,N_23961,N_20080);
xor U29320 (N_29320,N_20226,N_20016);
or U29321 (N_29321,N_20677,N_20233);
nor U29322 (N_29322,N_22957,N_24588);
nor U29323 (N_29323,N_24361,N_23307);
xnor U29324 (N_29324,N_22705,N_22126);
nand U29325 (N_29325,N_23946,N_20048);
and U29326 (N_29326,N_22173,N_22764);
nor U29327 (N_29327,N_21623,N_21306);
nor U29328 (N_29328,N_20988,N_21794);
nand U29329 (N_29329,N_21488,N_24252);
nand U29330 (N_29330,N_20963,N_21375);
xnor U29331 (N_29331,N_24316,N_24496);
or U29332 (N_29332,N_22392,N_23710);
or U29333 (N_29333,N_24684,N_20193);
xnor U29334 (N_29334,N_24361,N_24365);
and U29335 (N_29335,N_20914,N_24344);
or U29336 (N_29336,N_23256,N_23792);
or U29337 (N_29337,N_23719,N_20463);
nor U29338 (N_29338,N_20610,N_23153);
nor U29339 (N_29339,N_21823,N_23703);
and U29340 (N_29340,N_20506,N_21447);
or U29341 (N_29341,N_20368,N_21218);
nand U29342 (N_29342,N_22079,N_21492);
and U29343 (N_29343,N_24156,N_20343);
nor U29344 (N_29344,N_23901,N_21436);
and U29345 (N_29345,N_23881,N_20833);
and U29346 (N_29346,N_24713,N_24959);
xor U29347 (N_29347,N_23063,N_24984);
xor U29348 (N_29348,N_21655,N_23773);
nand U29349 (N_29349,N_24861,N_20392);
nor U29350 (N_29350,N_23186,N_21851);
nand U29351 (N_29351,N_22028,N_23246);
xnor U29352 (N_29352,N_20430,N_20562);
nor U29353 (N_29353,N_24322,N_20827);
nor U29354 (N_29354,N_22133,N_20283);
xnor U29355 (N_29355,N_20134,N_23880);
or U29356 (N_29356,N_22496,N_23601);
and U29357 (N_29357,N_22649,N_21109);
or U29358 (N_29358,N_22090,N_22888);
and U29359 (N_29359,N_20075,N_21653);
nand U29360 (N_29360,N_20256,N_20711);
or U29361 (N_29361,N_21754,N_23559);
and U29362 (N_29362,N_22915,N_22107);
nand U29363 (N_29363,N_23876,N_24327);
or U29364 (N_29364,N_20232,N_22202);
and U29365 (N_29365,N_21779,N_24536);
nor U29366 (N_29366,N_20259,N_24132);
nor U29367 (N_29367,N_22681,N_23878);
or U29368 (N_29368,N_22390,N_22532);
or U29369 (N_29369,N_22222,N_22126);
nand U29370 (N_29370,N_23827,N_22447);
nor U29371 (N_29371,N_23334,N_23843);
and U29372 (N_29372,N_24946,N_22991);
nand U29373 (N_29373,N_22019,N_20203);
nor U29374 (N_29374,N_23901,N_23037);
nand U29375 (N_29375,N_21378,N_22714);
xnor U29376 (N_29376,N_20950,N_22368);
nor U29377 (N_29377,N_20191,N_20740);
nor U29378 (N_29378,N_24722,N_24339);
nor U29379 (N_29379,N_21503,N_20384);
nor U29380 (N_29380,N_20134,N_20082);
and U29381 (N_29381,N_21378,N_22907);
nand U29382 (N_29382,N_22837,N_21773);
and U29383 (N_29383,N_23612,N_22686);
nand U29384 (N_29384,N_24007,N_22580);
xor U29385 (N_29385,N_23255,N_21777);
or U29386 (N_29386,N_23645,N_24349);
and U29387 (N_29387,N_20549,N_23222);
nand U29388 (N_29388,N_22771,N_20713);
xor U29389 (N_29389,N_20246,N_22580);
nor U29390 (N_29390,N_23853,N_24353);
or U29391 (N_29391,N_21726,N_22108);
xnor U29392 (N_29392,N_21066,N_22976);
nor U29393 (N_29393,N_24681,N_24061);
nand U29394 (N_29394,N_21051,N_23268);
nor U29395 (N_29395,N_20456,N_20360);
and U29396 (N_29396,N_20132,N_20154);
nand U29397 (N_29397,N_21135,N_20871);
and U29398 (N_29398,N_23349,N_23464);
and U29399 (N_29399,N_20652,N_21941);
nor U29400 (N_29400,N_20275,N_20311);
xnor U29401 (N_29401,N_23006,N_20142);
nand U29402 (N_29402,N_23367,N_23448);
nor U29403 (N_29403,N_22516,N_23386);
xnor U29404 (N_29404,N_20130,N_23264);
xnor U29405 (N_29405,N_24487,N_23367);
nor U29406 (N_29406,N_20155,N_23021);
nor U29407 (N_29407,N_20920,N_20248);
and U29408 (N_29408,N_20723,N_23208);
or U29409 (N_29409,N_23877,N_21768);
nor U29410 (N_29410,N_23899,N_24045);
or U29411 (N_29411,N_24866,N_22774);
and U29412 (N_29412,N_23027,N_21344);
nor U29413 (N_29413,N_21986,N_23354);
nand U29414 (N_29414,N_21380,N_24629);
and U29415 (N_29415,N_21834,N_20133);
and U29416 (N_29416,N_22114,N_23263);
xor U29417 (N_29417,N_24958,N_21177);
and U29418 (N_29418,N_22598,N_20107);
or U29419 (N_29419,N_23746,N_20463);
and U29420 (N_29420,N_20401,N_22869);
xnor U29421 (N_29421,N_24872,N_21933);
or U29422 (N_29422,N_24391,N_23547);
and U29423 (N_29423,N_23975,N_21589);
nor U29424 (N_29424,N_24193,N_23275);
nand U29425 (N_29425,N_20064,N_22919);
nor U29426 (N_29426,N_20175,N_21924);
or U29427 (N_29427,N_23461,N_24110);
xor U29428 (N_29428,N_23706,N_21089);
nand U29429 (N_29429,N_21961,N_21009);
nand U29430 (N_29430,N_24208,N_24058);
and U29431 (N_29431,N_22037,N_22088);
and U29432 (N_29432,N_24885,N_24787);
and U29433 (N_29433,N_23345,N_24428);
and U29434 (N_29434,N_23882,N_24657);
nor U29435 (N_29435,N_21490,N_21759);
xor U29436 (N_29436,N_23756,N_21228);
xor U29437 (N_29437,N_20994,N_23270);
nor U29438 (N_29438,N_24620,N_24656);
or U29439 (N_29439,N_20971,N_20609);
nor U29440 (N_29440,N_23295,N_21539);
or U29441 (N_29441,N_21341,N_24759);
nand U29442 (N_29442,N_23039,N_20722);
xnor U29443 (N_29443,N_24328,N_21737);
xor U29444 (N_29444,N_23593,N_23190);
and U29445 (N_29445,N_20172,N_23390);
or U29446 (N_29446,N_20389,N_20141);
nand U29447 (N_29447,N_21461,N_22740);
nand U29448 (N_29448,N_23084,N_22218);
nand U29449 (N_29449,N_22653,N_20296);
nand U29450 (N_29450,N_21894,N_23672);
or U29451 (N_29451,N_23787,N_21842);
or U29452 (N_29452,N_23230,N_22659);
or U29453 (N_29453,N_24439,N_21492);
nand U29454 (N_29454,N_21719,N_24779);
or U29455 (N_29455,N_23547,N_20797);
or U29456 (N_29456,N_24832,N_20419);
nand U29457 (N_29457,N_23805,N_22984);
and U29458 (N_29458,N_21156,N_20099);
nor U29459 (N_29459,N_20626,N_23918);
nor U29460 (N_29460,N_20097,N_23046);
or U29461 (N_29461,N_24368,N_24716);
nand U29462 (N_29462,N_20998,N_21934);
nand U29463 (N_29463,N_21543,N_20014);
nand U29464 (N_29464,N_21733,N_24185);
or U29465 (N_29465,N_22491,N_23782);
or U29466 (N_29466,N_21792,N_21060);
and U29467 (N_29467,N_23574,N_24637);
nor U29468 (N_29468,N_21583,N_21039);
nand U29469 (N_29469,N_23461,N_23899);
xnor U29470 (N_29470,N_20464,N_20725);
and U29471 (N_29471,N_22013,N_21183);
xnor U29472 (N_29472,N_20655,N_20947);
or U29473 (N_29473,N_24549,N_20983);
xor U29474 (N_29474,N_24503,N_21929);
and U29475 (N_29475,N_20120,N_21679);
xnor U29476 (N_29476,N_22751,N_22299);
or U29477 (N_29477,N_21537,N_21878);
nand U29478 (N_29478,N_22026,N_21359);
nand U29479 (N_29479,N_22236,N_22205);
nor U29480 (N_29480,N_23849,N_21843);
nand U29481 (N_29481,N_20116,N_21576);
and U29482 (N_29482,N_22977,N_20805);
and U29483 (N_29483,N_21809,N_20400);
nand U29484 (N_29484,N_24249,N_20127);
xnor U29485 (N_29485,N_21646,N_20905);
nand U29486 (N_29486,N_20093,N_23012);
nor U29487 (N_29487,N_24378,N_20400);
nand U29488 (N_29488,N_21860,N_20791);
nor U29489 (N_29489,N_24624,N_20878);
and U29490 (N_29490,N_20836,N_20973);
and U29491 (N_29491,N_22736,N_21108);
nand U29492 (N_29492,N_22119,N_21444);
or U29493 (N_29493,N_24421,N_20779);
nor U29494 (N_29494,N_21138,N_23380);
or U29495 (N_29495,N_23623,N_22157);
or U29496 (N_29496,N_23033,N_20247);
nor U29497 (N_29497,N_23505,N_21193);
and U29498 (N_29498,N_20039,N_24276);
xor U29499 (N_29499,N_24975,N_20207);
and U29500 (N_29500,N_22596,N_21298);
or U29501 (N_29501,N_21823,N_22529);
or U29502 (N_29502,N_22450,N_21406);
or U29503 (N_29503,N_21908,N_22792);
and U29504 (N_29504,N_23771,N_22778);
xor U29505 (N_29505,N_22812,N_24466);
nand U29506 (N_29506,N_20210,N_24455);
or U29507 (N_29507,N_22531,N_24395);
nand U29508 (N_29508,N_21560,N_20062);
xor U29509 (N_29509,N_20327,N_23102);
xnor U29510 (N_29510,N_20059,N_24892);
and U29511 (N_29511,N_22248,N_20327);
and U29512 (N_29512,N_20059,N_22727);
nor U29513 (N_29513,N_21496,N_20520);
xor U29514 (N_29514,N_21326,N_24351);
nand U29515 (N_29515,N_21334,N_23525);
xor U29516 (N_29516,N_22503,N_21251);
xor U29517 (N_29517,N_21071,N_24911);
xnor U29518 (N_29518,N_22980,N_20880);
nand U29519 (N_29519,N_21290,N_20886);
or U29520 (N_29520,N_23089,N_24149);
or U29521 (N_29521,N_21842,N_23033);
xor U29522 (N_29522,N_21897,N_22419);
or U29523 (N_29523,N_22069,N_20323);
or U29524 (N_29524,N_23373,N_22629);
nor U29525 (N_29525,N_20273,N_24773);
or U29526 (N_29526,N_21801,N_20857);
xnor U29527 (N_29527,N_24558,N_23648);
or U29528 (N_29528,N_24727,N_22998);
nor U29529 (N_29529,N_20567,N_22249);
or U29530 (N_29530,N_23154,N_21901);
nor U29531 (N_29531,N_21042,N_22465);
xor U29532 (N_29532,N_22845,N_21026);
nor U29533 (N_29533,N_22032,N_20349);
or U29534 (N_29534,N_24378,N_22189);
nand U29535 (N_29535,N_21331,N_22342);
nand U29536 (N_29536,N_24580,N_24343);
or U29537 (N_29537,N_20344,N_20932);
or U29538 (N_29538,N_20687,N_23111);
nand U29539 (N_29539,N_24220,N_22952);
and U29540 (N_29540,N_21874,N_20125);
or U29541 (N_29541,N_24730,N_21751);
xnor U29542 (N_29542,N_21414,N_23910);
nand U29543 (N_29543,N_21677,N_21208);
or U29544 (N_29544,N_21123,N_23570);
xor U29545 (N_29545,N_21854,N_23773);
xnor U29546 (N_29546,N_24947,N_23902);
xnor U29547 (N_29547,N_23825,N_20577);
or U29548 (N_29548,N_23278,N_23207);
and U29549 (N_29549,N_21543,N_21764);
and U29550 (N_29550,N_21565,N_22241);
and U29551 (N_29551,N_24677,N_21047);
xor U29552 (N_29552,N_24795,N_24363);
nor U29553 (N_29553,N_22316,N_24197);
xor U29554 (N_29554,N_21338,N_20831);
or U29555 (N_29555,N_21904,N_21603);
xnor U29556 (N_29556,N_22468,N_24481);
or U29557 (N_29557,N_24537,N_23556);
xnor U29558 (N_29558,N_22166,N_24010);
and U29559 (N_29559,N_24494,N_21808);
nor U29560 (N_29560,N_20522,N_22048);
nor U29561 (N_29561,N_20617,N_23105);
xnor U29562 (N_29562,N_24509,N_21128);
and U29563 (N_29563,N_20125,N_23042);
nand U29564 (N_29564,N_22075,N_20148);
xor U29565 (N_29565,N_22379,N_22403);
xor U29566 (N_29566,N_20936,N_21369);
and U29567 (N_29567,N_20697,N_20829);
xnor U29568 (N_29568,N_20401,N_20949);
or U29569 (N_29569,N_24268,N_21702);
and U29570 (N_29570,N_22884,N_20909);
nor U29571 (N_29571,N_23391,N_21953);
or U29572 (N_29572,N_20432,N_21414);
and U29573 (N_29573,N_21602,N_20782);
and U29574 (N_29574,N_23060,N_20243);
and U29575 (N_29575,N_22784,N_20918);
and U29576 (N_29576,N_23782,N_21288);
nand U29577 (N_29577,N_22545,N_21606);
xor U29578 (N_29578,N_20656,N_21203);
nand U29579 (N_29579,N_20934,N_21046);
or U29580 (N_29580,N_20080,N_20820);
or U29581 (N_29581,N_24669,N_22871);
nand U29582 (N_29582,N_22577,N_21904);
or U29583 (N_29583,N_21754,N_20024);
or U29584 (N_29584,N_24745,N_20547);
nor U29585 (N_29585,N_23850,N_23733);
and U29586 (N_29586,N_24098,N_23101);
nand U29587 (N_29587,N_24984,N_20841);
and U29588 (N_29588,N_21206,N_24333);
nand U29589 (N_29589,N_22407,N_22122);
or U29590 (N_29590,N_21340,N_22062);
xnor U29591 (N_29591,N_24165,N_22061);
or U29592 (N_29592,N_24688,N_21905);
xor U29593 (N_29593,N_23269,N_20526);
or U29594 (N_29594,N_22993,N_20576);
and U29595 (N_29595,N_20729,N_20513);
nor U29596 (N_29596,N_24560,N_21407);
or U29597 (N_29597,N_23485,N_20613);
or U29598 (N_29598,N_21123,N_21854);
xnor U29599 (N_29599,N_21360,N_21032);
or U29600 (N_29600,N_21449,N_22320);
xnor U29601 (N_29601,N_24290,N_20748);
xor U29602 (N_29602,N_22792,N_21327);
nor U29603 (N_29603,N_24868,N_20148);
and U29604 (N_29604,N_24609,N_22083);
or U29605 (N_29605,N_21808,N_24578);
or U29606 (N_29606,N_23549,N_22791);
nand U29607 (N_29607,N_23776,N_21659);
nor U29608 (N_29608,N_23012,N_24988);
nand U29609 (N_29609,N_21505,N_20652);
nand U29610 (N_29610,N_23856,N_21504);
or U29611 (N_29611,N_21250,N_21915);
and U29612 (N_29612,N_24656,N_23385);
and U29613 (N_29613,N_22687,N_23103);
or U29614 (N_29614,N_20864,N_24542);
and U29615 (N_29615,N_23778,N_22370);
and U29616 (N_29616,N_22511,N_23090);
nand U29617 (N_29617,N_22740,N_20843);
and U29618 (N_29618,N_23540,N_23546);
nor U29619 (N_29619,N_21527,N_23433);
nor U29620 (N_29620,N_22129,N_20376);
and U29621 (N_29621,N_21935,N_20355);
and U29622 (N_29622,N_23004,N_21664);
nand U29623 (N_29623,N_20290,N_24582);
and U29624 (N_29624,N_24224,N_20710);
xnor U29625 (N_29625,N_20836,N_22702);
or U29626 (N_29626,N_23946,N_24066);
or U29627 (N_29627,N_23869,N_20334);
and U29628 (N_29628,N_20813,N_23376);
and U29629 (N_29629,N_24980,N_23071);
and U29630 (N_29630,N_21936,N_20236);
and U29631 (N_29631,N_22062,N_21515);
xnor U29632 (N_29632,N_23278,N_24201);
xor U29633 (N_29633,N_24244,N_22213);
or U29634 (N_29634,N_24345,N_23622);
nand U29635 (N_29635,N_20061,N_21978);
and U29636 (N_29636,N_20544,N_23695);
xnor U29637 (N_29637,N_22317,N_20579);
nor U29638 (N_29638,N_22032,N_24217);
nand U29639 (N_29639,N_22932,N_24152);
nor U29640 (N_29640,N_20008,N_23054);
or U29641 (N_29641,N_23209,N_23471);
nand U29642 (N_29642,N_23108,N_21500);
nand U29643 (N_29643,N_22375,N_20680);
xor U29644 (N_29644,N_20432,N_23179);
xor U29645 (N_29645,N_23253,N_21996);
and U29646 (N_29646,N_20917,N_21428);
or U29647 (N_29647,N_23104,N_20964);
or U29648 (N_29648,N_20064,N_20944);
or U29649 (N_29649,N_23764,N_20766);
xor U29650 (N_29650,N_21009,N_24014);
nand U29651 (N_29651,N_20821,N_21688);
nand U29652 (N_29652,N_22832,N_22450);
nand U29653 (N_29653,N_23411,N_20965);
nand U29654 (N_29654,N_21285,N_24548);
nor U29655 (N_29655,N_23195,N_23161);
nor U29656 (N_29656,N_21353,N_24250);
or U29657 (N_29657,N_20634,N_23882);
or U29658 (N_29658,N_20450,N_21870);
xnor U29659 (N_29659,N_20389,N_20507);
and U29660 (N_29660,N_20925,N_23852);
xnor U29661 (N_29661,N_22494,N_21346);
xnor U29662 (N_29662,N_22395,N_24521);
nand U29663 (N_29663,N_20576,N_20550);
or U29664 (N_29664,N_20011,N_24945);
nand U29665 (N_29665,N_21992,N_24546);
nor U29666 (N_29666,N_23854,N_22733);
and U29667 (N_29667,N_22554,N_20901);
nand U29668 (N_29668,N_23355,N_24172);
nand U29669 (N_29669,N_21953,N_23570);
and U29670 (N_29670,N_21468,N_22115);
nor U29671 (N_29671,N_21397,N_21725);
nor U29672 (N_29672,N_20065,N_23898);
xor U29673 (N_29673,N_23712,N_20994);
or U29674 (N_29674,N_23368,N_23661);
and U29675 (N_29675,N_20134,N_24129);
and U29676 (N_29676,N_20565,N_24357);
and U29677 (N_29677,N_23550,N_20508);
or U29678 (N_29678,N_21080,N_21334);
nand U29679 (N_29679,N_23494,N_24653);
or U29680 (N_29680,N_24132,N_24670);
or U29681 (N_29681,N_20845,N_20774);
and U29682 (N_29682,N_24106,N_24217);
and U29683 (N_29683,N_22350,N_22622);
and U29684 (N_29684,N_21141,N_23704);
and U29685 (N_29685,N_24278,N_21939);
nand U29686 (N_29686,N_23168,N_23710);
xor U29687 (N_29687,N_23605,N_24845);
nor U29688 (N_29688,N_24086,N_23793);
nor U29689 (N_29689,N_20304,N_22095);
nor U29690 (N_29690,N_22233,N_24063);
nor U29691 (N_29691,N_20152,N_24608);
and U29692 (N_29692,N_23154,N_22472);
nor U29693 (N_29693,N_20027,N_23720);
xnor U29694 (N_29694,N_20791,N_22553);
and U29695 (N_29695,N_22309,N_22088);
nor U29696 (N_29696,N_22187,N_22018);
nor U29697 (N_29697,N_23427,N_22198);
nand U29698 (N_29698,N_21922,N_22629);
xnor U29699 (N_29699,N_24020,N_23621);
nor U29700 (N_29700,N_22465,N_22418);
nand U29701 (N_29701,N_22093,N_24895);
nand U29702 (N_29702,N_21812,N_21452);
or U29703 (N_29703,N_22479,N_23409);
nand U29704 (N_29704,N_24242,N_20058);
nand U29705 (N_29705,N_20613,N_20087);
or U29706 (N_29706,N_23792,N_20446);
or U29707 (N_29707,N_23189,N_21780);
nand U29708 (N_29708,N_23118,N_23528);
xor U29709 (N_29709,N_23290,N_23592);
xor U29710 (N_29710,N_21339,N_24566);
or U29711 (N_29711,N_21363,N_20925);
nand U29712 (N_29712,N_24758,N_24444);
nor U29713 (N_29713,N_22114,N_22931);
xnor U29714 (N_29714,N_20075,N_22948);
nor U29715 (N_29715,N_24049,N_20301);
and U29716 (N_29716,N_23295,N_24300);
and U29717 (N_29717,N_20731,N_21045);
nor U29718 (N_29718,N_22821,N_20394);
nand U29719 (N_29719,N_23936,N_23559);
nor U29720 (N_29720,N_23992,N_23017);
and U29721 (N_29721,N_20670,N_24884);
nand U29722 (N_29722,N_22560,N_21953);
nor U29723 (N_29723,N_23004,N_20200);
nor U29724 (N_29724,N_21182,N_22457);
xor U29725 (N_29725,N_22452,N_24516);
or U29726 (N_29726,N_23867,N_23152);
and U29727 (N_29727,N_22907,N_21051);
xnor U29728 (N_29728,N_20971,N_24214);
or U29729 (N_29729,N_20003,N_23655);
or U29730 (N_29730,N_20562,N_24901);
and U29731 (N_29731,N_20008,N_20085);
nor U29732 (N_29732,N_23611,N_22545);
and U29733 (N_29733,N_24390,N_20366);
xor U29734 (N_29734,N_21688,N_21300);
and U29735 (N_29735,N_24679,N_24174);
nand U29736 (N_29736,N_24916,N_24702);
or U29737 (N_29737,N_20910,N_24739);
nor U29738 (N_29738,N_23181,N_23903);
nand U29739 (N_29739,N_23330,N_21406);
xnor U29740 (N_29740,N_20149,N_22572);
nand U29741 (N_29741,N_20357,N_23761);
and U29742 (N_29742,N_23205,N_23117);
nand U29743 (N_29743,N_24349,N_20164);
or U29744 (N_29744,N_23231,N_21470);
or U29745 (N_29745,N_24212,N_24969);
xnor U29746 (N_29746,N_23565,N_24559);
nand U29747 (N_29747,N_21928,N_21330);
or U29748 (N_29748,N_22107,N_21753);
and U29749 (N_29749,N_20478,N_21297);
nand U29750 (N_29750,N_20646,N_23182);
nor U29751 (N_29751,N_24607,N_24652);
nor U29752 (N_29752,N_21607,N_23358);
nor U29753 (N_29753,N_20388,N_21266);
nand U29754 (N_29754,N_23660,N_24956);
xnor U29755 (N_29755,N_22124,N_23109);
xor U29756 (N_29756,N_21995,N_24526);
nor U29757 (N_29757,N_24362,N_21956);
xor U29758 (N_29758,N_22184,N_22004);
or U29759 (N_29759,N_22908,N_21032);
or U29760 (N_29760,N_22251,N_21892);
xor U29761 (N_29761,N_24850,N_20703);
and U29762 (N_29762,N_23676,N_22954);
nand U29763 (N_29763,N_23344,N_23504);
xnor U29764 (N_29764,N_24818,N_23893);
nand U29765 (N_29765,N_20018,N_24446);
nand U29766 (N_29766,N_20004,N_24494);
xnor U29767 (N_29767,N_22581,N_21562);
or U29768 (N_29768,N_20653,N_23177);
or U29769 (N_29769,N_23736,N_24750);
or U29770 (N_29770,N_24089,N_22172);
xnor U29771 (N_29771,N_24291,N_22525);
or U29772 (N_29772,N_23008,N_23152);
nor U29773 (N_29773,N_21487,N_22677);
nand U29774 (N_29774,N_23069,N_22435);
or U29775 (N_29775,N_22658,N_21711);
nand U29776 (N_29776,N_22944,N_22857);
or U29777 (N_29777,N_23971,N_24140);
xor U29778 (N_29778,N_21898,N_23391);
or U29779 (N_29779,N_22509,N_20484);
nand U29780 (N_29780,N_22590,N_22136);
nand U29781 (N_29781,N_24127,N_23561);
nor U29782 (N_29782,N_20707,N_24317);
nand U29783 (N_29783,N_21593,N_22025);
nor U29784 (N_29784,N_20041,N_21171);
nand U29785 (N_29785,N_22710,N_20573);
or U29786 (N_29786,N_23213,N_24227);
or U29787 (N_29787,N_23794,N_21919);
and U29788 (N_29788,N_20951,N_23457);
xor U29789 (N_29789,N_20942,N_23432);
or U29790 (N_29790,N_23882,N_22995);
and U29791 (N_29791,N_23023,N_20004);
and U29792 (N_29792,N_21128,N_21067);
and U29793 (N_29793,N_23334,N_23697);
or U29794 (N_29794,N_24346,N_24307);
and U29795 (N_29795,N_20012,N_23722);
nand U29796 (N_29796,N_21849,N_22002);
and U29797 (N_29797,N_21016,N_21533);
nand U29798 (N_29798,N_21474,N_23351);
or U29799 (N_29799,N_24994,N_22183);
and U29800 (N_29800,N_22692,N_21656);
and U29801 (N_29801,N_22071,N_24494);
or U29802 (N_29802,N_20539,N_22237);
nor U29803 (N_29803,N_20076,N_24318);
xnor U29804 (N_29804,N_21593,N_23318);
nand U29805 (N_29805,N_20257,N_20441);
nor U29806 (N_29806,N_21229,N_20474);
nor U29807 (N_29807,N_20816,N_21848);
nor U29808 (N_29808,N_24515,N_21913);
and U29809 (N_29809,N_20674,N_24950);
and U29810 (N_29810,N_24607,N_24413);
and U29811 (N_29811,N_23528,N_23763);
nor U29812 (N_29812,N_22246,N_20694);
nand U29813 (N_29813,N_20530,N_20140);
nor U29814 (N_29814,N_22347,N_24382);
nor U29815 (N_29815,N_22698,N_24548);
nor U29816 (N_29816,N_21783,N_23155);
and U29817 (N_29817,N_20902,N_21254);
or U29818 (N_29818,N_22603,N_20321);
and U29819 (N_29819,N_24072,N_23782);
nand U29820 (N_29820,N_24756,N_21322);
and U29821 (N_29821,N_24609,N_23618);
nor U29822 (N_29822,N_22998,N_23763);
and U29823 (N_29823,N_22883,N_22448);
or U29824 (N_29824,N_20098,N_24885);
nand U29825 (N_29825,N_22722,N_21193);
nor U29826 (N_29826,N_22806,N_24127);
nand U29827 (N_29827,N_23732,N_20979);
xor U29828 (N_29828,N_21659,N_20658);
or U29829 (N_29829,N_20508,N_23300);
or U29830 (N_29830,N_24248,N_23363);
nand U29831 (N_29831,N_23098,N_20097);
nand U29832 (N_29832,N_20665,N_23379);
nor U29833 (N_29833,N_21286,N_23039);
or U29834 (N_29834,N_24296,N_21906);
or U29835 (N_29835,N_22852,N_24134);
xor U29836 (N_29836,N_22578,N_23681);
or U29837 (N_29837,N_21333,N_21093);
and U29838 (N_29838,N_21478,N_21780);
and U29839 (N_29839,N_23959,N_20232);
or U29840 (N_29840,N_24495,N_23967);
nand U29841 (N_29841,N_21222,N_24298);
nor U29842 (N_29842,N_22493,N_22226);
xor U29843 (N_29843,N_20538,N_22312);
xnor U29844 (N_29844,N_20983,N_23070);
or U29845 (N_29845,N_20509,N_24490);
or U29846 (N_29846,N_22645,N_20372);
nor U29847 (N_29847,N_20222,N_21187);
nor U29848 (N_29848,N_20333,N_22348);
and U29849 (N_29849,N_21193,N_20441);
xor U29850 (N_29850,N_21665,N_23914);
xnor U29851 (N_29851,N_22581,N_20042);
xor U29852 (N_29852,N_24523,N_24363);
xnor U29853 (N_29853,N_24302,N_20749);
nor U29854 (N_29854,N_20968,N_20236);
nor U29855 (N_29855,N_20907,N_22101);
or U29856 (N_29856,N_24443,N_21539);
nor U29857 (N_29857,N_22178,N_24237);
nand U29858 (N_29858,N_21710,N_23059);
or U29859 (N_29859,N_24571,N_21058);
xnor U29860 (N_29860,N_23631,N_23377);
xnor U29861 (N_29861,N_21915,N_21684);
or U29862 (N_29862,N_22724,N_24195);
or U29863 (N_29863,N_20875,N_24881);
or U29864 (N_29864,N_20813,N_20103);
or U29865 (N_29865,N_21358,N_22636);
and U29866 (N_29866,N_20033,N_21679);
xnor U29867 (N_29867,N_21788,N_21464);
or U29868 (N_29868,N_24134,N_24080);
nor U29869 (N_29869,N_24636,N_24784);
nor U29870 (N_29870,N_22184,N_23173);
nand U29871 (N_29871,N_22355,N_24377);
nor U29872 (N_29872,N_24341,N_20155);
nor U29873 (N_29873,N_22248,N_21996);
nor U29874 (N_29874,N_22696,N_21457);
xnor U29875 (N_29875,N_22773,N_23200);
xnor U29876 (N_29876,N_20806,N_20060);
xor U29877 (N_29877,N_23357,N_24279);
or U29878 (N_29878,N_21496,N_21563);
nor U29879 (N_29879,N_24226,N_20206);
or U29880 (N_29880,N_23120,N_24982);
or U29881 (N_29881,N_20139,N_20024);
and U29882 (N_29882,N_24131,N_22912);
or U29883 (N_29883,N_22254,N_23674);
and U29884 (N_29884,N_20841,N_24340);
nor U29885 (N_29885,N_23837,N_24307);
and U29886 (N_29886,N_21968,N_24156);
and U29887 (N_29887,N_22641,N_23987);
and U29888 (N_29888,N_22657,N_24818);
xnor U29889 (N_29889,N_22928,N_23367);
nand U29890 (N_29890,N_23163,N_21805);
and U29891 (N_29891,N_23777,N_23900);
and U29892 (N_29892,N_24805,N_20033);
nand U29893 (N_29893,N_22717,N_20027);
or U29894 (N_29894,N_22101,N_23122);
or U29895 (N_29895,N_23623,N_23693);
nand U29896 (N_29896,N_23783,N_23585);
and U29897 (N_29897,N_23241,N_23781);
nand U29898 (N_29898,N_23058,N_20214);
or U29899 (N_29899,N_21558,N_20966);
nand U29900 (N_29900,N_22927,N_20079);
xor U29901 (N_29901,N_21930,N_21645);
xnor U29902 (N_29902,N_21174,N_23054);
and U29903 (N_29903,N_23033,N_22597);
xnor U29904 (N_29904,N_21100,N_22836);
nand U29905 (N_29905,N_23250,N_23977);
and U29906 (N_29906,N_21185,N_21841);
xor U29907 (N_29907,N_21291,N_20757);
and U29908 (N_29908,N_24331,N_22822);
nor U29909 (N_29909,N_20921,N_24975);
and U29910 (N_29910,N_23404,N_20987);
or U29911 (N_29911,N_24681,N_20965);
nor U29912 (N_29912,N_22003,N_21190);
nor U29913 (N_29913,N_22823,N_24816);
or U29914 (N_29914,N_23335,N_22554);
nand U29915 (N_29915,N_24095,N_23917);
xor U29916 (N_29916,N_20428,N_22982);
nand U29917 (N_29917,N_22243,N_24688);
or U29918 (N_29918,N_21780,N_20786);
nor U29919 (N_29919,N_22197,N_24534);
xnor U29920 (N_29920,N_20742,N_23561);
and U29921 (N_29921,N_24416,N_22785);
or U29922 (N_29922,N_22011,N_22728);
nor U29923 (N_29923,N_21106,N_22746);
or U29924 (N_29924,N_24261,N_24047);
and U29925 (N_29925,N_21022,N_20335);
or U29926 (N_29926,N_23665,N_24675);
and U29927 (N_29927,N_21520,N_24810);
and U29928 (N_29928,N_20753,N_21829);
and U29929 (N_29929,N_23878,N_21420);
and U29930 (N_29930,N_20629,N_24374);
or U29931 (N_29931,N_22594,N_22170);
nor U29932 (N_29932,N_24528,N_22725);
and U29933 (N_29933,N_24700,N_20212);
nor U29934 (N_29934,N_23541,N_24619);
or U29935 (N_29935,N_24072,N_23956);
or U29936 (N_29936,N_22711,N_21868);
and U29937 (N_29937,N_24799,N_23535);
or U29938 (N_29938,N_22758,N_20153);
and U29939 (N_29939,N_21091,N_20331);
or U29940 (N_29940,N_21255,N_21119);
or U29941 (N_29941,N_24323,N_21096);
and U29942 (N_29942,N_21950,N_23442);
xor U29943 (N_29943,N_23099,N_20079);
and U29944 (N_29944,N_23188,N_24489);
nor U29945 (N_29945,N_24307,N_22211);
nor U29946 (N_29946,N_23971,N_23427);
and U29947 (N_29947,N_20157,N_24935);
or U29948 (N_29948,N_20562,N_22483);
nand U29949 (N_29949,N_20597,N_20462);
nand U29950 (N_29950,N_22106,N_23462);
xnor U29951 (N_29951,N_23761,N_21043);
and U29952 (N_29952,N_24683,N_24571);
xor U29953 (N_29953,N_20624,N_21856);
nand U29954 (N_29954,N_24656,N_24016);
nor U29955 (N_29955,N_21443,N_24108);
and U29956 (N_29956,N_23478,N_21509);
or U29957 (N_29957,N_24794,N_24991);
nand U29958 (N_29958,N_22077,N_22544);
or U29959 (N_29959,N_20811,N_20386);
nand U29960 (N_29960,N_24171,N_20173);
and U29961 (N_29961,N_24762,N_23837);
nand U29962 (N_29962,N_21021,N_21342);
xnor U29963 (N_29963,N_20097,N_23612);
and U29964 (N_29964,N_24864,N_24764);
nor U29965 (N_29965,N_21398,N_24179);
and U29966 (N_29966,N_20649,N_22646);
nor U29967 (N_29967,N_21810,N_23138);
nor U29968 (N_29968,N_20197,N_22037);
nor U29969 (N_29969,N_20624,N_21752);
and U29970 (N_29970,N_20952,N_21053);
and U29971 (N_29971,N_24290,N_21285);
nor U29972 (N_29972,N_21661,N_23130);
and U29973 (N_29973,N_23444,N_24575);
or U29974 (N_29974,N_24585,N_21066);
xor U29975 (N_29975,N_21443,N_23962);
xor U29976 (N_29976,N_24558,N_21351);
xor U29977 (N_29977,N_24796,N_23807);
and U29978 (N_29978,N_22690,N_22743);
and U29979 (N_29979,N_24554,N_24559);
or U29980 (N_29980,N_24024,N_24942);
nand U29981 (N_29981,N_21028,N_23282);
xor U29982 (N_29982,N_22974,N_21891);
nand U29983 (N_29983,N_22706,N_20841);
nor U29984 (N_29984,N_22969,N_24393);
and U29985 (N_29985,N_23714,N_23339);
nor U29986 (N_29986,N_20735,N_24795);
nor U29987 (N_29987,N_21384,N_21349);
xnor U29988 (N_29988,N_20187,N_22906);
nor U29989 (N_29989,N_23564,N_24559);
and U29990 (N_29990,N_24590,N_24507);
and U29991 (N_29991,N_20143,N_21794);
xnor U29992 (N_29992,N_24028,N_23063);
nor U29993 (N_29993,N_21689,N_22933);
or U29994 (N_29994,N_20499,N_22170);
nand U29995 (N_29995,N_24913,N_23734);
xnor U29996 (N_29996,N_24953,N_24512);
xor U29997 (N_29997,N_22643,N_21574);
nor U29998 (N_29998,N_22631,N_21556);
nor U29999 (N_29999,N_24574,N_22874);
and U30000 (N_30000,N_26644,N_26735);
nand U30001 (N_30001,N_27969,N_27184);
xnor U30002 (N_30002,N_25259,N_28697);
xnor U30003 (N_30003,N_26740,N_28759);
nand U30004 (N_30004,N_29691,N_26446);
and U30005 (N_30005,N_29704,N_28483);
and U30006 (N_30006,N_26168,N_29282);
nand U30007 (N_30007,N_25842,N_28803);
xor U30008 (N_30008,N_28149,N_29042);
xor U30009 (N_30009,N_28201,N_25454);
nor U30010 (N_30010,N_28033,N_25283);
or U30011 (N_30011,N_27636,N_28061);
nor U30012 (N_30012,N_27803,N_25479);
or U30013 (N_30013,N_25351,N_25589);
and U30014 (N_30014,N_28006,N_26177);
nor U30015 (N_30015,N_26943,N_26607);
and U30016 (N_30016,N_29799,N_29026);
xnor U30017 (N_30017,N_27880,N_25230);
or U30018 (N_30018,N_26890,N_28053);
nor U30019 (N_30019,N_28262,N_28980);
nand U30020 (N_30020,N_28232,N_28545);
and U30021 (N_30021,N_29615,N_26901);
nor U30022 (N_30022,N_29394,N_25848);
or U30023 (N_30023,N_27532,N_27280);
or U30024 (N_30024,N_26143,N_25244);
or U30025 (N_30025,N_27894,N_29240);
and U30026 (N_30026,N_28255,N_25622);
and U30027 (N_30027,N_28625,N_28039);
or U30028 (N_30028,N_27930,N_25973);
xnor U30029 (N_30029,N_26090,N_29851);
and U30030 (N_30030,N_25167,N_26336);
nor U30031 (N_30031,N_26785,N_25046);
or U30032 (N_30032,N_27733,N_29739);
nand U30033 (N_30033,N_29253,N_28674);
or U30034 (N_30034,N_26438,N_25918);
nand U30035 (N_30035,N_27629,N_26338);
nand U30036 (N_30036,N_25724,N_26781);
or U30037 (N_30037,N_26236,N_27093);
nand U30038 (N_30038,N_28455,N_27654);
or U30039 (N_30039,N_28692,N_25541);
xnor U30040 (N_30040,N_29568,N_28351);
or U30041 (N_30041,N_27186,N_27888);
and U30042 (N_30042,N_29450,N_27463);
nand U30043 (N_30043,N_29660,N_25129);
nor U30044 (N_30044,N_26344,N_29608);
or U30045 (N_30045,N_28133,N_29297);
or U30046 (N_30046,N_27817,N_29538);
and U30047 (N_30047,N_29056,N_25568);
nand U30048 (N_30048,N_28067,N_28983);
nor U30049 (N_30049,N_26179,N_28636);
and U30050 (N_30050,N_27064,N_29333);
xor U30051 (N_30051,N_28044,N_26967);
xor U30052 (N_30052,N_26492,N_26816);
and U30053 (N_30053,N_29051,N_26082);
nor U30054 (N_30054,N_28872,N_28529);
or U30055 (N_30055,N_25159,N_27163);
xnor U30056 (N_30056,N_25470,N_25325);
nand U30057 (N_30057,N_29870,N_29134);
and U30058 (N_30058,N_28215,N_28181);
nor U30059 (N_30059,N_25047,N_28454);
or U30060 (N_30060,N_28820,N_28842);
and U30061 (N_30061,N_27649,N_29596);
nor U30062 (N_30062,N_26135,N_25988);
xnor U30063 (N_30063,N_25342,N_27558);
nor U30064 (N_30064,N_26960,N_27068);
or U30065 (N_30065,N_26511,N_26879);
xor U30066 (N_30066,N_26889,N_25874);
xor U30067 (N_30067,N_26963,N_29111);
or U30068 (N_30068,N_28762,N_28038);
nand U30069 (N_30069,N_26340,N_25496);
xor U30070 (N_30070,N_28008,N_25742);
nor U30071 (N_30071,N_27597,N_26124);
xnor U30072 (N_30072,N_29569,N_28861);
nor U30073 (N_30073,N_26353,N_25088);
and U30074 (N_30074,N_26581,N_26831);
nand U30075 (N_30075,N_25916,N_28802);
nand U30076 (N_30076,N_27840,N_25465);
nor U30077 (N_30077,N_29182,N_27360);
xor U30078 (N_30078,N_29611,N_25243);
nor U30079 (N_30079,N_27049,N_27039);
and U30080 (N_30080,N_28945,N_25741);
and U30081 (N_30081,N_27397,N_29590);
and U30082 (N_30082,N_29554,N_27435);
and U30083 (N_30083,N_28113,N_28275);
nor U30084 (N_30084,N_27772,N_28942);
or U30085 (N_30085,N_28894,N_28757);
and U30086 (N_30086,N_26727,N_29278);
and U30087 (N_30087,N_29945,N_25793);
xor U30088 (N_30088,N_27099,N_26391);
nand U30089 (N_30089,N_27715,N_26563);
xnor U30090 (N_30090,N_25068,N_27094);
xnor U30091 (N_30091,N_25921,N_29120);
and U30092 (N_30092,N_26545,N_26473);
nand U30093 (N_30093,N_27077,N_29874);
or U30094 (N_30094,N_28378,N_25640);
nor U30095 (N_30095,N_29458,N_25662);
nor U30096 (N_30096,N_28306,N_27819);
nand U30097 (N_30097,N_27417,N_29939);
or U30098 (N_30098,N_28731,N_27838);
nand U30099 (N_30099,N_28429,N_25947);
and U30100 (N_30100,N_29213,N_25367);
or U30101 (N_30101,N_27992,N_28463);
and U30102 (N_30102,N_27546,N_26404);
or U30103 (N_30103,N_27524,N_25987);
and U30104 (N_30104,N_25080,N_29839);
nor U30105 (N_30105,N_28702,N_29141);
and U30106 (N_30106,N_25048,N_29369);
or U30107 (N_30107,N_28755,N_27506);
nor U30108 (N_30108,N_29571,N_28583);
and U30109 (N_30109,N_29299,N_27828);
or U30110 (N_30110,N_27850,N_29152);
nor U30111 (N_30111,N_29639,N_28564);
xnor U30112 (N_30112,N_25019,N_28587);
xnor U30113 (N_30113,N_25978,N_28093);
xor U30114 (N_30114,N_26462,N_25743);
and U30115 (N_30115,N_27698,N_28089);
and U30116 (N_30116,N_27413,N_27353);
xor U30117 (N_30117,N_26379,N_26799);
or U30118 (N_30118,N_28348,N_28316);
or U30119 (N_30119,N_28254,N_25285);
nand U30120 (N_30120,N_25762,N_25786);
and U30121 (N_30121,N_26623,N_28882);
and U30122 (N_30122,N_29508,N_29577);
and U30123 (N_30123,N_28616,N_26695);
nand U30124 (N_30124,N_29789,N_25008);
nor U30125 (N_30125,N_28209,N_29835);
or U30126 (N_30126,N_27909,N_26037);
and U30127 (N_30127,N_25029,N_25893);
and U30128 (N_30128,N_26771,N_25677);
nand U30129 (N_30129,N_28270,N_29429);
or U30130 (N_30130,N_28419,N_26742);
or U30131 (N_30131,N_27374,N_28117);
and U30132 (N_30132,N_26915,N_29700);
xnor U30133 (N_30133,N_25946,N_27403);
and U30134 (N_30134,N_27202,N_29613);
nor U30135 (N_30135,N_29309,N_28237);
nand U30136 (N_30136,N_29673,N_29880);
xnor U30137 (N_30137,N_28175,N_25968);
nand U30138 (N_30138,N_27644,N_26280);
nand U30139 (N_30139,N_25766,N_25820);
nand U30140 (N_30140,N_26657,N_26957);
nor U30141 (N_30141,N_29295,N_26940);
and U30142 (N_30142,N_28612,N_27499);
xor U30143 (N_30143,N_28108,N_29514);
xor U30144 (N_30144,N_28396,N_29667);
nand U30145 (N_30145,N_27661,N_25193);
and U30146 (N_30146,N_28100,N_28105);
xnor U30147 (N_30147,N_28163,N_25588);
xnor U30148 (N_30148,N_25369,N_28077);
nand U30149 (N_30149,N_29886,N_28952);
and U30150 (N_30150,N_29178,N_29387);
xor U30151 (N_30151,N_29216,N_29267);
nor U30152 (N_30152,N_26906,N_26579);
or U30153 (N_30153,N_27680,N_27950);
nand U30154 (N_30154,N_29517,N_27052);
and U30155 (N_30155,N_25992,N_25431);
xor U30156 (N_30156,N_26712,N_25180);
nor U30157 (N_30157,N_26204,N_25513);
nor U30158 (N_30158,N_27712,N_28049);
or U30159 (N_30159,N_29265,N_29787);
xnor U30160 (N_30160,N_29550,N_25179);
xnor U30161 (N_30161,N_27199,N_27272);
nor U30162 (N_30162,N_26567,N_25931);
nor U30163 (N_30163,N_25516,N_28600);
xnor U30164 (N_30164,N_26898,N_26639);
or U30165 (N_30165,N_25170,N_26628);
or U30166 (N_30166,N_26158,N_29579);
xor U30167 (N_30167,N_26346,N_27694);
or U30168 (N_30168,N_29620,N_29435);
or U30169 (N_30169,N_27875,N_25328);
nor U30170 (N_30170,N_27300,N_27309);
xor U30171 (N_30171,N_29200,N_27014);
and U30172 (N_30172,N_28214,N_29015);
nand U30173 (N_30173,N_29832,N_28888);
and U30174 (N_30174,N_28732,N_28588);
xor U30175 (N_30175,N_29259,N_29012);
xor U30176 (N_30176,N_27588,N_29499);
xor U30177 (N_30177,N_27935,N_28667);
xnor U30178 (N_30178,N_26128,N_26034);
or U30179 (N_30179,N_28937,N_29980);
nor U30180 (N_30180,N_29487,N_26621);
nor U30181 (N_30181,N_28460,N_28317);
and U30182 (N_30182,N_26948,N_27291);
xnor U30183 (N_30183,N_28357,N_27387);
and U30184 (N_30184,N_28442,N_28934);
and U30185 (N_30185,N_29208,N_27748);
nand U30186 (N_30186,N_26994,N_26064);
xnor U30187 (N_30187,N_28760,N_26660);
or U30188 (N_30188,N_29247,N_29630);
nor U30189 (N_30189,N_25688,N_27503);
or U30190 (N_30190,N_27356,N_27135);
nor U30191 (N_30191,N_28481,N_29441);
and U30192 (N_30192,N_29105,N_29558);
xnor U30193 (N_30193,N_28260,N_25349);
xor U30194 (N_30194,N_26384,N_25203);
nor U30195 (N_30195,N_26383,N_27329);
and U30196 (N_30196,N_27181,N_25954);
xor U30197 (N_30197,N_29676,N_26427);
nand U30198 (N_30198,N_26864,N_29541);
nand U30199 (N_30199,N_28459,N_28989);
nor U30200 (N_30200,N_28405,N_28308);
and U30201 (N_30201,N_28522,N_26116);
nor U30202 (N_30202,N_25854,N_28095);
xor U30203 (N_30203,N_26171,N_29128);
nor U30204 (N_30204,N_29266,N_28694);
nor U30205 (N_30205,N_26471,N_28103);
or U30206 (N_30206,N_28070,N_26424);
xnor U30207 (N_30207,N_27316,N_26920);
or U30208 (N_30208,N_25627,N_28532);
and U30209 (N_30209,N_25265,N_25616);
nor U30210 (N_30210,N_29380,N_28230);
nand U30211 (N_30211,N_29258,N_26038);
or U30212 (N_30212,N_28791,N_29697);
xnor U30213 (N_30213,N_28121,N_25052);
nor U30214 (N_30214,N_29674,N_26531);
and U30215 (N_30215,N_29588,N_26538);
nor U30216 (N_30216,N_27053,N_28533);
nor U30217 (N_30217,N_29388,N_28805);
and U30218 (N_30218,N_29201,N_28110);
nor U30219 (N_30219,N_25464,N_26672);
and U30220 (N_30220,N_29603,N_29055);
xor U30221 (N_30221,N_29275,N_25785);
or U30222 (N_30222,N_25288,N_28960);
nor U30223 (N_30223,N_29456,N_27368);
nand U30224 (N_30224,N_26369,N_29931);
or U30225 (N_30225,N_25530,N_29332);
and U30226 (N_30226,N_27660,N_29447);
nor U30227 (N_30227,N_29101,N_29474);
xnor U30228 (N_30228,N_29032,N_25683);
nor U30229 (N_30229,N_29918,N_27713);
nand U30230 (N_30230,N_28680,N_26618);
or U30231 (N_30231,N_26333,N_25885);
nor U30232 (N_30232,N_25495,N_28000);
nand U30233 (N_30233,N_25700,N_28489);
or U30234 (N_30234,N_29280,N_27630);
and U30235 (N_30235,N_27254,N_25957);
xor U30236 (N_30236,N_26812,N_27301);
or U30237 (N_30237,N_26578,N_25849);
nand U30238 (N_30238,N_28373,N_28783);
nor U30239 (N_30239,N_27378,N_25754);
or U30240 (N_30240,N_25482,N_29251);
or U30241 (N_30241,N_29898,N_28347);
or U30242 (N_30242,N_27340,N_26190);
and U30243 (N_30243,N_27210,N_26653);
nand U30244 (N_30244,N_26127,N_26325);
and U30245 (N_30245,N_27986,N_25308);
and U30246 (N_30246,N_25756,N_27668);
and U30247 (N_30247,N_25281,N_27284);
or U30248 (N_30248,N_27354,N_27573);
or U30249 (N_30249,N_25561,N_27615);
and U30250 (N_30250,N_29567,N_29402);
and U30251 (N_30251,N_26169,N_29338);
xnor U30252 (N_30252,N_28106,N_26520);
xnor U30253 (N_30253,N_26592,N_26480);
nor U30254 (N_30254,N_26700,N_25360);
xnor U30255 (N_30255,N_25703,N_27515);
nor U30256 (N_30256,N_27142,N_28575);
nand U30257 (N_30257,N_27814,N_27307);
or U30258 (N_30258,N_26780,N_27032);
xnor U30259 (N_30259,N_28366,N_28509);
xor U30260 (N_30260,N_26375,N_28136);
and U30261 (N_30261,N_26376,N_27616);
and U30262 (N_30262,N_25296,N_29304);
and U30263 (N_30263,N_25544,N_25016);
and U30264 (N_30264,N_29320,N_29059);
xnor U30265 (N_30265,N_25924,N_29595);
nor U30266 (N_30266,N_25022,N_29719);
or U30267 (N_30267,N_27991,N_25608);
and U30268 (N_30268,N_28838,N_27115);
nor U30269 (N_30269,N_29661,N_29927);
and U30270 (N_30270,N_29840,N_25376);
nand U30271 (N_30271,N_25933,N_27275);
and U30272 (N_30272,N_28372,N_27504);
xnor U30273 (N_30273,N_27355,N_25166);
nand U30274 (N_30274,N_26434,N_28258);
nor U30275 (N_30275,N_26223,N_25459);
xnor U30276 (N_30276,N_27213,N_25996);
nor U30277 (N_30277,N_27683,N_29405);
nor U30278 (N_30278,N_29188,N_27623);
nor U30279 (N_30279,N_28458,N_26077);
nand U30280 (N_30280,N_27187,N_29262);
nor U30281 (N_30281,N_25878,N_27574);
nand U30282 (N_30282,N_25485,N_25930);
xnor U30283 (N_30283,N_28046,N_25876);
xor U30284 (N_30284,N_28556,N_28431);
or U30285 (N_30285,N_28764,N_25261);
nand U30286 (N_30286,N_27790,N_28182);
nand U30287 (N_30287,N_26288,N_25660);
or U30288 (N_30288,N_27951,N_29680);
or U30289 (N_30289,N_26709,N_29283);
and U30290 (N_30290,N_28603,N_26356);
or U30291 (N_30291,N_26374,N_29484);
nand U30292 (N_30292,N_29720,N_27312);
or U30293 (N_30293,N_25447,N_25292);
nand U30294 (N_30294,N_25553,N_29688);
xnor U30295 (N_30295,N_26468,N_27200);
nand U30296 (N_30296,N_29656,N_28825);
xor U30297 (N_30297,N_25679,N_27366);
or U30298 (N_30298,N_27605,N_28524);
and U30299 (N_30299,N_28997,N_28924);
and U30300 (N_30300,N_25634,N_26410);
nand U30301 (N_30301,N_28804,N_28280);
xor U30302 (N_30302,N_26686,N_27205);
xnor U30303 (N_30303,N_26928,N_25737);
or U30304 (N_30304,N_26448,N_25260);
nand U30305 (N_30305,N_26795,N_25250);
nor U30306 (N_30306,N_27454,N_25215);
nand U30307 (N_30307,N_26897,N_29504);
xor U30308 (N_30308,N_25391,N_25307);
nor U30309 (N_30309,N_29138,N_29029);
nor U30310 (N_30310,N_29627,N_27973);
or U30311 (N_30311,N_26377,N_28024);
nand U30312 (N_30312,N_28915,N_29800);
nand U30313 (N_30313,N_29129,N_25739);
nor U30314 (N_30314,N_27678,N_27942);
and U30315 (N_30315,N_26066,N_29760);
nand U30316 (N_30316,N_29916,N_25663);
or U30317 (N_30317,N_29731,N_27161);
nand U30318 (N_30318,N_29073,N_29601);
nand U30319 (N_30319,N_27538,N_27544);
or U30320 (N_30320,N_27507,N_26568);
xnor U30321 (N_30321,N_28059,N_25934);
nand U30322 (N_30322,N_26396,N_29766);
and U30323 (N_30323,N_29996,N_27062);
or U30324 (N_30324,N_27686,N_28464);
or U30325 (N_30325,N_27826,N_27883);
and U30326 (N_30326,N_25770,N_27578);
or U30327 (N_30327,N_26313,N_26634);
nand U30328 (N_30328,N_25382,N_29825);
xor U30329 (N_30329,N_27138,N_28475);
or U30330 (N_30330,N_25542,N_29862);
nor U30331 (N_30331,N_27236,N_25975);
nand U30332 (N_30332,N_27019,N_26632);
and U30333 (N_30333,N_28987,N_29727);
xnor U30334 (N_30334,N_26242,N_26437);
and U30335 (N_30335,N_25582,N_26667);
or U30336 (N_30336,N_27079,N_28752);
and U30337 (N_30337,N_25729,N_28869);
nor U30338 (N_30338,N_25566,N_27137);
nor U30339 (N_30339,N_28144,N_26865);
nor U30340 (N_30340,N_26663,N_27857);
xnor U30341 (N_30341,N_28146,N_25249);
xnor U30342 (N_30342,N_26167,N_26266);
and U30343 (N_30343,N_27624,N_26662);
xor U30344 (N_30344,N_28452,N_26454);
nor U30345 (N_30345,N_26231,N_25084);
xor U30346 (N_30346,N_25735,N_27260);
xor U30347 (N_30347,N_28526,N_27839);
nor U30348 (N_30348,N_25337,N_27907);
or U30349 (N_30349,N_25038,N_29088);
nand U30350 (N_30350,N_26389,N_27610);
and U30351 (N_30351,N_28893,N_26845);
and U30352 (N_30352,N_26359,N_26944);
or U30353 (N_30353,N_26074,N_27044);
or U30354 (N_30354,N_29962,N_28437);
nand U30355 (N_30355,N_27865,N_27171);
xor U30356 (N_30356,N_27448,N_26707);
nor U30357 (N_30357,N_26729,N_28718);
xnor U30358 (N_30358,N_29077,N_25574);
xnor U30359 (N_30359,N_29664,N_25161);
or U30360 (N_30360,N_29049,N_27095);
and U30361 (N_30361,N_29445,N_27509);
nand U30362 (N_30362,N_26899,N_27553);
nand U30363 (N_30363,N_26256,N_26835);
nor U30364 (N_30364,N_27145,N_25081);
nor U30365 (N_30365,N_26238,N_26401);
and U30366 (N_30366,N_27432,N_29810);
or U30367 (N_30367,N_28268,N_25158);
xor U30368 (N_30368,N_29586,N_26832);
nor U30369 (N_30369,N_27483,N_25590);
or U30370 (N_30370,N_27427,N_29254);
and U30371 (N_30371,N_29008,N_29838);
nor U30372 (N_30372,N_26725,N_25149);
nand U30373 (N_30373,N_27781,N_26748);
nor U30374 (N_30374,N_26875,N_27600);
and U30375 (N_30375,N_26051,N_27031);
and U30376 (N_30376,N_28474,N_27144);
and U30377 (N_30377,N_26788,N_27394);
xor U30378 (N_30378,N_25644,N_28969);
or U30379 (N_30379,N_29775,N_25486);
xor U30380 (N_30380,N_27856,N_26393);
nand U30381 (N_30381,N_25466,N_27916);
and U30382 (N_30382,N_29533,N_29378);
nand U30383 (N_30383,N_28862,N_25870);
or U30384 (N_30384,N_26499,N_27794);
or U30385 (N_30385,N_27552,N_25286);
and U30386 (N_30386,N_28523,N_29413);
nand U30387 (N_30387,N_25945,N_28758);
or U30388 (N_30388,N_29273,N_27050);
nor U30389 (N_30389,N_26230,N_28127);
nand U30390 (N_30390,N_29035,N_25936);
nor U30391 (N_30391,N_26429,N_29334);
or U30392 (N_30392,N_26552,N_28245);
or U30393 (N_30393,N_28834,N_29118);
xor U30394 (N_30394,N_27167,N_26909);
or U30395 (N_30395,N_27297,N_29048);
and U30396 (N_30396,N_28909,N_28074);
xnor U30397 (N_30397,N_27811,N_28343);
nand U30398 (N_30398,N_28015,N_25626);
or U30399 (N_30399,N_27899,N_28076);
nand U30400 (N_30400,N_29342,N_27268);
xnor U30401 (N_30401,N_27286,N_27179);
nand U30402 (N_30402,N_27861,N_26642);
and U30403 (N_30403,N_27412,N_29665);
nor U30404 (N_30404,N_28822,N_26409);
nor U30405 (N_30405,N_28620,N_29854);
nand U30406 (N_30406,N_25314,N_27190);
nor U30407 (N_30407,N_28951,N_27570);
and U30408 (N_30408,N_25552,N_29235);
or U30409 (N_30409,N_26752,N_29867);
nor U30410 (N_30410,N_29606,N_29140);
nand U30411 (N_30411,N_28148,N_27306);
xor U30412 (N_30412,N_29797,N_29506);
nor U30413 (N_30413,N_29988,N_28361);
xor U30414 (N_30414,N_29167,N_28473);
and U30415 (N_30415,N_27807,N_28957);
or U30416 (N_30416,N_25102,N_29881);
and U30417 (N_30417,N_28013,N_29845);
and U30418 (N_30418,N_27734,N_29168);
nor U30419 (N_30419,N_28837,N_26883);
and U30420 (N_30420,N_25809,N_27218);
nor U30421 (N_30421,N_28516,N_25071);
nor U30422 (N_30422,N_26041,N_28300);
xnor U30423 (N_30423,N_25007,N_27714);
and U30424 (N_30424,N_26108,N_27441);
and U30425 (N_30425,N_26650,N_28827);
nand U30426 (N_30426,N_28828,N_29022);
nor U30427 (N_30427,N_26905,N_27024);
xnor U30428 (N_30428,N_26371,N_29855);
nand U30429 (N_30429,N_29805,N_26229);
or U30430 (N_30430,N_27317,N_27896);
nand U30431 (N_30431,N_26061,N_27549);
xor U30432 (N_30432,N_27554,N_25025);
and U30433 (N_30433,N_26274,N_25110);
or U30434 (N_30434,N_25607,N_29084);
and U30435 (N_30435,N_28104,N_27869);
xnor U30436 (N_30436,N_25818,N_27939);
nor U30437 (N_30437,N_28075,N_25753);
and U30438 (N_30438,N_26365,N_27735);
and U30439 (N_30439,N_26711,N_27350);
nor U30440 (N_30440,N_28427,N_28644);
and U30441 (N_30441,N_29328,N_28188);
nand U30442 (N_30442,N_27513,N_26951);
xor U30443 (N_30443,N_27622,N_26014);
nor U30444 (N_30444,N_27932,N_28001);
and U30445 (N_30445,N_29065,N_29423);
or U30446 (N_30446,N_27620,N_28841);
nor U30447 (N_30447,N_28173,N_25977);
and U30448 (N_30448,N_28398,N_29221);
nor U30449 (N_30449,N_25771,N_25136);
and U30450 (N_30450,N_29752,N_29462);
or U30451 (N_30451,N_25504,N_25605);
and U30452 (N_30452,N_27727,N_26458);
and U30453 (N_30453,N_29636,N_25652);
xor U30454 (N_30454,N_26301,N_26465);
or U30455 (N_30455,N_29205,N_28277);
or U30456 (N_30456,N_26512,N_25557);
or U30457 (N_30457,N_29373,N_28714);
xnor U30458 (N_30458,N_25415,N_25103);
or U30459 (N_30459,N_26170,N_28567);
nand U30460 (N_30460,N_27274,N_27569);
or U30461 (N_30461,N_25144,N_26507);
and U30462 (N_30462,N_27671,N_29733);
and U30463 (N_30463,N_29637,N_29856);
nand U30464 (N_30464,N_29281,N_26011);
nor U30465 (N_30465,N_25816,N_25023);
xnor U30466 (N_30466,N_25377,N_27116);
or U30467 (N_30467,N_29311,N_29543);
or U30468 (N_30468,N_29677,N_29893);
or U30469 (N_30469,N_27055,N_25448);
nand U30470 (N_30470,N_25419,N_27197);
nand U30471 (N_30471,N_26503,N_26858);
nor U30472 (N_30472,N_26351,N_28723);
xnor U30473 (N_30473,N_27607,N_29994);
xor U30474 (N_30474,N_29875,N_26922);
nor U30475 (N_30475,N_26271,N_25295);
nor U30476 (N_30476,N_28978,N_27711);
and U30477 (N_30477,N_25759,N_27005);
nor U30478 (N_30478,N_26586,N_29829);
or U30479 (N_30479,N_29316,N_27363);
and U30480 (N_30480,N_25814,N_28979);
xnor U30481 (N_30481,N_28307,N_29806);
xnor U30482 (N_30482,N_27957,N_27259);
or U30483 (N_30483,N_27122,N_26009);
or U30484 (N_30484,N_26387,N_29274);
xnor U30485 (N_30485,N_28767,N_29317);
and U30486 (N_30486,N_29807,N_29908);
or U30487 (N_30487,N_28456,N_28335);
nor U30488 (N_30488,N_29990,N_26100);
xor U30489 (N_30489,N_27905,N_28010);
or U30490 (N_30490,N_25256,N_25411);
and U30491 (N_30491,N_29699,N_25837);
nand U30492 (N_30492,N_26232,N_27723);
nand U30493 (N_30493,N_25014,N_25300);
xor U30494 (N_30494,N_29385,N_28507);
and U30495 (N_30495,N_29446,N_29969);
nor U30496 (N_30496,N_28678,N_27121);
nor U30497 (N_30497,N_26398,N_26562);
nor U30498 (N_30498,N_27114,N_25851);
or U30499 (N_30499,N_28699,N_28851);
and U30500 (N_30500,N_27423,N_25383);
nand U30501 (N_30501,N_25789,N_29477);
xor U30502 (N_30502,N_27343,N_27471);
nand U30503 (N_30503,N_29549,N_29072);
and U30504 (N_30504,N_26099,N_28530);
xnor U30505 (N_30505,N_25344,N_28712);
nor U30506 (N_30506,N_26872,N_25248);
xnor U30507 (N_30507,N_28213,N_25498);
and U30508 (N_30508,N_29301,N_25709);
nand U30509 (N_30509,N_28330,N_28115);
nand U30510 (N_30510,N_28400,N_26267);
nand U30511 (N_30511,N_29286,N_28040);
xnor U30512 (N_30512,N_28988,N_27180);
xnor U30513 (N_30513,N_26605,N_25392);
nor U30514 (N_30514,N_29315,N_28698);
nand U30515 (N_30515,N_27467,N_27217);
and U30516 (N_30516,N_28420,N_27691);
nand U30517 (N_30517,N_29237,N_27108);
or U30518 (N_30518,N_26968,N_29545);
nand U30519 (N_30519,N_28168,N_28928);
nand U30520 (N_30520,N_25503,N_28964);
nor U30521 (N_30521,N_29837,N_25073);
and U30522 (N_30522,N_28547,N_26123);
nand U30523 (N_30523,N_28897,N_26215);
nor U30524 (N_30524,N_27917,N_29811);
and U30525 (N_30525,N_25241,N_28795);
and U30526 (N_30526,N_26715,N_28319);
and U30527 (N_30527,N_27501,N_28025);
nor U30528 (N_30528,N_29119,N_25266);
or U30529 (N_30529,N_29928,N_29580);
and U30530 (N_30530,N_29657,N_27706);
xnor U30531 (N_30531,N_29229,N_25133);
and U30532 (N_30532,N_29634,N_27288);
or U30533 (N_30533,N_28299,N_25686);
xor U30534 (N_30534,N_27146,N_27771);
nand U30535 (N_30535,N_26850,N_27729);
nand U30536 (N_30536,N_25546,N_29609);
or U30537 (N_30537,N_28401,N_26322);
nand U30538 (N_30538,N_27994,N_29973);
xnor U30539 (N_30539,N_25755,N_26705);
nor U30540 (N_30540,N_29798,N_27999);
or U30541 (N_30541,N_29562,N_25824);
xnor U30542 (N_30542,N_27789,N_25026);
nand U30543 (N_30543,N_29058,N_25775);
and U30544 (N_30544,N_27362,N_26924);
and U30545 (N_30545,N_27183,N_26330);
nor U30546 (N_30546,N_28505,N_28511);
xnor U30547 (N_30547,N_26060,N_25155);
and U30548 (N_30548,N_28131,N_29284);
and U30549 (N_30549,N_27273,N_25699);
xnor U30550 (N_30550,N_25333,N_25746);
xnor U30551 (N_30551,N_27398,N_27744);
or U30552 (N_30552,N_29420,N_29436);
nor U30553 (N_30553,N_27380,N_29268);
nand U30554 (N_30554,N_27703,N_28637);
xor U30555 (N_30555,N_25698,N_28211);
and U30556 (N_30556,N_27601,N_26962);
xnor U30557 (N_30557,N_26980,N_26796);
or U30558 (N_30558,N_28309,N_26174);
nor U30559 (N_30559,N_29820,N_28810);
xnor U30560 (N_30560,N_28064,N_25252);
xnor U30561 (N_30561,N_29658,N_27603);
nand U30562 (N_30562,N_27681,N_27670);
nand U30563 (N_30563,N_26484,N_26008);
xor U30564 (N_30564,N_28261,N_25917);
nor U30565 (N_30565,N_27007,N_27018);
nand U30566 (N_30566,N_26400,N_27192);
xnor U30567 (N_30567,N_28471,N_25997);
nor U30568 (N_30568,N_28298,N_28655);
xnor U30569 (N_30569,N_27245,N_29644);
nand U30570 (N_30570,N_27089,N_26934);
nor U30571 (N_30571,N_29175,N_29864);
or U30572 (N_30572,N_29062,N_28036);
nand U30573 (N_30573,N_28514,N_29210);
nor U30574 (N_30574,N_25638,N_28424);
xor U30575 (N_30575,N_28051,N_29495);
or U30576 (N_30576,N_28501,N_29046);
nor U30577 (N_30577,N_27255,N_25435);
or U30578 (N_30578,N_28005,N_26591);
or U30579 (N_30579,N_25003,N_28026);
nor U30580 (N_30580,N_28495,N_29399);
nand U30581 (N_30581,N_28664,N_29848);
xnor U30582 (N_30582,N_25358,N_27141);
xor U30583 (N_30583,N_29001,N_26609);
or U30584 (N_30584,N_29233,N_25779);
xnor U30585 (N_30585,N_26991,N_26680);
nor U30586 (N_30586,N_25811,N_29375);
or U30587 (N_30587,N_27863,N_29750);
or U30588 (N_30588,N_27673,N_29386);
xor U30589 (N_30589,N_28063,N_25421);
and U30590 (N_30590,N_28439,N_26272);
or U30591 (N_30591,N_27963,N_27525);
xnor U30592 (N_30592,N_29147,N_27281);
nand U30593 (N_30593,N_29785,N_25163);
xnor U30594 (N_30594,N_27296,N_27438);
xnor U30595 (N_30595,N_25579,N_26031);
or U30596 (N_30596,N_26133,N_29871);
xor U30597 (N_30597,N_27119,N_25063);
nand U30598 (N_30598,N_28072,N_26857);
or U30599 (N_30599,N_28435,N_28352);
or U30600 (N_30600,N_27303,N_28387);
and U30601 (N_30601,N_27402,N_28118);
xor U30602 (N_30602,N_28407,N_29542);
xor U30603 (N_30603,N_29471,N_29245);
nor U30604 (N_30604,N_27746,N_29024);
nor U30605 (N_30605,N_26150,N_29411);
nor U30606 (N_30606,N_25475,N_29076);
nand U30607 (N_30607,N_27773,N_26988);
nand U30608 (N_30608,N_27822,N_27648);
xnor U30609 (N_30609,N_28441,N_26829);
or U30610 (N_30610,N_26422,N_29438);
nand U30611 (N_30611,N_25706,N_29747);
nor U30612 (N_30612,N_25390,N_26192);
nor U30613 (N_30613,N_25444,N_26390);
nor U30614 (N_30614,N_26938,N_26493);
xnor U30615 (N_30615,N_28303,N_28327);
and U30616 (N_30616,N_28745,N_28949);
or U30617 (N_30617,N_26360,N_29594);
xnor U30618 (N_30618,N_28037,N_29426);
nand U30619 (N_30619,N_26992,N_26608);
nor U30620 (N_30620,N_28286,N_27252);
nor U30621 (N_30621,N_28034,N_27204);
or U30622 (N_30622,N_29536,N_25711);
and U30623 (N_30623,N_28968,N_26076);
and U30624 (N_30624,N_25013,N_26868);
nand U30625 (N_30625,N_25752,N_28333);
xor U30626 (N_30626,N_28640,N_29707);
and U30627 (N_30627,N_28071,N_28374);
and U30628 (N_30628,N_27872,N_28295);
and U30629 (N_30629,N_25736,N_28773);
xor U30630 (N_30630,N_29773,N_28786);
xnor U30631 (N_30631,N_25558,N_29011);
or U30632 (N_30632,N_25125,N_26691);
nor U30633 (N_30633,N_29080,N_26881);
and U30634 (N_30634,N_29872,N_28681);
and U30635 (N_30635,N_29428,N_25646);
xor U30636 (N_30636,N_29947,N_26372);
nand U30637 (N_30637,N_26891,N_25011);
nor U30638 (N_30638,N_25116,N_29721);
nor U30639 (N_30639,N_29414,N_28058);
nor U30640 (N_30640,N_28189,N_28740);
or U30641 (N_30641,N_25798,N_29419);
nor U30642 (N_30642,N_26739,N_27365);
nor U30643 (N_30643,N_25725,N_26576);
nand U30644 (N_30644,N_27693,N_27310);
nor U30645 (N_30645,N_28832,N_25320);
nand U30646 (N_30646,N_26794,N_26260);
nand U30647 (N_30647,N_29986,N_28138);
nor U30648 (N_30648,N_28056,N_27010);
nor U30649 (N_30649,N_26624,N_27737);
nand U30650 (N_30650,N_25536,N_29381);
nand U30651 (N_30651,N_27975,N_28153);
xor U30652 (N_30652,N_27912,N_27396);
xnor U30653 (N_30653,N_25330,N_28833);
xnor U30654 (N_30654,N_26258,N_29687);
and U30655 (N_30655,N_28627,N_27662);
nand U30656 (N_30656,N_27550,N_27250);
and U30657 (N_30657,N_28933,N_27690);
and U30658 (N_30658,N_29597,N_27801);
and U30659 (N_30659,N_25247,N_27477);
nor U30660 (N_30660,N_28014,N_25153);
xnor U30661 (N_30661,N_26114,N_25359);
and U30662 (N_30662,N_25919,N_27731);
nand U30663 (N_30663,N_27923,N_25716);
and U30664 (N_30664,N_29144,N_28598);
and U30665 (N_30665,N_26678,N_29925);
or U30666 (N_30666,N_29091,N_27359);
and U30667 (N_30667,N_25697,N_26860);
nand U30668 (N_30668,N_27315,N_29057);
and U30669 (N_30669,N_29082,N_28778);
nor U30670 (N_30670,N_26057,N_29863);
nor U30671 (N_30671,N_26109,N_28320);
or U30672 (N_30672,N_26839,N_29751);
or U30673 (N_30673,N_27945,N_29983);
nor U30674 (N_30674,N_28226,N_29575);
nand U30675 (N_30675,N_26030,N_27647);
and U30676 (N_30676,N_29292,N_25976);
nor U30677 (N_30677,N_29288,N_27791);
xor U30678 (N_30678,N_25750,N_28187);
nand U30679 (N_30679,N_27589,N_26151);
xor U30680 (N_30680,N_26896,N_29228);
or U30681 (N_30681,N_27533,N_26277);
and U30682 (N_30682,N_27070,N_27617);
nand U30683 (N_30683,N_26362,N_26297);
nand U30684 (N_30684,N_27023,N_29028);
nand U30685 (N_30685,N_26855,N_28356);
nand U30686 (N_30686,N_28470,N_28701);
and U30687 (N_30687,N_27977,N_29043);
nand U30688 (N_30688,N_28923,N_27433);
xor U30689 (N_30689,N_25587,N_27765);
nor U30690 (N_30690,N_29515,N_26931);
xor U30691 (N_30691,N_26787,N_27220);
nor U30692 (N_30692,N_25757,N_26689);
xnor U30693 (N_30693,N_27972,N_27700);
nand U30694 (N_30694,N_28339,N_25598);
and U30695 (N_30695,N_27572,N_28650);
and U30696 (N_30696,N_28568,N_26674);
nor U30697 (N_30697,N_27168,N_29972);
nor U30698 (N_30698,N_27152,N_26193);
and U30699 (N_30699,N_25491,N_28635);
nor U30700 (N_30700,N_26106,N_28938);
xor U30701 (N_30701,N_26085,N_29250);
xor U30702 (N_30702,N_28011,N_28479);
or U30703 (N_30703,N_25580,N_28601);
nand U30704 (N_30704,N_27392,N_25623);
and U30705 (N_30705,N_28592,N_26055);
xnor U30706 (N_30706,N_25044,N_27189);
and U30707 (N_30707,N_25426,N_29982);
or U30708 (N_30708,N_29298,N_26958);
and U30709 (N_30709,N_27777,N_28683);
nand U30710 (N_30710,N_27760,N_29884);
or U30711 (N_30711,N_25302,N_28354);
nand U30712 (N_30712,N_26261,N_28311);
nand U30713 (N_30713,N_27021,N_26886);
and U30714 (N_30714,N_27347,N_26320);
or U30715 (N_30715,N_28843,N_28112);
or U30716 (N_30716,N_29628,N_27514);
nand U30717 (N_30717,N_28162,N_29177);
nand U30718 (N_30718,N_28634,N_26959);
nor U30719 (N_30719,N_29761,N_29834);
xor U30720 (N_30720,N_27124,N_29600);
nand U30721 (N_30721,N_25543,N_28709);
xor U30722 (N_30722,N_25601,N_28857);
or U30723 (N_30723,N_29291,N_26572);
and U30724 (N_30724,N_25443,N_25667);
or U30725 (N_30725,N_28519,N_26276);
nor U30726 (N_30726,N_29126,N_27277);
nor U30727 (N_30727,N_29464,N_29941);
and U30728 (N_30728,N_28436,N_28515);
and U30729 (N_30729,N_27674,N_26540);
nand U30730 (N_30730,N_26433,N_28101);
nor U30731 (N_30731,N_29424,N_25985);
xor U30732 (N_30732,N_26306,N_25118);
nand U30733 (N_30733,N_25902,N_28184);
or U30734 (N_30734,N_29643,N_26139);
nand U30735 (N_30735,N_25319,N_29079);
and U30736 (N_30736,N_25188,N_29729);
nand U30737 (N_30737,N_29061,N_27964);
nand U30738 (N_30738,N_26841,N_27873);
nor U30739 (N_30739,N_27450,N_26048);
nand U30740 (N_30740,N_29070,N_26824);
or U30741 (N_30741,N_28941,N_27475);
or U30742 (N_30742,N_28597,N_25445);
nor U30743 (N_30743,N_29307,N_29757);
xnor U30744 (N_30744,N_26766,N_27046);
nand U30745 (N_30745,N_28349,N_25284);
and U30746 (N_30746,N_28007,N_27004);
nand U30747 (N_30747,N_27484,N_27320);
xor U30748 (N_30748,N_28318,N_29276);
nor U30749 (N_30749,N_28743,N_29005);
or U30750 (N_30750,N_25887,N_26595);
or U30751 (N_30751,N_29344,N_26091);
nand U30752 (N_30752,N_27370,N_29393);
nor U30753 (N_30753,N_27029,N_25723);
nand U30754 (N_30754,N_25331,N_25437);
nor U30755 (N_30755,N_27054,N_28573);
xor U30756 (N_30756,N_26533,N_25540);
nor U30757 (N_30757,N_26601,N_26825);
and U30758 (N_30758,N_27565,N_28248);
nand U30759 (N_30759,N_26286,N_25480);
nor U30760 (N_30760,N_29121,N_27929);
or U30761 (N_30761,N_25903,N_29546);
nand U30762 (N_30762,N_29869,N_27290);
or U30763 (N_30763,N_26876,N_27786);
or U30764 (N_30764,N_29849,N_29907);
nor U30765 (N_30765,N_25471,N_29249);
nor U30766 (N_30766,N_27871,N_26734);
and U30767 (N_30767,N_26443,N_25657);
or U30768 (N_30768,N_25304,N_26428);
nor U30769 (N_30769,N_29507,N_26202);
and U30770 (N_30770,N_28465,N_28484);
xnor U30771 (N_30771,N_27422,N_27792);
nand U30772 (N_30772,N_26939,N_27984);
nor U30773 (N_30773,N_25339,N_25093);
xnor U30774 (N_30774,N_28098,N_26494);
nand U30775 (N_30775,N_27747,N_29479);
xnor U30776 (N_30776,N_26370,N_26873);
and U30777 (N_30777,N_29778,N_25104);
and U30778 (N_30778,N_27389,N_27799);
or U30779 (N_30779,N_27540,N_28741);
nor U30780 (N_30780,N_25629,N_27824);
nand U30781 (N_30781,N_29584,N_29148);
nand U30782 (N_30782,N_26862,N_26341);
xnor U30783 (N_30783,N_28534,N_27762);
nor U30784 (N_30784,N_25593,N_25142);
nand U30785 (N_30785,N_27908,N_27188);
and U30786 (N_30786,N_27289,N_25922);
nor U30787 (N_30787,N_25907,N_25473);
or U30788 (N_30788,N_29942,N_29416);
or U30789 (N_30789,N_28331,N_25412);
nand U30790 (N_30790,N_25920,N_25335);
or U30791 (N_30791,N_27443,N_27103);
nand U30792 (N_30792,N_29192,N_29331);
nand U30793 (N_30793,N_26045,N_26923);
nor U30794 (N_30794,N_29553,N_26145);
nor U30795 (N_30795,N_28744,N_25141);
xor U30796 (N_30796,N_25317,N_29525);
or U30797 (N_30797,N_25615,N_27854);
or U30798 (N_30798,N_27906,N_28028);
nor U30799 (N_30799,N_25612,N_26050);
or U30800 (N_30800,N_29713,N_28648);
or U30801 (N_30801,N_26243,N_25056);
nand U30802 (N_30802,N_26765,N_27716);
nor U30803 (N_30803,N_28630,N_26853);
or U30804 (N_30804,N_25915,N_25050);
nor U30805 (N_30805,N_28030,N_29964);
xor U30806 (N_30806,N_25625,N_26852);
nand U30807 (N_30807,N_25108,N_26191);
xor U30808 (N_30808,N_27480,N_25474);
nand U30809 (N_30809,N_28898,N_28705);
and U30810 (N_30810,N_27710,N_27947);
and U30811 (N_30811,N_25855,N_27851);
nor U30812 (N_30812,N_27439,N_28614);
nor U30813 (N_30813,N_28687,N_26447);
xor U30814 (N_30814,N_25365,N_27655);
or U30815 (N_30815,N_29155,N_27314);
and U30816 (N_30816,N_26413,N_29570);
nand U30817 (N_30817,N_28571,N_27174);
nand U30818 (N_30818,N_29053,N_29696);
nand U30819 (N_30819,N_26355,N_26300);
xor U30820 (N_30820,N_25520,N_26289);
xnor U30821 (N_30821,N_26483,N_29768);
nor U30822 (N_30822,N_27372,N_25417);
nand U30823 (N_30823,N_25597,N_28297);
xnor U30824 (N_30824,N_27754,N_28658);
nand U30825 (N_30825,N_28961,N_25151);
nor U30826 (N_30826,N_28212,N_29762);
nand U30827 (N_30827,N_29374,N_26095);
nor U30828 (N_30828,N_28272,N_26324);
xnor U30829 (N_30829,N_27566,N_27720);
or U30830 (N_30830,N_29407,N_28932);
nand U30831 (N_30831,N_25935,N_26786);
xnor U30832 (N_30832,N_26436,N_29186);
xor U30833 (N_30833,N_26757,N_26815);
or U30834 (N_30834,N_25143,N_25150);
nand U30835 (N_30835,N_25669,N_27755);
and U30836 (N_30836,N_26637,N_26081);
and U30837 (N_30837,N_28443,N_29968);
nand U30838 (N_30838,N_26987,N_26509);
and U30839 (N_30839,N_26210,N_28027);
nor U30840 (N_30840,N_29003,N_29367);
xnor U30841 (N_30841,N_29455,N_29649);
and U30842 (N_30842,N_29965,N_26874);
nor U30843 (N_30843,N_27743,N_27575);
nor U30844 (N_30844,N_27222,N_27057);
or U30845 (N_30845,N_25272,N_25617);
nor U30846 (N_30846,N_25087,N_25653);
or U30847 (N_30847,N_28386,N_28581);
and U30848 (N_30848,N_27421,N_27842);
and U30849 (N_30849,N_27749,N_25406);
and U30850 (N_30850,N_25800,N_29777);
xnor U30851 (N_30851,N_27618,N_27692);
nor U30852 (N_30852,N_28881,N_27993);
nand U30853 (N_30853,N_28726,N_29009);
nand U30854 (N_30854,N_29725,N_26087);
nor U30855 (N_30855,N_28264,N_25363);
xnor U30856 (N_30856,N_25097,N_29626);
xnor U30857 (N_30857,N_28555,N_26200);
xnor U30858 (N_30858,N_29472,N_26183);
nand U30859 (N_30859,N_25943,N_28194);
or U30860 (N_30860,N_27913,N_25713);
xor U30861 (N_30861,N_26073,N_29345);
nand U30862 (N_30862,N_27976,N_29547);
xnor U30863 (N_30863,N_25461,N_28021);
xnor U30864 (N_30864,N_26016,N_26452);
xnor U30865 (N_30865,N_27379,N_29622);
and U30866 (N_30866,N_25511,N_29578);
nand U30867 (N_30867,N_26541,N_25324);
and U30868 (N_30868,N_28411,N_29544);
nand U30869 (N_30869,N_29503,N_28643);
nor U30870 (N_30870,N_26535,N_28346);
or U30871 (N_30871,N_28641,N_26933);
and U30872 (N_30872,N_27944,N_29842);
nor U30873 (N_30873,N_26088,N_28922);
nand U30874 (N_30874,N_28946,N_27891);
nand U30875 (N_30875,N_27949,N_29348);
and U30876 (N_30876,N_28416,N_29976);
nor U30877 (N_30877,N_29432,N_27830);
and U30878 (N_30878,N_29104,N_28780);
nand U30879 (N_30879,N_27383,N_27488);
or U30880 (N_30880,N_28735,N_29937);
or U30881 (N_30881,N_28904,N_29002);
or U30882 (N_30882,N_25280,N_28651);
nor U30883 (N_30883,N_27965,N_28700);
nor U30884 (N_30884,N_27160,N_28737);
and U30885 (N_30885,N_27322,N_29242);
and U30886 (N_30886,N_26803,N_25214);
or U30887 (N_30887,N_29623,N_27261);
or U30888 (N_30888,N_26665,N_26884);
xnor U30889 (N_30889,N_26626,N_27225);
and U30890 (N_30890,N_27640,N_25720);
and U30891 (N_30891,N_28563,N_26635);
nand U30892 (N_30892,N_25500,N_25705);
nand U30893 (N_30893,N_25940,N_26764);
xnor U30894 (N_30894,N_26806,N_29052);
or U30895 (N_30895,N_29075,N_26554);
and U30896 (N_30896,N_28130,N_27299);
nand U30897 (N_30897,N_28935,N_28242);
xnor U30898 (N_30898,N_28809,N_29710);
or U30899 (N_30899,N_28632,N_28608);
nor U30900 (N_30900,N_25956,N_26585);
and U30901 (N_30901,N_27669,N_25695);
xnor U30902 (N_30902,N_26759,N_25969);
nand U30903 (N_30903,N_26307,N_25010);
or U30904 (N_30904,N_25323,N_26062);
nand U30905 (N_30905,N_25210,N_27967);
nand U30906 (N_30906,N_26640,N_27495);
or U30907 (N_30907,N_26453,N_25949);
nand U30908 (N_30908,N_29183,N_25613);
nand U30909 (N_30909,N_27319,N_27282);
nor U30910 (N_30910,N_27983,N_27140);
nand U30911 (N_30911,N_29788,N_28180);
and U30912 (N_30912,N_28128,N_26756);
or U30913 (N_30913,N_25298,N_26187);
and U30914 (N_30914,N_28662,N_25032);
and U30915 (N_30915,N_28649,N_25501);
nor U30916 (N_30916,N_25184,N_25955);
and U30917 (N_30917,N_29173,N_26063);
nand U30918 (N_30918,N_28665,N_26791);
and U30919 (N_30919,N_29176,N_28369);
xor U30920 (N_30920,N_25195,N_27593);
nand U30921 (N_30921,N_26583,N_28457);
and U30922 (N_30922,N_25115,N_29277);
xor U30923 (N_30923,N_26137,N_27738);
xor U30924 (N_30924,N_28537,N_29793);
or U30925 (N_30925,N_28294,N_29502);
nand U30926 (N_30926,N_25747,N_29362);
xnor U30927 (N_30927,N_27173,N_29217);
or U30928 (N_30928,N_26357,N_29290);
nor U30929 (N_30929,N_27521,N_25092);
or U30930 (N_30930,N_29616,N_26012);
xor U30931 (N_30931,N_25374,N_28126);
xnor U30932 (N_30932,N_29404,N_27915);
nand U30933 (N_30933,N_25799,N_28596);
or U30934 (N_30934,N_29459,N_28375);
and U30935 (N_30935,N_29031,N_27453);
xor U30936 (N_30936,N_26826,N_26015);
or U30937 (N_30937,N_25594,N_27584);
nand U30938 (N_30938,N_25694,N_29532);
nor U30939 (N_30939,N_25575,N_26685);
nor U30940 (N_30940,N_25276,N_25439);
and U30941 (N_30941,N_26347,N_29654);
and U30942 (N_30942,N_26518,N_25453);
and U30943 (N_30943,N_26775,N_28761);
nand U30944 (N_30944,N_29748,N_26590);
nand U30945 (N_30945,N_28565,N_25661);
nand U30946 (N_30946,N_27555,N_29363);
xnor U30947 (N_30947,N_29439,N_26560);
xnor U30948 (N_30948,N_29199,N_29765);
nor U30949 (N_30949,N_25506,N_26440);
or U30950 (N_30950,N_29364,N_25847);
xnor U30951 (N_30951,N_25472,N_26040);
and U30952 (N_30952,N_27002,N_28642);
or U30953 (N_30953,N_28660,N_27757);
or U30954 (N_30954,N_29153,N_25291);
xnor U30955 (N_30955,N_26871,N_27881);
nor U30956 (N_30956,N_29561,N_28719);
or U30957 (N_30957,N_27219,N_25532);
nor U30958 (N_30958,N_29422,N_27581);
nor U30959 (N_30959,N_27808,N_28217);
xor U30960 (N_30960,N_29264,N_27591);
xor U30961 (N_30961,N_25578,N_25114);
and U30962 (N_30962,N_27332,N_27958);
or U30963 (N_30963,N_26054,N_28210);
and U30964 (N_30964,N_27292,N_29180);
nor U30965 (N_30965,N_29260,N_28677);
and U30966 (N_30966,N_26971,N_28769);
nand U30967 (N_30967,N_29564,N_26681);
or U30968 (N_30968,N_28956,N_29006);
or U30969 (N_30969,N_29071,N_25145);
and U30970 (N_30970,N_27472,N_29534);
xor U30971 (N_30971,N_29904,N_25487);
and U30972 (N_30972,N_27346,N_29675);
and U30973 (N_30973,N_27056,N_29212);
or U30974 (N_30974,N_29555,N_25378);
xnor U30975 (N_30975,N_25828,N_29163);
nand U30976 (N_30976,N_28273,N_29230);
xor U30977 (N_30977,N_26136,N_25024);
xnor U30978 (N_30978,N_27627,N_26487);
nor U30979 (N_30979,N_29802,N_29818);
xnor U30980 (N_30980,N_28925,N_29759);
and U30981 (N_30981,N_27086,N_29531);
and U30982 (N_30982,N_27326,N_28754);
and U30983 (N_30983,N_28382,N_26245);
xnor U30984 (N_30984,N_29470,N_28288);
and U30985 (N_30985,N_25321,N_25238);
nand U30986 (N_30986,N_29647,N_25299);
nor U30987 (N_30987,N_28498,N_29826);
nand U30988 (N_30988,N_27511,N_27568);
nand U30989 (N_30989,N_26597,N_28675);
nor U30990 (N_30990,N_25539,N_29137);
xnor U30991 (N_30991,N_28686,N_25883);
xnor U30992 (N_30992,N_25217,N_29844);
nor U30993 (N_30993,N_29158,N_29860);
nor U30994 (N_30994,N_26878,N_29852);
xnor U30995 (N_30995,N_29758,N_25704);
nand U30996 (N_30996,N_28151,N_27318);
xnor U30997 (N_30997,N_28233,N_29556);
or U30998 (N_30998,N_29497,N_27221);
or U30999 (N_30999,N_25869,N_27175);
and U31000 (N_31000,N_25373,N_25463);
or U31001 (N_31001,N_26309,N_26569);
or U31002 (N_31002,N_28388,N_28913);
nand U31003 (N_31003,N_26577,N_29901);
nand U31004 (N_31004,N_27416,N_28859);
nand U31005 (N_31005,N_25895,N_28972);
nor U31006 (N_31006,N_26003,N_27076);
and U31007 (N_31007,N_25614,N_25185);
or U31008 (N_31008,N_27265,N_25732);
or U31009 (N_31009,N_27845,N_28850);
nor U31010 (N_31010,N_28906,N_29734);
nor U31011 (N_31011,N_28304,N_26750);
xor U31012 (N_31012,N_26588,N_26761);
or U31013 (N_31013,N_29007,N_26270);
nor U31014 (N_31014,N_25730,N_26194);
nand U31015 (N_31015,N_25126,N_29511);
xor U31016 (N_31016,N_27742,N_29287);
or U31017 (N_31017,N_26698,N_26810);
nand U31018 (N_31018,N_25549,N_28165);
or U31019 (N_31019,N_26599,N_26559);
nor U31020 (N_31020,N_26439,N_28224);
and U31021 (N_31021,N_28191,N_25689);
or U31022 (N_31022,N_28315,N_27352);
nor U31023 (N_31023,N_29958,N_25168);
or U31024 (N_31024,N_25565,N_28976);
xor U31025 (N_31025,N_28055,N_29261);
and U31026 (N_31026,N_29598,N_29431);
nor U31027 (N_31027,N_26547,N_25131);
xnor U31028 (N_31028,N_28525,N_28018);
or U31029 (N_31029,N_25106,N_29081);
xnor U31030 (N_31030,N_26264,N_28503);
and U31031 (N_31031,N_28970,N_27836);
xnor U31032 (N_31032,N_27542,N_28394);
xor U31033 (N_31033,N_29631,N_26528);
or U31034 (N_31034,N_26932,N_25127);
nand U31035 (N_31035,N_29485,N_28559);
xnor U31036 (N_31036,N_28549,N_25676);
or U31037 (N_31037,N_26543,N_29489);
xnor U31038 (N_31038,N_28535,N_29368);
nor U31039 (N_31039,N_27635,N_28240);
xor U31040 (N_31040,N_26246,N_26582);
or U31041 (N_31041,N_28751,N_28445);
or U31042 (N_31042,N_25400,N_26373);
nor U31043 (N_31043,N_27904,N_27474);
and U31044 (N_31044,N_26273,N_25791);
nor U31045 (N_31045,N_25297,N_29984);
and U31046 (N_31046,N_26394,N_25821);
nand U31047 (N_31047,N_25316,N_29724);
or U31048 (N_31048,N_26488,N_26403);
nand U31049 (N_31049,N_26159,N_25122);
nand U31050 (N_31050,N_26500,N_25389);
or U31051 (N_31051,N_25422,N_25993);
or U31052 (N_31052,N_28541,N_27240);
or U31053 (N_31053,N_28283,N_29961);
xnor U31054 (N_31054,N_25687,N_28599);
xor U31055 (N_31055,N_29565,N_25960);
nor U31056 (N_31056,N_29231,N_26848);
nor U31057 (N_31057,N_26774,N_29382);
xnor U31058 (N_31058,N_26767,N_26821);
nor U31059 (N_31059,N_26070,N_25112);
and U31060 (N_31060,N_25424,N_29302);
nor U31061 (N_31061,N_29911,N_28003);
nor U31062 (N_31062,N_25031,N_27580);
xnor U31063 (N_31063,N_26762,N_26104);
nor U31064 (N_31064,N_28950,N_26046);
nand U31065 (N_31065,N_28080,N_29524);
or U31066 (N_31066,N_26047,N_29457);
xnor U31067 (N_31067,N_25733,N_27677);
or U31068 (N_31068,N_27809,N_29343);
and U31069 (N_31069,N_28943,N_27780);
and U31070 (N_31070,N_26112,N_25654);
nand U31071 (N_31071,N_27696,N_25803);
or U31072 (N_31072,N_27106,N_26334);
nor U31073 (N_31073,N_26703,N_25006);
xor U31074 (N_31074,N_25182,N_28875);
nor U31075 (N_31075,N_26161,N_29756);
nand U31076 (N_31076,N_25564,N_27704);
nor U31077 (N_31077,N_25051,N_26993);
xnor U31078 (N_31078,N_28707,N_25751);
and U31079 (N_31079,N_28340,N_26198);
nand U31080 (N_31080,N_26225,N_29529);
nor U31081 (N_31081,N_25066,N_28708);
and U31082 (N_31082,N_25176,N_27582);
nand U31083 (N_31083,N_27741,N_27996);
or U31084 (N_31084,N_26544,N_28012);
or U31085 (N_31085,N_29038,N_25229);
nand U31086 (N_31086,N_28205,N_25991);
xor U31087 (N_31087,N_25591,N_26702);
and U31088 (N_31088,N_26565,N_27015);
or U31089 (N_31089,N_27130,N_27264);
and U31090 (N_31090,N_28633,N_26203);
nand U31091 (N_31091,N_27249,N_27779);
or U31092 (N_31092,N_25618,N_26444);
xor U31093 (N_31093,N_27371,N_27242);
nand U31094 (N_31094,N_26949,N_27428);
and U31095 (N_31095,N_28812,N_27424);
and U31096 (N_31096,N_28561,N_25387);
nor U31097 (N_31097,N_28421,N_27980);
nand U31098 (N_31098,N_27464,N_26420);
nor U31099 (N_31099,N_25223,N_29746);
or U31100 (N_31100,N_25372,N_25226);
xnor U31101 (N_31101,N_26316,N_26275);
and U31102 (N_31102,N_29093,N_29563);
nor U31103 (N_31103,N_25727,N_26425);
nand U31104 (N_31104,N_28493,N_25191);
xnor U31105 (N_31105,N_27345,N_28392);
nor U31106 (N_31106,N_28231,N_26546);
nand U31107 (N_31107,N_25889,N_26804);
or U31108 (N_31108,N_26348,N_28995);
nor U31109 (N_31109,N_26807,N_26648);
and U31110 (N_31110,N_27892,N_25805);
or U31111 (N_31111,N_27736,N_29360);
or U31112 (N_31112,N_27682,N_25442);
nand U31113 (N_31113,N_26553,N_27498);
and U31114 (N_31114,N_28150,N_27726);
or U31115 (N_31115,N_25577,N_28787);
nor U31116 (N_31116,N_29113,N_25666);
xor U31117 (N_31117,N_25290,N_28155);
nor U31118 (N_31118,N_25624,N_29410);
xor U31119 (N_31119,N_25021,N_26455);
and U31120 (N_31120,N_29225,N_27890);
and U31121 (N_31121,N_27756,N_25483);
and U31122 (N_31122,N_27385,N_28434);
or U31123 (N_31123,N_25147,N_29913);
and U31124 (N_31124,N_25213,N_27596);
xnor U31125 (N_31125,N_29906,N_25986);
and U31126 (N_31126,N_25478,N_28926);
xnor U31127 (N_31127,N_26721,N_28917);
xor U31128 (N_31128,N_25524,N_28669);
and U31129 (N_31129,N_28779,N_27604);
and U31130 (N_31130,N_26737,N_28724);
and U31131 (N_31131,N_29635,N_27434);
and U31132 (N_31132,N_27695,N_26078);
or U31133 (N_31133,N_27061,N_26950);
xor U31134 (N_31134,N_28646,N_25364);
xor U31135 (N_31135,N_28123,N_27877);
nor U31136 (N_31136,N_25277,N_29125);
nand U31137 (N_31137,N_26141,N_26007);
nand U31138 (N_31138,N_25758,N_27800);
xnor U31139 (N_31139,N_27675,N_27098);
or U31140 (N_31140,N_26773,N_26910);
or U31141 (N_31141,N_29895,N_25875);
and U31142 (N_31142,N_28239,N_25585);
nor U31143 (N_31143,N_26318,N_27882);
nor U31144 (N_31144,N_29589,N_27020);
or U31145 (N_31145,N_26587,N_29841);
nor U31146 (N_31146,N_28876,N_28993);
or U31147 (N_31147,N_28808,N_26677);
xnor U31148 (N_31148,N_26984,N_25899);
or U31149 (N_31149,N_25682,N_28244);
or U31150 (N_31150,N_25109,N_27758);
and U31151 (N_31151,N_26432,N_25707);
nand U31152 (N_31152,N_27063,N_27928);
xor U31153 (N_31153,N_26321,N_25547);
or U31154 (N_31154,N_27833,N_26570);
and U31155 (N_31155,N_28661,N_26205);
nand U31156 (N_31156,N_28204,N_25722);
nor U31157 (N_31157,N_29786,N_27375);
or U31158 (N_31158,N_26122,N_29383);
xor U31159 (N_31159,N_27287,N_29858);
or U31160 (N_31160,N_29612,N_27941);
nand U31161 (N_31161,N_29496,N_25963);
xor U31162 (N_31162,N_29692,N_27341);
xnor U31163 (N_31163,N_25420,N_28880);
nand U31164 (N_31164,N_29823,N_26475);
xor U31165 (N_31165,N_27527,N_26813);
nor U31166 (N_31166,N_27369,N_26633);
nand U31167 (N_31167,N_25512,N_26305);
and U31168 (N_31168,N_28716,N_28878);
nor U31169 (N_31169,N_28595,N_29943);
and U31170 (N_31170,N_25018,N_29833);
and U31171 (N_31171,N_29572,N_29132);
nor U31172 (N_31172,N_25348,N_27599);
or U31173 (N_31173,N_28679,N_28579);
and U31174 (N_31174,N_27411,N_28984);
xor U31175 (N_31175,N_28418,N_28856);
nand U31176 (N_31176,N_27665,N_27585);
or U31177 (N_31177,N_25499,N_26147);
and U31178 (N_31178,N_29351,N_26697);
nand U31179 (N_31179,N_25091,N_29790);
nor U31180 (N_31180,N_29873,N_26854);
or U31181 (N_31181,N_27399,N_25132);
nor U31182 (N_31182,N_27058,N_29443);
nor U31183 (N_31183,N_29776,N_25278);
and U31184 (N_31184,N_27769,N_29741);
and U31185 (N_31185,N_26399,N_29678);
or U31186 (N_31186,N_28364,N_28826);
and U31187 (N_31187,N_29461,N_29108);
or U31188 (N_31188,N_28908,N_29979);
xor U31189 (N_31189,N_25456,N_27430);
and U31190 (N_31190,N_27974,N_27490);
and U31191 (N_31191,N_28141,N_26188);
nand U31192 (N_31192,N_25611,N_25990);
and U31193 (N_31193,N_28721,N_29668);
nand U31194 (N_31194,N_28611,N_29321);
and U31195 (N_31195,N_26701,N_29574);
xnor U31196 (N_31196,N_25356,N_26110);
nand U31197 (N_31197,N_25740,N_27798);
nand U31198 (N_31198,N_26990,N_28256);
xor U31199 (N_31199,N_27602,N_25815);
nor U31200 (N_31200,N_27216,N_25177);
or U31201 (N_31201,N_28433,N_29509);
nor U31202 (N_31202,N_27156,N_26838);
nand U31203 (N_31203,N_28771,N_27613);
and U31204 (N_31204,N_29679,N_26602);
nand U31205 (N_31205,N_28504,N_29551);
or U31206 (N_31206,N_28066,N_26975);
and U31207 (N_31207,N_26534,N_27446);
nand U31208 (N_31208,N_29891,N_28377);
nor U31209 (N_31209,N_29139,N_26522);
xnor U31210 (N_31210,N_25649,N_26255);
nor U31211 (N_31211,N_27386,N_28385);
and U31212 (N_31212,N_25015,N_28606);
nor U31213 (N_31213,N_25839,N_26751);
or U31214 (N_31214,N_27870,N_29530);
nand U31215 (N_31215,N_27619,N_27985);
nor U31216 (N_31216,N_25900,N_28654);
or U31217 (N_31217,N_28219,N_27926);
nand U31218 (N_31218,N_26925,N_29040);
nand U31219 (N_31219,N_26134,N_26331);
nor U31220 (N_31220,N_25827,N_25866);
nand U31221 (N_31221,N_25888,N_28874);
xor U31222 (N_31222,N_25525,N_28252);
xor U31223 (N_31223,N_28114,N_26052);
or U31224 (N_31224,N_26615,N_28999);
xor U31225 (N_31225,N_29083,N_29325);
xnor U31226 (N_31226,N_27164,N_26970);
nand U31227 (N_31227,N_25064,N_28032);
nor U31228 (N_31228,N_28276,N_29279);
nor U31229 (N_31229,N_29560,N_29819);
or U31230 (N_31230,N_29094,N_28328);
or U31231 (N_31231,N_27279,N_28570);
and U31232 (N_31232,N_29744,N_28520);
and U31233 (N_31233,N_25813,N_25251);
nor U31234 (N_31234,N_29483,N_26028);
nand U31235 (N_31235,N_29828,N_25645);
or U31236 (N_31236,N_27751,N_26733);
nor U31237 (N_31237,N_28365,N_28480);
and U31238 (N_31238,N_25418,N_25535);
or U31239 (N_31239,N_26589,N_25076);
and U31240 (N_31240,N_25562,N_25070);
xor U31241 (N_31241,N_26481,N_28855);
and U31242 (N_31242,N_25710,N_28982);
nor U31243 (N_31243,N_25332,N_29770);
nor U31244 (N_31244,N_25484,N_28543);
xor U31245 (N_31245,N_26102,N_25650);
xnor U31246 (N_31246,N_25979,N_26557);
xnor U31247 (N_31247,N_27793,N_29950);
or U31248 (N_31248,N_25892,N_25772);
nor U31249 (N_31249,N_26652,N_27110);
nor U31250 (N_31250,N_26973,N_26622);
and U31251 (N_31251,N_29535,N_26000);
nand U31252 (N_31252,N_25165,N_28914);
xnor U31253 (N_31253,N_28781,N_28353);
and U31254 (N_31254,N_29944,N_29406);
or U31255 (N_31255,N_25187,N_29415);
xor U31256 (N_31256,N_29218,N_29935);
and U31257 (N_31257,N_26335,N_29060);
nor U31258 (N_31258,N_27285,N_27111);
or U31259 (N_31259,N_25000,N_27404);
nor U31260 (N_31260,N_27128,N_25207);
and U31261 (N_31261,N_25749,N_27409);
and U31262 (N_31262,N_29593,N_27129);
nand U31263 (N_31263,N_29467,N_25637);
nor U31264 (N_31264,N_26747,N_26496);
or U31265 (N_31265,N_28497,N_25310);
xnor U31266 (N_31266,N_29671,N_25450);
xnor U31267 (N_31267,N_29460,N_25967);
or U31268 (N_31268,N_25164,N_26593);
nand U31269 (N_31269,N_27051,N_29822);
nor U31270 (N_31270,N_25428,N_27278);
nand U31271 (N_31271,N_27982,N_25432);
xor U31272 (N_31272,N_26946,N_25218);
xnor U31273 (N_31273,N_28954,N_28111);
nor U31274 (N_31274,N_28048,N_29468);
or U31275 (N_31275,N_28253,N_28147);
nand U31276 (N_31276,N_26421,N_26279);
and U31277 (N_31277,N_25181,N_28414);
and U31278 (N_31278,N_26817,N_25235);
xor U31279 (N_31279,N_27230,N_26699);
xor U31280 (N_31280,N_26779,N_25404);
xnor U31281 (N_31281,N_26079,N_26388);
nor U31282 (N_31282,N_27123,N_27535);
and U31283 (N_31283,N_26094,N_27834);
nand U31284 (N_31284,N_28393,N_29803);
and U31285 (N_31285,N_28236,N_29357);
nand U31286 (N_31286,N_28102,N_27571);
nand U31287 (N_31287,N_29526,N_25160);
xnor U31288 (N_31288,N_27223,N_26163);
nor U31289 (N_31289,N_28466,N_26929);
and U31290 (N_31290,N_27238,N_28207);
nand U31291 (N_31291,N_29449,N_28250);
or U31292 (N_31292,N_25085,N_27829);
or U31293 (N_31293,N_27959,N_29149);
or U31294 (N_31294,N_27096,N_27666);
or U31295 (N_31295,N_27539,N_28296);
xnor U31296 (N_31296,N_26029,N_29926);
nor U31297 (N_31297,N_27821,N_26326);
nor U31298 (N_31298,N_26178,N_29683);
nand U31299 (N_31299,N_27784,N_25830);
xor U31300 (N_31300,N_26176,N_26117);
and U31301 (N_31301,N_25861,N_25079);
xor U31302 (N_31302,N_28527,N_26498);
nor U31303 (N_31303,N_25228,N_28586);
and U31304 (N_31304,N_28860,N_26527);
or U31305 (N_31305,N_25303,N_27672);
or U31306 (N_31306,N_29993,N_29463);
or U31307 (N_31307,N_28107,N_25477);
or U31308 (N_31308,N_25844,N_26361);
xnor U31309 (N_31309,N_27783,N_25877);
nand U31310 (N_31310,N_27088,N_29753);
and U31311 (N_31311,N_25556,N_26596);
nor U31312 (N_31312,N_28510,N_29041);
xor U31313 (N_31313,N_27026,N_29136);
and U31314 (N_31314,N_26416,N_28593);
xor U31315 (N_31315,N_29241,N_27276);
or U31316 (N_31316,N_28817,N_29095);
nor U31317 (N_31317,N_28866,N_28367);
xor U31318 (N_31318,N_28412,N_29505);
xnor U31319 (N_31319,N_26730,N_29064);
xor U31320 (N_31320,N_25647,N_27782);
and U31321 (N_31321,N_29066,N_27775);
xnor U31322 (N_31322,N_26688,N_25951);
nor U31323 (N_31323,N_25041,N_25884);
and U31324 (N_31324,N_25401,N_25734);
nor U31325 (N_31325,N_25961,N_28799);
xor U31326 (N_31326,N_26160,N_29619);
or U31327 (N_31327,N_25769,N_26919);
or U31328 (N_31328,N_29184,N_29256);
or U31329 (N_31329,N_28770,N_28506);
or U31330 (N_31330,N_27717,N_28462);
xor U31331 (N_31331,N_28167,N_26184);
xor U31332 (N_31332,N_29706,N_29949);
xnor U31333 (N_31333,N_25192,N_29189);
nor U31334 (N_31334,N_28301,N_25595);
and U31335 (N_31335,N_26329,N_29581);
xor U31336 (N_31336,N_28814,N_28886);
xor U31337 (N_31337,N_25551,N_29151);
nand U31338 (N_31338,N_26113,N_26490);
nand U31339 (N_31339,N_25846,N_26972);
nor U31340 (N_31340,N_27961,N_28449);
or U31341 (N_31341,N_26743,N_29641);
xor U31342 (N_31342,N_26319,N_25206);
and U31343 (N_31343,N_29648,N_28792);
nor U31344 (N_31344,N_29607,N_25531);
or U31345 (N_31345,N_25570,N_25656);
or U31346 (N_31346,N_28122,N_27406);
nor U31347 (N_31347,N_29194,N_29159);
xnor U31348 (N_31348,N_27813,N_28746);
xnor U31349 (N_31349,N_27447,N_26426);
nor U31350 (N_31350,N_27889,N_25355);
and U31351 (N_31351,N_28727,N_28944);
or U31352 (N_31352,N_25908,N_29701);
xnor U31353 (N_31353,N_27331,N_27159);
and U31354 (N_31354,N_26892,N_27001);
or U31355 (N_31355,N_25274,N_28806);
xnor U31356 (N_31356,N_27536,N_28087);
or U31357 (N_31357,N_27445,N_25178);
nand U31358 (N_31358,N_29723,N_25077);
and U31359 (N_31359,N_27528,N_29179);
and U31360 (N_31360,N_25095,N_29978);
and U31361 (N_31361,N_28196,N_25264);
xor U31362 (N_31362,N_26182,N_29602);
xnor U31363 (N_31363,N_26366,N_28513);
and U31364 (N_31364,N_29488,N_27455);
nand U31365 (N_31365,N_27853,N_27866);
or U31366 (N_31366,N_28129,N_28602);
xor U31367 (N_31367,N_28734,N_29164);
nor U31368 (N_31368,N_26284,N_27642);
xor U31369 (N_31369,N_28607,N_28800);
or U31370 (N_31370,N_25642,N_25829);
and U31371 (N_31371,N_26887,N_27810);
and U31372 (N_31372,N_26119,N_27377);
or U31373 (N_31373,N_26478,N_27494);
nor U31374 (N_31374,N_27583,N_25675);
or U31375 (N_31375,N_25836,N_26291);
nor U31376 (N_31376,N_28550,N_25891);
or U31377 (N_31377,N_29882,N_26148);
nand U31378 (N_31378,N_26263,N_26523);
or U31379 (N_31379,N_28499,N_25246);
nand U31380 (N_31380,N_27943,N_25045);
nor U31381 (N_31381,N_27646,N_26604);
xnor U31382 (N_31382,N_28830,N_27466);
xor U31383 (N_31383,N_26842,N_28220);
nand U31384 (N_31384,N_29754,N_28623);
xnor U31385 (N_31385,N_29078,N_25287);
xor U31386 (N_31386,N_25438,N_26186);
nor U31387 (N_31387,N_26402,N_25490);
and U31388 (N_31388,N_27764,N_27017);
nor U31389 (N_31389,N_28363,N_25005);
nand U31390 (N_31390,N_26822,N_26684);
nand U31391 (N_31391,N_28312,N_26154);
xor U31392 (N_31392,N_29246,N_26075);
nand U31393 (N_31393,N_25911,N_26783);
nor U31394 (N_31394,N_26658,N_28613);
and U31395 (N_31395,N_29716,N_28895);
nor U31396 (N_31396,N_26718,N_25510);
or U31397 (N_31397,N_25001,N_26996);
or U31398 (N_31398,N_29359,N_29592);
nand U31399 (N_31399,N_28553,N_25405);
and U31400 (N_31400,N_28444,N_26798);
or U31401 (N_31401,N_27770,N_27069);
and U31402 (N_31402,N_28671,N_27305);
nor U31403 (N_31403,N_25146,N_26530);
nand U31404 (N_31404,N_25950,N_26467);
nand U31405 (N_31405,N_25345,N_27937);
xnor U31406 (N_31406,N_25731,N_26129);
xor U31407 (N_31407,N_26647,N_28195);
nand U31408 (N_31408,N_26671,N_28417);
or U31409 (N_31409,N_27587,N_27656);
or U31410 (N_31410,N_27479,N_27653);
nand U31411 (N_31411,N_25099,N_26669);
nand U31412 (N_31412,N_29621,N_28689);
nor U31413 (N_31413,N_25493,N_25172);
or U31414 (N_31414,N_25926,N_28912);
and U31415 (N_31415,N_28161,N_28358);
nor U31416 (N_31416,N_25995,N_27611);
nand U31417 (N_31417,N_27505,N_26978);
xnor U31418 (N_31418,N_28574,N_29518);
or U31419 (N_31419,N_26278,N_27632);
nand U31420 (N_31420,N_29133,N_26625);
or U31421 (N_31421,N_26310,N_29528);
xor U31422 (N_31422,N_29004,N_27083);
or U31423 (N_31423,N_29646,N_27832);
nor U31424 (N_31424,N_27657,N_26019);
or U31425 (N_31425,N_29824,N_29143);
xor U31426 (N_31426,N_25999,N_29255);
nand U31427 (N_31427,N_29728,N_27022);
nand U31428 (N_31428,N_29587,N_29349);
xnor U31429 (N_31429,N_26843,N_26708);
nand U31430 (N_31430,N_25641,N_29122);
or U31431 (N_31431,N_27150,N_28345);
nand U31432 (N_31432,N_25932,N_27688);
nor U31433 (N_31433,N_26172,N_26693);
nand U31434 (N_31434,N_28410,N_26013);
or U31435 (N_31435,N_26466,N_27788);
nand U31436 (N_31436,N_26555,N_29963);
nor U31437 (N_31437,N_25596,N_27232);
nand U31438 (N_31438,N_28695,N_28035);
nor U31439 (N_31439,N_27258,N_27625);
and U31440 (N_31440,N_28798,N_26659);
nor U31441 (N_31441,N_27954,N_29894);
xor U31442 (N_31442,N_28415,N_26024);
xnor U31443 (N_31443,N_27719,N_29774);
xnor U31444 (N_31444,N_29865,N_28531);
and U31445 (N_31445,N_29391,N_29917);
nor U31446 (N_31446,N_27531,N_27321);
or U31447 (N_31447,N_26130,N_29888);
nand U31448 (N_31448,N_28763,N_27308);
nand U31449 (N_31449,N_28083,N_28447);
nor U31450 (N_31450,N_27239,N_26226);
nand U31451 (N_31451,N_27522,N_25833);
xnor U31452 (N_31452,N_28137,N_28305);
and U31453 (N_31453,N_29521,N_27071);
xor U31454 (N_31454,N_28948,N_25481);
and U31455 (N_31455,N_27966,N_28494);
nand U31456 (N_31456,N_28440,N_26612);
or U31457 (N_31457,N_27512,N_28930);
xnor U31458 (N_31458,N_28722,N_28140);
or U31459 (N_31459,N_29087,N_25685);
nor U31460 (N_31460,N_26283,N_26069);
and U31461 (N_31461,N_25691,N_27126);
nor U31462 (N_31462,N_29512,N_28060);
and U31463 (N_31463,N_29610,N_28241);
nand U31464 (N_31464,N_26989,N_28371);
nor U31465 (N_31465,N_25427,N_28085);
or U31466 (N_31466,N_29308,N_25403);
or U31467 (N_31467,N_29197,N_27011);
nand U31468 (N_31468,N_29998,N_26800);
and U31469 (N_31469,N_29482,N_25610);
nor U31470 (N_31470,N_26521,N_28487);
xnor U31471 (N_31471,N_27132,N_28221);
nor U31472 (N_31472,N_25668,N_28218);
nand U31473 (N_31473,N_25831,N_29745);
nand U31474 (N_31474,N_27795,N_26720);
nand U31475 (N_31475,N_28461,N_25371);
or U31476 (N_31476,N_29063,N_27827);
and U31477 (N_31477,N_29659,N_27722);
and U31478 (N_31478,N_25409,N_28774);
or U31479 (N_31479,N_27725,N_25468);
nor U31480 (N_31480,N_26723,N_28263);
nand U31481 (N_31481,N_28145,N_29694);
nor U31482 (N_31482,N_29997,N_25684);
or U31483 (N_31483,N_26979,N_27048);
or U31484 (N_31484,N_27902,N_25867);
nor U31485 (N_31485,N_28360,N_28257);
and U31486 (N_31486,N_27328,N_27267);
and U31487 (N_31487,N_29319,N_25835);
and U31488 (N_31488,N_27815,N_27849);
nor U31489 (N_31489,N_26574,N_25559);
nand U31490 (N_31490,N_26851,N_26036);
or U31491 (N_31491,N_29115,N_28622);
and U31492 (N_31492,N_26736,N_26913);
nor U31493 (N_31493,N_28617,N_26244);
nor U31494 (N_31494,N_29130,N_28631);
or U31495 (N_31495,N_25289,N_26580);
nand U31496 (N_31496,N_25385,N_25592);
nor U31497 (N_31497,N_25279,N_28736);
or U31498 (N_31498,N_26731,N_27548);
and U31499 (N_31499,N_26302,N_29645);
or U31500 (N_31500,N_27878,N_28871);
xnor U31501 (N_31501,N_29146,N_27997);
xor U31502 (N_31502,N_26086,N_26636);
xor U31503 (N_31503,N_25726,N_28673);
nand U31504 (N_31504,N_29672,N_29036);
or U31505 (N_31505,N_28931,N_27516);
nor U31506 (N_31506,N_27702,N_28069);
or U31507 (N_31507,N_25782,N_26616);
xor U31508 (N_31508,N_27911,N_27038);
nor U31509 (N_31509,N_25529,N_25202);
xor U31510 (N_31510,N_25602,N_26630);
xor U31511 (N_31511,N_25693,N_28584);
or U31512 (N_31512,N_25599,N_29573);
xor U31513 (N_31513,N_29145,N_25433);
nand U31514 (N_31514,N_27410,N_25402);
and U31515 (N_31515,N_25965,N_26655);
nor U31516 (N_31516,N_28172,N_25457);
or U31517 (N_31517,N_29795,N_29131);
and U31518 (N_31518,N_28920,N_29327);
or U31519 (N_31519,N_29473,N_28042);
and U31520 (N_31520,N_29020,N_27253);
nor U31521 (N_31521,N_27149,N_29039);
nor U31522 (N_31522,N_29951,N_25135);
or U31523 (N_31523,N_27330,N_25196);
nor U31524 (N_31524,N_25350,N_27006);
nor U31525 (N_31525,N_28023,N_25807);
or U31526 (N_31526,N_25254,N_26877);
nand U31527 (N_31527,N_28666,N_28546);
xor U31528 (N_31528,N_25859,N_26250);
and U31529 (N_31529,N_28994,N_26227);
nand U31530 (N_31530,N_25370,N_29106);
or U31531 (N_31531,N_25882,N_26772);
or U31532 (N_31532,N_29303,N_27025);
nor U31533 (N_31533,N_26033,N_25062);
nor U31534 (N_31534,N_27523,N_27458);
xor U31535 (N_31535,N_26770,N_27847);
nand U31536 (N_31536,N_26519,N_27169);
or U31537 (N_31537,N_25174,N_29527);
or U31538 (N_31538,N_25393,N_27469);
and U31539 (N_31539,N_28645,N_28890);
or U31540 (N_31540,N_27699,N_27541);
or U31541 (N_31541,N_26819,N_26212);
nor U31542 (N_31542,N_25620,N_29625);
nand U31543 (N_31543,N_26945,N_25808);
and U31544 (N_31544,N_28896,N_29540);
nor U31545 (N_31545,N_26827,N_27886);
nor U31546 (N_31546,N_25072,N_26380);
nand U31547 (N_31547,N_28482,N_29971);
or U31548 (N_31548,N_28831,N_25545);
xnor U31549 (N_31549,N_25794,N_27739);
and U31550 (N_31550,N_28390,N_29478);
nor U31551 (N_31551,N_29599,N_25205);
xnor U31552 (N_31552,N_29909,N_25233);
nand U31553 (N_31553,N_29632,N_26156);
and U31554 (N_31554,N_27485,N_27721);
and U31555 (N_31555,N_29992,N_25928);
nor U31556 (N_31556,N_29252,N_27893);
nand U31557 (N_31557,N_28086,N_27257);
nor U31558 (N_31558,N_25211,N_29486);
xor U31559 (N_31559,N_27041,N_29412);
and U31560 (N_31560,N_26209,N_29185);
or U31561 (N_31561,N_27576,N_29232);
nand U31562 (N_31562,N_27224,N_27468);
and U31563 (N_31563,N_29902,N_27925);
xnor U31564 (N_31564,N_25923,N_28016);
or U31565 (N_31565,N_25311,N_27987);
or U31566 (N_31566,N_29861,N_25763);
nor U31567 (N_31567,N_28247,N_27960);
nand U31568 (N_31568,N_25343,N_27030);
or U31569 (N_31569,N_29705,N_26575);
or U31570 (N_31570,N_27283,N_26392);
nand U31571 (N_31571,N_25232,N_26213);
nand U31572 (N_31572,N_25628,N_25362);
xnor U31573 (N_31573,N_26673,N_25982);
nand U31574 (N_31574,N_27785,N_27388);
or U31575 (N_31575,N_29034,N_28384);
or U31576 (N_31576,N_27806,N_25154);
nand U31577 (N_31577,N_25306,N_28706);
nor U31578 (N_31578,N_25670,N_28490);
and U31579 (N_31579,N_26237,N_28785);
xor U31580 (N_31580,N_25665,N_26997);
nand U31581 (N_31581,N_26502,N_27311);
nor U31582 (N_31582,N_25009,N_27766);
or U31583 (N_31583,N_29605,N_29099);
or U31584 (N_31584,N_25055,N_28202);
nor U31585 (N_31585,N_25639,N_29209);
or U31586 (N_31586,N_26442,N_27165);
xor U31587 (N_31587,N_25236,N_28609);
nand U31588 (N_31588,N_25492,N_28652);
nor U31589 (N_31589,N_25873,N_25856);
nand U31590 (N_31590,N_26749,N_27970);
nor U31591 (N_31591,N_25826,N_28159);
and U31592 (N_31592,N_28747,N_26744);
nor U31593 (N_31593,N_28821,N_27650);
or U31594 (N_31594,N_28918,N_28084);
nor U31595 (N_31595,N_25386,N_26224);
and U31596 (N_31596,N_29453,N_27556);
nor U31597 (N_31597,N_28682,N_28099);
nor U31598 (N_31598,N_25792,N_29801);
nor U31599 (N_31599,N_26189,N_25476);
nor U31600 (N_31600,N_25137,N_26603);
or U31601 (N_31601,N_28279,N_29938);
xnor U31602 (N_31602,N_25864,N_26349);
nor U31603 (N_31603,N_25326,N_29624);
nor U31604 (N_31604,N_28109,N_29987);
xor U31605 (N_31605,N_26235,N_26917);
nand U31606 (N_31606,N_28200,N_28551);
xor U31607 (N_31607,N_25305,N_27707);
xor U31608 (N_31608,N_25678,N_26491);
nand U31609 (N_31609,N_29480,N_27493);
or U31610 (N_31610,N_27460,N_25216);
or U31611 (N_31611,N_27451,N_25966);
xnor U31612 (N_31612,N_25043,N_29715);
nor U31613 (N_31613,N_29174,N_27860);
and U31614 (N_31614,N_28998,N_28733);
nor U31615 (N_31615,N_29737,N_29110);
or U31616 (N_31616,N_27381,N_25413);
or U31617 (N_31617,N_28179,N_25718);
nand U31618 (N_31618,N_28756,N_29306);
nor U31619 (N_31619,N_25057,N_26641);
nand U31620 (N_31620,N_25327,N_29476);
xor U31621 (N_31621,N_25958,N_28397);
nor U31622 (N_31622,N_29878,N_27621);
or U31623 (N_31623,N_26269,N_25255);
nor U31624 (N_31624,N_29771,N_27651);
nor U31625 (N_31625,N_27293,N_27449);
nand U31626 (N_31626,N_29050,N_28560);
xor U31627 (N_31627,N_26317,N_27091);
nor U31628 (N_31628,N_25200,N_28742);
nand U31629 (N_31629,N_27579,N_27701);
and U31630 (N_31630,N_25715,N_29932);
nor U31631 (N_31631,N_25942,N_26252);
xnor U31632 (N_31632,N_28703,N_28738);
xnor U31633 (N_31633,N_29940,N_25728);
nor U31634 (N_31634,N_26281,N_25905);
or U31635 (N_31635,N_27687,N_27226);
nand U31636 (N_31636,N_25027,N_25845);
and U31637 (N_31637,N_26801,N_27510);
or U31638 (N_31638,N_25171,N_29236);
nand U31639 (N_31639,N_27112,N_29559);
and U31640 (N_31640,N_29355,N_27101);
nor U31641 (N_31641,N_25322,N_27400);
xnor U31642 (N_31642,N_27774,N_27728);
xor U31643 (N_31643,N_28120,N_29392);
or U31644 (N_31644,N_27887,N_26352);
xnor U31645 (N_31645,N_28610,N_25812);
and U31646 (N_31646,N_25863,N_26513);
xnor U31647 (N_31647,N_28119,N_25537);
nor U31648 (N_31648,N_26614,N_29903);
nor U31649 (N_31649,N_28815,N_26023);
xor U31650 (N_31650,N_25082,N_29347);
nand U31651 (N_31651,N_26312,N_25534);
or U31652 (N_31652,N_29537,N_25858);
xor U31653 (N_31653,N_27709,N_27927);
nor U31654 (N_31654,N_27125,N_26248);
nand U31655 (N_31655,N_25788,N_27302);
nand U31656 (N_31656,N_27796,N_26646);
nor U31657 (N_31657,N_25060,N_29516);
nor U31658 (N_31658,N_27903,N_28193);
and U31659 (N_31659,N_27502,N_25209);
xor U31660 (N_31660,N_28868,N_25270);
or U31661 (N_31661,N_27562,N_26311);
or U31662 (N_31662,N_27962,N_25175);
and U31663 (N_31663,N_29030,N_27195);
and U31664 (N_31664,N_28322,N_29326);
nor U31665 (N_31665,N_26456,N_26823);
nor U31666 (N_31666,N_29866,N_27373);
xnor U31667 (N_31667,N_25139,N_28289);
nand U31668 (N_31668,N_26412,N_29977);
or U31669 (N_31669,N_25555,N_29985);
and U31670 (N_31670,N_29092,N_28004);
and U31671 (N_31671,N_27155,N_27075);
nand U31672 (N_31672,N_26668,N_28325);
or U31673 (N_31673,N_26619,N_25446);
nor U31674 (N_31674,N_29689,N_26474);
xnor U31675 (N_31675,N_28884,N_29068);
or U31676 (N_31676,N_29617,N_29466);
xnor U31677 (N_31677,N_26617,N_26414);
xnor U31678 (N_31678,N_25197,N_26895);
nand U31679 (N_31679,N_25430,N_25801);
xor U31680 (N_31680,N_25275,N_29019);
xor U31681 (N_31681,N_27837,N_26696);
and U31682 (N_31682,N_28899,N_27191);
and U31683 (N_31683,N_29566,N_28170);
nor U31684 (N_31684,N_26830,N_29717);
nor U31685 (N_31685,N_27763,N_29156);
nand U31686 (N_31686,N_26354,N_29821);
nor U31687 (N_31687,N_27269,N_25458);
and U31688 (N_31688,N_25227,N_27000);
nand U31689 (N_31689,N_25257,N_25655);
or U31690 (N_31690,N_25972,N_25234);
nor U31691 (N_31691,N_27109,N_26863);
or U31692 (N_31692,N_26539,N_28990);
xor U31693 (N_31693,N_26111,N_26566);
nor U31694 (N_31694,N_25384,N_28748);
and U31695 (N_31695,N_29103,N_28776);
or U31696 (N_31696,N_25231,N_26921);
nor U31697 (N_31697,N_27045,N_26902);
nand U31698 (N_31698,N_26856,N_28313);
or U31699 (N_31699,N_29490,N_28684);
xor U31700 (N_31700,N_28845,N_27491);
nand U31701 (N_31701,N_28380,N_26449);
xor U31702 (N_31702,N_25156,N_25658);
nand U31703 (N_31703,N_25157,N_26185);
nor U31704 (N_31704,N_25049,N_26327);
nor U31705 (N_31705,N_25239,N_26999);
nand U31706 (N_31706,N_26121,N_29929);
or U31707 (N_31707,N_29633,N_26097);
nand U31708 (N_31708,N_27358,N_26916);
nand U31709 (N_31709,N_29684,N_28438);
xnor U31710 (N_31710,N_25100,N_26303);
nor U31711 (N_31711,N_26760,N_29905);
and U31712 (N_31712,N_29305,N_28502);
xor U31713 (N_31713,N_27113,N_25834);
xnor U31714 (N_31714,N_25065,N_29045);
or U31715 (N_31715,N_26207,N_29135);
nand U31716 (N_31716,N_28653,N_27294);
or U31717 (N_31717,N_26407,N_28562);
xnor U31718 (N_31718,N_28959,N_25488);
or U31719 (N_31719,N_25347,N_27858);
nor U31720 (N_31720,N_25449,N_28225);
nand U31721 (N_31721,N_26584,N_27910);
or U31722 (N_31722,N_25381,N_26482);
nand U31723 (N_31723,N_26532,N_27952);
nor U31724 (N_31724,N_28905,N_26966);
xor U31725 (N_31725,N_25263,N_26704);
and U31726 (N_31726,N_28801,N_28381);
and U31727 (N_31727,N_28688,N_29850);
nor U31728 (N_31728,N_28164,N_27820);
nand U31729 (N_31729,N_25240,N_27855);
nand U31730 (N_31730,N_25984,N_29195);
and U31731 (N_31731,N_28078,N_26638);
nor U31732 (N_31732,N_26144,N_26337);
nand U31733 (N_31733,N_26620,N_28422);
or U31734 (N_31734,N_26900,N_25105);
or U31735 (N_31735,N_29981,N_28870);
xor U31736 (N_31736,N_28402,N_26406);
nor U31737 (N_31737,N_27335,N_27931);
nand U31738 (N_31738,N_28670,N_28626);
and U31739 (N_31739,N_28267,N_29366);
xor U31740 (N_31740,N_28190,N_26461);
nand U31741 (N_31741,N_28590,N_26594);
or U31742 (N_31742,N_26247,N_27408);
nor U31743 (N_31743,N_27752,N_25282);
and U31744 (N_31744,N_26385,N_28569);
nor U31745 (N_31745,N_27178,N_27831);
nor U31746 (N_31746,N_28847,N_26035);
nand U31747 (N_31747,N_29582,N_25059);
and U31748 (N_31748,N_25778,N_25571);
nand U31749 (N_31749,N_29248,N_29726);
nor U31750 (N_31750,N_25341,N_25904);
xnor U31751 (N_31751,N_29014,N_28376);
xor U31752 (N_31752,N_29936,N_26253);
xor U31753 (N_31753,N_25120,N_28073);
xor U31754 (N_31754,N_29890,N_26018);
or U31755 (N_31755,N_28029,N_26942);
xor U31756 (N_31756,N_25981,N_26976);
or U31757 (N_31757,N_26367,N_28578);
and U31758 (N_31758,N_26687,N_28576);
and U31759 (N_31759,N_28720,N_25635);
nand U31760 (N_31760,N_25819,N_26907);
or U31761 (N_31761,N_26926,N_29172);
or U31762 (N_31762,N_29074,N_28391);
nand U31763 (N_31763,N_26131,N_27304);
nand U31764 (N_31764,N_25140,N_25455);
or U31765 (N_31765,N_26769,N_26157);
or U31766 (N_31766,N_27689,N_26445);
or U31767 (N_31767,N_28359,N_25604);
nand U31768 (N_31768,N_29451,N_27382);
and U31769 (N_31769,N_29418,N_27229);
nand U31770 (N_31770,N_26430,N_29781);
nand U31771 (N_31771,N_29974,N_29792);
or U31772 (N_31772,N_28088,N_27405);
xor U31773 (N_31773,N_29827,N_27900);
xor U31774 (N_31774,N_29742,N_27436);
nand U31775 (N_31775,N_28469,N_25569);
xor U31776 (N_31776,N_26083,N_28002);
nor U31777 (N_31777,N_29730,N_29892);
xnor U31778 (N_31778,N_29377,N_27638);
nand U31779 (N_31779,N_25194,N_28310);
nor U31780 (N_31780,N_26840,N_28542);
or U31781 (N_31781,N_27172,N_28496);
nor U31782 (N_31782,N_25690,N_28730);
nand U31783 (N_31783,N_25078,N_26894);
nand U31784 (N_31784,N_26717,N_29539);
xor U31785 (N_31785,N_29166,N_25929);
and U31786 (N_31786,N_26105,N_29879);
and U31787 (N_31787,N_29090,N_26710);
nor U31788 (N_31788,N_28448,N_28134);
nor U31789 (N_31789,N_29712,N_27920);
nor U31790 (N_31790,N_26600,N_25494);
nor U31791 (N_31791,N_27482,N_29920);
and U31792 (N_31792,N_28739,N_29492);
xnor U31793 (N_31793,N_29843,N_29033);
or U31794 (N_31794,N_28020,N_29202);
and U31795 (N_31795,N_26006,N_29021);
nor U31796 (N_31796,N_26022,N_26268);
xor U31797 (N_31797,N_27348,N_27134);
or U31798 (N_31798,N_28321,N_25862);
and U31799 (N_31799,N_28657,N_27936);
and U31800 (N_31800,N_28334,N_26216);
or U31801 (N_31801,N_27489,N_29966);
or U31802 (N_31802,N_26645,N_29604);
nor U31803 (N_31803,N_28605,N_29323);
nand U31804 (N_31804,N_28963,N_25212);
or U31805 (N_31805,N_28068,N_26363);
nor U31806 (N_31806,N_27897,N_29772);
and U31807 (N_31807,N_26977,N_26732);
and U31808 (N_31808,N_26457,N_29112);
xnor U31809 (N_31809,N_26405,N_25425);
nand U31810 (N_31810,N_26649,N_28271);
or U31811 (N_31811,N_26524,N_28824);
or U31812 (N_31812,N_25554,N_26165);
xnor U31813 (N_31813,N_27390,N_26954);
nor U31814 (N_31814,N_25020,N_28818);
or U31815 (N_31815,N_28154,N_25366);
or U31816 (N_31816,N_28081,N_27956);
nor U31817 (N_31817,N_29732,N_26259);
or U31818 (N_31818,N_28591,N_25436);
nor U31819 (N_31819,N_27590,N_25522);
or U31820 (N_31820,N_27133,N_27198);
nand U31821 (N_31821,N_28885,N_25042);
nor U31822 (N_31822,N_27684,N_28350);
or U31823 (N_31823,N_28711,N_28621);
xor U31824 (N_31824,N_26713,N_25012);
xor U31825 (N_31825,N_26558,N_29591);
and U31826 (N_31826,N_29957,N_29154);
nor U31827 (N_31827,N_27659,N_25225);
nand U31828 (N_31828,N_28274,N_29722);
nand U31829 (N_31829,N_29027,N_28750);
xor U31830 (N_31830,N_27818,N_26809);
xor U31831 (N_31831,N_25672,N_26670);
nor U31832 (N_31832,N_28615,N_29791);
xnor U31833 (N_31833,N_25262,N_28156);
nor U31834 (N_31834,N_28807,N_28022);
nor U31835 (N_31835,N_27979,N_26726);
xnor U31836 (N_31836,N_28500,N_29223);
and U31837 (N_31837,N_29384,N_29329);
xor U31838 (N_31838,N_27327,N_27251);
nor U31839 (N_31839,N_25183,N_29812);
nand U31840 (N_31840,N_26241,N_28975);
nand U31841 (N_31841,N_27414,N_25221);
xnor U31842 (N_31842,N_27235,N_25964);
nand U31843 (N_31843,N_26784,N_28395);
xor U31844 (N_31844,N_29954,N_28775);
and U31845 (N_31845,N_26536,N_27517);
nand U31846 (N_31846,N_28285,N_29693);
or U31847 (N_31847,N_25774,N_27212);
and U31848 (N_31848,N_25914,N_25939);
and U31849 (N_31849,N_28096,N_25817);
nor U31850 (N_31850,N_26716,N_26792);
nand U31851 (N_31851,N_29640,N_27563);
and U31852 (N_31852,N_28249,N_26676);
or U31853 (N_31853,N_26285,N_25721);
nor U31854 (N_31854,N_29169,N_27805);
or U31855 (N_31855,N_28728,N_25408);
nand U31856 (N_31856,N_29782,N_27248);
or U31857 (N_31857,N_26292,N_28835);
and U31858 (N_31858,N_25912,N_29206);
xor U31859 (N_31859,N_26510,N_27497);
nor U31860 (N_31860,N_29257,N_25113);
nand U31861 (N_31861,N_25696,N_27990);
or U31862 (N_31862,N_26629,N_28362);
xor U31863 (N_31863,N_27339,N_27092);
or U31864 (N_31864,N_25037,N_27823);
or U31865 (N_31865,N_27263,N_29653);
or U31866 (N_31866,N_26197,N_28566);
xnor U31867 (N_31867,N_28552,N_28955);
xnor U31868 (N_31868,N_25361,N_26811);
nor U31869 (N_31869,N_28183,N_28985);
and U31870 (N_31870,N_27645,N_28765);
and U31871 (N_31871,N_26866,N_28142);
nand U31872 (N_31872,N_27118,N_27595);
or U31873 (N_31873,N_29372,N_27384);
and U31874 (N_31874,N_27415,N_28485);
or U31875 (N_31875,N_27028,N_25806);
or U31876 (N_31876,N_25237,N_26265);
and U31877 (N_31877,N_25002,N_25822);
xnor U31878 (N_31878,N_27233,N_29318);
xor U31879 (N_31879,N_25101,N_26793);
and U31880 (N_31880,N_29960,N_27065);
nor U31881 (N_31881,N_28528,N_28991);
nand U31882 (N_31882,N_29421,N_27357);
nand U31883 (N_31883,N_29769,N_27918);
xor U31884 (N_31884,N_26397,N_25340);
xnor U31885 (N_31885,N_27333,N_29520);
nand U31886 (N_31886,N_28409,N_27724);
nand U31887 (N_31887,N_28166,N_25505);
nand U31888 (N_31888,N_29970,N_27708);
and U31889 (N_31889,N_29322,N_28428);
or U31890 (N_31890,N_25550,N_28668);
xnor U31891 (N_31891,N_28858,N_29868);
or U31892 (N_31892,N_26561,N_26495);
or U31893 (N_31893,N_29294,N_26947);
nand U31894 (N_31894,N_27919,N_28676);
nand U31895 (N_31895,N_26955,N_29395);
or U31896 (N_31896,N_26814,N_29272);
and U31897 (N_31897,N_25572,N_27080);
and U31898 (N_31898,N_26930,N_26836);
nor U31899 (N_31899,N_26146,N_26441);
or U31900 (N_31900,N_27995,N_26084);
and U31901 (N_31901,N_28197,N_28548);
xnor U31902 (N_31902,N_27778,N_27008);
xnor U31903 (N_31903,N_28370,N_26706);
or U31904 (N_31904,N_27431,N_28811);
or U31905 (N_31905,N_27560,N_28185);
nor U31906 (N_31906,N_25028,N_26005);
nor U31907 (N_31907,N_26556,N_29669);
nor U31908 (N_31908,N_27626,N_25204);
and U31909 (N_31909,N_27520,N_26956);
nand U31910 (N_31910,N_29681,N_25271);
and U31911 (N_31911,N_25962,N_26776);
and U31912 (N_31912,N_28539,N_28768);
and U31913 (N_31913,N_27035,N_26417);
nor U31914 (N_31914,N_27085,N_25198);
and U31915 (N_31915,N_25659,N_25781);
or U31916 (N_31916,N_25294,N_27136);
nor U31917 (N_31917,N_29013,N_27342);
xor U31918 (N_31918,N_25039,N_28887);
xnor U31919 (N_31919,N_28717,N_26199);
xor U31920 (N_31920,N_29967,N_28491);
xor U31921 (N_31921,N_27148,N_25054);
nor U31922 (N_31922,N_26464,N_27492);
nand U31923 (N_31923,N_27867,N_25760);
or U31924 (N_31924,N_28794,N_25925);
nor U31925 (N_31925,N_29813,N_29089);
nor U31926 (N_31926,N_29475,N_29501);
or U31927 (N_31927,N_26517,N_25989);
or U31928 (N_31928,N_29638,N_25379);
nor U31929 (N_31929,N_27998,N_27162);
nor U31930 (N_31930,N_29222,N_29444);
and U31931 (N_31931,N_26314,N_27066);
nand U31932 (N_31932,N_26021,N_26692);
nor U31933 (N_31933,N_28222,N_28468);
nor U31934 (N_31934,N_29350,N_29975);
or U31935 (N_31935,N_29740,N_27843);
and U31936 (N_31936,N_25489,N_27087);
or U31937 (N_31937,N_25224,N_27196);
or U31938 (N_31938,N_26964,N_28050);
nor U31939 (N_31939,N_26132,N_25396);
and U31940 (N_31940,N_26758,N_28192);
and U31941 (N_31941,N_29238,N_27577);
nand U31942 (N_31942,N_28430,N_27170);
xor U31943 (N_31943,N_26952,N_28169);
and U31944 (N_31944,N_27868,N_29914);
and U31945 (N_31945,N_28704,N_26294);
and U31946 (N_31946,N_29999,N_27922);
and U31947 (N_31947,N_26651,N_27862);
and U31948 (N_31948,N_26981,N_25796);
and U31949 (N_31949,N_27594,N_29389);
nand U31950 (N_31950,N_28819,N_26995);
or U31951 (N_31951,N_26542,N_29836);
nor U31952 (N_31952,N_26068,N_28413);
nor U31953 (N_31953,N_29263,N_26118);
or U31954 (N_31954,N_26722,N_27104);
nor U31955 (N_31955,N_25301,N_27802);
and U31956 (N_31956,N_27885,N_25567);
xor U31957 (N_31957,N_27153,N_28324);
xor U31958 (N_31958,N_29767,N_25090);
and U31959 (N_31959,N_29662,N_26058);
xor U31960 (N_31960,N_26149,N_28082);
nand U31961 (N_31961,N_28939,N_27633);
or U31962 (N_31962,N_28246,N_25094);
and U31963 (N_31963,N_27564,N_25407);
or U31964 (N_31964,N_27117,N_25879);
or U31965 (N_31965,N_25069,N_25868);
nand U31966 (N_31966,N_28696,N_28157);
nor U31967 (N_31967,N_26459,N_29150);
and U31968 (N_31968,N_26833,N_27194);
nor U31969 (N_31969,N_27978,N_26096);
nor U31970 (N_31970,N_27074,N_29023);
or U31971 (N_31971,N_26287,N_27420);
xor U31972 (N_31972,N_28691,N_26986);
nor U31973 (N_31973,N_27841,N_29500);
or U31974 (N_31974,N_26882,N_28618);
xor U31975 (N_31975,N_28536,N_26195);
nor U31976 (N_31976,N_29191,N_26777);
nand U31977 (N_31977,N_25719,N_26719);
or U31978 (N_31978,N_27298,N_29576);
nand U31979 (N_31979,N_26152,N_28092);
or U31980 (N_31980,N_29877,N_27097);
or U31981 (N_31981,N_29086,N_25631);
and U31982 (N_31982,N_26044,N_27750);
nor U31983 (N_31983,N_28017,N_28797);
or U31984 (N_31984,N_29069,N_29814);
nand U31985 (N_31985,N_25245,N_28790);
xnor U31986 (N_31986,N_25030,N_27598);
or U31987 (N_31987,N_26497,N_27537);
nor U31988 (N_31988,N_27459,N_26342);
nor U31989 (N_31989,N_28753,N_26485);
xor U31990 (N_31990,N_26598,N_25515);
and U31991 (N_31991,N_26368,N_27037);
xor U31992 (N_31992,N_29370,N_26666);
and U31993 (N_31993,N_25507,N_29165);
and U31994 (N_31994,N_27003,N_29123);
and U31995 (N_31995,N_27879,N_28796);
nor U31996 (N_31996,N_28638,N_25397);
nor U31997 (N_31997,N_29698,N_26904);
or U31998 (N_31998,N_26257,N_26515);
or U31999 (N_31999,N_28582,N_27614);
and U32000 (N_32000,N_29085,N_25312);
xor U32001 (N_32001,N_25201,N_28235);
nand U32002 (N_32002,N_29708,N_25309);
and U32003 (N_32003,N_29915,N_28326);
or U32004 (N_32004,N_25452,N_26820);
nor U32005 (N_32005,N_28125,N_26643);
xor U32006 (N_32006,N_27639,N_29017);
xor U32007 (N_32007,N_26211,N_26166);
xor U32008 (N_32008,N_26364,N_28135);
nor U32009 (N_32009,N_25423,N_27419);
xnor U32010 (N_32010,N_28585,N_27211);
nor U32011 (N_32011,N_27462,N_27586);
or U32012 (N_32012,N_27102,N_27718);
and U32013 (N_32013,N_25852,N_27496);
or U32014 (N_32014,N_26181,N_29702);
or U32015 (N_32015,N_28143,N_29491);
and U32016 (N_32016,N_27084,N_28472);
and U32017 (N_32017,N_29948,N_28302);
nor U32018 (N_32018,N_28902,N_27338);
nor U32019 (N_32019,N_26098,N_29067);
or U32020 (N_32020,N_27203,N_29830);
or U32021 (N_32021,N_25497,N_28266);
or U32022 (N_32022,N_26423,N_26918);
and U32023 (N_32023,N_29187,N_25941);
xnor U32024 (N_32024,N_27812,N_26328);
xnor U32025 (N_32025,N_26613,N_29171);
nor U32026 (N_32026,N_26529,N_29494);
nor U32027 (N_32027,N_29614,N_28788);
and U32028 (N_32028,N_28323,N_28849);
or U32029 (N_32029,N_26763,N_27182);
nor U32030 (N_32030,N_25434,N_27612);
and U32031 (N_32031,N_27072,N_25514);
or U32032 (N_32032,N_28965,N_28517);
or U32033 (N_32033,N_27664,N_25944);
or U32034 (N_32034,N_29804,N_25651);
xnor U32035 (N_32035,N_27027,N_26343);
xor U32036 (N_32036,N_28558,N_25744);
or U32037 (N_32037,N_28782,N_28019);
xnor U32038 (N_32038,N_29244,N_27606);
and U32039 (N_32039,N_29847,N_28203);
nor U32040 (N_32040,N_27228,N_27679);
xnor U32041 (N_32041,N_28628,N_27470);
and U32042 (N_32042,N_25913,N_26571);
nor U32043 (N_32043,N_28091,N_29269);
and U32044 (N_32044,N_26982,N_29682);
and U32045 (N_32045,N_25134,N_26435);
or U32046 (N_32046,N_29227,N_28045);
nand U32047 (N_32047,N_26753,N_25909);
and U32048 (N_32048,N_27247,N_25823);
nor U32049 (N_32049,N_27631,N_25315);
and U32050 (N_32050,N_28873,N_26115);
xor U32051 (N_32051,N_26846,N_29371);
nand U32052 (N_32052,N_29448,N_29425);
and U32053 (N_32053,N_26381,N_26103);
nor U32054 (N_32054,N_29102,N_25034);
nand U32055 (N_32055,N_26339,N_25508);
nor U32056 (N_32056,N_29234,N_27835);
xor U32057 (N_32057,N_28554,N_28336);
and U32058 (N_32058,N_26138,N_28477);
nor U32059 (N_32059,N_28423,N_26071);
and U32060 (N_32060,N_25573,N_28967);
and U32061 (N_32061,N_25398,N_26551);
xor U32062 (N_32062,N_26315,N_26220);
or U32063 (N_32063,N_26378,N_27500);
nor U32064 (N_32064,N_29203,N_27349);
nand U32065 (N_32065,N_26745,N_26027);
xnor U32066 (N_32066,N_29239,N_25004);
nor U32067 (N_32067,N_26162,N_27295);
nor U32068 (N_32068,N_29162,N_27561);
nor U32069 (N_32069,N_27013,N_29098);
nor U32070 (N_32070,N_25441,N_28094);
nor U32071 (N_32071,N_29923,N_29300);
xor U32072 (N_32072,N_25517,N_28052);
xnor U32073 (N_32073,N_29764,N_25346);
nor U32074 (N_32074,N_27177,N_28344);
or U32075 (N_32075,N_25680,N_27478);
nor U32076 (N_32076,N_28426,N_25083);
nor U32077 (N_32077,N_28425,N_25538);
nor U32078 (N_32078,N_25586,N_27768);
nand U32079 (N_32079,N_27081,N_26526);
nor U32080 (N_32080,N_26828,N_26564);
and U32081 (N_32081,N_28973,N_27214);
or U32082 (N_32082,N_29271,N_26017);
nor U32083 (N_32083,N_25526,N_27898);
xnor U32084 (N_32084,N_27016,N_25974);
xnor U32085 (N_32085,N_28921,N_29207);
nor U32086 (N_32086,N_27193,N_25633);
or U32087 (N_32087,N_25380,N_28848);
or U32088 (N_32088,N_26548,N_27641);
xnor U32089 (N_32089,N_26032,N_25765);
xnor U32090 (N_32090,N_25117,N_28342);
xor U32091 (N_32091,N_25606,N_28453);
and U32092 (N_32092,N_26789,N_26941);
and U32093 (N_32093,N_27776,N_26738);
xnor U32094 (N_32094,N_25293,N_29709);
or U32095 (N_32095,N_25061,N_26611);
nor U32096 (N_32096,N_28234,N_27244);
xor U32097 (N_32097,N_25841,N_29409);
xnor U32098 (N_32098,N_26228,N_25460);
nor U32099 (N_32099,N_29995,N_27767);
xnor U32100 (N_32100,N_26610,N_26778);
nand U32101 (N_32101,N_25162,N_29181);
xor U32102 (N_32102,N_27948,N_25609);
or U32103 (N_32103,N_28823,N_25632);
and U32104 (N_32104,N_27009,N_29454);
xnor U32105 (N_32105,N_29686,N_28863);
or U32106 (N_32106,N_25764,N_29831);
nor U32107 (N_32107,N_27033,N_27989);
and U32108 (N_32108,N_26479,N_28158);
nor U32109 (N_32109,N_27334,N_28854);
or U32110 (N_32110,N_28243,N_25843);
nor U32111 (N_32111,N_28892,N_25777);
or U32112 (N_32112,N_25910,N_25898);
nand U32113 (N_32113,N_25576,N_27457);
xor U32114 (N_32114,N_28974,N_27090);
nor U32115 (N_32115,N_28629,N_26020);
and U32116 (N_32116,N_27185,N_27921);
nand U32117 (N_32117,N_26885,N_27914);
nand U32118 (N_32118,N_27444,N_25894);
and U32119 (N_32119,N_28043,N_25128);
and U32120 (N_32120,N_26239,N_27147);
nor U32121 (N_32121,N_26415,N_29557);
and U32122 (N_32122,N_29703,N_27060);
nor U32123 (N_32123,N_28940,N_26549);
and U32124 (N_32124,N_26631,N_29817);
xor U32125 (N_32125,N_26472,N_25469);
nand U32126 (N_32126,N_28508,N_29735);
nor U32127 (N_32127,N_25107,N_28903);
xor U32128 (N_32128,N_26754,N_27628);
nor U32129 (N_32129,N_29481,N_27059);
and U32130 (N_32130,N_27073,N_28992);
or U32131 (N_32131,N_25267,N_29896);
nor U32132 (N_32132,N_25643,N_25890);
or U32133 (N_32133,N_28057,N_28877);
nor U32134 (N_32134,N_28793,N_29685);
or U32135 (N_32135,N_25857,N_28953);
nand U32136 (N_32136,N_25086,N_29956);
and U32137 (N_32137,N_28647,N_28292);
nand U32138 (N_32138,N_26254,N_26460);
nand U32139 (N_32139,N_25354,N_26175);
or U32140 (N_32140,N_27241,N_27658);
nand U32141 (N_32141,N_26240,N_26664);
nand U32142 (N_32142,N_25357,N_28379);
nor U32143 (N_32143,N_28659,N_25664);
nand U32144 (N_32144,N_28171,N_29109);
and U32145 (N_32145,N_25111,N_25523);
nor U32146 (N_32146,N_29224,N_29897);
or U32147 (N_32147,N_27036,N_28329);
and U32148 (N_32148,N_28399,N_26304);
or U32149 (N_32149,N_28341,N_29037);
or U32150 (N_32150,N_26039,N_27047);
nor U32151 (N_32151,N_27442,N_29666);
xor U32152 (N_32152,N_25440,N_27262);
nor U32153 (N_32153,N_25881,N_27940);
nand U32154 (N_32154,N_25783,N_26936);
nand U32155 (N_32155,N_28478,N_26196);
nand U32156 (N_32156,N_25952,N_26869);
nand U32157 (N_32157,N_27753,N_27592);
and U32158 (N_32158,N_25702,N_26965);
nor U32159 (N_32159,N_28054,N_27324);
xor U32160 (N_32160,N_26790,N_29408);
nor U32161 (N_32161,N_26293,N_29352);
nor U32162 (N_32162,N_27559,N_29417);
nor U32163 (N_32163,N_28772,N_27761);
nand U32164 (N_32164,N_25528,N_27859);
nor U32165 (N_32165,N_27452,N_29398);
nor U32166 (N_32166,N_25784,N_28725);
nand U32167 (N_32167,N_28291,N_29047);
and U32168 (N_32168,N_29749,N_29493);
and U32169 (N_32169,N_27545,N_25850);
or U32170 (N_32170,N_26125,N_29743);
nor U32171 (N_32171,N_26880,N_29853);
or U32172 (N_32172,N_29220,N_25152);
nor U32173 (N_32173,N_27486,N_26859);
nor U32174 (N_32174,N_26080,N_29427);
nand U32175 (N_32175,N_26682,N_28041);
xnor U32176 (N_32176,N_28177,N_26249);
and U32177 (N_32177,N_27529,N_26797);
nor U32178 (N_32178,N_28604,N_27323);
nand U32179 (N_32179,N_28900,N_28293);
xnor U32180 (N_32180,N_25872,N_25692);
or U32181 (N_32181,N_26101,N_28451);
nor U32182 (N_32182,N_25787,N_27473);
xor U32183 (N_32183,N_25780,N_25313);
and U32184 (N_32184,N_25563,N_29955);
nand U32185 (N_32185,N_27440,N_28097);
and U32186 (N_32186,N_27924,N_29190);
xnor U32187 (N_32187,N_27237,N_28337);
and U32188 (N_32188,N_27895,N_28174);
and U32189 (N_32189,N_28777,N_29346);
xnor U32190 (N_32190,N_27270,N_26308);
or U32191 (N_32191,N_28432,N_29100);
and U32192 (N_32192,N_25840,N_29922);
nor U32193 (N_32193,N_28132,N_26323);
xor U32194 (N_32194,N_25983,N_29211);
xnor U32195 (N_32195,N_29289,N_29469);
nand U32196 (N_32196,N_29054,N_25560);
nor U32197 (N_32197,N_26683,N_27227);
nand U32198 (N_32198,N_27067,N_27634);
and U32199 (N_32199,N_25190,N_29044);
and U32200 (N_32200,N_28947,N_28521);
or U32201 (N_32201,N_27266,N_27407);
or U32202 (N_32202,N_25795,N_25773);
or U32203 (N_32203,N_28685,N_27534);
or U32204 (N_32204,N_28883,N_29214);
xnor U32205 (N_32205,N_29763,N_28538);
nor U32206 (N_32206,N_28047,N_26072);
nand U32207 (N_32207,N_29243,N_27344);
nor U32208 (N_32208,N_25804,N_25040);
and U32209 (N_32209,N_25648,N_26262);
nor U32210 (N_32210,N_29430,N_26219);
xor U32211 (N_32211,N_28208,N_29736);
and U32212 (N_32212,N_27543,N_25738);
nand U32213 (N_32213,N_28996,N_29376);
and U32214 (N_32214,N_25717,N_25761);
xor U32215 (N_32215,N_25671,N_25334);
and U32216 (N_32216,N_26155,N_27968);
nor U32217 (N_32217,N_26408,N_25219);
nor U32218 (N_32218,N_29160,N_26506);
nor U32219 (N_32219,N_26107,N_26222);
nor U32220 (N_32220,N_28624,N_27401);
or U32221 (N_32221,N_25375,N_26514);
xnor U32222 (N_32222,N_25394,N_27557);
or U32223 (N_32223,N_27429,N_29522);
and U32224 (N_32224,N_25927,N_25748);
xnor U32225 (N_32225,N_28846,N_25353);
nand U32226 (N_32226,N_27325,N_26332);
nand U32227 (N_32227,N_28966,N_28176);
nor U32228 (N_32228,N_28467,N_25825);
or U32229 (N_32229,N_28816,N_29629);
nand U32230 (N_32230,N_26295,N_29816);
xor U32231 (N_32231,N_29815,N_26450);
nor U32232 (N_32232,N_29226,N_29887);
xnor U32233 (N_32233,N_28062,N_29196);
and U32234 (N_32234,N_26714,N_29341);
and U32235 (N_32235,N_29452,N_27864);
or U32236 (N_32236,N_28715,N_28269);
nand U32237 (N_32237,N_26927,N_29117);
xor U32238 (N_32238,N_25075,N_25329);
and U32239 (N_32239,N_26724,N_26059);
nand U32240 (N_32240,N_27848,N_28090);
nor U32241 (N_32241,N_28160,N_27391);
xnor U32242 (N_32242,N_27231,N_26654);
or U32243 (N_32243,N_27376,N_28789);
xnor U32244 (N_32244,N_29335,N_25518);
or U32245 (N_32245,N_26201,N_28867);
or U32246 (N_32246,N_25948,N_26089);
and U32247 (N_32247,N_25681,N_27139);
nand U32248 (N_32248,N_29193,N_25810);
xor U32249 (N_32249,N_29738,N_27105);
nor U32250 (N_32250,N_27361,N_29755);
and U32251 (N_32251,N_28749,N_29876);
nand U32252 (N_32252,N_29114,N_25714);
nor U32253 (N_32253,N_27206,N_29379);
nand U32254 (N_32254,N_28986,N_26525);
nor U32255 (N_32255,N_27884,N_26893);
nand U32256 (N_32256,N_27157,N_28844);
and U32257 (N_32257,N_29910,N_28594);
and U32258 (N_32258,N_25673,N_26298);
xor U32259 (N_32259,N_29663,N_25603);
nand U32260 (N_32260,N_25521,N_28829);
and U32261 (N_32261,N_28839,N_28690);
xnor U32262 (N_32262,N_29016,N_29296);
and U32263 (N_32263,N_26606,N_29285);
nor U32264 (N_32264,N_28901,N_25138);
and U32265 (N_32265,N_26550,N_25838);
and U32266 (N_32266,N_28282,N_29358);
xor U32267 (N_32267,N_26469,N_27988);
or U32268 (N_32268,N_27981,N_28124);
and U32269 (N_32269,N_26675,N_29018);
and U32270 (N_32270,N_29900,N_26358);
or U32271 (N_32271,N_28919,N_25880);
or U32272 (N_32272,N_26065,N_26049);
and U32273 (N_32273,N_29337,N_28766);
or U32274 (N_32274,N_25636,N_27166);
nor U32275 (N_32275,N_28206,N_28476);
xor U32276 (N_32276,N_28139,N_28853);
nor U32277 (N_32277,N_26961,N_25701);
or U32278 (N_32278,N_28852,N_27143);
or U32279 (N_32279,N_26911,N_26501);
xor U32280 (N_32280,N_29437,N_29959);
and U32281 (N_32281,N_28488,N_27337);
nand U32282 (N_32282,N_25033,N_27530);
nand U32283 (N_32283,N_27816,N_26233);
and U32284 (N_32284,N_25853,N_29340);
xnor U32285 (N_32285,N_25519,N_26296);
xnor U32286 (N_32286,N_25548,N_25096);
nand U32287 (N_32287,N_28031,N_25414);
and U32288 (N_32288,N_28403,N_27100);
and U32289 (N_32289,N_28713,N_25871);
xor U32290 (N_32290,N_28962,N_27364);
or U32291 (N_32291,N_25121,N_26818);
nand U32292 (N_32292,N_28540,N_25186);
or U32293 (N_32293,N_26908,N_29330);
nor U32294 (N_32294,N_28251,N_28265);
nand U32295 (N_32295,N_29690,N_27336);
and U32296 (N_32296,N_26573,N_27797);
and U32297 (N_32297,N_27740,N_25035);
or U32298 (N_32298,N_26746,N_29585);
or U32299 (N_32299,N_25119,N_28865);
and U32300 (N_32300,N_29670,N_29899);
nand U32301 (N_32301,N_27425,N_26411);
nor U32302 (N_32302,N_27971,N_27437);
xor U32303 (N_32303,N_27676,N_25937);
and U32304 (N_32304,N_28544,N_27082);
and U32305 (N_32305,N_25509,N_28840);
and U32306 (N_32306,N_28486,N_27351);
nor U32307 (N_32307,N_27208,N_27395);
and U32308 (N_32308,N_26419,N_26489);
xor U32309 (N_32309,N_28864,N_26208);
nor U32310 (N_32310,N_28227,N_28284);
or U32311 (N_32311,N_27901,N_26290);
nor U32312 (N_32312,N_25998,N_27643);
and U32313 (N_32313,N_29403,N_28580);
nor U32314 (N_32314,N_29846,N_29519);
nor U32315 (N_32315,N_26043,N_27876);
and U32316 (N_32316,N_27176,N_27519);
and U32317 (N_32317,N_26395,N_25462);
nand U32318 (N_32318,N_25994,N_25067);
or U32319 (N_32319,N_27043,N_27685);
xnor U32320 (N_32320,N_25970,N_26234);
nor U32321 (N_32321,N_25036,N_29953);
and U32322 (N_32322,N_29293,N_25776);
xnor U32323 (N_32323,N_25790,N_26126);
xnor U32324 (N_32324,N_27215,N_28889);
nand U32325 (N_32325,N_26768,N_27393);
nor U32326 (N_32326,N_25242,N_26463);
nor U32327 (N_32327,N_29433,N_26656);
xnor U32328 (N_32328,N_25388,N_29946);
nand U32329 (N_32329,N_25395,N_26470);
xor U32330 (N_32330,N_25399,N_26486);
xor U32331 (N_32331,N_28368,N_27874);
and U32332 (N_32332,N_25938,N_29921);
xnor U32333 (N_32333,N_28408,N_26728);
nand U32334 (N_32334,N_27012,N_28238);
or U32335 (N_32335,N_27201,N_28589);
and U32336 (N_32336,N_25410,N_27243);
and U32337 (N_32337,N_28152,N_29650);
nor U32338 (N_32338,N_27426,N_25258);
or U32339 (N_32339,N_28927,N_29642);
nand U32340 (N_32340,N_26627,N_29107);
nor U32341 (N_32341,N_29324,N_29952);
or U32342 (N_32342,N_29270,N_29989);
or U32343 (N_32343,N_28656,N_26755);
xor U32344 (N_32344,N_29779,N_26282);
nand U32345 (N_32345,N_25017,N_27608);
xor U32346 (N_32346,N_28278,N_26477);
nor U32347 (N_32347,N_28198,N_29142);
xnor U32348 (N_32348,N_27846,N_26042);
nand U32349 (N_32349,N_25222,N_25797);
nand U32350 (N_32350,N_27955,N_25416);
nor U32351 (N_32351,N_27487,N_28907);
xnor U32352 (N_32352,N_29401,N_25581);
and U32353 (N_32353,N_25630,N_27107);
or U32354 (N_32354,N_26504,N_29354);
nand U32355 (N_32355,N_26888,N_29465);
or U32356 (N_32356,N_29930,N_28879);
xnor U32357 (N_32357,N_29204,N_27663);
xnor U32358 (N_32358,N_25352,N_26382);
nand U32359 (N_32359,N_26026,N_29390);
nor U32360 (N_32360,N_28710,N_27609);
or U32361 (N_32361,N_25199,N_27120);
xnor U32362 (N_32362,N_26912,N_26505);
nor U32363 (N_32363,N_26953,N_25089);
nor U32364 (N_32364,N_29934,N_27825);
and U32365 (N_32365,N_25971,N_28338);
or U32366 (N_32366,N_26010,N_25098);
nand U32367 (N_32367,N_27040,N_28971);
or U32368 (N_32368,N_26694,N_27759);
or U32369 (N_32369,N_25901,N_27246);
nand U32370 (N_32370,N_29510,N_29552);
xor U32371 (N_32371,N_29714,N_28572);
and U32372 (N_32372,N_27127,N_29361);
nor U32373 (N_32373,N_25074,N_29912);
and U32374 (N_32374,N_28450,N_29718);
xor U32375 (N_32375,N_27207,N_25745);
nand U32376 (N_32376,N_26173,N_25502);
xor U32377 (N_32377,N_25336,N_25906);
and U32378 (N_32378,N_29314,N_25708);
xor U32379 (N_32379,N_26870,N_26782);
xor U32380 (N_32380,N_29651,N_27042);
nand U32381 (N_32381,N_26431,N_28178);
nor U32382 (N_32382,N_25148,N_27526);
nand U32383 (N_32383,N_27209,N_28891);
and U32384 (N_32384,N_27131,N_26164);
or U32385 (N_32385,N_29313,N_29498);
nand U32386 (N_32386,N_29336,N_28223);
nand U32387 (N_32387,N_25767,N_26802);
or U32388 (N_32388,N_25220,N_26251);
and U32389 (N_32389,N_29353,N_26985);
nand U32390 (N_32390,N_26056,N_29808);
xnor U32391 (N_32391,N_29695,N_29548);
nand U32392 (N_32392,N_25058,N_26969);
xor U32393 (N_32393,N_27418,N_29365);
nor U32394 (N_32394,N_26451,N_29883);
xnor U32395 (N_32395,N_27804,N_26418);
xor U32396 (N_32396,N_26844,N_25253);
xnor U32397 (N_32397,N_26004,N_27461);
xor U32398 (N_32398,N_28332,N_25124);
or U32399 (N_32399,N_25368,N_26741);
nor U32400 (N_32400,N_25318,N_26805);
xor U32401 (N_32401,N_28404,N_26935);
and U32402 (N_32402,N_26386,N_25621);
nand U32403 (N_32403,N_26218,N_27234);
nand U32404 (N_32404,N_29924,N_26345);
or U32405 (N_32405,N_29991,N_25865);
or U32406 (N_32406,N_27481,N_25269);
xor U32407 (N_32407,N_25189,N_26837);
xor U32408 (N_32408,N_28672,N_26914);
nor U32409 (N_32409,N_26053,N_25173);
nor U32410 (N_32410,N_25169,N_27508);
nor U32411 (N_32411,N_29780,N_27367);
or U32412 (N_32412,N_27154,N_28936);
xor U32413 (N_32413,N_25619,N_25832);
xnor U32414 (N_32414,N_25584,N_27567);
or U32415 (N_32415,N_25860,N_28639);
or U32416 (N_32416,N_28065,N_26153);
or U32417 (N_32417,N_29025,N_28229);
xor U32418 (N_32418,N_29583,N_25768);
and U32419 (N_32419,N_28929,N_28446);
nand U32420 (N_32420,N_28557,N_26002);
xnor U32421 (N_32421,N_26092,N_29397);
or U32422 (N_32422,N_27745,N_26937);
or U32423 (N_32423,N_25953,N_27652);
nor U32424 (N_32424,N_25959,N_29356);
and U32425 (N_32425,N_28009,N_27667);
or U32426 (N_32426,N_28813,N_25802);
and U32427 (N_32427,N_26180,N_26847);
and U32428 (N_32428,N_27933,N_25053);
or U32429 (N_32429,N_26903,N_29000);
xnor U32430 (N_32430,N_26849,N_27551);
and U32431 (N_32431,N_25583,N_29618);
nand U32432 (N_32432,N_26808,N_26983);
nand U32433 (N_32433,N_29096,N_27518);
xor U32434 (N_32434,N_29796,N_26025);
and U32435 (N_32435,N_29312,N_29513);
or U32436 (N_32436,N_25429,N_29219);
nand U32437 (N_32437,N_28693,N_28492);
xnor U32438 (N_32438,N_29523,N_28911);
nor U32439 (N_32439,N_29310,N_26142);
or U32440 (N_32440,N_29097,N_29783);
nor U32441 (N_32441,N_29157,N_28228);
xor U32442 (N_32442,N_26221,N_28916);
and U32443 (N_32443,N_26661,N_29784);
xor U32444 (N_32444,N_27476,N_29170);
or U32445 (N_32445,N_28199,N_27078);
nor U32446 (N_32446,N_27465,N_29857);
and U32447 (N_32447,N_25268,N_29885);
or U32448 (N_32448,N_27151,N_26679);
or U32449 (N_32449,N_28977,N_28663);
or U32450 (N_32450,N_29339,N_25208);
nor U32451 (N_32451,N_29859,N_29127);
and U32452 (N_32452,N_27730,N_28512);
and U32453 (N_32453,N_28216,N_28910);
or U32454 (N_32454,N_28355,N_26690);
or U32455 (N_32455,N_29161,N_27938);
or U32456 (N_32456,N_27034,N_27456);
nor U32457 (N_32457,N_26206,N_28729);
or U32458 (N_32458,N_26861,N_28406);
nor U32459 (N_32459,N_26217,N_28784);
or U32460 (N_32460,N_29124,N_29794);
and U32461 (N_32461,N_29933,N_26867);
xnor U32462 (N_32462,N_28577,N_29652);
and U32463 (N_32463,N_28281,N_28186);
nand U32464 (N_32464,N_26067,N_29010);
nor U32465 (N_32465,N_25896,N_27256);
nor U32466 (N_32466,N_27946,N_27852);
nand U32467 (N_32467,N_25886,N_29655);
and U32468 (N_32468,N_25451,N_25712);
nor U32469 (N_32469,N_29116,N_25130);
xor U32470 (N_32470,N_29215,N_28981);
nor U32471 (N_32471,N_26476,N_26350);
xor U32472 (N_32472,N_27313,N_29434);
nor U32473 (N_32473,N_26974,N_29809);
nand U32474 (N_32474,N_29198,N_27953);
nand U32475 (N_32475,N_25897,N_28383);
nand U32476 (N_32476,N_28290,N_27844);
nand U32477 (N_32477,N_27271,N_29400);
xor U32478 (N_32478,N_29889,N_28314);
or U32479 (N_32479,N_26516,N_27732);
nand U32480 (N_32480,N_25338,N_25527);
nor U32481 (N_32481,N_27547,N_27705);
and U32482 (N_32482,N_26998,N_26508);
xor U32483 (N_32483,N_29396,N_26299);
and U32484 (N_32484,N_28958,N_27934);
nand U32485 (N_32485,N_29442,N_27158);
nor U32486 (N_32486,N_28287,N_28389);
nand U32487 (N_32487,N_28079,N_27637);
nand U32488 (N_32488,N_29711,N_26120);
nand U32489 (N_32489,N_25123,N_28116);
or U32490 (N_32490,N_28518,N_26093);
xor U32491 (N_32491,N_25600,N_26537);
or U32492 (N_32492,N_27697,N_26140);
or U32493 (N_32493,N_28836,N_25467);
and U32494 (N_32494,N_25533,N_29440);
nor U32495 (N_32495,N_26834,N_26001);
nand U32496 (N_32496,N_27787,N_28259);
xnor U32497 (N_32497,N_25980,N_25273);
xor U32498 (N_32498,N_26214,N_25674);
nand U32499 (N_32499,N_28619,N_29919);
nand U32500 (N_32500,N_27529,N_25908);
and U32501 (N_32501,N_28126,N_29621);
or U32502 (N_32502,N_29358,N_29295);
and U32503 (N_32503,N_26133,N_26168);
and U32504 (N_32504,N_28563,N_26814);
and U32505 (N_32505,N_28416,N_27489);
nand U32506 (N_32506,N_26206,N_25387);
or U32507 (N_32507,N_25925,N_26551);
nand U32508 (N_32508,N_25179,N_27118);
or U32509 (N_32509,N_25488,N_25384);
or U32510 (N_32510,N_28214,N_25338);
and U32511 (N_32511,N_25519,N_29329);
nand U32512 (N_32512,N_27065,N_25811);
nor U32513 (N_32513,N_26995,N_27306);
or U32514 (N_32514,N_25567,N_29214);
and U32515 (N_32515,N_28043,N_28285);
and U32516 (N_32516,N_29997,N_26682);
nand U32517 (N_32517,N_29811,N_29784);
and U32518 (N_32518,N_28750,N_28635);
and U32519 (N_32519,N_26107,N_26332);
nor U32520 (N_32520,N_29176,N_27043);
xnor U32521 (N_32521,N_25628,N_25730);
or U32522 (N_32522,N_26812,N_27311);
nand U32523 (N_32523,N_26793,N_26679);
or U32524 (N_32524,N_28674,N_25874);
nand U32525 (N_32525,N_26734,N_27106);
nor U32526 (N_32526,N_26581,N_27678);
nand U32527 (N_32527,N_29129,N_27202);
or U32528 (N_32528,N_25706,N_25505);
or U32529 (N_32529,N_28836,N_26084);
xnor U32530 (N_32530,N_26306,N_25230);
xnor U32531 (N_32531,N_26536,N_29649);
and U32532 (N_32532,N_29853,N_25183);
or U32533 (N_32533,N_26141,N_25927);
nor U32534 (N_32534,N_25159,N_28812);
nand U32535 (N_32535,N_25724,N_25324);
and U32536 (N_32536,N_29863,N_29258);
xor U32537 (N_32537,N_26325,N_29844);
or U32538 (N_32538,N_25011,N_27026);
xor U32539 (N_32539,N_25251,N_26960);
and U32540 (N_32540,N_27639,N_29717);
nand U32541 (N_32541,N_26610,N_26884);
or U32542 (N_32542,N_29714,N_25084);
nor U32543 (N_32543,N_29624,N_26539);
and U32544 (N_32544,N_27384,N_26997);
nor U32545 (N_32545,N_28552,N_26408);
and U32546 (N_32546,N_28671,N_26122);
and U32547 (N_32547,N_29551,N_25415);
xor U32548 (N_32548,N_27612,N_29595);
nand U32549 (N_32549,N_25947,N_27468);
nor U32550 (N_32550,N_25770,N_28403);
xnor U32551 (N_32551,N_27567,N_28927);
and U32552 (N_32552,N_25200,N_29492);
nand U32553 (N_32553,N_27801,N_25232);
or U32554 (N_32554,N_27836,N_29360);
and U32555 (N_32555,N_29549,N_27335);
and U32556 (N_32556,N_25774,N_28596);
xor U32557 (N_32557,N_27128,N_26283);
or U32558 (N_32558,N_29623,N_29157);
or U32559 (N_32559,N_25323,N_26339);
and U32560 (N_32560,N_25639,N_27353);
nor U32561 (N_32561,N_25405,N_26758);
nand U32562 (N_32562,N_27879,N_26949);
or U32563 (N_32563,N_29142,N_27279);
nand U32564 (N_32564,N_25253,N_28450);
or U32565 (N_32565,N_25347,N_28762);
nand U32566 (N_32566,N_28794,N_28556);
and U32567 (N_32567,N_27519,N_27552);
xor U32568 (N_32568,N_28511,N_29290);
nor U32569 (N_32569,N_26712,N_27240);
or U32570 (N_32570,N_25678,N_26201);
or U32571 (N_32571,N_27357,N_28331);
nor U32572 (N_32572,N_27081,N_27583);
xor U32573 (N_32573,N_29011,N_28537);
and U32574 (N_32574,N_29503,N_27660);
nand U32575 (N_32575,N_27836,N_28353);
xor U32576 (N_32576,N_27220,N_27334);
xnor U32577 (N_32577,N_28322,N_28425);
xor U32578 (N_32578,N_27479,N_28685);
and U32579 (N_32579,N_26858,N_26521);
nor U32580 (N_32580,N_28047,N_29583);
and U32581 (N_32581,N_28433,N_29436);
xor U32582 (N_32582,N_29793,N_26539);
and U32583 (N_32583,N_25192,N_25801);
xor U32584 (N_32584,N_26626,N_29005);
or U32585 (N_32585,N_29674,N_27372);
nor U32586 (N_32586,N_29001,N_28839);
nor U32587 (N_32587,N_25761,N_25953);
xor U32588 (N_32588,N_25492,N_29972);
or U32589 (N_32589,N_25850,N_26115);
nand U32590 (N_32590,N_29435,N_26622);
nand U32591 (N_32591,N_27768,N_28901);
nor U32592 (N_32592,N_27879,N_28343);
and U32593 (N_32593,N_25693,N_28270);
or U32594 (N_32594,N_26517,N_25938);
xnor U32595 (N_32595,N_25741,N_25517);
and U32596 (N_32596,N_27679,N_27006);
nor U32597 (N_32597,N_28287,N_26748);
and U32598 (N_32598,N_27984,N_27005);
nor U32599 (N_32599,N_26074,N_26064);
or U32600 (N_32600,N_29936,N_27337);
and U32601 (N_32601,N_28606,N_27751);
xnor U32602 (N_32602,N_29005,N_29198);
and U32603 (N_32603,N_25298,N_25764);
nor U32604 (N_32604,N_25836,N_29278);
nor U32605 (N_32605,N_27294,N_28783);
and U32606 (N_32606,N_28100,N_26460);
xnor U32607 (N_32607,N_29555,N_27490);
nand U32608 (N_32608,N_27509,N_29676);
nand U32609 (N_32609,N_28286,N_29501);
and U32610 (N_32610,N_28233,N_29501);
nor U32611 (N_32611,N_29075,N_27207);
and U32612 (N_32612,N_28139,N_26296);
xnor U32613 (N_32613,N_28752,N_28943);
and U32614 (N_32614,N_27680,N_29880);
and U32615 (N_32615,N_26926,N_25060);
xnor U32616 (N_32616,N_27015,N_28870);
and U32617 (N_32617,N_26997,N_29689);
or U32618 (N_32618,N_28056,N_26281);
xnor U32619 (N_32619,N_25605,N_29345);
nand U32620 (N_32620,N_28348,N_25348);
nor U32621 (N_32621,N_26233,N_29703);
or U32622 (N_32622,N_28042,N_27486);
and U32623 (N_32623,N_27733,N_29712);
xor U32624 (N_32624,N_26122,N_29509);
or U32625 (N_32625,N_29561,N_26941);
xor U32626 (N_32626,N_29540,N_25219);
or U32627 (N_32627,N_26327,N_28639);
and U32628 (N_32628,N_29941,N_25795);
or U32629 (N_32629,N_25662,N_29439);
and U32630 (N_32630,N_26735,N_29548);
nand U32631 (N_32631,N_26829,N_29442);
nor U32632 (N_32632,N_29499,N_25587);
xnor U32633 (N_32633,N_26972,N_25219);
nand U32634 (N_32634,N_26424,N_25832);
nand U32635 (N_32635,N_26216,N_27760);
or U32636 (N_32636,N_25509,N_27167);
xor U32637 (N_32637,N_26837,N_29586);
and U32638 (N_32638,N_28810,N_27533);
or U32639 (N_32639,N_29429,N_26417);
nand U32640 (N_32640,N_29059,N_27432);
xnor U32641 (N_32641,N_29219,N_26298);
and U32642 (N_32642,N_28809,N_25252);
and U32643 (N_32643,N_26915,N_25526);
xor U32644 (N_32644,N_28777,N_25194);
and U32645 (N_32645,N_25467,N_28163);
nor U32646 (N_32646,N_26415,N_26387);
nor U32647 (N_32647,N_26435,N_25678);
nand U32648 (N_32648,N_29598,N_26948);
nor U32649 (N_32649,N_25593,N_28636);
and U32650 (N_32650,N_25069,N_28425);
xnor U32651 (N_32651,N_27837,N_27556);
or U32652 (N_32652,N_28009,N_25954);
or U32653 (N_32653,N_28726,N_25128);
or U32654 (N_32654,N_29512,N_25864);
nand U32655 (N_32655,N_27144,N_29303);
xnor U32656 (N_32656,N_29684,N_29149);
xor U32657 (N_32657,N_27477,N_28645);
nand U32658 (N_32658,N_29248,N_27513);
and U32659 (N_32659,N_28623,N_27660);
nand U32660 (N_32660,N_27839,N_26777);
or U32661 (N_32661,N_26889,N_27745);
nor U32662 (N_32662,N_28559,N_25676);
and U32663 (N_32663,N_29839,N_26380);
nor U32664 (N_32664,N_28834,N_25456);
nand U32665 (N_32665,N_29255,N_27159);
xor U32666 (N_32666,N_25260,N_25198);
or U32667 (N_32667,N_26949,N_25805);
xor U32668 (N_32668,N_27494,N_26782);
or U32669 (N_32669,N_25193,N_25840);
nor U32670 (N_32670,N_27001,N_29552);
and U32671 (N_32671,N_25359,N_25695);
nand U32672 (N_32672,N_28278,N_28255);
nor U32673 (N_32673,N_27321,N_26548);
or U32674 (N_32674,N_28950,N_27548);
xnor U32675 (N_32675,N_26630,N_25687);
nand U32676 (N_32676,N_28155,N_28396);
or U32677 (N_32677,N_25218,N_26399);
nand U32678 (N_32678,N_27626,N_29159);
nand U32679 (N_32679,N_28790,N_29639);
and U32680 (N_32680,N_28784,N_25410);
xnor U32681 (N_32681,N_27550,N_25005);
nor U32682 (N_32682,N_27331,N_26940);
and U32683 (N_32683,N_25469,N_28695);
xnor U32684 (N_32684,N_27295,N_25617);
xor U32685 (N_32685,N_29943,N_26623);
nand U32686 (N_32686,N_25531,N_29804);
nand U32687 (N_32687,N_28183,N_29525);
and U32688 (N_32688,N_27551,N_25082);
nor U32689 (N_32689,N_27418,N_26026);
nand U32690 (N_32690,N_27835,N_26349);
or U32691 (N_32691,N_25496,N_28440);
xor U32692 (N_32692,N_25559,N_26577);
nand U32693 (N_32693,N_28067,N_29652);
and U32694 (N_32694,N_26448,N_27266);
and U32695 (N_32695,N_29859,N_26603);
nand U32696 (N_32696,N_28640,N_26878);
xnor U32697 (N_32697,N_27882,N_29161);
and U32698 (N_32698,N_25303,N_28432);
nand U32699 (N_32699,N_27314,N_27409);
or U32700 (N_32700,N_29560,N_27219);
nand U32701 (N_32701,N_29900,N_25519);
and U32702 (N_32702,N_25873,N_27055);
xnor U32703 (N_32703,N_29256,N_28808);
nand U32704 (N_32704,N_29644,N_28165);
or U32705 (N_32705,N_29866,N_25794);
and U32706 (N_32706,N_25647,N_29050);
nand U32707 (N_32707,N_28381,N_26487);
nand U32708 (N_32708,N_26466,N_26985);
nor U32709 (N_32709,N_27011,N_25009);
and U32710 (N_32710,N_25032,N_28605);
xor U32711 (N_32711,N_27474,N_26480);
and U32712 (N_32712,N_28411,N_26320);
nand U32713 (N_32713,N_26546,N_29540);
nor U32714 (N_32714,N_26639,N_29921);
nor U32715 (N_32715,N_25586,N_25536);
nor U32716 (N_32716,N_27208,N_25371);
nand U32717 (N_32717,N_28808,N_28834);
or U32718 (N_32718,N_25633,N_28278);
nor U32719 (N_32719,N_28603,N_26491);
and U32720 (N_32720,N_29232,N_26812);
and U32721 (N_32721,N_26734,N_29091);
nor U32722 (N_32722,N_28769,N_28465);
xor U32723 (N_32723,N_28182,N_28214);
and U32724 (N_32724,N_25696,N_27796);
nand U32725 (N_32725,N_25636,N_25067);
nor U32726 (N_32726,N_28360,N_25178);
xor U32727 (N_32727,N_26545,N_25237);
and U32728 (N_32728,N_29929,N_29094);
or U32729 (N_32729,N_28253,N_28812);
and U32730 (N_32730,N_25353,N_28993);
and U32731 (N_32731,N_27720,N_28530);
or U32732 (N_32732,N_28904,N_25966);
or U32733 (N_32733,N_27593,N_25718);
xor U32734 (N_32734,N_25739,N_28686);
or U32735 (N_32735,N_28422,N_27187);
and U32736 (N_32736,N_25638,N_29520);
or U32737 (N_32737,N_28178,N_27151);
nand U32738 (N_32738,N_27559,N_28700);
nand U32739 (N_32739,N_27200,N_28546);
xnor U32740 (N_32740,N_26102,N_29850);
or U32741 (N_32741,N_29793,N_27844);
xor U32742 (N_32742,N_27269,N_28992);
or U32743 (N_32743,N_29946,N_25585);
or U32744 (N_32744,N_25294,N_28383);
or U32745 (N_32745,N_25838,N_27307);
or U32746 (N_32746,N_25759,N_27699);
or U32747 (N_32747,N_29321,N_27120);
nor U32748 (N_32748,N_29261,N_26121);
nor U32749 (N_32749,N_28110,N_28834);
nand U32750 (N_32750,N_28892,N_27787);
xnor U32751 (N_32751,N_27042,N_28841);
nand U32752 (N_32752,N_26277,N_29073);
nor U32753 (N_32753,N_27839,N_26358);
and U32754 (N_32754,N_25688,N_25005);
xnor U32755 (N_32755,N_27756,N_27506);
nor U32756 (N_32756,N_25857,N_28148);
and U32757 (N_32757,N_27212,N_26670);
or U32758 (N_32758,N_27579,N_26794);
nor U32759 (N_32759,N_25669,N_29439);
nor U32760 (N_32760,N_28943,N_28306);
xnor U32761 (N_32761,N_25276,N_27648);
nand U32762 (N_32762,N_26708,N_28637);
nor U32763 (N_32763,N_28216,N_25425);
nor U32764 (N_32764,N_25532,N_26399);
or U32765 (N_32765,N_25012,N_29761);
nor U32766 (N_32766,N_25731,N_28685);
nand U32767 (N_32767,N_26314,N_28111);
and U32768 (N_32768,N_27468,N_29250);
nand U32769 (N_32769,N_29933,N_29418);
xnor U32770 (N_32770,N_27051,N_25252);
nor U32771 (N_32771,N_26412,N_27464);
nor U32772 (N_32772,N_29116,N_26530);
nand U32773 (N_32773,N_27666,N_27333);
or U32774 (N_32774,N_28052,N_25521);
nand U32775 (N_32775,N_26995,N_26159);
nand U32776 (N_32776,N_27525,N_25617);
nand U32777 (N_32777,N_25439,N_25284);
nand U32778 (N_32778,N_26483,N_27574);
xor U32779 (N_32779,N_27804,N_29044);
and U32780 (N_32780,N_25325,N_27193);
nand U32781 (N_32781,N_27900,N_29095);
and U32782 (N_32782,N_27984,N_28158);
xnor U32783 (N_32783,N_28295,N_29463);
xnor U32784 (N_32784,N_26613,N_27867);
nor U32785 (N_32785,N_29852,N_28140);
or U32786 (N_32786,N_27025,N_28889);
or U32787 (N_32787,N_28152,N_25614);
nand U32788 (N_32788,N_27925,N_25160);
nor U32789 (N_32789,N_26310,N_27719);
nor U32790 (N_32790,N_25198,N_28033);
nor U32791 (N_32791,N_25308,N_28906);
or U32792 (N_32792,N_28610,N_29433);
or U32793 (N_32793,N_25528,N_27636);
nor U32794 (N_32794,N_29816,N_26846);
and U32795 (N_32795,N_25626,N_28944);
or U32796 (N_32796,N_28452,N_27977);
nand U32797 (N_32797,N_28657,N_29612);
or U32798 (N_32798,N_25957,N_28230);
nor U32799 (N_32799,N_25488,N_25257);
nand U32800 (N_32800,N_27804,N_29437);
xnor U32801 (N_32801,N_29794,N_25162);
and U32802 (N_32802,N_28749,N_26601);
xnor U32803 (N_32803,N_28674,N_28253);
nand U32804 (N_32804,N_28190,N_27258);
nand U32805 (N_32805,N_26207,N_29273);
nand U32806 (N_32806,N_29991,N_28015);
nand U32807 (N_32807,N_25854,N_27795);
and U32808 (N_32808,N_29744,N_28173);
nand U32809 (N_32809,N_29247,N_28128);
nand U32810 (N_32810,N_26092,N_25883);
nor U32811 (N_32811,N_25570,N_29322);
or U32812 (N_32812,N_27814,N_29418);
nor U32813 (N_32813,N_27742,N_29129);
nand U32814 (N_32814,N_26973,N_29228);
nand U32815 (N_32815,N_28342,N_25266);
nand U32816 (N_32816,N_25002,N_26539);
or U32817 (N_32817,N_25492,N_28319);
and U32818 (N_32818,N_26806,N_29209);
or U32819 (N_32819,N_26177,N_26348);
or U32820 (N_32820,N_29611,N_26344);
or U32821 (N_32821,N_28159,N_25658);
xnor U32822 (N_32822,N_25593,N_27746);
nor U32823 (N_32823,N_27626,N_29907);
xnor U32824 (N_32824,N_25333,N_27947);
nand U32825 (N_32825,N_27867,N_26978);
xor U32826 (N_32826,N_29019,N_28196);
xor U32827 (N_32827,N_26686,N_28732);
or U32828 (N_32828,N_26912,N_25942);
or U32829 (N_32829,N_26998,N_29056);
and U32830 (N_32830,N_26736,N_27525);
nand U32831 (N_32831,N_26029,N_29234);
nor U32832 (N_32832,N_28157,N_26601);
xnor U32833 (N_32833,N_27537,N_25996);
xnor U32834 (N_32834,N_25219,N_25678);
xnor U32835 (N_32835,N_25604,N_25960);
or U32836 (N_32836,N_26003,N_28238);
nand U32837 (N_32837,N_29121,N_25007);
nor U32838 (N_32838,N_28672,N_25629);
xnor U32839 (N_32839,N_25094,N_25130);
and U32840 (N_32840,N_25481,N_26066);
nor U32841 (N_32841,N_26606,N_27619);
xor U32842 (N_32842,N_29741,N_29573);
nor U32843 (N_32843,N_27040,N_29138);
and U32844 (N_32844,N_27982,N_25122);
nand U32845 (N_32845,N_27821,N_27372);
xor U32846 (N_32846,N_27594,N_26336);
nand U32847 (N_32847,N_29362,N_27628);
nand U32848 (N_32848,N_28889,N_27471);
and U32849 (N_32849,N_26315,N_28878);
nand U32850 (N_32850,N_27446,N_25911);
and U32851 (N_32851,N_25914,N_29888);
xor U32852 (N_32852,N_27875,N_29027);
nand U32853 (N_32853,N_28410,N_28692);
nand U32854 (N_32854,N_27707,N_29399);
or U32855 (N_32855,N_29440,N_27321);
nor U32856 (N_32856,N_25490,N_28354);
and U32857 (N_32857,N_29412,N_29218);
xor U32858 (N_32858,N_28370,N_25248);
or U32859 (N_32859,N_26714,N_25170);
xnor U32860 (N_32860,N_28786,N_27298);
nand U32861 (N_32861,N_29597,N_27240);
nor U32862 (N_32862,N_27573,N_26920);
nand U32863 (N_32863,N_25242,N_28415);
nor U32864 (N_32864,N_27156,N_26239);
nor U32865 (N_32865,N_26355,N_27905);
xnor U32866 (N_32866,N_28537,N_27714);
xnor U32867 (N_32867,N_28065,N_28290);
and U32868 (N_32868,N_29479,N_26605);
and U32869 (N_32869,N_28306,N_27303);
nand U32870 (N_32870,N_29573,N_25910);
nor U32871 (N_32871,N_27093,N_28644);
or U32872 (N_32872,N_28236,N_28375);
and U32873 (N_32873,N_28281,N_29781);
xnor U32874 (N_32874,N_27962,N_27914);
and U32875 (N_32875,N_25170,N_28129);
and U32876 (N_32876,N_25857,N_26562);
nand U32877 (N_32877,N_26621,N_28775);
nor U32878 (N_32878,N_28229,N_28437);
nor U32879 (N_32879,N_28777,N_29278);
nor U32880 (N_32880,N_27212,N_27642);
and U32881 (N_32881,N_26115,N_25694);
nor U32882 (N_32882,N_26957,N_27464);
nand U32883 (N_32883,N_29790,N_25957);
nor U32884 (N_32884,N_26914,N_27478);
nor U32885 (N_32885,N_25197,N_29317);
nor U32886 (N_32886,N_29072,N_28448);
xnor U32887 (N_32887,N_29072,N_26635);
nor U32888 (N_32888,N_29251,N_25013);
or U32889 (N_32889,N_29616,N_26098);
and U32890 (N_32890,N_28082,N_25820);
nor U32891 (N_32891,N_28852,N_27159);
nor U32892 (N_32892,N_26562,N_26610);
nand U32893 (N_32893,N_27201,N_28430);
xor U32894 (N_32894,N_27881,N_29499);
nor U32895 (N_32895,N_29920,N_27804);
and U32896 (N_32896,N_29675,N_29966);
xnor U32897 (N_32897,N_27267,N_27898);
nor U32898 (N_32898,N_28571,N_29298);
nand U32899 (N_32899,N_25303,N_26449);
or U32900 (N_32900,N_29381,N_26993);
xor U32901 (N_32901,N_26131,N_27528);
xnor U32902 (N_32902,N_29325,N_28340);
nand U32903 (N_32903,N_25863,N_27008);
nor U32904 (N_32904,N_25753,N_26855);
nand U32905 (N_32905,N_25836,N_29201);
nand U32906 (N_32906,N_27930,N_26152);
and U32907 (N_32907,N_26218,N_25835);
or U32908 (N_32908,N_26378,N_28412);
or U32909 (N_32909,N_29084,N_29106);
nand U32910 (N_32910,N_25658,N_26514);
nor U32911 (N_32911,N_26684,N_29038);
and U32912 (N_32912,N_28234,N_27677);
xnor U32913 (N_32913,N_25297,N_27539);
xnor U32914 (N_32914,N_26897,N_26467);
nor U32915 (N_32915,N_26385,N_29125);
nand U32916 (N_32916,N_28095,N_25056);
or U32917 (N_32917,N_27241,N_28783);
nand U32918 (N_32918,N_28125,N_25889);
nor U32919 (N_32919,N_26868,N_29110);
nor U32920 (N_32920,N_25618,N_25594);
nand U32921 (N_32921,N_27343,N_28554);
and U32922 (N_32922,N_29908,N_26691);
nor U32923 (N_32923,N_25436,N_26213);
xnor U32924 (N_32924,N_27767,N_29412);
and U32925 (N_32925,N_27594,N_29628);
xnor U32926 (N_32926,N_26452,N_29051);
xnor U32927 (N_32927,N_29267,N_26591);
nand U32928 (N_32928,N_27731,N_29156);
nand U32929 (N_32929,N_27241,N_25769);
nand U32930 (N_32930,N_25212,N_29957);
nand U32931 (N_32931,N_28847,N_29920);
nor U32932 (N_32932,N_25269,N_25572);
xnor U32933 (N_32933,N_26150,N_27040);
or U32934 (N_32934,N_29464,N_28917);
and U32935 (N_32935,N_27450,N_26179);
and U32936 (N_32936,N_26134,N_26014);
nor U32937 (N_32937,N_25953,N_28868);
and U32938 (N_32938,N_25078,N_25836);
or U32939 (N_32939,N_29855,N_29822);
nor U32940 (N_32940,N_28604,N_29864);
nand U32941 (N_32941,N_26307,N_25262);
nand U32942 (N_32942,N_27621,N_28618);
xor U32943 (N_32943,N_29994,N_29707);
and U32944 (N_32944,N_29500,N_29994);
xor U32945 (N_32945,N_29614,N_27777);
nor U32946 (N_32946,N_26594,N_27165);
xor U32947 (N_32947,N_28896,N_28886);
or U32948 (N_32948,N_29695,N_25425);
xor U32949 (N_32949,N_25416,N_28585);
nand U32950 (N_32950,N_27477,N_26449);
xnor U32951 (N_32951,N_28775,N_29219);
and U32952 (N_32952,N_28075,N_29399);
nand U32953 (N_32953,N_27206,N_26833);
nor U32954 (N_32954,N_27483,N_29980);
nor U32955 (N_32955,N_28314,N_29724);
xnor U32956 (N_32956,N_27584,N_27692);
or U32957 (N_32957,N_27351,N_25485);
nand U32958 (N_32958,N_29596,N_28137);
nand U32959 (N_32959,N_26113,N_27116);
or U32960 (N_32960,N_27247,N_28884);
and U32961 (N_32961,N_25611,N_28925);
nand U32962 (N_32962,N_26360,N_28878);
or U32963 (N_32963,N_27919,N_28295);
xnor U32964 (N_32964,N_26650,N_26275);
xnor U32965 (N_32965,N_28076,N_25272);
or U32966 (N_32966,N_29191,N_25877);
xor U32967 (N_32967,N_25832,N_28069);
and U32968 (N_32968,N_26096,N_25814);
nor U32969 (N_32969,N_29046,N_25861);
xnor U32970 (N_32970,N_28808,N_27480);
xor U32971 (N_32971,N_25520,N_27705);
or U32972 (N_32972,N_28853,N_27185);
or U32973 (N_32973,N_29894,N_26255);
nor U32974 (N_32974,N_29019,N_26239);
and U32975 (N_32975,N_29440,N_29579);
nand U32976 (N_32976,N_25281,N_26732);
nor U32977 (N_32977,N_27296,N_26061);
nor U32978 (N_32978,N_28127,N_27538);
and U32979 (N_32979,N_26034,N_27602);
nor U32980 (N_32980,N_25038,N_29702);
or U32981 (N_32981,N_25789,N_29242);
and U32982 (N_32982,N_28718,N_26213);
and U32983 (N_32983,N_27730,N_26742);
and U32984 (N_32984,N_29959,N_26610);
nor U32985 (N_32985,N_25291,N_28974);
xor U32986 (N_32986,N_25279,N_28101);
xor U32987 (N_32987,N_26476,N_27703);
nor U32988 (N_32988,N_29643,N_29516);
nand U32989 (N_32989,N_27010,N_25026);
xor U32990 (N_32990,N_25878,N_27338);
and U32991 (N_32991,N_26384,N_27596);
and U32992 (N_32992,N_25662,N_29010);
nand U32993 (N_32993,N_28196,N_28534);
nand U32994 (N_32994,N_27984,N_25311);
nand U32995 (N_32995,N_28502,N_27591);
or U32996 (N_32996,N_25954,N_27597);
nand U32997 (N_32997,N_25907,N_28624);
or U32998 (N_32998,N_29063,N_25148);
xnor U32999 (N_32999,N_27033,N_29926);
and U33000 (N_33000,N_28353,N_25323);
or U33001 (N_33001,N_29835,N_25956);
nor U33002 (N_33002,N_28055,N_27307);
and U33003 (N_33003,N_27641,N_25594);
nand U33004 (N_33004,N_27302,N_26498);
and U33005 (N_33005,N_27880,N_27043);
and U33006 (N_33006,N_25971,N_25827);
nor U33007 (N_33007,N_25811,N_27860);
and U33008 (N_33008,N_25512,N_26391);
and U33009 (N_33009,N_29498,N_28515);
nor U33010 (N_33010,N_26320,N_25689);
or U33011 (N_33011,N_25801,N_28049);
xnor U33012 (N_33012,N_28089,N_28378);
and U33013 (N_33013,N_26353,N_25624);
xor U33014 (N_33014,N_29776,N_29530);
xnor U33015 (N_33015,N_28829,N_26063);
xor U33016 (N_33016,N_27767,N_25506);
xor U33017 (N_33017,N_25881,N_28479);
nor U33018 (N_33018,N_27554,N_26865);
xor U33019 (N_33019,N_25136,N_26163);
and U33020 (N_33020,N_25338,N_25774);
and U33021 (N_33021,N_27965,N_27263);
and U33022 (N_33022,N_26578,N_29612);
and U33023 (N_33023,N_25934,N_26287);
or U33024 (N_33024,N_28659,N_25226);
xor U33025 (N_33025,N_26498,N_26533);
nand U33026 (N_33026,N_26123,N_27268);
nor U33027 (N_33027,N_26302,N_25745);
nor U33028 (N_33028,N_25358,N_27509);
xnor U33029 (N_33029,N_29023,N_28447);
xnor U33030 (N_33030,N_26691,N_26457);
xor U33031 (N_33031,N_25538,N_28637);
nand U33032 (N_33032,N_25191,N_26080);
nand U33033 (N_33033,N_28256,N_29767);
xor U33034 (N_33034,N_27536,N_28925);
xor U33035 (N_33035,N_29242,N_26317);
nand U33036 (N_33036,N_28130,N_26820);
or U33037 (N_33037,N_28067,N_28657);
or U33038 (N_33038,N_29981,N_27747);
nand U33039 (N_33039,N_27043,N_26308);
and U33040 (N_33040,N_29072,N_26208);
or U33041 (N_33041,N_25158,N_26532);
or U33042 (N_33042,N_29141,N_25315);
or U33043 (N_33043,N_26591,N_28358);
or U33044 (N_33044,N_27109,N_28150);
nor U33045 (N_33045,N_28222,N_29098);
or U33046 (N_33046,N_26686,N_28114);
nor U33047 (N_33047,N_25356,N_29307);
nor U33048 (N_33048,N_28545,N_25507);
nand U33049 (N_33049,N_26823,N_27275);
and U33050 (N_33050,N_26165,N_25242);
nor U33051 (N_33051,N_25192,N_29617);
and U33052 (N_33052,N_27346,N_25884);
xnor U33053 (N_33053,N_26378,N_25007);
nand U33054 (N_33054,N_25393,N_26108);
xor U33055 (N_33055,N_27992,N_29755);
and U33056 (N_33056,N_25782,N_29837);
nand U33057 (N_33057,N_26761,N_28675);
nor U33058 (N_33058,N_28985,N_28808);
nor U33059 (N_33059,N_25479,N_28144);
nor U33060 (N_33060,N_29413,N_29869);
nand U33061 (N_33061,N_25706,N_26006);
or U33062 (N_33062,N_26461,N_28615);
or U33063 (N_33063,N_29844,N_26885);
or U33064 (N_33064,N_26762,N_25260);
nand U33065 (N_33065,N_28394,N_29353);
or U33066 (N_33066,N_29465,N_29140);
nand U33067 (N_33067,N_25634,N_26444);
xor U33068 (N_33068,N_25871,N_28449);
nor U33069 (N_33069,N_26877,N_29599);
nor U33070 (N_33070,N_25087,N_29067);
nor U33071 (N_33071,N_26718,N_29217);
nor U33072 (N_33072,N_27975,N_25936);
and U33073 (N_33073,N_25317,N_25446);
and U33074 (N_33074,N_27076,N_29124);
or U33075 (N_33075,N_25495,N_28700);
nor U33076 (N_33076,N_26541,N_29895);
nand U33077 (N_33077,N_27786,N_29118);
nor U33078 (N_33078,N_27883,N_25687);
xor U33079 (N_33079,N_27281,N_28590);
nand U33080 (N_33080,N_25491,N_29647);
nand U33081 (N_33081,N_28065,N_27959);
nand U33082 (N_33082,N_26580,N_27851);
or U33083 (N_33083,N_28194,N_25152);
or U33084 (N_33084,N_26051,N_28761);
and U33085 (N_33085,N_25790,N_25594);
or U33086 (N_33086,N_28663,N_26223);
or U33087 (N_33087,N_29666,N_26418);
nand U33088 (N_33088,N_27297,N_25574);
and U33089 (N_33089,N_27961,N_27991);
and U33090 (N_33090,N_29536,N_27333);
and U33091 (N_33091,N_26474,N_29279);
and U33092 (N_33092,N_25942,N_29883);
nor U33093 (N_33093,N_27254,N_26729);
nand U33094 (N_33094,N_25724,N_29683);
nand U33095 (N_33095,N_25689,N_29430);
nor U33096 (N_33096,N_27359,N_25760);
nor U33097 (N_33097,N_27226,N_29684);
nor U33098 (N_33098,N_25368,N_26775);
nand U33099 (N_33099,N_29612,N_25401);
nand U33100 (N_33100,N_29251,N_28375);
xor U33101 (N_33101,N_28896,N_27140);
xnor U33102 (N_33102,N_25804,N_28386);
or U33103 (N_33103,N_28781,N_27348);
or U33104 (N_33104,N_27624,N_28114);
or U33105 (N_33105,N_27405,N_27744);
and U33106 (N_33106,N_29649,N_26056);
nor U33107 (N_33107,N_25396,N_27123);
and U33108 (N_33108,N_27635,N_27399);
and U33109 (N_33109,N_28766,N_29257);
nand U33110 (N_33110,N_25118,N_25576);
nor U33111 (N_33111,N_29536,N_27491);
and U33112 (N_33112,N_27183,N_27185);
nand U33113 (N_33113,N_28952,N_27844);
nand U33114 (N_33114,N_26785,N_27849);
nor U33115 (N_33115,N_27106,N_26441);
nand U33116 (N_33116,N_25913,N_29485);
or U33117 (N_33117,N_26360,N_29521);
and U33118 (N_33118,N_26941,N_26450);
nor U33119 (N_33119,N_28687,N_29118);
nand U33120 (N_33120,N_27582,N_29443);
nand U33121 (N_33121,N_25270,N_25931);
or U33122 (N_33122,N_29833,N_28026);
or U33123 (N_33123,N_27304,N_29214);
or U33124 (N_33124,N_25550,N_29520);
nor U33125 (N_33125,N_28289,N_26299);
and U33126 (N_33126,N_26927,N_26775);
and U33127 (N_33127,N_26723,N_25265);
or U33128 (N_33128,N_26886,N_27294);
or U33129 (N_33129,N_29916,N_29642);
xnor U33130 (N_33130,N_27124,N_26029);
nand U33131 (N_33131,N_28137,N_25665);
nand U33132 (N_33132,N_27354,N_27607);
nor U33133 (N_33133,N_29727,N_28928);
and U33134 (N_33134,N_26956,N_27933);
or U33135 (N_33135,N_25107,N_26024);
and U33136 (N_33136,N_28087,N_27344);
and U33137 (N_33137,N_26585,N_27570);
or U33138 (N_33138,N_28558,N_29677);
nand U33139 (N_33139,N_29028,N_27932);
and U33140 (N_33140,N_25308,N_26615);
xor U33141 (N_33141,N_25545,N_25183);
nand U33142 (N_33142,N_27570,N_25804);
and U33143 (N_33143,N_27615,N_25487);
and U33144 (N_33144,N_26536,N_27793);
and U33145 (N_33145,N_25773,N_26649);
and U33146 (N_33146,N_26550,N_29106);
and U33147 (N_33147,N_26756,N_29139);
nor U33148 (N_33148,N_29270,N_25432);
nor U33149 (N_33149,N_28197,N_28817);
nand U33150 (N_33150,N_25416,N_29982);
nand U33151 (N_33151,N_26170,N_28736);
nand U33152 (N_33152,N_25025,N_28531);
nor U33153 (N_33153,N_29937,N_28027);
xor U33154 (N_33154,N_25459,N_28560);
and U33155 (N_33155,N_27040,N_26064);
nand U33156 (N_33156,N_26045,N_29653);
or U33157 (N_33157,N_25261,N_25547);
xor U33158 (N_33158,N_28430,N_25954);
nor U33159 (N_33159,N_28229,N_26959);
or U33160 (N_33160,N_26861,N_25809);
nor U33161 (N_33161,N_27298,N_25671);
or U33162 (N_33162,N_28767,N_26947);
and U33163 (N_33163,N_29951,N_26722);
or U33164 (N_33164,N_27816,N_29325);
or U33165 (N_33165,N_26269,N_25166);
nor U33166 (N_33166,N_26302,N_25224);
xor U33167 (N_33167,N_27698,N_28436);
or U33168 (N_33168,N_28965,N_29368);
and U33169 (N_33169,N_28322,N_27690);
and U33170 (N_33170,N_26088,N_25085);
xor U33171 (N_33171,N_29030,N_27367);
xor U33172 (N_33172,N_27039,N_25395);
nand U33173 (N_33173,N_26453,N_26258);
xor U33174 (N_33174,N_25264,N_29572);
and U33175 (N_33175,N_25453,N_29319);
and U33176 (N_33176,N_29204,N_26800);
nand U33177 (N_33177,N_27629,N_29031);
nor U33178 (N_33178,N_29204,N_26918);
nand U33179 (N_33179,N_26784,N_29207);
nor U33180 (N_33180,N_27634,N_28897);
nand U33181 (N_33181,N_27287,N_28883);
xnor U33182 (N_33182,N_29444,N_26511);
xor U33183 (N_33183,N_27630,N_25603);
or U33184 (N_33184,N_25397,N_26689);
and U33185 (N_33185,N_28473,N_26048);
and U33186 (N_33186,N_26070,N_27212);
xnor U33187 (N_33187,N_28866,N_27619);
or U33188 (N_33188,N_28325,N_29308);
nor U33189 (N_33189,N_26877,N_29123);
and U33190 (N_33190,N_28666,N_26850);
xor U33191 (N_33191,N_27727,N_27579);
and U33192 (N_33192,N_27706,N_26541);
nand U33193 (N_33193,N_28369,N_27113);
nand U33194 (N_33194,N_26886,N_26457);
and U33195 (N_33195,N_27744,N_29280);
xor U33196 (N_33196,N_28310,N_25482);
xor U33197 (N_33197,N_25063,N_29602);
nor U33198 (N_33198,N_25570,N_29015);
xor U33199 (N_33199,N_28752,N_25025);
or U33200 (N_33200,N_27978,N_27675);
xor U33201 (N_33201,N_28842,N_25255);
and U33202 (N_33202,N_28971,N_27460);
nor U33203 (N_33203,N_25248,N_26950);
xnor U33204 (N_33204,N_28038,N_28366);
nand U33205 (N_33205,N_29648,N_29960);
nand U33206 (N_33206,N_27665,N_28401);
xor U33207 (N_33207,N_25506,N_28171);
xor U33208 (N_33208,N_29140,N_27019);
nand U33209 (N_33209,N_26457,N_27211);
nor U33210 (N_33210,N_26730,N_28487);
nand U33211 (N_33211,N_26496,N_29795);
nor U33212 (N_33212,N_25967,N_29572);
xor U33213 (N_33213,N_28328,N_28873);
nand U33214 (N_33214,N_29594,N_25280);
nand U33215 (N_33215,N_28740,N_27686);
nand U33216 (N_33216,N_25803,N_26993);
and U33217 (N_33217,N_25445,N_26424);
xor U33218 (N_33218,N_28938,N_27731);
xor U33219 (N_33219,N_27290,N_27120);
or U33220 (N_33220,N_25757,N_25387);
or U33221 (N_33221,N_27430,N_27158);
nor U33222 (N_33222,N_29911,N_28069);
nand U33223 (N_33223,N_27440,N_27845);
or U33224 (N_33224,N_27790,N_27732);
nand U33225 (N_33225,N_27999,N_28340);
xnor U33226 (N_33226,N_27223,N_26333);
nor U33227 (N_33227,N_27728,N_29208);
nor U33228 (N_33228,N_26410,N_28478);
or U33229 (N_33229,N_27719,N_26003);
or U33230 (N_33230,N_25889,N_29075);
xor U33231 (N_33231,N_28519,N_27796);
or U33232 (N_33232,N_28470,N_26317);
or U33233 (N_33233,N_27964,N_29593);
and U33234 (N_33234,N_29231,N_25762);
xnor U33235 (N_33235,N_25483,N_29694);
or U33236 (N_33236,N_29108,N_26000);
nor U33237 (N_33237,N_27783,N_26240);
and U33238 (N_33238,N_29171,N_25571);
nand U33239 (N_33239,N_25275,N_26852);
xnor U33240 (N_33240,N_28155,N_25901);
or U33241 (N_33241,N_26261,N_29672);
xor U33242 (N_33242,N_29511,N_25900);
nand U33243 (N_33243,N_27294,N_29310);
nor U33244 (N_33244,N_29288,N_27913);
nand U33245 (N_33245,N_27660,N_29603);
and U33246 (N_33246,N_29992,N_26301);
or U33247 (N_33247,N_25519,N_28950);
xnor U33248 (N_33248,N_28004,N_29074);
and U33249 (N_33249,N_27225,N_29551);
or U33250 (N_33250,N_28320,N_26132);
nand U33251 (N_33251,N_27070,N_28511);
or U33252 (N_33252,N_26569,N_28806);
nand U33253 (N_33253,N_25243,N_27365);
and U33254 (N_33254,N_27575,N_25332);
or U33255 (N_33255,N_27918,N_27437);
nor U33256 (N_33256,N_26109,N_25971);
xor U33257 (N_33257,N_26869,N_28791);
or U33258 (N_33258,N_29475,N_26010);
nor U33259 (N_33259,N_28512,N_25276);
or U33260 (N_33260,N_25922,N_25378);
nand U33261 (N_33261,N_26938,N_28465);
and U33262 (N_33262,N_25199,N_27868);
nand U33263 (N_33263,N_29213,N_28370);
nand U33264 (N_33264,N_26351,N_28683);
nor U33265 (N_33265,N_29247,N_27498);
xnor U33266 (N_33266,N_26757,N_26333);
nand U33267 (N_33267,N_28331,N_26754);
or U33268 (N_33268,N_25523,N_26286);
nor U33269 (N_33269,N_25265,N_28289);
nand U33270 (N_33270,N_29647,N_26827);
and U33271 (N_33271,N_29480,N_26289);
or U33272 (N_33272,N_27146,N_26849);
nor U33273 (N_33273,N_27226,N_29789);
or U33274 (N_33274,N_29403,N_28735);
xnor U33275 (N_33275,N_29849,N_29427);
xor U33276 (N_33276,N_27855,N_28113);
or U33277 (N_33277,N_26131,N_26435);
nand U33278 (N_33278,N_27708,N_26326);
or U33279 (N_33279,N_28761,N_29294);
or U33280 (N_33280,N_26244,N_26164);
and U33281 (N_33281,N_29434,N_28599);
nor U33282 (N_33282,N_25727,N_27678);
xnor U33283 (N_33283,N_29677,N_29745);
or U33284 (N_33284,N_25310,N_27163);
nand U33285 (N_33285,N_26631,N_27557);
nand U33286 (N_33286,N_27791,N_27944);
and U33287 (N_33287,N_29263,N_25016);
or U33288 (N_33288,N_28138,N_27672);
nor U33289 (N_33289,N_26440,N_29717);
xor U33290 (N_33290,N_29343,N_25773);
and U33291 (N_33291,N_28856,N_25635);
xnor U33292 (N_33292,N_26306,N_29626);
xnor U33293 (N_33293,N_29155,N_27642);
nand U33294 (N_33294,N_28497,N_25023);
xor U33295 (N_33295,N_28311,N_28927);
or U33296 (N_33296,N_25124,N_27879);
nor U33297 (N_33297,N_28952,N_27875);
nand U33298 (N_33298,N_27251,N_25218);
or U33299 (N_33299,N_25007,N_29376);
and U33300 (N_33300,N_28633,N_26905);
and U33301 (N_33301,N_27044,N_28416);
and U33302 (N_33302,N_29105,N_27310);
nor U33303 (N_33303,N_26200,N_29405);
and U33304 (N_33304,N_27303,N_28085);
or U33305 (N_33305,N_29116,N_28029);
xnor U33306 (N_33306,N_26211,N_26583);
xnor U33307 (N_33307,N_29139,N_28683);
and U33308 (N_33308,N_27855,N_28255);
nand U33309 (N_33309,N_29281,N_27872);
nand U33310 (N_33310,N_25136,N_29092);
and U33311 (N_33311,N_27642,N_28382);
or U33312 (N_33312,N_29885,N_29479);
nand U33313 (N_33313,N_27174,N_28311);
nor U33314 (N_33314,N_25857,N_29475);
nand U33315 (N_33315,N_29235,N_26034);
or U33316 (N_33316,N_25991,N_26756);
xor U33317 (N_33317,N_28005,N_29266);
nand U33318 (N_33318,N_27080,N_26242);
or U33319 (N_33319,N_25558,N_25180);
nor U33320 (N_33320,N_26248,N_25910);
nand U33321 (N_33321,N_28769,N_27742);
and U33322 (N_33322,N_25778,N_28102);
nand U33323 (N_33323,N_25585,N_26048);
nand U33324 (N_33324,N_27765,N_29793);
and U33325 (N_33325,N_29225,N_25145);
and U33326 (N_33326,N_27547,N_26190);
and U33327 (N_33327,N_29894,N_27703);
and U33328 (N_33328,N_25420,N_28894);
nand U33329 (N_33329,N_27342,N_26019);
nand U33330 (N_33330,N_28460,N_25948);
nand U33331 (N_33331,N_29131,N_26949);
nor U33332 (N_33332,N_27109,N_28208);
and U33333 (N_33333,N_28061,N_29377);
or U33334 (N_33334,N_27642,N_28069);
and U33335 (N_33335,N_28195,N_27073);
and U33336 (N_33336,N_25045,N_26817);
xnor U33337 (N_33337,N_28404,N_26888);
and U33338 (N_33338,N_25433,N_29864);
and U33339 (N_33339,N_27642,N_25766);
nor U33340 (N_33340,N_29692,N_27033);
and U33341 (N_33341,N_28717,N_29505);
nor U33342 (N_33342,N_27284,N_25635);
and U33343 (N_33343,N_29334,N_28177);
nand U33344 (N_33344,N_28534,N_25785);
xor U33345 (N_33345,N_28120,N_29013);
or U33346 (N_33346,N_29474,N_28769);
nand U33347 (N_33347,N_26070,N_26112);
or U33348 (N_33348,N_29542,N_26433);
and U33349 (N_33349,N_29850,N_29187);
nor U33350 (N_33350,N_26153,N_28600);
and U33351 (N_33351,N_29685,N_26686);
and U33352 (N_33352,N_27980,N_26931);
xnor U33353 (N_33353,N_27091,N_27671);
and U33354 (N_33354,N_25817,N_29648);
nand U33355 (N_33355,N_29803,N_25300);
or U33356 (N_33356,N_29011,N_29333);
nor U33357 (N_33357,N_27794,N_29437);
nand U33358 (N_33358,N_25269,N_27350);
nand U33359 (N_33359,N_29948,N_27267);
or U33360 (N_33360,N_25357,N_28279);
nor U33361 (N_33361,N_29950,N_27696);
or U33362 (N_33362,N_29595,N_28340);
nor U33363 (N_33363,N_28523,N_28894);
and U33364 (N_33364,N_29829,N_29313);
or U33365 (N_33365,N_28933,N_27168);
nand U33366 (N_33366,N_27028,N_28252);
or U33367 (N_33367,N_28370,N_28246);
or U33368 (N_33368,N_28238,N_25352);
nand U33369 (N_33369,N_28916,N_26349);
and U33370 (N_33370,N_26123,N_28307);
or U33371 (N_33371,N_27525,N_27078);
or U33372 (N_33372,N_29352,N_29473);
nand U33373 (N_33373,N_28998,N_25286);
nand U33374 (N_33374,N_29382,N_26514);
or U33375 (N_33375,N_28066,N_25172);
and U33376 (N_33376,N_25212,N_26285);
or U33377 (N_33377,N_29328,N_29788);
or U33378 (N_33378,N_26105,N_27855);
nor U33379 (N_33379,N_27535,N_27946);
xor U33380 (N_33380,N_27773,N_26042);
nand U33381 (N_33381,N_27346,N_27369);
nand U33382 (N_33382,N_26613,N_27505);
nor U33383 (N_33383,N_26390,N_28968);
xnor U33384 (N_33384,N_27120,N_29067);
xor U33385 (N_33385,N_25754,N_27804);
xnor U33386 (N_33386,N_27292,N_27471);
nor U33387 (N_33387,N_26774,N_28411);
nand U33388 (N_33388,N_28310,N_26645);
xor U33389 (N_33389,N_27519,N_26879);
nor U33390 (N_33390,N_26624,N_28764);
and U33391 (N_33391,N_27445,N_26767);
nor U33392 (N_33392,N_28608,N_25818);
nor U33393 (N_33393,N_26760,N_25600);
nor U33394 (N_33394,N_28233,N_26141);
nand U33395 (N_33395,N_27902,N_29678);
nor U33396 (N_33396,N_25985,N_29712);
and U33397 (N_33397,N_26731,N_25285);
nor U33398 (N_33398,N_26507,N_26371);
or U33399 (N_33399,N_25613,N_29654);
nor U33400 (N_33400,N_28339,N_27259);
or U33401 (N_33401,N_27185,N_26775);
nand U33402 (N_33402,N_27059,N_28757);
and U33403 (N_33403,N_29741,N_28199);
or U33404 (N_33404,N_26314,N_26188);
nand U33405 (N_33405,N_25565,N_27676);
and U33406 (N_33406,N_29065,N_29076);
and U33407 (N_33407,N_29017,N_29131);
xor U33408 (N_33408,N_26693,N_28649);
xnor U33409 (N_33409,N_25325,N_25764);
and U33410 (N_33410,N_29825,N_27593);
xnor U33411 (N_33411,N_26783,N_26811);
and U33412 (N_33412,N_27224,N_28420);
nor U33413 (N_33413,N_25636,N_29554);
nand U33414 (N_33414,N_26954,N_26415);
and U33415 (N_33415,N_27135,N_28215);
and U33416 (N_33416,N_27324,N_29698);
or U33417 (N_33417,N_29973,N_29603);
xnor U33418 (N_33418,N_27668,N_26269);
nor U33419 (N_33419,N_27224,N_29883);
xnor U33420 (N_33420,N_26339,N_25445);
xnor U33421 (N_33421,N_27393,N_26312);
nor U33422 (N_33422,N_29187,N_25028);
and U33423 (N_33423,N_27884,N_28658);
nand U33424 (N_33424,N_28672,N_26479);
xnor U33425 (N_33425,N_27030,N_26072);
nand U33426 (N_33426,N_28837,N_25992);
nand U33427 (N_33427,N_27247,N_26619);
and U33428 (N_33428,N_26167,N_25381);
nor U33429 (N_33429,N_29526,N_26688);
xnor U33430 (N_33430,N_26433,N_28876);
nor U33431 (N_33431,N_25652,N_27373);
xor U33432 (N_33432,N_28366,N_25036);
xor U33433 (N_33433,N_29523,N_28860);
nand U33434 (N_33434,N_28274,N_26323);
or U33435 (N_33435,N_28241,N_26474);
or U33436 (N_33436,N_29358,N_29293);
and U33437 (N_33437,N_29082,N_27232);
nand U33438 (N_33438,N_27391,N_29768);
nand U33439 (N_33439,N_29307,N_29225);
nor U33440 (N_33440,N_25087,N_27984);
or U33441 (N_33441,N_27799,N_25365);
nand U33442 (N_33442,N_25205,N_25936);
nor U33443 (N_33443,N_25170,N_25946);
nor U33444 (N_33444,N_28786,N_28864);
nand U33445 (N_33445,N_29914,N_29354);
xor U33446 (N_33446,N_26899,N_25978);
and U33447 (N_33447,N_25205,N_28843);
nand U33448 (N_33448,N_29635,N_27528);
xnor U33449 (N_33449,N_26661,N_27596);
xnor U33450 (N_33450,N_26320,N_25982);
and U33451 (N_33451,N_28827,N_29345);
nand U33452 (N_33452,N_27557,N_26170);
xor U33453 (N_33453,N_28704,N_25686);
nand U33454 (N_33454,N_26106,N_28791);
nor U33455 (N_33455,N_26114,N_25658);
and U33456 (N_33456,N_25771,N_26602);
or U33457 (N_33457,N_26381,N_26632);
or U33458 (N_33458,N_28479,N_29866);
and U33459 (N_33459,N_27300,N_26748);
nand U33460 (N_33460,N_28538,N_27594);
nand U33461 (N_33461,N_28528,N_28922);
or U33462 (N_33462,N_27790,N_28512);
or U33463 (N_33463,N_26690,N_29838);
nand U33464 (N_33464,N_28778,N_29858);
nor U33465 (N_33465,N_27415,N_26469);
xor U33466 (N_33466,N_29137,N_27851);
nand U33467 (N_33467,N_29611,N_28164);
and U33468 (N_33468,N_29632,N_29096);
and U33469 (N_33469,N_26801,N_25480);
and U33470 (N_33470,N_26079,N_28085);
or U33471 (N_33471,N_25787,N_28076);
xnor U33472 (N_33472,N_25811,N_27681);
nand U33473 (N_33473,N_28602,N_29540);
and U33474 (N_33474,N_26772,N_29496);
nand U33475 (N_33475,N_27338,N_28832);
nand U33476 (N_33476,N_28679,N_29654);
nand U33477 (N_33477,N_25543,N_27536);
nand U33478 (N_33478,N_25717,N_27431);
xor U33479 (N_33479,N_26478,N_28733);
or U33480 (N_33480,N_27859,N_26420);
nor U33481 (N_33481,N_27124,N_29315);
or U33482 (N_33482,N_28772,N_28839);
nor U33483 (N_33483,N_26439,N_29855);
nand U33484 (N_33484,N_27288,N_25106);
nand U33485 (N_33485,N_27619,N_25490);
nand U33486 (N_33486,N_25215,N_27435);
nand U33487 (N_33487,N_28133,N_25559);
xor U33488 (N_33488,N_25020,N_28200);
or U33489 (N_33489,N_29412,N_28984);
xor U33490 (N_33490,N_25510,N_25646);
nand U33491 (N_33491,N_26757,N_26820);
nand U33492 (N_33492,N_26779,N_26609);
or U33493 (N_33493,N_26022,N_29948);
nand U33494 (N_33494,N_29929,N_25520);
nand U33495 (N_33495,N_28649,N_26071);
or U33496 (N_33496,N_26764,N_29382);
nor U33497 (N_33497,N_27591,N_26119);
or U33498 (N_33498,N_25242,N_29463);
or U33499 (N_33499,N_27718,N_25756);
nand U33500 (N_33500,N_28055,N_25237);
xor U33501 (N_33501,N_26898,N_27270);
nand U33502 (N_33502,N_29923,N_26838);
xnor U33503 (N_33503,N_29925,N_29015);
xor U33504 (N_33504,N_25437,N_25749);
nor U33505 (N_33505,N_27215,N_28876);
nor U33506 (N_33506,N_29191,N_26126);
and U33507 (N_33507,N_26045,N_26430);
nor U33508 (N_33508,N_25480,N_28273);
or U33509 (N_33509,N_25882,N_27003);
xnor U33510 (N_33510,N_29379,N_29725);
or U33511 (N_33511,N_25147,N_25008);
nor U33512 (N_33512,N_28793,N_28110);
or U33513 (N_33513,N_27286,N_26943);
nor U33514 (N_33514,N_27488,N_25350);
nor U33515 (N_33515,N_25012,N_27182);
or U33516 (N_33516,N_27927,N_27313);
nor U33517 (N_33517,N_26408,N_29863);
or U33518 (N_33518,N_26739,N_29322);
nand U33519 (N_33519,N_27563,N_28205);
or U33520 (N_33520,N_29207,N_27533);
xnor U33521 (N_33521,N_29314,N_26963);
xor U33522 (N_33522,N_26713,N_26732);
nand U33523 (N_33523,N_25477,N_28091);
and U33524 (N_33524,N_27231,N_29431);
xor U33525 (N_33525,N_28846,N_26485);
and U33526 (N_33526,N_27866,N_26030);
xnor U33527 (N_33527,N_28138,N_28817);
and U33528 (N_33528,N_25670,N_26694);
nor U33529 (N_33529,N_27093,N_29100);
nor U33530 (N_33530,N_26157,N_27654);
nor U33531 (N_33531,N_29825,N_27401);
xnor U33532 (N_33532,N_25824,N_29398);
nand U33533 (N_33533,N_28617,N_29301);
and U33534 (N_33534,N_29075,N_26226);
nor U33535 (N_33535,N_27928,N_27937);
and U33536 (N_33536,N_26303,N_27691);
xnor U33537 (N_33537,N_28444,N_25717);
or U33538 (N_33538,N_28659,N_27210);
xor U33539 (N_33539,N_27790,N_26780);
nor U33540 (N_33540,N_25187,N_28859);
or U33541 (N_33541,N_28096,N_28696);
and U33542 (N_33542,N_28322,N_29177);
nand U33543 (N_33543,N_27868,N_29248);
or U33544 (N_33544,N_28446,N_26486);
and U33545 (N_33545,N_28135,N_25193);
and U33546 (N_33546,N_25446,N_28011);
and U33547 (N_33547,N_25388,N_28757);
nand U33548 (N_33548,N_25690,N_29140);
nor U33549 (N_33549,N_28127,N_26271);
nand U33550 (N_33550,N_25992,N_26823);
or U33551 (N_33551,N_27033,N_29663);
or U33552 (N_33552,N_28978,N_28243);
xnor U33553 (N_33553,N_27159,N_29446);
nand U33554 (N_33554,N_26286,N_29251);
nor U33555 (N_33555,N_28103,N_26356);
nor U33556 (N_33556,N_29988,N_26859);
nand U33557 (N_33557,N_29197,N_29369);
xor U33558 (N_33558,N_26942,N_25879);
or U33559 (N_33559,N_27205,N_27042);
xor U33560 (N_33560,N_26101,N_28968);
nor U33561 (N_33561,N_29004,N_29990);
nor U33562 (N_33562,N_27239,N_29690);
xor U33563 (N_33563,N_27656,N_29203);
nor U33564 (N_33564,N_28674,N_27056);
nor U33565 (N_33565,N_26475,N_25865);
nand U33566 (N_33566,N_29414,N_25004);
nor U33567 (N_33567,N_28402,N_27108);
xor U33568 (N_33568,N_28490,N_29030);
xnor U33569 (N_33569,N_25190,N_28149);
xnor U33570 (N_33570,N_29843,N_28646);
nor U33571 (N_33571,N_29525,N_28903);
or U33572 (N_33572,N_25783,N_26979);
nor U33573 (N_33573,N_28407,N_27601);
or U33574 (N_33574,N_28207,N_26956);
xnor U33575 (N_33575,N_28798,N_27881);
and U33576 (N_33576,N_29628,N_28936);
nand U33577 (N_33577,N_27033,N_25867);
or U33578 (N_33578,N_29211,N_27711);
nor U33579 (N_33579,N_25362,N_27391);
nor U33580 (N_33580,N_28919,N_25490);
and U33581 (N_33581,N_26153,N_28077);
nor U33582 (N_33582,N_25371,N_25522);
or U33583 (N_33583,N_27847,N_25081);
xnor U33584 (N_33584,N_26362,N_28308);
xor U33585 (N_33585,N_25286,N_28922);
and U33586 (N_33586,N_26580,N_27316);
and U33587 (N_33587,N_28156,N_25537);
nor U33588 (N_33588,N_28620,N_25645);
xnor U33589 (N_33589,N_25026,N_26876);
or U33590 (N_33590,N_26636,N_28484);
or U33591 (N_33591,N_29513,N_29314);
nand U33592 (N_33592,N_28197,N_25122);
and U33593 (N_33593,N_26887,N_28792);
and U33594 (N_33594,N_26799,N_28002);
or U33595 (N_33595,N_28723,N_29795);
or U33596 (N_33596,N_28579,N_25757);
xnor U33597 (N_33597,N_29793,N_26510);
or U33598 (N_33598,N_29746,N_27988);
xor U33599 (N_33599,N_25201,N_25320);
or U33600 (N_33600,N_26271,N_26176);
nor U33601 (N_33601,N_29032,N_27781);
nand U33602 (N_33602,N_25129,N_29594);
nand U33603 (N_33603,N_29291,N_28609);
or U33604 (N_33604,N_26219,N_26062);
nor U33605 (N_33605,N_25112,N_26456);
xor U33606 (N_33606,N_26839,N_29274);
xnor U33607 (N_33607,N_26103,N_25193);
xor U33608 (N_33608,N_28190,N_28553);
nand U33609 (N_33609,N_25372,N_25990);
xnor U33610 (N_33610,N_28830,N_25067);
and U33611 (N_33611,N_29139,N_28479);
xor U33612 (N_33612,N_29095,N_28270);
nand U33613 (N_33613,N_27383,N_29893);
nand U33614 (N_33614,N_29941,N_29316);
and U33615 (N_33615,N_29820,N_25227);
nor U33616 (N_33616,N_29025,N_26620);
and U33617 (N_33617,N_26561,N_26765);
nor U33618 (N_33618,N_27870,N_28582);
and U33619 (N_33619,N_27563,N_29231);
nor U33620 (N_33620,N_26181,N_27561);
and U33621 (N_33621,N_27266,N_29141);
or U33622 (N_33622,N_27645,N_26380);
and U33623 (N_33623,N_27907,N_28707);
or U33624 (N_33624,N_29077,N_29852);
nor U33625 (N_33625,N_27199,N_28853);
nand U33626 (N_33626,N_26924,N_27999);
or U33627 (N_33627,N_27696,N_26230);
nand U33628 (N_33628,N_27026,N_26816);
nor U33629 (N_33629,N_27493,N_28289);
or U33630 (N_33630,N_28302,N_27447);
and U33631 (N_33631,N_29059,N_27233);
xnor U33632 (N_33632,N_26344,N_25447);
nor U33633 (N_33633,N_26227,N_26271);
or U33634 (N_33634,N_26708,N_28696);
or U33635 (N_33635,N_26041,N_28647);
and U33636 (N_33636,N_29114,N_25506);
and U33637 (N_33637,N_26945,N_28571);
and U33638 (N_33638,N_28387,N_25195);
or U33639 (N_33639,N_28870,N_26854);
nor U33640 (N_33640,N_28305,N_28670);
and U33641 (N_33641,N_26649,N_27971);
or U33642 (N_33642,N_25188,N_26783);
nor U33643 (N_33643,N_29754,N_26755);
or U33644 (N_33644,N_26627,N_28086);
and U33645 (N_33645,N_28505,N_26579);
nor U33646 (N_33646,N_25606,N_26036);
and U33647 (N_33647,N_27955,N_27721);
nand U33648 (N_33648,N_27380,N_27024);
nor U33649 (N_33649,N_25556,N_29014);
and U33650 (N_33650,N_29797,N_28505);
xor U33651 (N_33651,N_25562,N_28763);
or U33652 (N_33652,N_28174,N_27437);
or U33653 (N_33653,N_27990,N_28418);
nor U33654 (N_33654,N_29325,N_27720);
xor U33655 (N_33655,N_25983,N_25409);
xor U33656 (N_33656,N_27721,N_25399);
nor U33657 (N_33657,N_27926,N_26786);
or U33658 (N_33658,N_28708,N_29755);
and U33659 (N_33659,N_29735,N_27298);
and U33660 (N_33660,N_27875,N_29911);
and U33661 (N_33661,N_26060,N_27050);
or U33662 (N_33662,N_29264,N_25813);
nor U33663 (N_33663,N_25300,N_29265);
nor U33664 (N_33664,N_26654,N_28469);
and U33665 (N_33665,N_27417,N_28685);
xnor U33666 (N_33666,N_25233,N_27854);
xor U33667 (N_33667,N_29510,N_26779);
and U33668 (N_33668,N_29033,N_28187);
or U33669 (N_33669,N_26551,N_28863);
nor U33670 (N_33670,N_29784,N_25126);
nand U33671 (N_33671,N_27094,N_28916);
or U33672 (N_33672,N_28484,N_25169);
nor U33673 (N_33673,N_29859,N_27155);
nor U33674 (N_33674,N_27969,N_29327);
xor U33675 (N_33675,N_29990,N_27139);
xor U33676 (N_33676,N_27084,N_28938);
nand U33677 (N_33677,N_25538,N_25783);
xnor U33678 (N_33678,N_29180,N_26616);
nor U33679 (N_33679,N_26402,N_28376);
nand U33680 (N_33680,N_26364,N_26327);
and U33681 (N_33681,N_26973,N_29790);
and U33682 (N_33682,N_29295,N_27009);
nand U33683 (N_33683,N_28760,N_28466);
xor U33684 (N_33684,N_28340,N_27681);
or U33685 (N_33685,N_27589,N_26810);
or U33686 (N_33686,N_26320,N_27534);
or U33687 (N_33687,N_28609,N_27185);
nand U33688 (N_33688,N_25149,N_26424);
nand U33689 (N_33689,N_25655,N_29452);
nand U33690 (N_33690,N_25435,N_27995);
xor U33691 (N_33691,N_25458,N_29815);
nand U33692 (N_33692,N_28326,N_25360);
and U33693 (N_33693,N_27167,N_26398);
xor U33694 (N_33694,N_27074,N_27759);
and U33695 (N_33695,N_27241,N_29206);
and U33696 (N_33696,N_28389,N_25345);
or U33697 (N_33697,N_29334,N_25620);
xnor U33698 (N_33698,N_25034,N_28804);
xnor U33699 (N_33699,N_25756,N_28141);
and U33700 (N_33700,N_26216,N_27725);
nor U33701 (N_33701,N_28307,N_26248);
xnor U33702 (N_33702,N_28545,N_27972);
nand U33703 (N_33703,N_27289,N_27950);
nor U33704 (N_33704,N_26473,N_26108);
or U33705 (N_33705,N_27337,N_28100);
and U33706 (N_33706,N_26640,N_25035);
nand U33707 (N_33707,N_28012,N_28240);
and U33708 (N_33708,N_26821,N_27395);
xor U33709 (N_33709,N_27760,N_25415);
nor U33710 (N_33710,N_29047,N_27691);
or U33711 (N_33711,N_25775,N_25789);
or U33712 (N_33712,N_25938,N_26715);
and U33713 (N_33713,N_25568,N_26204);
nor U33714 (N_33714,N_25958,N_28487);
or U33715 (N_33715,N_27925,N_27130);
xor U33716 (N_33716,N_27299,N_29860);
nor U33717 (N_33717,N_26293,N_25868);
or U33718 (N_33718,N_25439,N_25609);
and U33719 (N_33719,N_29061,N_25819);
and U33720 (N_33720,N_28542,N_25725);
xor U33721 (N_33721,N_26733,N_29667);
nor U33722 (N_33722,N_25814,N_26948);
and U33723 (N_33723,N_29728,N_27758);
or U33724 (N_33724,N_25662,N_28610);
nand U33725 (N_33725,N_26180,N_29504);
or U33726 (N_33726,N_26230,N_29679);
nand U33727 (N_33727,N_27588,N_29753);
nand U33728 (N_33728,N_29038,N_29666);
nand U33729 (N_33729,N_26685,N_25925);
xor U33730 (N_33730,N_27320,N_26998);
and U33731 (N_33731,N_28150,N_28814);
xnor U33732 (N_33732,N_25115,N_25288);
or U33733 (N_33733,N_26124,N_26372);
and U33734 (N_33734,N_27818,N_28744);
or U33735 (N_33735,N_25539,N_27445);
nand U33736 (N_33736,N_29572,N_29443);
nand U33737 (N_33737,N_28166,N_28533);
xor U33738 (N_33738,N_29028,N_28675);
nor U33739 (N_33739,N_28557,N_28812);
or U33740 (N_33740,N_25562,N_27547);
and U33741 (N_33741,N_26591,N_25219);
nand U33742 (N_33742,N_27548,N_29271);
nor U33743 (N_33743,N_25355,N_29274);
nand U33744 (N_33744,N_28754,N_26182);
nor U33745 (N_33745,N_28361,N_25292);
nor U33746 (N_33746,N_27610,N_27895);
nand U33747 (N_33747,N_28665,N_26856);
and U33748 (N_33748,N_28376,N_29246);
nand U33749 (N_33749,N_28828,N_28442);
or U33750 (N_33750,N_27696,N_27078);
and U33751 (N_33751,N_26939,N_26793);
nand U33752 (N_33752,N_28820,N_26393);
xor U33753 (N_33753,N_28629,N_26428);
or U33754 (N_33754,N_28388,N_27208);
and U33755 (N_33755,N_25926,N_26578);
xor U33756 (N_33756,N_27156,N_29921);
or U33757 (N_33757,N_25160,N_26667);
nor U33758 (N_33758,N_27115,N_25055);
xor U33759 (N_33759,N_27811,N_25895);
or U33760 (N_33760,N_29871,N_27857);
nand U33761 (N_33761,N_25900,N_27969);
and U33762 (N_33762,N_25450,N_29666);
xor U33763 (N_33763,N_28165,N_26919);
nand U33764 (N_33764,N_28393,N_28329);
nor U33765 (N_33765,N_26525,N_25279);
or U33766 (N_33766,N_27635,N_27581);
or U33767 (N_33767,N_29402,N_29111);
xor U33768 (N_33768,N_28052,N_29883);
nand U33769 (N_33769,N_27078,N_29903);
xnor U33770 (N_33770,N_26382,N_29926);
and U33771 (N_33771,N_26313,N_29377);
and U33772 (N_33772,N_29066,N_28205);
nand U33773 (N_33773,N_29621,N_26402);
and U33774 (N_33774,N_27580,N_26895);
xnor U33775 (N_33775,N_29811,N_25666);
xor U33776 (N_33776,N_28457,N_28276);
xor U33777 (N_33777,N_25019,N_27196);
xor U33778 (N_33778,N_26919,N_25698);
or U33779 (N_33779,N_29181,N_25954);
nand U33780 (N_33780,N_25430,N_26353);
nor U33781 (N_33781,N_25180,N_27350);
xor U33782 (N_33782,N_25058,N_26524);
nor U33783 (N_33783,N_27343,N_26424);
xor U33784 (N_33784,N_26998,N_25897);
nand U33785 (N_33785,N_27827,N_25108);
xor U33786 (N_33786,N_25895,N_29236);
nand U33787 (N_33787,N_29744,N_26744);
and U33788 (N_33788,N_26335,N_28902);
xnor U33789 (N_33789,N_27458,N_25058);
nor U33790 (N_33790,N_29212,N_25654);
xor U33791 (N_33791,N_26999,N_26320);
xor U33792 (N_33792,N_25270,N_28760);
or U33793 (N_33793,N_27274,N_26974);
nor U33794 (N_33794,N_27659,N_29035);
nand U33795 (N_33795,N_26398,N_27541);
or U33796 (N_33796,N_26083,N_28774);
nand U33797 (N_33797,N_26998,N_27347);
and U33798 (N_33798,N_27342,N_27305);
nand U33799 (N_33799,N_27802,N_25249);
nand U33800 (N_33800,N_26351,N_29058);
or U33801 (N_33801,N_28718,N_28348);
xnor U33802 (N_33802,N_29916,N_25389);
or U33803 (N_33803,N_26172,N_26243);
nor U33804 (N_33804,N_25494,N_26641);
xor U33805 (N_33805,N_25097,N_27423);
nor U33806 (N_33806,N_26012,N_26455);
and U33807 (N_33807,N_29382,N_26469);
nand U33808 (N_33808,N_29909,N_27558);
xnor U33809 (N_33809,N_28528,N_25337);
nor U33810 (N_33810,N_27229,N_29702);
and U33811 (N_33811,N_26707,N_29834);
and U33812 (N_33812,N_28346,N_29911);
nand U33813 (N_33813,N_25160,N_28024);
or U33814 (N_33814,N_29823,N_25569);
and U33815 (N_33815,N_27887,N_25977);
xnor U33816 (N_33816,N_26418,N_28605);
nor U33817 (N_33817,N_27664,N_29835);
nor U33818 (N_33818,N_29422,N_26988);
nor U33819 (N_33819,N_28083,N_27319);
nand U33820 (N_33820,N_27048,N_28212);
and U33821 (N_33821,N_27541,N_28208);
and U33822 (N_33822,N_25548,N_29000);
nand U33823 (N_33823,N_28899,N_26089);
and U33824 (N_33824,N_29579,N_29175);
nor U33825 (N_33825,N_28424,N_28837);
or U33826 (N_33826,N_28796,N_25999);
xnor U33827 (N_33827,N_29050,N_28409);
nand U33828 (N_33828,N_27517,N_25950);
nor U33829 (N_33829,N_28962,N_27781);
nand U33830 (N_33830,N_29197,N_29038);
xor U33831 (N_33831,N_27639,N_29279);
and U33832 (N_33832,N_26098,N_26197);
and U33833 (N_33833,N_26126,N_26251);
nor U33834 (N_33834,N_29552,N_28142);
nor U33835 (N_33835,N_27813,N_29001);
nand U33836 (N_33836,N_29177,N_27643);
and U33837 (N_33837,N_26504,N_26286);
and U33838 (N_33838,N_25421,N_27327);
xor U33839 (N_33839,N_26377,N_27972);
or U33840 (N_33840,N_28214,N_25733);
and U33841 (N_33841,N_26085,N_27416);
nand U33842 (N_33842,N_26054,N_25131);
xnor U33843 (N_33843,N_28798,N_28521);
xnor U33844 (N_33844,N_29662,N_28003);
and U33845 (N_33845,N_26726,N_25362);
nand U33846 (N_33846,N_27052,N_29740);
nand U33847 (N_33847,N_28211,N_27654);
xor U33848 (N_33848,N_25019,N_25420);
nor U33849 (N_33849,N_25051,N_29656);
nor U33850 (N_33850,N_28922,N_29972);
and U33851 (N_33851,N_29589,N_29074);
nand U33852 (N_33852,N_25035,N_26997);
or U33853 (N_33853,N_26842,N_27395);
or U33854 (N_33854,N_25760,N_26215);
xor U33855 (N_33855,N_25780,N_29893);
nand U33856 (N_33856,N_27033,N_29094);
or U33857 (N_33857,N_25085,N_29174);
or U33858 (N_33858,N_25913,N_29860);
and U33859 (N_33859,N_25561,N_25372);
or U33860 (N_33860,N_26128,N_26330);
nor U33861 (N_33861,N_26837,N_26274);
nand U33862 (N_33862,N_29619,N_26598);
xor U33863 (N_33863,N_29766,N_29997);
xor U33864 (N_33864,N_27273,N_25526);
nand U33865 (N_33865,N_25892,N_29843);
nor U33866 (N_33866,N_29134,N_28627);
nand U33867 (N_33867,N_29335,N_29110);
xor U33868 (N_33868,N_28709,N_25404);
or U33869 (N_33869,N_26543,N_27551);
nor U33870 (N_33870,N_27635,N_25709);
nand U33871 (N_33871,N_27938,N_25417);
or U33872 (N_33872,N_29718,N_28555);
nand U33873 (N_33873,N_28621,N_27426);
nor U33874 (N_33874,N_29753,N_29669);
nor U33875 (N_33875,N_26784,N_25887);
and U33876 (N_33876,N_28053,N_25225);
nand U33877 (N_33877,N_27833,N_26558);
xor U33878 (N_33878,N_29082,N_27863);
nand U33879 (N_33879,N_28227,N_27677);
nand U33880 (N_33880,N_25316,N_25538);
and U33881 (N_33881,N_27293,N_29467);
nor U33882 (N_33882,N_28824,N_26936);
nor U33883 (N_33883,N_27969,N_27904);
xnor U33884 (N_33884,N_26666,N_27380);
and U33885 (N_33885,N_25387,N_27050);
nor U33886 (N_33886,N_26916,N_27935);
nand U33887 (N_33887,N_25099,N_28746);
nand U33888 (N_33888,N_25895,N_26502);
xor U33889 (N_33889,N_29363,N_26573);
nor U33890 (N_33890,N_25036,N_28886);
nor U33891 (N_33891,N_27518,N_29291);
nand U33892 (N_33892,N_28602,N_26384);
nor U33893 (N_33893,N_28473,N_26867);
nor U33894 (N_33894,N_29776,N_25700);
nand U33895 (N_33895,N_26372,N_25121);
nand U33896 (N_33896,N_27298,N_26635);
xor U33897 (N_33897,N_29468,N_28536);
or U33898 (N_33898,N_25006,N_29356);
and U33899 (N_33899,N_26650,N_27708);
nor U33900 (N_33900,N_29485,N_25194);
nand U33901 (N_33901,N_29040,N_26739);
or U33902 (N_33902,N_25755,N_25774);
xnor U33903 (N_33903,N_26433,N_27294);
nor U33904 (N_33904,N_26316,N_26859);
xnor U33905 (N_33905,N_26045,N_27709);
xor U33906 (N_33906,N_25459,N_26358);
nor U33907 (N_33907,N_26822,N_25091);
xor U33908 (N_33908,N_25601,N_25958);
or U33909 (N_33909,N_25165,N_28884);
nor U33910 (N_33910,N_25583,N_26269);
and U33911 (N_33911,N_26027,N_29185);
xor U33912 (N_33912,N_28093,N_26077);
nand U33913 (N_33913,N_28227,N_26398);
nand U33914 (N_33914,N_25142,N_27788);
or U33915 (N_33915,N_25773,N_27633);
and U33916 (N_33916,N_28964,N_29758);
and U33917 (N_33917,N_29752,N_26272);
nor U33918 (N_33918,N_28661,N_27780);
nor U33919 (N_33919,N_29065,N_27581);
nor U33920 (N_33920,N_27811,N_29380);
nor U33921 (N_33921,N_29396,N_25878);
nor U33922 (N_33922,N_25569,N_26740);
nor U33923 (N_33923,N_26111,N_25785);
nor U33924 (N_33924,N_25707,N_28469);
or U33925 (N_33925,N_27168,N_26910);
nand U33926 (N_33926,N_28821,N_25506);
or U33927 (N_33927,N_29436,N_29676);
or U33928 (N_33928,N_28708,N_25467);
nor U33929 (N_33929,N_28508,N_25705);
and U33930 (N_33930,N_28353,N_27806);
nand U33931 (N_33931,N_26734,N_29762);
nor U33932 (N_33932,N_25371,N_26014);
and U33933 (N_33933,N_29257,N_29573);
and U33934 (N_33934,N_25516,N_25729);
nand U33935 (N_33935,N_28115,N_29923);
or U33936 (N_33936,N_27298,N_26739);
nor U33937 (N_33937,N_25179,N_25547);
and U33938 (N_33938,N_29965,N_28387);
nand U33939 (N_33939,N_25277,N_26684);
xor U33940 (N_33940,N_29230,N_25520);
and U33941 (N_33941,N_26924,N_28384);
and U33942 (N_33942,N_25588,N_28846);
xor U33943 (N_33943,N_28702,N_29977);
or U33944 (N_33944,N_27213,N_27850);
or U33945 (N_33945,N_26436,N_25705);
or U33946 (N_33946,N_27449,N_26624);
and U33947 (N_33947,N_27021,N_26584);
and U33948 (N_33948,N_29209,N_26192);
xnor U33949 (N_33949,N_29552,N_28857);
xnor U33950 (N_33950,N_27056,N_25566);
and U33951 (N_33951,N_28739,N_29114);
or U33952 (N_33952,N_29196,N_25364);
and U33953 (N_33953,N_27920,N_25856);
or U33954 (N_33954,N_29285,N_25093);
nor U33955 (N_33955,N_28528,N_25404);
and U33956 (N_33956,N_27343,N_27827);
or U33957 (N_33957,N_26580,N_25325);
nand U33958 (N_33958,N_28816,N_28148);
nor U33959 (N_33959,N_26936,N_25176);
and U33960 (N_33960,N_26878,N_27187);
or U33961 (N_33961,N_26033,N_28771);
xor U33962 (N_33962,N_26738,N_29188);
or U33963 (N_33963,N_27969,N_28847);
or U33964 (N_33964,N_27132,N_25032);
and U33965 (N_33965,N_29030,N_29764);
nand U33966 (N_33966,N_29923,N_29221);
nand U33967 (N_33967,N_25860,N_27433);
xor U33968 (N_33968,N_26496,N_28352);
nor U33969 (N_33969,N_29161,N_27811);
and U33970 (N_33970,N_25463,N_25093);
or U33971 (N_33971,N_25005,N_29045);
nor U33972 (N_33972,N_25951,N_25526);
nand U33973 (N_33973,N_25204,N_27051);
and U33974 (N_33974,N_28444,N_25770);
xor U33975 (N_33975,N_27433,N_29573);
nand U33976 (N_33976,N_28811,N_25303);
or U33977 (N_33977,N_29277,N_25256);
or U33978 (N_33978,N_26343,N_29775);
nand U33979 (N_33979,N_28720,N_27390);
and U33980 (N_33980,N_29885,N_28540);
and U33981 (N_33981,N_26213,N_25609);
or U33982 (N_33982,N_25404,N_28397);
xor U33983 (N_33983,N_26801,N_26697);
or U33984 (N_33984,N_25636,N_25100);
and U33985 (N_33985,N_25272,N_29575);
or U33986 (N_33986,N_27197,N_29102);
xnor U33987 (N_33987,N_27124,N_25524);
nor U33988 (N_33988,N_25647,N_26567);
nand U33989 (N_33989,N_26024,N_26551);
or U33990 (N_33990,N_26400,N_29450);
nand U33991 (N_33991,N_25105,N_27130);
xor U33992 (N_33992,N_28112,N_29709);
xor U33993 (N_33993,N_27533,N_28544);
xnor U33994 (N_33994,N_26521,N_25616);
or U33995 (N_33995,N_28057,N_29501);
or U33996 (N_33996,N_25531,N_25843);
nand U33997 (N_33997,N_28685,N_27577);
xnor U33998 (N_33998,N_29339,N_29220);
or U33999 (N_33999,N_25806,N_28344);
nand U34000 (N_34000,N_28845,N_26609);
or U34001 (N_34001,N_28291,N_25427);
nand U34002 (N_34002,N_29235,N_29939);
and U34003 (N_34003,N_25148,N_27719);
or U34004 (N_34004,N_26109,N_29621);
xnor U34005 (N_34005,N_27285,N_27392);
and U34006 (N_34006,N_27327,N_27367);
and U34007 (N_34007,N_29242,N_26414);
and U34008 (N_34008,N_29049,N_28164);
nor U34009 (N_34009,N_26605,N_26602);
and U34010 (N_34010,N_26389,N_28554);
xnor U34011 (N_34011,N_25246,N_28221);
nand U34012 (N_34012,N_27821,N_26470);
nand U34013 (N_34013,N_26112,N_25281);
or U34014 (N_34014,N_25115,N_28932);
nand U34015 (N_34015,N_29425,N_27108);
nand U34016 (N_34016,N_25299,N_29330);
and U34017 (N_34017,N_29966,N_29395);
or U34018 (N_34018,N_27893,N_28870);
nor U34019 (N_34019,N_29365,N_28630);
or U34020 (N_34020,N_25367,N_29601);
and U34021 (N_34021,N_27677,N_26393);
and U34022 (N_34022,N_27687,N_28026);
nand U34023 (N_34023,N_27090,N_25469);
xor U34024 (N_34024,N_27071,N_27480);
nor U34025 (N_34025,N_28251,N_27709);
xor U34026 (N_34026,N_27087,N_28466);
and U34027 (N_34027,N_28874,N_27856);
or U34028 (N_34028,N_27111,N_26546);
xor U34029 (N_34029,N_25354,N_28502);
nor U34030 (N_34030,N_27018,N_25734);
and U34031 (N_34031,N_29172,N_28011);
nor U34032 (N_34032,N_29661,N_27231);
xor U34033 (N_34033,N_27226,N_28374);
nor U34034 (N_34034,N_29167,N_26876);
and U34035 (N_34035,N_27227,N_26277);
nand U34036 (N_34036,N_26353,N_27475);
xnor U34037 (N_34037,N_27456,N_28520);
xnor U34038 (N_34038,N_28634,N_28534);
xnor U34039 (N_34039,N_26308,N_29068);
nor U34040 (N_34040,N_26502,N_29869);
and U34041 (N_34041,N_28963,N_28862);
xnor U34042 (N_34042,N_27743,N_26157);
or U34043 (N_34043,N_25254,N_25528);
or U34044 (N_34044,N_27720,N_29857);
nor U34045 (N_34045,N_26085,N_29102);
xor U34046 (N_34046,N_28102,N_26611);
or U34047 (N_34047,N_28882,N_29146);
and U34048 (N_34048,N_25428,N_26730);
or U34049 (N_34049,N_25094,N_26696);
and U34050 (N_34050,N_28580,N_29016);
nor U34051 (N_34051,N_26494,N_25779);
nand U34052 (N_34052,N_28789,N_25609);
nor U34053 (N_34053,N_29616,N_25752);
nand U34054 (N_34054,N_28997,N_25616);
xor U34055 (N_34055,N_27849,N_29135);
nand U34056 (N_34056,N_29132,N_26271);
and U34057 (N_34057,N_25219,N_25982);
nor U34058 (N_34058,N_27143,N_28299);
nand U34059 (N_34059,N_25604,N_26897);
or U34060 (N_34060,N_27927,N_26011);
and U34061 (N_34061,N_29804,N_25000);
nor U34062 (N_34062,N_26820,N_29735);
nand U34063 (N_34063,N_29218,N_25246);
nor U34064 (N_34064,N_29198,N_28072);
and U34065 (N_34065,N_25359,N_29798);
or U34066 (N_34066,N_28554,N_28975);
nor U34067 (N_34067,N_27915,N_28736);
nor U34068 (N_34068,N_28175,N_28538);
nand U34069 (N_34069,N_26342,N_25280);
xnor U34070 (N_34070,N_27970,N_28995);
nand U34071 (N_34071,N_28278,N_29539);
or U34072 (N_34072,N_29177,N_26654);
or U34073 (N_34073,N_25102,N_29356);
nor U34074 (N_34074,N_25879,N_26104);
and U34075 (N_34075,N_25532,N_27716);
xor U34076 (N_34076,N_28691,N_26258);
nor U34077 (N_34077,N_27666,N_27473);
or U34078 (N_34078,N_26253,N_26666);
xor U34079 (N_34079,N_29242,N_27946);
nor U34080 (N_34080,N_28892,N_27879);
nor U34081 (N_34081,N_28967,N_28637);
and U34082 (N_34082,N_27513,N_29971);
nor U34083 (N_34083,N_29776,N_27643);
xnor U34084 (N_34084,N_26126,N_26371);
xor U34085 (N_34085,N_25503,N_25521);
or U34086 (N_34086,N_25393,N_29238);
xnor U34087 (N_34087,N_27815,N_28787);
and U34088 (N_34088,N_25856,N_27043);
or U34089 (N_34089,N_29044,N_28382);
and U34090 (N_34090,N_26658,N_26919);
or U34091 (N_34091,N_26445,N_25691);
and U34092 (N_34092,N_25375,N_27298);
nor U34093 (N_34093,N_27334,N_28883);
nand U34094 (N_34094,N_28879,N_27552);
xor U34095 (N_34095,N_26263,N_28319);
xnor U34096 (N_34096,N_27208,N_27944);
and U34097 (N_34097,N_25330,N_26338);
and U34098 (N_34098,N_26709,N_28497);
nand U34099 (N_34099,N_26044,N_26235);
xnor U34100 (N_34100,N_27799,N_28157);
nand U34101 (N_34101,N_29134,N_26695);
nor U34102 (N_34102,N_28359,N_27239);
and U34103 (N_34103,N_26299,N_25719);
nand U34104 (N_34104,N_28277,N_27895);
and U34105 (N_34105,N_27943,N_26913);
or U34106 (N_34106,N_27557,N_28417);
nor U34107 (N_34107,N_29088,N_26645);
nor U34108 (N_34108,N_26412,N_28717);
or U34109 (N_34109,N_27489,N_27646);
nor U34110 (N_34110,N_25826,N_29583);
nor U34111 (N_34111,N_26703,N_27227);
and U34112 (N_34112,N_28607,N_26134);
xnor U34113 (N_34113,N_29725,N_26710);
and U34114 (N_34114,N_28009,N_26845);
or U34115 (N_34115,N_29061,N_25147);
and U34116 (N_34116,N_27821,N_25316);
or U34117 (N_34117,N_25955,N_28109);
or U34118 (N_34118,N_28461,N_27303);
xor U34119 (N_34119,N_27934,N_26583);
and U34120 (N_34120,N_25109,N_29199);
xnor U34121 (N_34121,N_27819,N_29317);
nand U34122 (N_34122,N_29120,N_26004);
xor U34123 (N_34123,N_28155,N_29543);
nor U34124 (N_34124,N_26420,N_25124);
nand U34125 (N_34125,N_26723,N_25797);
or U34126 (N_34126,N_29631,N_25004);
or U34127 (N_34127,N_29350,N_28140);
nor U34128 (N_34128,N_27483,N_26773);
xnor U34129 (N_34129,N_26083,N_29517);
nor U34130 (N_34130,N_29420,N_27095);
nand U34131 (N_34131,N_25992,N_29096);
or U34132 (N_34132,N_26841,N_27092);
and U34133 (N_34133,N_27171,N_28180);
nand U34134 (N_34134,N_29589,N_25614);
xnor U34135 (N_34135,N_26253,N_25987);
or U34136 (N_34136,N_27170,N_29533);
xor U34137 (N_34137,N_27442,N_25862);
nand U34138 (N_34138,N_28732,N_28771);
and U34139 (N_34139,N_29866,N_27955);
nor U34140 (N_34140,N_25624,N_25531);
or U34141 (N_34141,N_29536,N_27682);
nand U34142 (N_34142,N_26647,N_25027);
nor U34143 (N_34143,N_29512,N_27244);
and U34144 (N_34144,N_26213,N_26277);
or U34145 (N_34145,N_25840,N_25907);
nand U34146 (N_34146,N_28721,N_28679);
and U34147 (N_34147,N_29527,N_29093);
nand U34148 (N_34148,N_27818,N_25816);
nand U34149 (N_34149,N_27081,N_29413);
xnor U34150 (N_34150,N_26354,N_26090);
nand U34151 (N_34151,N_29744,N_25001);
or U34152 (N_34152,N_26577,N_29793);
and U34153 (N_34153,N_26047,N_29531);
nand U34154 (N_34154,N_27775,N_27871);
and U34155 (N_34155,N_29376,N_29196);
nand U34156 (N_34156,N_28091,N_27279);
or U34157 (N_34157,N_27124,N_29817);
xnor U34158 (N_34158,N_27914,N_28984);
nor U34159 (N_34159,N_27680,N_28915);
xnor U34160 (N_34160,N_25666,N_28009);
nor U34161 (N_34161,N_26270,N_29649);
or U34162 (N_34162,N_28202,N_26230);
nor U34163 (N_34163,N_27175,N_29062);
xnor U34164 (N_34164,N_28006,N_27461);
nor U34165 (N_34165,N_26964,N_27403);
and U34166 (N_34166,N_25262,N_29970);
nand U34167 (N_34167,N_28372,N_27987);
or U34168 (N_34168,N_27305,N_26031);
or U34169 (N_34169,N_26745,N_25021);
and U34170 (N_34170,N_27919,N_25740);
nor U34171 (N_34171,N_26843,N_25515);
and U34172 (N_34172,N_27272,N_26045);
or U34173 (N_34173,N_25195,N_28805);
or U34174 (N_34174,N_25808,N_25992);
xor U34175 (N_34175,N_29939,N_27011);
nor U34176 (N_34176,N_27790,N_28784);
xnor U34177 (N_34177,N_29134,N_29079);
nor U34178 (N_34178,N_28455,N_29576);
nand U34179 (N_34179,N_28121,N_27337);
and U34180 (N_34180,N_26469,N_29803);
nor U34181 (N_34181,N_29257,N_26797);
and U34182 (N_34182,N_28108,N_26235);
and U34183 (N_34183,N_25521,N_25476);
nor U34184 (N_34184,N_25946,N_27165);
and U34185 (N_34185,N_29022,N_25645);
and U34186 (N_34186,N_29708,N_26811);
nor U34187 (N_34187,N_26090,N_25753);
or U34188 (N_34188,N_26376,N_29813);
and U34189 (N_34189,N_25304,N_28722);
and U34190 (N_34190,N_27768,N_28152);
xor U34191 (N_34191,N_25571,N_28565);
or U34192 (N_34192,N_27791,N_28136);
or U34193 (N_34193,N_27192,N_25098);
nor U34194 (N_34194,N_27761,N_25751);
nand U34195 (N_34195,N_26006,N_27910);
and U34196 (N_34196,N_25351,N_27282);
and U34197 (N_34197,N_28157,N_27636);
nand U34198 (N_34198,N_25697,N_27961);
and U34199 (N_34199,N_25339,N_26395);
or U34200 (N_34200,N_27581,N_27252);
nor U34201 (N_34201,N_27380,N_28973);
nand U34202 (N_34202,N_26015,N_26796);
and U34203 (N_34203,N_29231,N_25261);
or U34204 (N_34204,N_29480,N_29940);
xnor U34205 (N_34205,N_26878,N_25446);
nor U34206 (N_34206,N_28530,N_29463);
or U34207 (N_34207,N_25227,N_28145);
nor U34208 (N_34208,N_27581,N_25935);
and U34209 (N_34209,N_27383,N_29597);
or U34210 (N_34210,N_25109,N_29494);
and U34211 (N_34211,N_26227,N_26797);
nand U34212 (N_34212,N_25914,N_26724);
xnor U34213 (N_34213,N_26382,N_29804);
xnor U34214 (N_34214,N_26650,N_25830);
nor U34215 (N_34215,N_26378,N_28659);
and U34216 (N_34216,N_26613,N_25377);
nor U34217 (N_34217,N_29411,N_27761);
nand U34218 (N_34218,N_29152,N_26443);
nand U34219 (N_34219,N_25741,N_27114);
or U34220 (N_34220,N_27270,N_25639);
xnor U34221 (N_34221,N_25000,N_25346);
or U34222 (N_34222,N_28558,N_25365);
and U34223 (N_34223,N_26098,N_28288);
and U34224 (N_34224,N_29121,N_26665);
and U34225 (N_34225,N_27572,N_27740);
or U34226 (N_34226,N_25816,N_27701);
xor U34227 (N_34227,N_29745,N_26047);
nand U34228 (N_34228,N_25784,N_26869);
or U34229 (N_34229,N_28944,N_29008);
and U34230 (N_34230,N_29779,N_25846);
nor U34231 (N_34231,N_28230,N_25685);
nand U34232 (N_34232,N_28341,N_25311);
xor U34233 (N_34233,N_29834,N_26963);
nor U34234 (N_34234,N_26576,N_27421);
nor U34235 (N_34235,N_25336,N_28981);
and U34236 (N_34236,N_25452,N_28269);
nor U34237 (N_34237,N_29145,N_29625);
nor U34238 (N_34238,N_27057,N_25451);
or U34239 (N_34239,N_25773,N_26845);
and U34240 (N_34240,N_27667,N_29691);
nand U34241 (N_34241,N_29678,N_25425);
nor U34242 (N_34242,N_29560,N_27729);
nand U34243 (N_34243,N_27380,N_29715);
or U34244 (N_34244,N_26505,N_29725);
or U34245 (N_34245,N_26834,N_26462);
or U34246 (N_34246,N_27469,N_26773);
or U34247 (N_34247,N_29901,N_26494);
nor U34248 (N_34248,N_29681,N_28101);
nand U34249 (N_34249,N_26206,N_27500);
nor U34250 (N_34250,N_29021,N_26595);
nand U34251 (N_34251,N_26578,N_28403);
and U34252 (N_34252,N_25678,N_25384);
or U34253 (N_34253,N_25179,N_28334);
or U34254 (N_34254,N_25061,N_27401);
xnor U34255 (N_34255,N_28355,N_25829);
xor U34256 (N_34256,N_25887,N_29657);
or U34257 (N_34257,N_27104,N_28001);
nor U34258 (N_34258,N_27927,N_28426);
xor U34259 (N_34259,N_28420,N_26393);
xor U34260 (N_34260,N_29462,N_27177);
or U34261 (N_34261,N_29488,N_25038);
or U34262 (N_34262,N_27554,N_26044);
xor U34263 (N_34263,N_26305,N_25702);
or U34264 (N_34264,N_26703,N_25950);
or U34265 (N_34265,N_29013,N_25779);
nand U34266 (N_34266,N_29471,N_29758);
xor U34267 (N_34267,N_28779,N_28946);
or U34268 (N_34268,N_25609,N_26888);
nor U34269 (N_34269,N_28948,N_25006);
and U34270 (N_34270,N_29378,N_25696);
or U34271 (N_34271,N_26924,N_28100);
xnor U34272 (N_34272,N_26649,N_26642);
nand U34273 (N_34273,N_29512,N_27574);
nand U34274 (N_34274,N_29187,N_27798);
nor U34275 (N_34275,N_29318,N_27591);
nor U34276 (N_34276,N_26614,N_28384);
nor U34277 (N_34277,N_25530,N_27121);
and U34278 (N_34278,N_28072,N_26983);
nor U34279 (N_34279,N_28598,N_26567);
and U34280 (N_34280,N_25865,N_29045);
and U34281 (N_34281,N_26677,N_25919);
or U34282 (N_34282,N_25845,N_28590);
or U34283 (N_34283,N_28468,N_27463);
xor U34284 (N_34284,N_26067,N_28001);
nor U34285 (N_34285,N_26547,N_26811);
nand U34286 (N_34286,N_27279,N_28817);
nor U34287 (N_34287,N_29237,N_28487);
nand U34288 (N_34288,N_28572,N_28771);
and U34289 (N_34289,N_26916,N_26541);
nand U34290 (N_34290,N_28240,N_29513);
nor U34291 (N_34291,N_27593,N_28316);
and U34292 (N_34292,N_28175,N_26986);
and U34293 (N_34293,N_25405,N_26938);
nor U34294 (N_34294,N_25498,N_25984);
or U34295 (N_34295,N_26371,N_27125);
xor U34296 (N_34296,N_29597,N_29131);
xnor U34297 (N_34297,N_26427,N_27984);
nor U34298 (N_34298,N_28066,N_25146);
nand U34299 (N_34299,N_25122,N_29023);
xor U34300 (N_34300,N_29403,N_28509);
and U34301 (N_34301,N_27151,N_27923);
nor U34302 (N_34302,N_29711,N_27425);
nand U34303 (N_34303,N_29585,N_26116);
xnor U34304 (N_34304,N_28841,N_25512);
and U34305 (N_34305,N_29195,N_26700);
nor U34306 (N_34306,N_26928,N_26053);
and U34307 (N_34307,N_27713,N_28094);
xor U34308 (N_34308,N_27174,N_25252);
nand U34309 (N_34309,N_26936,N_29773);
or U34310 (N_34310,N_28336,N_27481);
and U34311 (N_34311,N_25052,N_29356);
nor U34312 (N_34312,N_26598,N_29641);
xor U34313 (N_34313,N_28315,N_27277);
and U34314 (N_34314,N_26378,N_25699);
nand U34315 (N_34315,N_27441,N_29738);
and U34316 (N_34316,N_28015,N_27949);
nand U34317 (N_34317,N_26319,N_25843);
nor U34318 (N_34318,N_29171,N_27670);
xnor U34319 (N_34319,N_25774,N_28637);
nor U34320 (N_34320,N_26409,N_27025);
and U34321 (N_34321,N_27759,N_28259);
or U34322 (N_34322,N_27566,N_28349);
nand U34323 (N_34323,N_29655,N_26084);
nand U34324 (N_34324,N_28169,N_29951);
or U34325 (N_34325,N_26209,N_26155);
nand U34326 (N_34326,N_28795,N_26639);
nand U34327 (N_34327,N_28932,N_28490);
nor U34328 (N_34328,N_25813,N_27307);
or U34329 (N_34329,N_25988,N_26336);
and U34330 (N_34330,N_28759,N_29238);
and U34331 (N_34331,N_29926,N_26162);
or U34332 (N_34332,N_29436,N_27429);
nor U34333 (N_34333,N_26974,N_25887);
xor U34334 (N_34334,N_28217,N_28430);
xor U34335 (N_34335,N_25545,N_28604);
nor U34336 (N_34336,N_25546,N_29459);
xor U34337 (N_34337,N_27285,N_29343);
nand U34338 (N_34338,N_29326,N_29473);
and U34339 (N_34339,N_27871,N_27609);
and U34340 (N_34340,N_29335,N_26290);
nand U34341 (N_34341,N_27976,N_28162);
and U34342 (N_34342,N_27533,N_25195);
nor U34343 (N_34343,N_25662,N_27248);
xnor U34344 (N_34344,N_25126,N_29781);
xnor U34345 (N_34345,N_28402,N_26876);
or U34346 (N_34346,N_25542,N_27936);
nor U34347 (N_34347,N_25224,N_29218);
nor U34348 (N_34348,N_26201,N_25473);
nor U34349 (N_34349,N_29811,N_25369);
or U34350 (N_34350,N_29098,N_28928);
nand U34351 (N_34351,N_26623,N_25592);
xnor U34352 (N_34352,N_25234,N_25004);
xnor U34353 (N_34353,N_25439,N_28371);
xor U34354 (N_34354,N_28208,N_29708);
nand U34355 (N_34355,N_27503,N_28398);
and U34356 (N_34356,N_27699,N_27472);
or U34357 (N_34357,N_26753,N_25652);
and U34358 (N_34358,N_27604,N_29974);
nor U34359 (N_34359,N_25058,N_27574);
nor U34360 (N_34360,N_29310,N_26326);
or U34361 (N_34361,N_25751,N_25788);
or U34362 (N_34362,N_25194,N_26441);
and U34363 (N_34363,N_26431,N_25498);
and U34364 (N_34364,N_26726,N_26692);
nand U34365 (N_34365,N_26978,N_27124);
xnor U34366 (N_34366,N_26668,N_28080);
nand U34367 (N_34367,N_29347,N_26301);
nor U34368 (N_34368,N_29106,N_28175);
or U34369 (N_34369,N_26809,N_28347);
xnor U34370 (N_34370,N_28420,N_27958);
xor U34371 (N_34371,N_28649,N_29996);
and U34372 (N_34372,N_27475,N_25826);
and U34373 (N_34373,N_28881,N_25110);
xor U34374 (N_34374,N_27700,N_25261);
xor U34375 (N_34375,N_27526,N_26262);
nand U34376 (N_34376,N_26349,N_28428);
and U34377 (N_34377,N_29050,N_29537);
and U34378 (N_34378,N_25110,N_29559);
nor U34379 (N_34379,N_28714,N_27332);
nor U34380 (N_34380,N_26529,N_28111);
nand U34381 (N_34381,N_26490,N_28169);
xor U34382 (N_34382,N_29150,N_28250);
and U34383 (N_34383,N_29999,N_25662);
and U34384 (N_34384,N_29761,N_29003);
xor U34385 (N_34385,N_27075,N_28455);
nor U34386 (N_34386,N_29448,N_28809);
and U34387 (N_34387,N_25740,N_28461);
nand U34388 (N_34388,N_27122,N_25786);
nor U34389 (N_34389,N_29430,N_25711);
nand U34390 (N_34390,N_29893,N_25938);
or U34391 (N_34391,N_25806,N_25397);
and U34392 (N_34392,N_27906,N_28334);
nor U34393 (N_34393,N_28734,N_27389);
xor U34394 (N_34394,N_28210,N_27030);
nor U34395 (N_34395,N_26412,N_27096);
xor U34396 (N_34396,N_28977,N_27926);
nor U34397 (N_34397,N_27833,N_26042);
nand U34398 (N_34398,N_29083,N_28695);
and U34399 (N_34399,N_27027,N_29156);
nand U34400 (N_34400,N_28262,N_28736);
nor U34401 (N_34401,N_29653,N_27288);
or U34402 (N_34402,N_28940,N_28989);
nor U34403 (N_34403,N_26953,N_25345);
nor U34404 (N_34404,N_28802,N_29208);
nor U34405 (N_34405,N_25176,N_29420);
nand U34406 (N_34406,N_28238,N_27336);
nand U34407 (N_34407,N_29463,N_29471);
or U34408 (N_34408,N_29223,N_28091);
xor U34409 (N_34409,N_28080,N_27147);
nor U34410 (N_34410,N_26617,N_27808);
nor U34411 (N_34411,N_27013,N_27182);
xnor U34412 (N_34412,N_27947,N_28666);
nand U34413 (N_34413,N_29055,N_28203);
nor U34414 (N_34414,N_26713,N_29985);
xor U34415 (N_34415,N_29526,N_26462);
xnor U34416 (N_34416,N_27227,N_27046);
or U34417 (N_34417,N_29687,N_27659);
or U34418 (N_34418,N_25848,N_28113);
or U34419 (N_34419,N_26419,N_29934);
nor U34420 (N_34420,N_27513,N_29684);
xor U34421 (N_34421,N_27445,N_26889);
nand U34422 (N_34422,N_26670,N_25086);
nand U34423 (N_34423,N_27519,N_28262);
and U34424 (N_34424,N_29419,N_26978);
nand U34425 (N_34425,N_29510,N_25693);
xnor U34426 (N_34426,N_29398,N_29090);
nor U34427 (N_34427,N_29683,N_26977);
or U34428 (N_34428,N_25083,N_26409);
nor U34429 (N_34429,N_27245,N_27398);
xnor U34430 (N_34430,N_25949,N_27038);
nor U34431 (N_34431,N_29255,N_27911);
nand U34432 (N_34432,N_29153,N_25129);
nand U34433 (N_34433,N_25575,N_28224);
nand U34434 (N_34434,N_25286,N_29514);
nand U34435 (N_34435,N_27097,N_25430);
nor U34436 (N_34436,N_25887,N_26958);
nand U34437 (N_34437,N_27018,N_29888);
nor U34438 (N_34438,N_25598,N_26878);
and U34439 (N_34439,N_25415,N_25265);
and U34440 (N_34440,N_27297,N_25099);
xor U34441 (N_34441,N_28634,N_28453);
nor U34442 (N_34442,N_28362,N_29722);
nor U34443 (N_34443,N_25788,N_27936);
and U34444 (N_34444,N_29830,N_26531);
nand U34445 (N_34445,N_25080,N_26910);
and U34446 (N_34446,N_29311,N_27356);
xor U34447 (N_34447,N_28448,N_25247);
nor U34448 (N_34448,N_26830,N_27901);
nand U34449 (N_34449,N_28908,N_26923);
or U34450 (N_34450,N_28488,N_25978);
and U34451 (N_34451,N_29621,N_27717);
nand U34452 (N_34452,N_27969,N_29373);
xnor U34453 (N_34453,N_25956,N_25019);
nand U34454 (N_34454,N_25793,N_25667);
and U34455 (N_34455,N_27679,N_25179);
nand U34456 (N_34456,N_26311,N_28231);
nor U34457 (N_34457,N_26482,N_25610);
nand U34458 (N_34458,N_25969,N_28549);
and U34459 (N_34459,N_27928,N_28151);
nor U34460 (N_34460,N_29119,N_25574);
nand U34461 (N_34461,N_25305,N_26572);
or U34462 (N_34462,N_26894,N_27362);
or U34463 (N_34463,N_28211,N_26266);
nand U34464 (N_34464,N_28475,N_27240);
and U34465 (N_34465,N_27759,N_28884);
and U34466 (N_34466,N_27260,N_26760);
nand U34467 (N_34467,N_29182,N_28892);
and U34468 (N_34468,N_28913,N_27829);
xor U34469 (N_34469,N_25317,N_28510);
and U34470 (N_34470,N_26103,N_29673);
xnor U34471 (N_34471,N_25730,N_26427);
and U34472 (N_34472,N_27379,N_28386);
xnor U34473 (N_34473,N_25855,N_29876);
xor U34474 (N_34474,N_27015,N_27268);
xnor U34475 (N_34475,N_26804,N_25723);
nand U34476 (N_34476,N_26818,N_25846);
xor U34477 (N_34477,N_26205,N_29980);
nand U34478 (N_34478,N_27134,N_26749);
or U34479 (N_34479,N_29866,N_28778);
and U34480 (N_34480,N_29004,N_27475);
and U34481 (N_34481,N_28968,N_27468);
and U34482 (N_34482,N_29448,N_26591);
or U34483 (N_34483,N_25842,N_25450);
nand U34484 (N_34484,N_28666,N_28218);
nor U34485 (N_34485,N_28455,N_25194);
nor U34486 (N_34486,N_27315,N_28085);
nand U34487 (N_34487,N_25090,N_25184);
and U34488 (N_34488,N_29260,N_26967);
nor U34489 (N_34489,N_25046,N_28945);
and U34490 (N_34490,N_27920,N_27554);
nand U34491 (N_34491,N_29814,N_26471);
nand U34492 (N_34492,N_27877,N_26783);
and U34493 (N_34493,N_25466,N_25295);
nand U34494 (N_34494,N_28329,N_29538);
and U34495 (N_34495,N_29242,N_27512);
and U34496 (N_34496,N_29710,N_28836);
and U34497 (N_34497,N_28832,N_29316);
or U34498 (N_34498,N_25959,N_29401);
nor U34499 (N_34499,N_27929,N_27054);
nand U34500 (N_34500,N_28602,N_27473);
nor U34501 (N_34501,N_26712,N_28333);
nand U34502 (N_34502,N_27713,N_26994);
nand U34503 (N_34503,N_27911,N_26526);
nor U34504 (N_34504,N_29235,N_29277);
nor U34505 (N_34505,N_27498,N_27337);
nor U34506 (N_34506,N_29196,N_26129);
nor U34507 (N_34507,N_29455,N_28356);
or U34508 (N_34508,N_25408,N_28413);
xor U34509 (N_34509,N_27961,N_27891);
or U34510 (N_34510,N_27855,N_28960);
nand U34511 (N_34511,N_27409,N_28721);
or U34512 (N_34512,N_26551,N_29452);
and U34513 (N_34513,N_26844,N_27114);
nand U34514 (N_34514,N_29345,N_28091);
and U34515 (N_34515,N_27547,N_25978);
xor U34516 (N_34516,N_27617,N_27039);
and U34517 (N_34517,N_27600,N_25995);
xor U34518 (N_34518,N_26987,N_26480);
and U34519 (N_34519,N_27050,N_26197);
nor U34520 (N_34520,N_27282,N_26834);
nor U34521 (N_34521,N_27166,N_26643);
nand U34522 (N_34522,N_26855,N_28982);
and U34523 (N_34523,N_27764,N_29627);
and U34524 (N_34524,N_26465,N_27153);
xnor U34525 (N_34525,N_29149,N_28951);
nor U34526 (N_34526,N_25190,N_28497);
nand U34527 (N_34527,N_27286,N_26558);
nor U34528 (N_34528,N_29060,N_26839);
xnor U34529 (N_34529,N_28193,N_25480);
and U34530 (N_34530,N_29708,N_29801);
and U34531 (N_34531,N_25834,N_27623);
or U34532 (N_34532,N_29803,N_29501);
or U34533 (N_34533,N_26445,N_29649);
or U34534 (N_34534,N_25425,N_28665);
nor U34535 (N_34535,N_25027,N_28041);
xor U34536 (N_34536,N_27246,N_29447);
nor U34537 (N_34537,N_29533,N_29643);
or U34538 (N_34538,N_28412,N_27376);
and U34539 (N_34539,N_28204,N_25029);
and U34540 (N_34540,N_27821,N_25617);
nor U34541 (N_34541,N_29071,N_29816);
or U34542 (N_34542,N_29768,N_29200);
nand U34543 (N_34543,N_26932,N_28978);
and U34544 (N_34544,N_25066,N_29522);
xor U34545 (N_34545,N_26023,N_27069);
or U34546 (N_34546,N_26701,N_25730);
or U34547 (N_34547,N_29430,N_25847);
nor U34548 (N_34548,N_29847,N_26034);
nor U34549 (N_34549,N_29664,N_27554);
or U34550 (N_34550,N_27649,N_27053);
or U34551 (N_34551,N_26722,N_25882);
and U34552 (N_34552,N_29303,N_27356);
xor U34553 (N_34553,N_29512,N_26723);
nor U34554 (N_34554,N_25775,N_29953);
and U34555 (N_34555,N_27909,N_26911);
nand U34556 (N_34556,N_29304,N_29475);
nand U34557 (N_34557,N_25562,N_28527);
nor U34558 (N_34558,N_29725,N_28618);
xnor U34559 (N_34559,N_26395,N_28177);
nor U34560 (N_34560,N_28161,N_26248);
xnor U34561 (N_34561,N_27474,N_26291);
nor U34562 (N_34562,N_26073,N_25366);
nand U34563 (N_34563,N_29440,N_25765);
nor U34564 (N_34564,N_29821,N_26703);
or U34565 (N_34565,N_26992,N_26027);
nand U34566 (N_34566,N_25551,N_28695);
xnor U34567 (N_34567,N_27727,N_27393);
xor U34568 (N_34568,N_26705,N_27396);
xnor U34569 (N_34569,N_27357,N_28978);
nand U34570 (N_34570,N_28171,N_26444);
nor U34571 (N_34571,N_29739,N_26002);
nand U34572 (N_34572,N_25549,N_25307);
and U34573 (N_34573,N_25412,N_29596);
or U34574 (N_34574,N_26687,N_27005);
nor U34575 (N_34575,N_27266,N_27753);
nor U34576 (N_34576,N_28382,N_29326);
and U34577 (N_34577,N_26859,N_28233);
nand U34578 (N_34578,N_26840,N_26940);
or U34579 (N_34579,N_25630,N_28098);
nor U34580 (N_34580,N_28533,N_28332);
or U34581 (N_34581,N_25873,N_27257);
or U34582 (N_34582,N_27736,N_28735);
nor U34583 (N_34583,N_26156,N_25332);
and U34584 (N_34584,N_26269,N_27928);
and U34585 (N_34585,N_26522,N_28072);
or U34586 (N_34586,N_29607,N_28337);
and U34587 (N_34587,N_29889,N_28054);
xor U34588 (N_34588,N_27410,N_29053);
and U34589 (N_34589,N_25605,N_25025);
nor U34590 (N_34590,N_27304,N_25145);
or U34591 (N_34591,N_28126,N_25664);
or U34592 (N_34592,N_27740,N_29757);
or U34593 (N_34593,N_29904,N_26156);
xor U34594 (N_34594,N_29449,N_27664);
xor U34595 (N_34595,N_28876,N_25077);
xor U34596 (N_34596,N_29634,N_25249);
nor U34597 (N_34597,N_27216,N_27044);
and U34598 (N_34598,N_28525,N_28225);
nand U34599 (N_34599,N_26581,N_26245);
nand U34600 (N_34600,N_29984,N_29649);
nand U34601 (N_34601,N_28025,N_28454);
nand U34602 (N_34602,N_27850,N_27402);
nand U34603 (N_34603,N_27390,N_25126);
nor U34604 (N_34604,N_28556,N_28691);
and U34605 (N_34605,N_25941,N_29120);
nor U34606 (N_34606,N_25003,N_25207);
or U34607 (N_34607,N_28846,N_25013);
nand U34608 (N_34608,N_25249,N_26422);
xnor U34609 (N_34609,N_28383,N_27358);
nand U34610 (N_34610,N_27997,N_26359);
nand U34611 (N_34611,N_26052,N_25495);
nand U34612 (N_34612,N_29015,N_28147);
and U34613 (N_34613,N_27707,N_26837);
nand U34614 (N_34614,N_28316,N_27668);
or U34615 (N_34615,N_26503,N_28873);
nand U34616 (N_34616,N_29546,N_27594);
nand U34617 (N_34617,N_26093,N_28020);
nor U34618 (N_34618,N_27468,N_26865);
nor U34619 (N_34619,N_25931,N_29065);
nand U34620 (N_34620,N_29651,N_26484);
nand U34621 (N_34621,N_26652,N_27405);
xnor U34622 (N_34622,N_26274,N_29394);
nor U34623 (N_34623,N_25160,N_25731);
or U34624 (N_34624,N_26921,N_27325);
nand U34625 (N_34625,N_29299,N_25959);
and U34626 (N_34626,N_26839,N_29110);
nand U34627 (N_34627,N_27116,N_29339);
nor U34628 (N_34628,N_27664,N_27062);
nor U34629 (N_34629,N_29725,N_28671);
and U34630 (N_34630,N_26824,N_26220);
nand U34631 (N_34631,N_28791,N_28656);
nor U34632 (N_34632,N_26294,N_27094);
and U34633 (N_34633,N_25427,N_28801);
or U34634 (N_34634,N_27573,N_27135);
xor U34635 (N_34635,N_26020,N_28408);
xnor U34636 (N_34636,N_29129,N_29361);
nand U34637 (N_34637,N_29964,N_25348);
xor U34638 (N_34638,N_28096,N_25849);
and U34639 (N_34639,N_29594,N_25607);
or U34640 (N_34640,N_29698,N_29332);
xor U34641 (N_34641,N_25694,N_26695);
xor U34642 (N_34642,N_28143,N_25862);
or U34643 (N_34643,N_28740,N_28073);
and U34644 (N_34644,N_28445,N_26197);
nor U34645 (N_34645,N_28940,N_26843);
nand U34646 (N_34646,N_29503,N_29361);
or U34647 (N_34647,N_25115,N_25760);
or U34648 (N_34648,N_29438,N_26351);
nor U34649 (N_34649,N_27929,N_28607);
and U34650 (N_34650,N_26925,N_29086);
or U34651 (N_34651,N_29361,N_26120);
and U34652 (N_34652,N_27775,N_26166);
nand U34653 (N_34653,N_29949,N_29241);
or U34654 (N_34654,N_25404,N_25800);
and U34655 (N_34655,N_26910,N_26299);
xnor U34656 (N_34656,N_29673,N_25194);
or U34657 (N_34657,N_28195,N_29982);
and U34658 (N_34658,N_27019,N_29404);
nor U34659 (N_34659,N_28484,N_27770);
xor U34660 (N_34660,N_29912,N_27237);
nand U34661 (N_34661,N_29354,N_26482);
nor U34662 (N_34662,N_26666,N_29539);
nor U34663 (N_34663,N_29490,N_28846);
and U34664 (N_34664,N_27399,N_27201);
nand U34665 (N_34665,N_27905,N_26406);
xnor U34666 (N_34666,N_25098,N_28295);
nor U34667 (N_34667,N_27424,N_28361);
and U34668 (N_34668,N_26374,N_28117);
or U34669 (N_34669,N_29162,N_26489);
nand U34670 (N_34670,N_29186,N_29944);
nor U34671 (N_34671,N_26354,N_25623);
nor U34672 (N_34672,N_26881,N_27738);
or U34673 (N_34673,N_26258,N_27439);
and U34674 (N_34674,N_28366,N_27721);
nor U34675 (N_34675,N_25308,N_27707);
and U34676 (N_34676,N_29630,N_25130);
nor U34677 (N_34677,N_29328,N_29236);
xnor U34678 (N_34678,N_29309,N_27539);
xor U34679 (N_34679,N_27287,N_27397);
nand U34680 (N_34680,N_26550,N_27735);
xnor U34681 (N_34681,N_28159,N_28265);
xnor U34682 (N_34682,N_26057,N_28556);
nand U34683 (N_34683,N_27853,N_25973);
nand U34684 (N_34684,N_25163,N_26205);
nand U34685 (N_34685,N_26159,N_26127);
nor U34686 (N_34686,N_28694,N_26278);
and U34687 (N_34687,N_25689,N_25005);
xnor U34688 (N_34688,N_29649,N_26217);
xor U34689 (N_34689,N_27725,N_28170);
nor U34690 (N_34690,N_29172,N_26383);
nor U34691 (N_34691,N_28424,N_26052);
nor U34692 (N_34692,N_26521,N_29000);
and U34693 (N_34693,N_26527,N_26234);
xor U34694 (N_34694,N_26625,N_25629);
xnor U34695 (N_34695,N_26735,N_26020);
xor U34696 (N_34696,N_29464,N_29317);
nand U34697 (N_34697,N_29309,N_28557);
nand U34698 (N_34698,N_29444,N_27599);
xnor U34699 (N_34699,N_26662,N_28567);
and U34700 (N_34700,N_26668,N_27014);
xor U34701 (N_34701,N_28553,N_28277);
xor U34702 (N_34702,N_28162,N_27167);
nand U34703 (N_34703,N_27696,N_28766);
xnor U34704 (N_34704,N_27529,N_26682);
nand U34705 (N_34705,N_25050,N_28805);
nand U34706 (N_34706,N_28240,N_29217);
nand U34707 (N_34707,N_25414,N_28006);
or U34708 (N_34708,N_26868,N_26611);
nand U34709 (N_34709,N_26018,N_25928);
xnor U34710 (N_34710,N_26277,N_28448);
or U34711 (N_34711,N_27031,N_29615);
nor U34712 (N_34712,N_27816,N_29596);
nor U34713 (N_34713,N_27229,N_28703);
nor U34714 (N_34714,N_27475,N_28870);
xor U34715 (N_34715,N_29053,N_27851);
nor U34716 (N_34716,N_26023,N_26920);
nand U34717 (N_34717,N_27332,N_28877);
nor U34718 (N_34718,N_25755,N_25260);
nor U34719 (N_34719,N_28865,N_29151);
and U34720 (N_34720,N_26439,N_27760);
or U34721 (N_34721,N_26786,N_26574);
or U34722 (N_34722,N_29650,N_26799);
xor U34723 (N_34723,N_27639,N_27728);
or U34724 (N_34724,N_28973,N_25552);
nor U34725 (N_34725,N_26340,N_27896);
or U34726 (N_34726,N_28360,N_28246);
xnor U34727 (N_34727,N_27564,N_29075);
and U34728 (N_34728,N_28709,N_26426);
nand U34729 (N_34729,N_29063,N_28469);
xnor U34730 (N_34730,N_26463,N_25815);
or U34731 (N_34731,N_29276,N_25448);
nand U34732 (N_34732,N_29035,N_28542);
nand U34733 (N_34733,N_28885,N_29898);
nand U34734 (N_34734,N_27781,N_29668);
xor U34735 (N_34735,N_27763,N_27543);
xor U34736 (N_34736,N_29471,N_27419);
xor U34737 (N_34737,N_28434,N_26010);
or U34738 (N_34738,N_26391,N_26494);
and U34739 (N_34739,N_29012,N_29667);
or U34740 (N_34740,N_26829,N_29905);
and U34741 (N_34741,N_26518,N_26716);
xnor U34742 (N_34742,N_25215,N_25151);
xnor U34743 (N_34743,N_26282,N_26176);
xor U34744 (N_34744,N_26149,N_28572);
xnor U34745 (N_34745,N_29513,N_26845);
xnor U34746 (N_34746,N_25817,N_25881);
nor U34747 (N_34747,N_28339,N_25639);
xor U34748 (N_34748,N_26167,N_26054);
nor U34749 (N_34749,N_27827,N_28077);
nor U34750 (N_34750,N_29435,N_28158);
xnor U34751 (N_34751,N_29452,N_27111);
nand U34752 (N_34752,N_29006,N_26672);
xor U34753 (N_34753,N_28251,N_27872);
nor U34754 (N_34754,N_25310,N_26410);
nor U34755 (N_34755,N_26664,N_26164);
or U34756 (N_34756,N_28352,N_27795);
or U34757 (N_34757,N_29110,N_29982);
nand U34758 (N_34758,N_29422,N_26705);
or U34759 (N_34759,N_26349,N_25447);
or U34760 (N_34760,N_26361,N_25669);
nor U34761 (N_34761,N_27963,N_29392);
nor U34762 (N_34762,N_29000,N_29772);
nand U34763 (N_34763,N_26410,N_26968);
xnor U34764 (N_34764,N_28778,N_26743);
xor U34765 (N_34765,N_28959,N_29835);
or U34766 (N_34766,N_29715,N_25973);
xnor U34767 (N_34767,N_29823,N_26152);
xor U34768 (N_34768,N_29329,N_28269);
or U34769 (N_34769,N_27760,N_26351);
nor U34770 (N_34770,N_29282,N_25803);
nor U34771 (N_34771,N_26496,N_29330);
or U34772 (N_34772,N_28109,N_27640);
and U34773 (N_34773,N_26924,N_25850);
nor U34774 (N_34774,N_27041,N_29838);
and U34775 (N_34775,N_28478,N_26661);
and U34776 (N_34776,N_26705,N_25430);
nand U34777 (N_34777,N_26452,N_26194);
nand U34778 (N_34778,N_26854,N_26786);
and U34779 (N_34779,N_27691,N_28250);
or U34780 (N_34780,N_26840,N_25405);
nand U34781 (N_34781,N_29303,N_29728);
and U34782 (N_34782,N_25108,N_26860);
or U34783 (N_34783,N_25508,N_28156);
nor U34784 (N_34784,N_29371,N_28363);
or U34785 (N_34785,N_29087,N_29376);
or U34786 (N_34786,N_27826,N_28448);
xor U34787 (N_34787,N_29608,N_27849);
and U34788 (N_34788,N_27550,N_26598);
or U34789 (N_34789,N_29687,N_29796);
xor U34790 (N_34790,N_25263,N_29726);
or U34791 (N_34791,N_29915,N_28928);
or U34792 (N_34792,N_26003,N_28957);
nor U34793 (N_34793,N_27403,N_26805);
and U34794 (N_34794,N_26708,N_25910);
xnor U34795 (N_34795,N_26422,N_28987);
xnor U34796 (N_34796,N_28011,N_25267);
nand U34797 (N_34797,N_28023,N_26515);
nand U34798 (N_34798,N_25743,N_25571);
nor U34799 (N_34799,N_28365,N_26748);
and U34800 (N_34800,N_25093,N_25398);
nor U34801 (N_34801,N_28247,N_28500);
xnor U34802 (N_34802,N_28857,N_29504);
nor U34803 (N_34803,N_28852,N_26927);
nand U34804 (N_34804,N_27763,N_29366);
nand U34805 (N_34805,N_28572,N_29602);
and U34806 (N_34806,N_28776,N_26854);
nand U34807 (N_34807,N_29272,N_29205);
xor U34808 (N_34808,N_26093,N_25137);
xnor U34809 (N_34809,N_28355,N_26982);
nor U34810 (N_34810,N_28670,N_25496);
nor U34811 (N_34811,N_26933,N_26351);
nor U34812 (N_34812,N_25548,N_26035);
nor U34813 (N_34813,N_27890,N_27190);
or U34814 (N_34814,N_28531,N_25356);
nand U34815 (N_34815,N_27987,N_26609);
nor U34816 (N_34816,N_29804,N_26881);
or U34817 (N_34817,N_28370,N_25057);
xor U34818 (N_34818,N_27965,N_29030);
or U34819 (N_34819,N_26394,N_25058);
xor U34820 (N_34820,N_26280,N_26455);
xnor U34821 (N_34821,N_26237,N_25229);
nor U34822 (N_34822,N_29585,N_25639);
or U34823 (N_34823,N_25797,N_27481);
or U34824 (N_34824,N_28240,N_28694);
and U34825 (N_34825,N_26866,N_25956);
xor U34826 (N_34826,N_28157,N_29808);
xnor U34827 (N_34827,N_29111,N_27385);
xor U34828 (N_34828,N_28929,N_28033);
nand U34829 (N_34829,N_28546,N_28345);
xor U34830 (N_34830,N_27264,N_28241);
xor U34831 (N_34831,N_27055,N_26548);
nand U34832 (N_34832,N_28894,N_29048);
nand U34833 (N_34833,N_25483,N_26597);
nand U34834 (N_34834,N_27569,N_26372);
and U34835 (N_34835,N_26281,N_25381);
nand U34836 (N_34836,N_25248,N_27703);
and U34837 (N_34837,N_29184,N_28853);
or U34838 (N_34838,N_28089,N_29711);
and U34839 (N_34839,N_29321,N_29263);
and U34840 (N_34840,N_28226,N_26915);
xnor U34841 (N_34841,N_27818,N_27506);
xnor U34842 (N_34842,N_28135,N_25633);
or U34843 (N_34843,N_28830,N_27273);
and U34844 (N_34844,N_26328,N_27428);
xor U34845 (N_34845,N_29112,N_28465);
or U34846 (N_34846,N_29500,N_28692);
nor U34847 (N_34847,N_26966,N_25580);
and U34848 (N_34848,N_29282,N_26056);
nor U34849 (N_34849,N_29599,N_28496);
or U34850 (N_34850,N_29699,N_28724);
nor U34851 (N_34851,N_26996,N_26840);
and U34852 (N_34852,N_25826,N_25340);
or U34853 (N_34853,N_28704,N_28220);
nand U34854 (N_34854,N_26881,N_25882);
xor U34855 (N_34855,N_29697,N_26722);
and U34856 (N_34856,N_29241,N_28580);
or U34857 (N_34857,N_28172,N_25107);
or U34858 (N_34858,N_25431,N_27113);
nor U34859 (N_34859,N_26441,N_27012);
and U34860 (N_34860,N_25969,N_25297);
nor U34861 (N_34861,N_26983,N_26276);
xor U34862 (N_34862,N_28517,N_27905);
or U34863 (N_34863,N_25724,N_25406);
or U34864 (N_34864,N_28853,N_29529);
nor U34865 (N_34865,N_25091,N_27039);
xnor U34866 (N_34866,N_25626,N_27112);
and U34867 (N_34867,N_25607,N_26768);
and U34868 (N_34868,N_29241,N_25227);
or U34869 (N_34869,N_25203,N_25054);
and U34870 (N_34870,N_28540,N_28325);
nor U34871 (N_34871,N_26913,N_27579);
nand U34872 (N_34872,N_29622,N_27113);
or U34873 (N_34873,N_25936,N_28319);
xor U34874 (N_34874,N_26525,N_25708);
nand U34875 (N_34875,N_27216,N_25144);
nor U34876 (N_34876,N_26576,N_29694);
or U34877 (N_34877,N_26903,N_26779);
nor U34878 (N_34878,N_28650,N_27413);
nand U34879 (N_34879,N_27059,N_27551);
nand U34880 (N_34880,N_29192,N_25854);
nor U34881 (N_34881,N_26519,N_26124);
xor U34882 (N_34882,N_29378,N_27122);
nand U34883 (N_34883,N_27321,N_26182);
and U34884 (N_34884,N_27629,N_25338);
nor U34885 (N_34885,N_26411,N_27797);
and U34886 (N_34886,N_27298,N_25613);
nor U34887 (N_34887,N_27078,N_25172);
nor U34888 (N_34888,N_28069,N_29984);
xor U34889 (N_34889,N_28957,N_26847);
and U34890 (N_34890,N_29997,N_26298);
nand U34891 (N_34891,N_28505,N_28762);
nand U34892 (N_34892,N_26993,N_29313);
nand U34893 (N_34893,N_25469,N_28037);
or U34894 (N_34894,N_28522,N_26286);
nor U34895 (N_34895,N_27969,N_28377);
nand U34896 (N_34896,N_27253,N_28753);
xor U34897 (N_34897,N_29751,N_29134);
xor U34898 (N_34898,N_25980,N_26268);
xnor U34899 (N_34899,N_27266,N_26394);
nor U34900 (N_34900,N_27974,N_27325);
nand U34901 (N_34901,N_26709,N_26342);
nand U34902 (N_34902,N_29646,N_25746);
or U34903 (N_34903,N_28806,N_27843);
nor U34904 (N_34904,N_26762,N_29882);
or U34905 (N_34905,N_27014,N_29761);
xor U34906 (N_34906,N_25981,N_26307);
nand U34907 (N_34907,N_29216,N_26544);
nor U34908 (N_34908,N_25371,N_27034);
nor U34909 (N_34909,N_26043,N_26003);
nor U34910 (N_34910,N_27986,N_25936);
and U34911 (N_34911,N_29782,N_26930);
or U34912 (N_34912,N_29666,N_29035);
nor U34913 (N_34913,N_26244,N_29989);
nand U34914 (N_34914,N_29969,N_29614);
nor U34915 (N_34915,N_26596,N_25661);
nand U34916 (N_34916,N_27621,N_29330);
nor U34917 (N_34917,N_28373,N_25520);
xor U34918 (N_34918,N_26508,N_25056);
xnor U34919 (N_34919,N_25890,N_26492);
nor U34920 (N_34920,N_25888,N_28879);
nand U34921 (N_34921,N_26984,N_25247);
nand U34922 (N_34922,N_29574,N_29528);
xor U34923 (N_34923,N_27581,N_26304);
nand U34924 (N_34924,N_29056,N_28623);
and U34925 (N_34925,N_25025,N_28308);
nand U34926 (N_34926,N_28987,N_28874);
nor U34927 (N_34927,N_27254,N_28215);
and U34928 (N_34928,N_29402,N_25515);
xnor U34929 (N_34929,N_27515,N_29224);
and U34930 (N_34930,N_26140,N_26868);
and U34931 (N_34931,N_29284,N_27332);
and U34932 (N_34932,N_26074,N_26990);
xnor U34933 (N_34933,N_27166,N_29301);
nand U34934 (N_34934,N_27094,N_29706);
nand U34935 (N_34935,N_26437,N_28363);
and U34936 (N_34936,N_29965,N_27980);
or U34937 (N_34937,N_25252,N_28417);
nor U34938 (N_34938,N_26545,N_28854);
xor U34939 (N_34939,N_25218,N_28767);
xor U34940 (N_34940,N_28247,N_26418);
and U34941 (N_34941,N_27861,N_25180);
xor U34942 (N_34942,N_25128,N_28958);
and U34943 (N_34943,N_27573,N_27068);
xor U34944 (N_34944,N_29304,N_25777);
or U34945 (N_34945,N_29149,N_25022);
nand U34946 (N_34946,N_26852,N_28941);
nand U34947 (N_34947,N_25273,N_29635);
or U34948 (N_34948,N_29650,N_29329);
nand U34949 (N_34949,N_27499,N_27646);
nand U34950 (N_34950,N_26455,N_28084);
or U34951 (N_34951,N_27135,N_26651);
and U34952 (N_34952,N_27451,N_29929);
nor U34953 (N_34953,N_25983,N_26434);
nor U34954 (N_34954,N_28644,N_26600);
and U34955 (N_34955,N_29045,N_25512);
nand U34956 (N_34956,N_27196,N_25079);
or U34957 (N_34957,N_26375,N_27077);
nand U34958 (N_34958,N_26154,N_29289);
nand U34959 (N_34959,N_26356,N_25874);
nand U34960 (N_34960,N_29344,N_25993);
xor U34961 (N_34961,N_29168,N_27646);
or U34962 (N_34962,N_29649,N_27820);
nor U34963 (N_34963,N_27988,N_27370);
nand U34964 (N_34964,N_25635,N_27697);
xnor U34965 (N_34965,N_28229,N_29995);
or U34966 (N_34966,N_29959,N_28317);
or U34967 (N_34967,N_28971,N_27751);
xor U34968 (N_34968,N_29325,N_29612);
and U34969 (N_34969,N_25769,N_25202);
nand U34970 (N_34970,N_26669,N_27205);
xnor U34971 (N_34971,N_27329,N_26983);
nor U34972 (N_34972,N_29880,N_29988);
nand U34973 (N_34973,N_25352,N_28835);
xor U34974 (N_34974,N_29122,N_25612);
or U34975 (N_34975,N_29697,N_26737);
nor U34976 (N_34976,N_27916,N_27686);
and U34977 (N_34977,N_26499,N_28297);
nand U34978 (N_34978,N_29292,N_29413);
xnor U34979 (N_34979,N_29017,N_25348);
nor U34980 (N_34980,N_27594,N_26645);
xor U34981 (N_34981,N_25781,N_28647);
nor U34982 (N_34982,N_29669,N_28238);
nor U34983 (N_34983,N_27782,N_28192);
and U34984 (N_34984,N_27663,N_28418);
or U34985 (N_34985,N_27024,N_29432);
and U34986 (N_34986,N_26387,N_27169);
or U34987 (N_34987,N_26243,N_26317);
nand U34988 (N_34988,N_29020,N_29249);
nor U34989 (N_34989,N_26324,N_29630);
or U34990 (N_34990,N_25968,N_26537);
nand U34991 (N_34991,N_28683,N_29543);
nand U34992 (N_34992,N_27365,N_25687);
or U34993 (N_34993,N_25505,N_27863);
and U34994 (N_34994,N_27344,N_25333);
nor U34995 (N_34995,N_28078,N_27805);
xnor U34996 (N_34996,N_25435,N_27101);
nand U34997 (N_34997,N_26687,N_28085);
xnor U34998 (N_34998,N_25821,N_27472);
nand U34999 (N_34999,N_28624,N_28952);
nand U35000 (N_35000,N_34954,N_34363);
xnor U35001 (N_35001,N_30581,N_34928);
and U35002 (N_35002,N_31900,N_34721);
nor U35003 (N_35003,N_30746,N_31409);
and U35004 (N_35004,N_34916,N_34979);
or U35005 (N_35005,N_30562,N_32298);
nor U35006 (N_35006,N_30007,N_34115);
and U35007 (N_35007,N_31803,N_32071);
nand U35008 (N_35008,N_31408,N_32973);
xor U35009 (N_35009,N_34658,N_32295);
nor U35010 (N_35010,N_31319,N_31637);
nand U35011 (N_35011,N_30878,N_31283);
and U35012 (N_35012,N_31556,N_33572);
nor U35013 (N_35013,N_31433,N_30870);
nor U35014 (N_35014,N_34023,N_30865);
xor U35015 (N_35015,N_33560,N_32429);
nor U35016 (N_35016,N_31581,N_33435);
nor U35017 (N_35017,N_31591,N_30180);
nand U35018 (N_35018,N_30088,N_33353);
nor U35019 (N_35019,N_31702,N_31429);
xnor U35020 (N_35020,N_32277,N_33437);
or U35021 (N_35021,N_30809,N_32190);
nand U35022 (N_35022,N_30889,N_31589);
xor U35023 (N_35023,N_31576,N_34564);
or U35024 (N_35024,N_31382,N_32212);
nor U35025 (N_35025,N_33331,N_30300);
and U35026 (N_35026,N_31874,N_31389);
or U35027 (N_35027,N_34615,N_34887);
or U35028 (N_35028,N_32644,N_34290);
nand U35029 (N_35029,N_30165,N_31437);
xnor U35030 (N_35030,N_32886,N_33381);
and U35031 (N_35031,N_30532,N_32284);
and U35032 (N_35032,N_33406,N_34538);
and U35033 (N_35033,N_33957,N_34071);
nand U35034 (N_35034,N_33279,N_30525);
nand U35035 (N_35035,N_31942,N_31203);
nor U35036 (N_35036,N_34265,N_31905);
and U35037 (N_35037,N_30254,N_34473);
or U35038 (N_35038,N_34902,N_31765);
xnor U35039 (N_35039,N_30908,N_31199);
nand U35040 (N_35040,N_31695,N_31582);
nor U35041 (N_35041,N_30716,N_30071);
nor U35042 (N_35042,N_32697,N_34355);
and U35043 (N_35043,N_33045,N_32322);
and U35044 (N_35044,N_33697,N_33388);
xnor U35045 (N_35045,N_30591,N_33173);
or U35046 (N_35046,N_32752,N_34974);
or U35047 (N_35047,N_34406,N_33681);
or U35048 (N_35048,N_31760,N_30329);
and U35049 (N_35049,N_32801,N_30319);
or U35050 (N_35050,N_34193,N_32845);
and U35051 (N_35051,N_34848,N_31420);
or U35052 (N_35052,N_34818,N_31109);
xnor U35053 (N_35053,N_32063,N_33981);
nand U35054 (N_35054,N_30008,N_33880);
and U35055 (N_35055,N_32565,N_33618);
or U35056 (N_35056,N_33079,N_30172);
or U35057 (N_35057,N_30408,N_34184);
nand U35058 (N_35058,N_34268,N_32596);
xor U35059 (N_35059,N_33531,N_34388);
nor U35060 (N_35060,N_32229,N_34311);
or U35061 (N_35061,N_30712,N_31662);
and U35062 (N_35062,N_30406,N_30139);
or U35063 (N_35063,N_34202,N_33204);
or U35064 (N_35064,N_33649,N_31691);
nand U35065 (N_35065,N_30346,N_33202);
nand U35066 (N_35066,N_32986,N_33899);
nor U35067 (N_35067,N_30484,N_34965);
xor U35068 (N_35068,N_30128,N_31643);
xnor U35069 (N_35069,N_32869,N_32529);
nor U35070 (N_35070,N_31380,N_33281);
or U35071 (N_35071,N_31128,N_31371);
nor U35072 (N_35072,N_32274,N_31031);
xor U35073 (N_35073,N_31627,N_33501);
nor U35074 (N_35074,N_30205,N_30987);
nor U35075 (N_35075,N_31796,N_33087);
nand U35076 (N_35076,N_33042,N_33772);
and U35077 (N_35077,N_33952,N_33360);
or U35078 (N_35078,N_31293,N_30174);
and U35079 (N_35079,N_32953,N_34940);
and U35080 (N_35080,N_30785,N_30695);
nand U35081 (N_35081,N_30850,N_32200);
nand U35082 (N_35082,N_32877,N_31344);
xor U35083 (N_35083,N_34240,N_33873);
or U35084 (N_35084,N_31879,N_33332);
nand U35085 (N_35085,N_31431,N_32416);
xor U35086 (N_35086,N_34671,N_30732);
or U35087 (N_35087,N_34936,N_32810);
and U35088 (N_35088,N_32796,N_34574);
nand U35089 (N_35089,N_31148,N_30937);
nand U35090 (N_35090,N_31041,N_31374);
nand U35091 (N_35091,N_33917,N_30125);
nand U35092 (N_35092,N_30580,N_32285);
nor U35093 (N_35093,N_30653,N_31728);
nand U35094 (N_35094,N_33194,N_32292);
nand U35095 (N_35095,N_34162,N_30586);
xnor U35096 (N_35096,N_31514,N_30787);
nor U35097 (N_35097,N_32572,N_30237);
and U35098 (N_35098,N_30980,N_34725);
or U35099 (N_35099,N_34672,N_30768);
nand U35100 (N_35100,N_30020,N_33887);
xnor U35101 (N_35101,N_31625,N_32034);
and U35102 (N_35102,N_34906,N_32121);
and U35103 (N_35103,N_31384,N_31926);
and U35104 (N_35104,N_33432,N_31354);
nor U35105 (N_35105,N_31010,N_33668);
or U35106 (N_35106,N_33518,N_32512);
and U35107 (N_35107,N_30110,N_31676);
nand U35108 (N_35108,N_32922,N_32041);
and U35109 (N_35109,N_33716,N_32882);
nor U35110 (N_35110,N_32148,N_34116);
or U35111 (N_35111,N_32055,N_31516);
nor U35112 (N_35112,N_30806,N_30799);
xnor U35113 (N_35113,N_32773,N_31217);
nand U35114 (N_35114,N_33617,N_33174);
nand U35115 (N_35115,N_31809,N_32413);
and U35116 (N_35116,N_31457,N_32770);
and U35117 (N_35117,N_30642,N_34398);
nand U35118 (N_35118,N_30881,N_30348);
nand U35119 (N_35119,N_31822,N_31648);
xnor U35120 (N_35120,N_31274,N_33236);
xnor U35121 (N_35121,N_32219,N_32974);
xnor U35122 (N_35122,N_31546,N_33597);
nor U35123 (N_35123,N_32500,N_31321);
xnor U35124 (N_35124,N_31739,N_32851);
or U35125 (N_35125,N_33163,N_32156);
and U35126 (N_35126,N_32318,N_31520);
or U35127 (N_35127,N_30207,N_30802);
xor U35128 (N_35128,N_32736,N_33551);
nand U35129 (N_35129,N_32996,N_34100);
nand U35130 (N_35130,N_31222,N_34846);
nand U35131 (N_35131,N_34352,N_33536);
nor U35132 (N_35132,N_34263,N_34409);
nand U35133 (N_35133,N_33116,N_30113);
or U35134 (N_35134,N_31945,N_34572);
nor U35135 (N_35135,N_34925,N_33034);
xnor U35136 (N_35136,N_30234,N_30480);
xnor U35137 (N_35137,N_34862,N_33591);
xnor U35138 (N_35138,N_32338,N_33914);
nand U35139 (N_35139,N_34700,N_30986);
or U35140 (N_35140,N_30855,N_33064);
nor U35141 (N_35141,N_30773,N_32852);
nor U35142 (N_35142,N_32023,N_30517);
and U35143 (N_35143,N_33569,N_30013);
and U35144 (N_35144,N_31503,N_34990);
xor U35145 (N_35145,N_32758,N_32369);
nor U35146 (N_35146,N_34179,N_30817);
nand U35147 (N_35147,N_30310,N_31071);
nand U35148 (N_35148,N_30301,N_33254);
nor U35149 (N_35149,N_33966,N_30116);
nand U35150 (N_35150,N_33639,N_32392);
nor U35151 (N_35151,N_31564,N_30616);
or U35152 (N_35152,N_31294,N_30371);
nor U35153 (N_35153,N_30612,N_34085);
nor U35154 (N_35154,N_31435,N_30068);
nand U35155 (N_35155,N_34086,N_31350);
nand U35156 (N_35156,N_33809,N_34093);
nand U35157 (N_35157,N_34771,N_31020);
or U35158 (N_35158,N_32164,N_32283);
nor U35159 (N_35159,N_30527,N_34946);
nand U35160 (N_35160,N_33260,N_34987);
or U35161 (N_35161,N_34767,N_33679);
xnor U35162 (N_35162,N_30705,N_33990);
nor U35163 (N_35163,N_34063,N_33315);
or U35164 (N_35164,N_30416,N_31745);
or U35165 (N_35165,N_32998,N_33152);
xor U35166 (N_35166,N_34644,N_32630);
nor U35167 (N_35167,N_33578,N_30968);
and U35168 (N_35168,N_31453,N_32811);
or U35169 (N_35169,N_30660,N_31779);
or U35170 (N_35170,N_34831,N_31061);
nor U35171 (N_35171,N_34981,N_31596);
and U35172 (N_35172,N_30085,N_31708);
or U35173 (N_35173,N_32123,N_32395);
xor U35174 (N_35174,N_30361,N_30436);
and U35175 (N_35175,N_30495,N_31527);
nor U35176 (N_35176,N_31507,N_32891);
xor U35177 (N_35177,N_34647,N_32965);
nor U35178 (N_35178,N_30141,N_31718);
nor U35179 (N_35179,N_30485,N_34960);
nand U35180 (N_35180,N_32401,N_30123);
and U35181 (N_35181,N_30339,N_34578);
xnor U35182 (N_35182,N_34806,N_31309);
nand U35183 (N_35183,N_30331,N_31894);
xnor U35184 (N_35184,N_33658,N_33935);
or U35185 (N_35185,N_32550,N_31163);
and U35186 (N_35186,N_33888,N_34429);
nand U35187 (N_35187,N_30282,N_30269);
xnor U35188 (N_35188,N_33166,N_33909);
nand U35189 (N_35189,N_33655,N_30720);
nor U35190 (N_35190,N_33594,N_33377);
nor U35191 (N_35191,N_34762,N_31143);
nand U35192 (N_35192,N_30906,N_31144);
xor U35193 (N_35193,N_31583,N_30506);
nor U35194 (N_35194,N_32586,N_34764);
or U35195 (N_35195,N_33013,N_34749);
nand U35196 (N_35196,N_33960,N_32211);
nor U35197 (N_35197,N_34356,N_34383);
nand U35198 (N_35198,N_34674,N_30019);
or U35199 (N_35199,N_32836,N_34339);
and U35200 (N_35200,N_31373,N_30613);
xnor U35201 (N_35201,N_30455,N_31855);
nand U35202 (N_35202,N_30468,N_34747);
nor U35203 (N_35203,N_33803,N_33024);
nand U35204 (N_35204,N_31614,N_30884);
or U35205 (N_35205,N_30121,N_30132);
nand U35206 (N_35206,N_33904,N_34114);
xnor U35207 (N_35207,N_34607,N_32091);
nor U35208 (N_35208,N_31050,N_33153);
and U35209 (N_35209,N_33155,N_32600);
or U35210 (N_35210,N_32964,N_30089);
nor U35211 (N_35211,N_34204,N_33656);
nand U35212 (N_35212,N_30335,N_32983);
nor U35213 (N_35213,N_31258,N_30062);
and U35214 (N_35214,N_34938,N_31290);
nor U35215 (N_35215,N_30907,N_31447);
xor U35216 (N_35216,N_33477,N_32070);
and U35217 (N_35217,N_31463,N_31553);
nand U35218 (N_35218,N_30771,N_33211);
or U35219 (N_35219,N_30425,N_33728);
nand U35220 (N_35220,N_32994,N_32124);
nor U35221 (N_35221,N_32393,N_31386);
nor U35222 (N_35222,N_32590,N_33417);
nor U35223 (N_35223,N_33647,N_32976);
xor U35224 (N_35224,N_33256,N_33409);
and U35225 (N_35225,N_34611,N_33036);
nand U35226 (N_35226,N_33158,N_31667);
and U35227 (N_35227,N_32405,N_31072);
xnor U35228 (N_35228,N_30553,N_30398);
and U35229 (N_35229,N_30904,N_33176);
nor U35230 (N_35230,N_30198,N_30251);
xor U35231 (N_35231,N_33644,N_32927);
xnor U35232 (N_35232,N_33747,N_33587);
nor U35233 (N_35233,N_33453,N_31248);
xor U35234 (N_35234,N_30411,N_34982);
nand U35235 (N_35235,N_32303,N_31103);
xor U35236 (N_35236,N_32737,N_31829);
or U35237 (N_35237,N_31366,N_31058);
xnor U35238 (N_35238,N_34354,N_33422);
nor U35239 (N_35239,N_30211,N_32892);
nand U35240 (N_35240,N_31873,N_33930);
and U35241 (N_35241,N_31774,N_32286);
nor U35242 (N_35242,N_34142,N_32247);
xor U35243 (N_35243,N_31000,N_34481);
nand U35244 (N_35244,N_31494,N_34408);
nand U35245 (N_35245,N_33666,N_32635);
nor U35246 (N_35246,N_34652,N_32198);
xor U35247 (N_35247,N_34673,N_30001);
and U35248 (N_35248,N_31339,N_34293);
xnor U35249 (N_35249,N_32439,N_31489);
xnor U35250 (N_35250,N_34817,N_30738);
nand U35251 (N_35251,N_34453,N_30639);
and U35252 (N_35252,N_30684,N_34335);
or U35253 (N_35253,N_34988,N_31152);
xor U35254 (N_35254,N_31915,N_34183);
and U35255 (N_35255,N_34504,N_34274);
and U35256 (N_35256,N_32033,N_34851);
nand U35257 (N_35257,N_31473,N_31198);
nand U35258 (N_35258,N_32833,N_31817);
or U35259 (N_35259,N_34560,N_34750);
nand U35260 (N_35260,N_31015,N_34103);
xnor U35261 (N_35261,N_34546,N_34048);
xnor U35262 (N_35262,N_32014,N_33600);
nand U35263 (N_35263,N_30432,N_31299);
nor U35264 (N_35264,N_30973,N_34096);
or U35265 (N_35265,N_34272,N_34108);
nand U35266 (N_35266,N_34455,N_33439);
nand U35267 (N_35267,N_32008,N_33817);
nor U35268 (N_35268,N_34963,N_31320);
nand U35269 (N_35269,N_33703,N_32116);
nand U35270 (N_35270,N_33942,N_34238);
xnor U35271 (N_35271,N_31977,N_34181);
nand U35272 (N_35272,N_33088,N_34182);
and U35273 (N_35273,N_32766,N_33227);
xnor U35274 (N_35274,N_34068,N_34614);
nor U35275 (N_35275,N_31726,N_30972);
and U35276 (N_35276,N_34235,N_31327);
nor U35277 (N_35277,N_31295,N_32088);
xor U35278 (N_35278,N_31452,N_34681);
nor U35279 (N_35279,N_33581,N_32784);
and U35280 (N_35280,N_32161,N_31095);
nor U35281 (N_35281,N_30831,N_33179);
nor U35282 (N_35282,N_31207,N_33623);
nand U35283 (N_35283,N_33225,N_33091);
xor U35284 (N_35284,N_31399,N_31037);
nor U35285 (N_35285,N_34878,N_34723);
and U35286 (N_35286,N_34402,N_31009);
nand U35287 (N_35287,N_33903,N_33702);
nand U35288 (N_35288,N_30084,N_32243);
and U35289 (N_35289,N_34378,N_33208);
nand U35290 (N_35290,N_30340,N_34853);
xnor U35291 (N_35291,N_30465,N_30325);
and U35292 (N_35292,N_34178,N_33740);
nand U35293 (N_35293,N_33418,N_34440);
or U35294 (N_35294,N_32954,N_34867);
nand U35295 (N_35295,N_30288,N_31690);
and U35296 (N_35296,N_33165,N_33607);
nand U35297 (N_35297,N_32856,N_30547);
nor U35298 (N_35298,N_33764,N_31303);
nor U35299 (N_35299,N_32263,N_33685);
or U35300 (N_35300,N_30775,N_32181);
or U35301 (N_35301,N_30515,N_30876);
or U35302 (N_35302,N_33533,N_32629);
and U35303 (N_35303,N_30015,N_31963);
xor U35304 (N_35304,N_32147,N_33508);
and U35305 (N_35305,N_32829,N_34168);
or U35306 (N_35306,N_30430,N_31785);
nor U35307 (N_35307,N_33854,N_33277);
nand U35308 (N_35308,N_34483,N_30063);
and U35309 (N_35309,N_30531,N_33366);
and U35310 (N_35310,N_33121,N_32020);
nor U35311 (N_35311,N_30192,N_34368);
nor U35312 (N_35312,N_32583,N_33449);
nor U35313 (N_35313,N_32894,N_31916);
xnor U35314 (N_35314,N_30588,N_34591);
nand U35315 (N_35315,N_33539,N_31574);
and U35316 (N_35316,N_32839,N_33057);
or U35317 (N_35317,N_34643,N_30179);
nand U35318 (N_35318,N_34194,N_33498);
nand U35319 (N_35319,N_31812,N_30112);
nor U35320 (N_35320,N_33312,N_32835);
xnor U35321 (N_35321,N_34242,N_33513);
and U35322 (N_35322,N_34506,N_31961);
or U35323 (N_35323,N_30471,N_32660);
or U35324 (N_35324,N_31467,N_32302);
xor U35325 (N_35325,N_34915,N_32577);
nor U35326 (N_35326,N_34474,N_31766);
and U35327 (N_35327,N_34195,N_32783);
or U35328 (N_35328,N_33995,N_34215);
and U35329 (N_35329,N_33721,N_33805);
nand U35330 (N_35330,N_34371,N_30208);
nor U35331 (N_35331,N_33185,N_31558);
and U35332 (N_35332,N_34733,N_30392);
and U35333 (N_35333,N_34002,N_30417);
xnor U35334 (N_35334,N_34830,N_31629);
or U35335 (N_35335,N_30434,N_30009);
xor U35336 (N_35336,N_32726,N_32676);
and U35337 (N_35337,N_33575,N_32472);
and U35338 (N_35338,N_33828,N_32978);
xnor U35339 (N_35339,N_30364,N_34797);
nand U35340 (N_35340,N_33813,N_33310);
nand U35341 (N_35341,N_31570,N_32196);
or U35342 (N_35342,N_33855,N_30841);
and U35343 (N_35343,N_31995,N_33124);
nor U35344 (N_35344,N_30628,N_31710);
xor U35345 (N_35345,N_33089,N_33856);
xor U35346 (N_35346,N_33577,N_34629);
nand U35347 (N_35347,N_31806,N_34230);
nor U35348 (N_35348,N_31657,N_31688);
nand U35349 (N_35349,N_33924,N_34174);
and U35350 (N_35350,N_34610,N_30136);
nand U35351 (N_35351,N_33654,N_33199);
and U35352 (N_35352,N_32499,N_33674);
nor U35353 (N_35353,N_30118,N_33328);
xnor U35354 (N_35354,N_30308,N_31665);
and U35355 (N_35355,N_30801,N_32666);
nor U35356 (N_35356,N_33457,N_31263);
and U35357 (N_35357,N_30691,N_33223);
nor U35358 (N_35358,N_30999,N_30663);
xor U35359 (N_35359,N_31707,N_31700);
xnor U35360 (N_35360,N_34985,N_33706);
nand U35361 (N_35361,N_33612,N_30885);
or U35362 (N_35362,N_31715,N_30212);
or U35363 (N_35363,N_33720,N_33290);
or U35364 (N_35364,N_34291,N_34296);
xnor U35365 (N_35365,N_31169,N_30679);
nor U35366 (N_35366,N_33000,N_34947);
or U35367 (N_35367,N_34734,N_32032);
and U35368 (N_35368,N_33992,N_32380);
and U35369 (N_35369,N_30444,N_31851);
or U35370 (N_35370,N_32645,N_34122);
nor U35371 (N_35371,N_31084,N_31981);
nand U35372 (N_35372,N_30038,N_32524);
nor U35373 (N_35373,N_33763,N_34869);
nand U35374 (N_35374,N_30776,N_34521);
or U35375 (N_35375,N_31150,N_33530);
nor U35376 (N_35376,N_33375,N_34881);
nand U35377 (N_35377,N_32937,N_34967);
nand U35378 (N_35378,N_31114,N_31346);
nand U35379 (N_35379,N_31156,N_32721);
nor U35380 (N_35380,N_30795,N_31846);
nor U35381 (N_35381,N_33120,N_31615);
or U35382 (N_35382,N_30095,N_30382);
or U35383 (N_35383,N_32001,N_32323);
nor U35384 (N_35384,N_33818,N_34285);
nand U35385 (N_35385,N_32554,N_30912);
or U35386 (N_35386,N_31862,N_30403);
xnor U35387 (N_35387,N_31027,N_31598);
or U35388 (N_35388,N_33963,N_32634);
nand U35389 (N_35389,N_34394,N_31278);
nor U35390 (N_35390,N_31039,N_34316);
nand U35391 (N_35391,N_32878,N_34787);
nand U35392 (N_35392,N_34860,N_32089);
and U35393 (N_35393,N_32804,N_33743);
nor U35394 (N_35394,N_33511,N_34101);
or U35395 (N_35395,N_34469,N_34702);
or U35396 (N_35396,N_32240,N_30175);
nor U35397 (N_35397,N_32368,N_34432);
and U35398 (N_35398,N_34426,N_34527);
and U35399 (N_35399,N_30466,N_32601);
nor U35400 (N_35400,N_30315,N_34739);
and U35401 (N_35401,N_31901,N_32970);
xor U35402 (N_35402,N_30291,N_34562);
nand U35403 (N_35403,N_33380,N_30094);
and U35404 (N_35404,N_31094,N_32188);
nand U35405 (N_35405,N_32742,N_34111);
nand U35406 (N_35406,N_33414,N_32867);
nor U35407 (N_35407,N_34328,N_33445);
nor U35408 (N_35408,N_33683,N_30564);
and U35409 (N_35409,N_31335,N_31651);
nand U35410 (N_35410,N_33500,N_34135);
nor U35411 (N_35411,N_33402,N_32534);
xor U35412 (N_35412,N_30263,N_34661);
or U35413 (N_35413,N_34015,N_32074);
nor U35414 (N_35414,N_31481,N_32604);
xnor U35415 (N_35415,N_32667,N_33460);
and U35416 (N_35416,N_34471,N_32253);
nor U35417 (N_35417,N_33907,N_30034);
and U35418 (N_35418,N_30213,N_33912);
or U35419 (N_35419,N_34510,N_32677);
nand U35420 (N_35420,N_34708,N_32987);
or U35421 (N_35421,N_33136,N_31940);
nand U35422 (N_35422,N_33020,N_34211);
nand U35423 (N_35423,N_30848,N_32636);
xnor U35424 (N_35424,N_33603,N_31815);
nor U35425 (N_35425,N_34253,N_32487);
and U35426 (N_35426,N_31750,N_32308);
or U35427 (N_35427,N_31045,N_34465);
and U35428 (N_35428,N_34698,N_33037);
and U35429 (N_35429,N_33363,N_34310);
nor U35430 (N_35430,N_32037,N_34978);
and U35431 (N_35431,N_32790,N_32771);
and U35432 (N_35432,N_34348,N_33394);
and U35433 (N_35433,N_31585,N_31983);
or U35434 (N_35434,N_32703,N_32704);
nor U35435 (N_35435,N_33219,N_32431);
nand U35436 (N_35436,N_34791,N_32481);
xor U35437 (N_35437,N_30488,N_30561);
xor U35438 (N_35438,N_32406,N_33985);
nand U35439 (N_35439,N_30701,N_30719);
nand U35440 (N_35440,N_31395,N_32426);
and U35441 (N_35441,N_33811,N_34013);
xor U35442 (N_35442,N_30276,N_30017);
and U35443 (N_35443,N_32767,N_31364);
and U35444 (N_35444,N_34199,N_30552);
xor U35445 (N_35445,N_34414,N_31017);
and U35446 (N_35446,N_31264,N_33301);
or U35447 (N_35447,N_32364,N_30459);
nand U35448 (N_35448,N_31259,N_30909);
xor U35449 (N_35449,N_30736,N_32933);
xnor U35450 (N_35450,N_34619,N_34294);
xor U35451 (N_35451,N_30900,N_32700);
or U35452 (N_35452,N_30474,N_34119);
xnor U35453 (N_35453,N_31459,N_30054);
and U35454 (N_35454,N_34362,N_31683);
and U35455 (N_35455,N_30750,N_31763);
xnor U35456 (N_35456,N_32238,N_34795);
or U35457 (N_35457,N_34456,N_31442);
nor U35458 (N_35458,N_33776,N_34950);
and U35459 (N_35459,N_34109,N_31099);
and U35460 (N_35460,N_32705,N_30565);
and U35461 (N_35461,N_30222,N_31405);
nor U35462 (N_35462,N_30400,N_33570);
xor U35463 (N_35463,N_30615,N_32476);
and U35464 (N_35464,N_32866,N_34924);
nand U35465 (N_35465,N_32496,N_31049);
nor U35466 (N_35466,N_34430,N_31110);
xnor U35467 (N_35467,N_34998,N_30717);
and U35468 (N_35468,N_33611,N_34569);
nand U35469 (N_35469,N_34609,N_33922);
xor U35470 (N_35470,N_34382,N_32419);
and U35471 (N_35471,N_33344,N_32789);
and U35472 (N_35472,N_34143,N_30862);
or U35473 (N_35473,N_30114,N_30933);
xor U35474 (N_35474,N_32776,N_33029);
nand U35475 (N_35475,N_34492,N_30209);
nor U35476 (N_35476,N_30693,N_31539);
nand U35477 (N_35477,N_32691,N_33780);
and U35478 (N_35478,N_34716,N_33172);
nor U35479 (N_35479,N_32669,N_34229);
nor U35480 (N_35480,N_33096,N_30818);
xnor U35481 (N_35481,N_30760,N_31853);
or U35482 (N_35482,N_33359,N_30868);
xor U35483 (N_35483,N_34177,N_30916);
nor U35484 (N_35484,N_33267,N_33845);
nand U35485 (N_35485,N_32265,N_33017);
or U35486 (N_35486,N_32077,N_34088);
nand U35487 (N_35487,N_34016,N_33040);
nor U35488 (N_35488,N_34014,N_32608);
nand U35489 (N_35489,N_34123,N_32919);
xnor U35490 (N_35490,N_30847,N_31474);
or U35491 (N_35491,N_32480,N_32174);
nand U35492 (N_35492,N_32528,N_31191);
or U35493 (N_35493,N_31944,N_34962);
nor U35494 (N_35494,N_30500,N_32162);
nor U35495 (N_35495,N_33693,N_32111);
or U35496 (N_35496,N_30169,N_30670);
xnor U35497 (N_35497,N_31559,N_33181);
or U35498 (N_35498,N_32735,N_30232);
nor U35499 (N_35499,N_33145,N_34668);
and U35500 (N_35500,N_34528,N_33392);
xnor U35501 (N_35501,N_33526,N_31286);
xor U35502 (N_35502,N_30835,N_31820);
nand U35503 (N_35503,N_32706,N_30934);
and U35504 (N_35504,N_32185,N_30388);
or U35505 (N_35505,N_34638,N_33291);
nand U35506 (N_35506,N_32548,N_31220);
and U35507 (N_35507,N_30477,N_31610);
and U35508 (N_35508,N_34582,N_34892);
nor U35509 (N_35509,N_32769,N_30324);
and U35510 (N_35510,N_34876,N_34137);
or U35511 (N_35511,N_33627,N_32026);
nor U35512 (N_35512,N_33565,N_33401);
nand U35513 (N_35513,N_32984,N_31550);
nand U35514 (N_35514,N_33475,N_34208);
or U35515 (N_35515,N_34520,N_30033);
and U35516 (N_35516,N_30600,N_32172);
and U35517 (N_35517,N_34872,N_30482);
or U35518 (N_35518,N_31795,N_34011);
nor U35519 (N_35519,N_32445,N_30077);
xnor U35520 (N_35520,N_31046,N_32837);
or U35521 (N_35521,N_34214,N_32307);
nor U35522 (N_35522,N_32873,N_33007);
nand U35523 (N_35523,N_31769,N_32948);
nor U35524 (N_35524,N_34247,N_32913);
or U35525 (N_35525,N_30936,N_32421);
nor U35526 (N_35526,N_33241,N_30772);
xor U35527 (N_35527,N_30022,N_31289);
nand U35528 (N_35528,N_34251,N_32202);
and U35529 (N_35529,N_33968,N_30953);
or U35530 (N_35530,N_30861,N_33258);
nand U35531 (N_35531,N_31390,N_33420);
and U35532 (N_35532,N_33791,N_34811);
and U35533 (N_35533,N_32112,N_34084);
nor U35534 (N_35534,N_33421,N_34000);
xor U35535 (N_35535,N_33848,N_31266);
nor U35536 (N_35536,N_34968,N_33978);
nor U35537 (N_35537,N_32025,N_33505);
nor U35538 (N_35538,N_33770,N_30437);
nand U35539 (N_35539,N_33188,N_30041);
nor U35540 (N_35540,N_34684,N_30740);
nor U35541 (N_35541,N_30607,N_32180);
xnor U35542 (N_35542,N_31880,N_33516);
and U35543 (N_35543,N_31348,N_32808);
xnor U35544 (N_35544,N_31954,N_31313);
xor U35545 (N_35545,N_34536,N_32661);
xor U35546 (N_35546,N_31256,N_30921);
or U35547 (N_35547,N_31361,N_33523);
and U35548 (N_35548,N_34841,N_31016);
or U35549 (N_35549,N_32201,N_32781);
or U35550 (N_35550,N_33846,N_32612);
and U35551 (N_35551,N_32093,N_32688);
xnor U35552 (N_35552,N_32567,N_31654);
xor U35553 (N_35553,N_34283,N_31560);
xor U35554 (N_35554,N_31407,N_33956);
nor U35555 (N_35555,N_34820,N_34566);
xnor U35556 (N_35556,N_33461,N_34544);
or U35557 (N_35557,N_34590,N_34167);
or U35558 (N_35558,N_30322,N_34255);
nand U35559 (N_35559,N_30568,N_30229);
or U35560 (N_35560,N_31599,N_31552);
xnor U35561 (N_35561,N_32598,N_32828);
nand U35562 (N_35562,N_33872,N_30521);
and U35563 (N_35563,N_31644,N_32969);
nand U35564 (N_35564,N_34326,N_30636);
or U35565 (N_35565,N_31077,N_31918);
nand U35566 (N_35566,N_33857,N_33387);
nand U35567 (N_35567,N_30035,N_33356);
or U35568 (N_35568,N_31404,N_33050);
and U35569 (N_35569,N_34252,N_32021);
and U35570 (N_35570,N_30306,N_33970);
nor U35571 (N_35571,N_31669,N_32379);
and U35572 (N_35572,N_34046,N_32489);
and U35573 (N_35573,N_32105,N_30592);
nand U35574 (N_35574,N_32078,N_33514);
nand U35575 (N_35575,N_30111,N_31907);
nor U35576 (N_35576,N_34152,N_33115);
and U35577 (N_35577,N_31336,N_30287);
xor U35578 (N_35578,N_34017,N_33370);
and U35579 (N_35579,N_31813,N_30744);
or U35580 (N_35580,N_33502,N_32786);
nand U35581 (N_35581,N_30487,N_33230);
nor U35582 (N_35582,N_33537,N_31768);
or U35583 (N_35583,N_31968,N_32324);
nor U35584 (N_35584,N_32017,N_34415);
nand U35585 (N_35585,N_30185,N_31764);
xor U35586 (N_35586,N_34508,N_30284);
nand U35587 (N_35587,N_32351,N_34006);
xnor U35588 (N_35588,N_34232,N_31419);
nand U35589 (N_35589,N_34439,N_34069);
nand U35590 (N_35590,N_33167,N_31003);
xor U35591 (N_35591,N_30014,N_34844);
nand U35592 (N_35592,N_34948,N_30181);
or U35593 (N_35593,N_31623,N_30991);
xnor U35594 (N_35594,N_31701,N_31048);
or U35595 (N_35595,N_30368,N_33519);
and U35596 (N_35596,N_32754,N_30573);
or U35597 (N_35597,N_32573,N_32119);
xnor U35598 (N_35598,N_32458,N_31311);
and U35599 (N_35599,N_34903,N_34443);
and U35600 (N_35600,N_34479,N_31092);
nand U35601 (N_35601,N_34212,N_32226);
or U35602 (N_35602,N_33795,N_32231);
nand U35603 (N_35603,N_33598,N_33060);
or U35604 (N_35604,N_33018,N_30575);
xor U35605 (N_35605,N_32215,N_32639);
nor U35606 (N_35606,N_33335,N_30313);
nand U35607 (N_35607,N_34956,N_30596);
and U35608 (N_35608,N_30641,N_34542);
or U35609 (N_35609,N_31988,N_32907);
nor U35610 (N_35610,N_32950,N_33682);
and U35611 (N_35611,N_33337,N_33562);
xnor U35612 (N_35612,N_33786,N_30273);
nor U35613 (N_35613,N_30714,N_31670);
nor U35614 (N_35614,N_30189,N_34838);
xor U35615 (N_35615,N_31328,N_31345);
nor U35616 (N_35616,N_30924,N_32287);
or U35617 (N_35617,N_31115,N_32407);
and U35618 (N_35618,N_31030,N_34337);
or U35619 (N_35619,N_30537,N_33512);
and U35620 (N_35620,N_30039,N_34980);
nand U35621 (N_35621,N_34269,N_30252);
xor U35622 (N_35622,N_32847,N_33014);
nor U35623 (N_35623,N_31171,N_30096);
and U35624 (N_35624,N_34038,N_34080);
nor U35625 (N_35625,N_33146,N_34450);
and U35626 (N_35626,N_34736,N_32755);
nand U35627 (N_35627,N_31960,N_34447);
xnor U35628 (N_35628,N_34390,N_30122);
and U35629 (N_35629,N_34540,N_31951);
nand U35630 (N_35630,N_30599,N_34117);
nand U35631 (N_35631,N_31857,N_31859);
nand U35632 (N_35632,N_30543,N_30621);
or U35633 (N_35633,N_31557,N_30275);
nor U35634 (N_35634,N_33792,N_33149);
or U35635 (N_35635,N_31436,N_31860);
or U35636 (N_35636,N_33474,N_32129);
and U35637 (N_35637,N_30117,N_30901);
or U35638 (N_35638,N_33712,N_32076);
nand U35639 (N_35639,N_33235,N_32578);
nor U35640 (N_35640,N_32291,N_32346);
xnor U35641 (N_35641,N_32497,N_31943);
xor U35642 (N_35642,N_30357,N_33454);
xnor U35643 (N_35643,N_33126,N_31751);
or U35644 (N_35644,N_32360,N_32473);
nor U35645 (N_35645,N_32544,N_34271);
or U35646 (N_35646,N_33999,N_31465);
and U35647 (N_35647,N_31786,N_34266);
nor U35648 (N_35648,N_32068,N_34670);
nand U35649 (N_35649,N_31979,N_34951);
or U35650 (N_35650,N_34320,N_33074);
nor U35651 (N_35651,N_32732,N_31160);
or U35652 (N_35652,N_30431,N_31424);
nand U35653 (N_35653,N_32424,N_32146);
or U35654 (N_35654,N_33710,N_30872);
and U35655 (N_35655,N_30511,N_31211);
or U35656 (N_35656,N_33098,N_32382);
nor U35657 (N_35657,N_34880,N_33285);
or U35658 (N_35658,N_31675,N_33698);
nor U35659 (N_35659,N_30704,N_33216);
and U35660 (N_35660,N_31931,N_31090);
nand U35661 (N_35661,N_32383,N_34989);
and U35662 (N_35662,N_32296,N_31650);
xnor U35663 (N_35663,N_31235,N_33299);
xor U35664 (N_35664,N_30332,N_30290);
or U35665 (N_35665,N_33419,N_32002);
and U35666 (N_35666,N_30808,N_34514);
xnor U35667 (N_35667,N_32814,N_30837);
nand U35668 (N_35668,N_31107,N_32988);
nand U35669 (N_35669,N_34267,N_33065);
nor U35670 (N_35670,N_33305,N_31370);
and U35671 (N_35671,N_34176,N_33503);
xnor U35672 (N_35672,N_31734,N_33396);
nand U35673 (N_35673,N_32535,N_34735);
nor U35674 (N_35674,N_33664,N_31261);
xnor U35675 (N_35675,N_32649,N_34417);
nor U35676 (N_35676,N_30302,N_33920);
xnor U35677 (N_35677,N_31306,N_31540);
xor U35678 (N_35678,N_31388,N_33535);
nand U35679 (N_35679,N_32515,N_34972);
xnor U35680 (N_35680,N_33362,N_33883);
nand U35681 (N_35681,N_30046,N_33642);
and U35682 (N_35682,N_34391,N_30522);
xnor U35683 (N_35683,N_31522,N_31976);
nor U35684 (N_35684,N_33247,N_30195);
nand U35685 (N_35685,N_31492,N_32222);
and U35686 (N_35686,N_33035,N_33183);
xor U35687 (N_35687,N_30097,N_32339);
or U35688 (N_35688,N_30938,N_33918);
and U35689 (N_35689,N_31555,N_32047);
xnor U35690 (N_35690,N_33651,N_32232);
or U35691 (N_35691,N_34323,N_31485);
xor U35692 (N_35692,N_31578,N_32605);
or U35693 (N_35693,N_34236,N_30093);
and U35694 (N_35694,N_30204,N_33885);
or U35695 (N_35695,N_32158,N_30354);
nand U35696 (N_35696,N_34125,N_31511);
nor U35697 (N_35697,N_33661,N_30066);
and U35698 (N_35698,N_34149,N_32144);
and U35699 (N_35699,N_33019,N_34387);
or U35700 (N_35700,N_31579,N_31875);
nand U35701 (N_35701,N_32641,N_31421);
xor U35702 (N_35702,N_30105,N_32513);
nor U35703 (N_35703,N_34489,N_34726);
nand U35704 (N_35704,N_31626,N_31930);
nor U35705 (N_35705,N_31638,N_30619);
or U35706 (N_35706,N_31797,N_30246);
xnor U35707 (N_35707,N_30268,N_34675);
nor U35708 (N_35708,N_30472,N_33033);
and U35709 (N_35709,N_30460,N_32761);
or U35710 (N_35710,N_34032,N_31087);
xor U35711 (N_35711,N_33774,N_33425);
nand U35712 (N_35712,N_32106,N_33933);
or U35713 (N_35713,N_31377,N_32991);
nor U35714 (N_35714,N_32084,N_32627);
nor U35715 (N_35715,N_33964,N_32224);
or U35716 (N_35716,N_31312,N_34003);
nor U35717 (N_35717,N_30629,N_33364);
or U35718 (N_35718,N_33708,N_31210);
nor U35719 (N_35719,N_33988,N_30554);
and U35720 (N_35720,N_32013,N_31450);
nand U35721 (N_35721,N_31997,N_30021);
nor U35722 (N_35722,N_31089,N_31323);
and U35723 (N_35723,N_31439,N_32367);
nor U35724 (N_35724,N_33972,N_32447);
and U35725 (N_35725,N_34778,N_31416);
xnor U35726 (N_35726,N_30752,N_32681);
nand U35727 (N_35727,N_31911,N_33605);
or U35728 (N_35728,N_32280,N_31184);
xnor U35729 (N_35729,N_30832,N_31518);
or U35730 (N_35730,N_34107,N_31254);
nand U35731 (N_35731,N_34669,N_33806);
nand U35732 (N_35732,N_32462,N_32207);
nor U35733 (N_35733,N_31508,N_34106);
nand U35734 (N_35734,N_31529,N_33379);
nand U35735 (N_35735,N_32505,N_32275);
xor U35736 (N_35736,N_34154,N_32571);
or U35737 (N_35737,N_33191,N_34319);
and U35738 (N_35738,N_33900,N_33713);
or U35739 (N_35739,N_33576,N_32532);
and U35740 (N_35740,N_33984,N_31592);
nand U35741 (N_35741,N_34602,N_34295);
xnor U35742 (N_35742,N_33411,N_31932);
nand U35743 (N_35743,N_32398,N_32155);
or U35744 (N_35744,N_34136,N_33015);
nand U35745 (N_35745,N_32936,N_30206);
nor U35746 (N_35746,N_31515,N_31561);
nor U35747 (N_35747,N_30373,N_30955);
or U35748 (N_35748,N_31532,N_32849);
or U35749 (N_35749,N_31839,N_30218);
and U35750 (N_35750,N_34513,N_31925);
nand U35751 (N_35751,N_30138,N_33117);
nor U35752 (N_35752,N_30215,N_31063);
nand U35753 (N_35753,N_34922,N_30721);
nand U35754 (N_35754,N_34009,N_30050);
or U35755 (N_35755,N_30974,N_33870);
or U35756 (N_35756,N_31136,N_30419);
and U35757 (N_35757,N_33424,N_34185);
and U35758 (N_35758,N_34970,N_33529);
or U35759 (N_35759,N_30700,N_33443);
or U35760 (N_35760,N_32173,N_30784);
nor U35761 (N_35761,N_30099,N_30966);
or U35762 (N_35762,N_32043,N_31133);
xnor U35763 (N_35763,N_31569,N_32132);
or U35764 (N_35764,N_32261,N_30957);
or U35765 (N_35765,N_34451,N_33341);
xnor U35766 (N_35766,N_31251,N_33160);
xor U35767 (N_35767,N_30076,N_33444);
xor U35768 (N_35768,N_34534,N_34343);
nor U35769 (N_35769,N_33292,N_34454);
nand U35770 (N_35770,N_32985,N_34040);
and U35771 (N_35771,N_33692,N_30260);
and U35772 (N_35772,N_31721,N_30669);
and U35773 (N_35773,N_30654,N_33090);
nand U35774 (N_35774,N_30632,N_30314);
or U35775 (N_35775,N_33571,N_33150);
or U35776 (N_35776,N_30450,N_34420);
nand U35777 (N_35777,N_32425,N_33351);
nand U35778 (N_35778,N_34418,N_32402);
or U35779 (N_35779,N_34931,N_31060);
nor U35780 (N_35780,N_34089,N_34507);
or U35781 (N_35781,N_34709,N_30871);
nor U35782 (N_35782,N_33525,N_34104);
nand U35783 (N_35783,N_33361,N_32582);
and U35784 (N_35784,N_31057,N_31018);
nor U35785 (N_35785,N_31281,N_34863);
or U35786 (N_35786,N_30000,N_32874);
nand U35787 (N_35787,N_31237,N_30798);
nand U35788 (N_35788,N_34834,N_30196);
nor U35789 (N_35789,N_31454,N_31186);
nor U35790 (N_35790,N_31257,N_33507);
xnor U35791 (N_35791,N_32945,N_31906);
nand U35792 (N_35792,N_32453,N_30086);
xnor U35793 (N_35793,N_33671,N_31677);
xor U35794 (N_35794,N_30969,N_32831);
and U35795 (N_35795,N_33808,N_34598);
or U35796 (N_35796,N_30372,N_34436);
and U35797 (N_35797,N_32918,N_33755);
xor U35798 (N_35798,N_34485,N_30800);
and U35799 (N_35799,N_32731,N_32748);
or U35800 (N_35800,N_34074,N_34784);
nand U35801 (N_35801,N_30984,N_33403);
or U35802 (N_35802,N_30739,N_31201);
nor U35803 (N_35803,N_30622,N_31491);
and U35804 (N_35804,N_30311,N_33601);
nor U35805 (N_35805,N_32536,N_33853);
nand U35806 (N_35806,N_30982,N_34498);
nand U35807 (N_35807,N_32166,N_31332);
and U35808 (N_35808,N_30741,N_32670);
or U35809 (N_35809,N_31028,N_32170);
nand U35810 (N_35810,N_31008,N_34871);
nor U35811 (N_35811,N_34225,N_30725);
or U35812 (N_35812,N_33249,N_33544);
or U35813 (N_35813,N_31272,N_34145);
nor U35814 (N_35814,N_34347,N_31711);
and U35815 (N_35815,N_31004,N_34503);
nand U35816 (N_35816,N_32809,N_31526);
xor U35817 (N_35817,N_34307,N_32038);
and U35818 (N_35818,N_33510,N_34034);
and U35819 (N_35819,N_32979,N_34132);
or U35820 (N_35820,N_34597,N_30520);
xnor U35821 (N_35821,N_31633,N_31032);
and U35822 (N_35822,N_30627,N_34761);
and U35823 (N_35823,N_34874,N_33787);
and U35824 (N_35824,N_32363,N_32625);
xnor U35825 (N_35825,N_33369,N_32744);
and U35826 (N_35826,N_32720,N_33358);
nor U35827 (N_35827,N_32273,N_32655);
or U35828 (N_35828,N_32067,N_31805);
or U35829 (N_35829,N_30389,N_32951);
nand U35830 (N_35830,N_33055,N_33404);
or U35831 (N_35831,N_31227,N_33031);
or U35832 (N_35832,N_31712,N_30281);
nor U35833 (N_35833,N_32603,N_30626);
xnor U35834 (N_35834,N_32659,N_33761);
nand U35835 (N_35835,N_31528,N_32467);
or U35836 (N_35836,N_31013,N_31819);
or U35837 (N_35837,N_32349,N_34688);
xor U35838 (N_35838,N_31922,N_32494);
and U35839 (N_35839,N_32819,N_31098);
nor U35840 (N_35840,N_34623,N_33971);
nand U35841 (N_35841,N_33592,N_30186);
nor U35842 (N_35842,N_33108,N_34091);
or U35843 (N_35843,N_30047,N_34911);
xor U35844 (N_35844,N_33038,N_33610);
nor U35845 (N_35845,N_33066,N_32062);
nor U35846 (N_35846,N_33428,N_34571);
xnor U35847 (N_35847,N_34551,N_30856);
nor U35848 (N_35848,N_31938,N_30454);
or U35849 (N_35849,N_32384,N_34711);
nand U35850 (N_35850,N_34303,N_30441);
nor U35851 (N_35851,N_32004,N_32355);
xor U35852 (N_35852,N_30271,N_33941);
and U35853 (N_35853,N_34497,N_32036);
or U35854 (N_35854,N_30692,N_30917);
xor U35855 (N_35855,N_33287,N_33874);
nor U35856 (N_35856,N_30226,N_34129);
or U35857 (N_35857,N_34741,N_34237);
xor U35858 (N_35858,N_31608,N_34188);
xor U35859 (N_35859,N_34786,N_30409);
nand U35860 (N_35860,N_31166,N_32250);
xor U35861 (N_35861,N_33459,N_34554);
xor U35862 (N_35862,N_33550,N_32225);
xor U35863 (N_35863,N_31800,N_33399);
nor U35864 (N_35864,N_34466,N_31652);
and U35865 (N_35865,N_30397,N_34836);
nand U35866 (N_35866,N_31342,N_34478);
or U35867 (N_35867,N_31267,N_31470);
nor U35868 (N_35868,N_30248,N_30699);
and U35869 (N_35869,N_31300,N_32484);
or U35870 (N_35870,N_30976,N_32335);
or U35871 (N_35871,N_30843,N_31367);
and U35872 (N_35872,N_34908,N_34877);
nor U35873 (N_35873,N_31921,N_33180);
xnor U35874 (N_35874,N_32685,N_32415);
or U35875 (N_35875,N_33481,N_33645);
xnor U35876 (N_35876,N_32566,N_31838);
nand U35877 (N_35877,N_30242,N_32103);
nor U35878 (N_35878,N_31804,N_30747);
nor U35879 (N_35879,N_31966,N_31139);
xor U35880 (N_35880,N_30620,N_34993);
nor U35881 (N_35881,N_33252,N_31268);
or U35882 (N_35882,N_34568,N_30778);
nor U35883 (N_35883,N_30223,N_34302);
or U35884 (N_35884,N_32827,N_33491);
nand U35885 (N_35885,N_30598,N_32632);
nor U35886 (N_35886,N_32518,N_34712);
xor U35887 (N_35887,N_33768,N_33168);
nor U35888 (N_35888,N_34099,N_34927);
nand U35889 (N_35889,N_31043,N_33925);
xor U35890 (N_35890,N_32297,N_31679);
xnor U35891 (N_35891,N_33324,N_33224);
or U35892 (N_35892,N_31537,N_32378);
xnor U35893 (N_35893,N_33296,N_31126);
nand U35894 (N_35894,N_34896,N_34662);
xnor U35895 (N_35895,N_33760,N_31239);
and U35896 (N_35896,N_33636,N_33892);
and U35897 (N_35897,N_34827,N_30298);
xor U35898 (N_35898,N_31044,N_30967);
nand U35899 (N_35899,N_31757,N_32656);
nor U35900 (N_35900,N_34943,N_34789);
nor U35901 (N_35901,N_34516,N_32187);
or U35902 (N_35902,N_32621,N_33906);
nand U35903 (N_35903,N_33450,N_31232);
xnor U35904 (N_35904,N_34539,N_30231);
or U35905 (N_35905,N_33083,N_32780);
and U35906 (N_35906,N_31912,N_32289);
or U35907 (N_35907,N_30142,N_34216);
or U35908 (N_35908,N_30493,N_30104);
nor U35909 (N_35909,N_33346,N_32079);
and U35910 (N_35910,N_34829,N_34163);
xnor U35911 (N_35911,N_34062,N_32785);
nor U35912 (N_35912,N_32968,N_34376);
nand U35913 (N_35913,N_34330,N_32024);
and U35914 (N_35914,N_33641,N_31502);
or U35915 (N_35915,N_34745,N_33415);
nand U35916 (N_35916,N_34150,N_30073);
nor U35917 (N_35917,N_33276,N_34024);
nor U35918 (N_35918,N_34861,N_30927);
or U35919 (N_35919,N_32876,N_34769);
and U35920 (N_35920,N_30366,N_31051);
xnor U35921 (N_35921,N_31939,N_30960);
nor U35922 (N_35922,N_34833,N_31024);
and U35923 (N_35923,N_34847,N_33833);
nand U35924 (N_35924,N_33723,N_34901);
and U35925 (N_35925,N_31113,N_32189);
nor U35926 (N_35926,N_32509,N_34939);
xor U35927 (N_35927,N_30059,N_30225);
xor U35928 (N_35928,N_34575,N_33100);
xor U35929 (N_35929,N_34545,N_32059);
nand U35930 (N_35930,N_33186,N_30556);
nor U35931 (N_35931,N_34777,N_32684);
nor U35932 (N_35932,N_30905,N_32353);
or U35933 (N_35933,N_31985,N_30935);
or U35934 (N_35934,N_34832,N_32657);
or U35935 (N_35935,N_33561,N_31192);
xor U35936 (N_35936,N_30582,N_30279);
xor U35937 (N_35937,N_34631,N_34913);
and U35938 (N_35938,N_32570,N_30749);
and U35939 (N_35939,N_32599,N_33549);
nand U35940 (N_35940,N_30178,N_31787);
or U35941 (N_35941,N_32561,N_31275);
nand U35942 (N_35942,N_31284,N_32589);
nor U35943 (N_35943,N_31243,N_30780);
or U35944 (N_35944,N_34315,N_32678);
or U35945 (N_35945,N_31206,N_32883);
nor U35946 (N_35946,N_30266,N_34190);
or U35947 (N_35947,N_34385,N_31112);
and U35948 (N_35948,N_33118,N_32643);
or U35949 (N_35949,N_34530,N_34775);
or U35950 (N_35950,N_33866,N_32197);
nand U35951 (N_35951,N_31767,N_34487);
nor U35952 (N_35952,N_33068,N_32179);
or U35953 (N_35953,N_33987,N_32908);
nand U35954 (N_35954,N_34217,N_33718);
or U35955 (N_35955,N_31040,N_33266);
or U35956 (N_35956,N_32714,N_32082);
nor U35957 (N_35957,N_31219,N_30894);
xor U35958 (N_35958,N_31488,N_34656);
and U35959 (N_35959,N_32693,N_34824);
nor U35960 (N_35960,N_33473,N_33973);
nor U35961 (N_35961,N_34025,N_33143);
and U35962 (N_35962,N_32136,N_32160);
or U35963 (N_35963,N_32167,N_33717);
xor U35964 (N_35964,N_30091,N_31920);
or U35965 (N_35965,N_30595,N_33197);
and U35966 (N_35966,N_30723,N_30623);
xor U35967 (N_35967,N_32348,N_32186);
and U35968 (N_35968,N_32482,N_34593);
and U35969 (N_35969,N_34585,N_33861);
nor U35970 (N_35970,N_33466,N_33470);
xor U35971 (N_35971,N_31130,N_34036);
nand U35972 (N_35972,N_31571,N_32097);
nand U35973 (N_35973,N_33727,N_31987);
nor U35974 (N_35974,N_31269,N_30353);
nor U35975 (N_35975,N_32654,N_30587);
nand U35976 (N_35976,N_33255,N_31432);
xor U35977 (N_35977,N_32734,N_31612);
and U35978 (N_35978,N_30563,N_30135);
and U35979 (N_35979,N_31562,N_32941);
or U35980 (N_35980,N_32503,N_34637);
xor U35981 (N_35981,N_32768,N_34626);
or U35982 (N_35982,N_30680,N_31542);
nand U35983 (N_35983,N_30731,N_34288);
nand U35984 (N_35984,N_31108,N_33590);
nand U35985 (N_35985,N_30697,N_31814);
nand U35986 (N_35986,N_32519,N_30386);
and U35987 (N_35987,N_32321,N_30931);
and U35988 (N_35988,N_32072,N_32728);
or U35989 (N_35989,N_32278,N_30708);
or U35990 (N_35990,N_33837,N_33558);
or U35991 (N_35991,N_33130,N_34092);
and U35992 (N_35992,N_32816,N_34687);
and U35993 (N_35993,N_32370,N_34366);
nand U35994 (N_35994,N_30662,N_34206);
xor U35995 (N_35995,N_34118,N_31741);
nor U35996 (N_35996,N_33119,N_33251);
or U35997 (N_35997,N_30951,N_30363);
nand U35998 (N_35998,N_32227,N_31890);
nand U35999 (N_35999,N_30814,N_32330);
nor U36000 (N_36000,N_32687,N_34961);
nor U36001 (N_36001,N_32863,N_32879);
xor U36002 (N_36002,N_32264,N_30737);
nand U36003 (N_36003,N_34792,N_32490);
or U36004 (N_36004,N_34097,N_30323);
nor U36005 (N_36005,N_31847,N_33733);
and U36006 (N_36006,N_34312,N_30558);
and U36007 (N_36007,N_32580,N_34810);
or U36008 (N_36008,N_31047,N_30249);
nor U36009 (N_36009,N_32889,N_34799);
and U36010 (N_36010,N_32410,N_34286);
or U36011 (N_36011,N_33412,N_32581);
or U36012 (N_36012,N_30236,N_32739);
or U36013 (N_36013,N_30959,N_32812);
or U36014 (N_36014,N_34393,N_31858);
nor U36015 (N_36015,N_34049,N_31881);
nor U36016 (N_36016,N_32165,N_32210);
nand U36017 (N_36017,N_31996,N_31825);
xnor U36018 (N_36018,N_32631,N_30519);
or U36019 (N_36019,N_34541,N_32995);
or U36020 (N_36020,N_33954,N_33729);
and U36021 (N_36021,N_33075,N_31120);
or U36022 (N_36022,N_31400,N_30645);
and U36023 (N_36023,N_30689,N_34297);
xor U36024 (N_36024,N_30140,N_34798);
and U36025 (N_36025,N_32971,N_31713);
xnor U36026 (N_36026,N_34054,N_30002);
nand U36027 (N_36027,N_34278,N_33814);
or U36028 (N_36028,N_31903,N_34133);
nor U36029 (N_36029,N_31310,N_32585);
nor U36030 (N_36030,N_33495,N_34580);
or U36031 (N_36031,N_32798,N_31141);
and U36032 (N_36032,N_30792,N_34796);
xnor U36033 (N_36033,N_33011,N_31178);
and U36034 (N_36034,N_33371,N_31196);
nor U36035 (N_36035,N_30637,N_33840);
or U36036 (N_36036,N_30915,N_32861);
nand U36037 (N_36037,N_30024,N_30709);
xnor U36038 (N_36038,N_33742,N_33901);
and U36039 (N_36039,N_32388,N_30274);
and U36040 (N_36040,N_34357,N_31709);
nand U36041 (N_36041,N_31189,N_31755);
nand U36042 (N_36042,N_30447,N_30952);
xnor U36043 (N_36043,N_31716,N_32525);
nor U36044 (N_36044,N_30404,N_30648);
xnor U36045 (N_36045,N_31005,N_34891);
and U36046 (N_36046,N_32329,N_33758);
and U36047 (N_36047,N_33884,N_31869);
nand U36048 (N_36048,N_30442,N_33711);
nand U36049 (N_36049,N_34694,N_34589);
xor U36050 (N_36050,N_32150,N_33735);
xnor U36051 (N_36051,N_32343,N_33297);
or U36052 (N_36052,N_34547,N_30548);
nor U36053 (N_36053,N_32797,N_33239);
and U36054 (N_36054,N_32018,N_30401);
nor U36055 (N_36055,N_30794,N_33916);
xnor U36056 (N_36056,N_32233,N_34992);
or U36057 (N_36057,N_34121,N_34373);
nor U36058 (N_36058,N_34030,N_30702);
or U36059 (N_36059,N_30793,N_31316);
nor U36060 (N_36060,N_33701,N_32841);
or U36061 (N_36061,N_34052,N_34813);
or U36062 (N_36062,N_31607,N_32775);
or U36063 (N_36063,N_32690,N_34139);
nor U36064 (N_36064,N_32375,N_34588);
and U36065 (N_36065,N_34917,N_30473);
xor U36066 (N_36066,N_31867,N_32747);
nand U36067 (N_36067,N_30829,N_32868);
nand U36068 (N_36068,N_32763,N_33939);
or U36069 (N_36069,N_30421,N_33739);
and U36070 (N_36070,N_32902,N_32299);
nand U36071 (N_36071,N_32795,N_33940);
nand U36072 (N_36072,N_34120,N_33556);
nor U36073 (N_36073,N_30075,N_30745);
nor U36074 (N_36074,N_31451,N_33433);
or U36075 (N_36075,N_34535,N_31426);
or U36076 (N_36076,N_34077,N_34642);
nand U36077 (N_36077,N_34160,N_32750);
nand U36078 (N_36078,N_34164,N_31414);
or U36079 (N_36079,N_31601,N_31205);
xor U36080 (N_36080,N_34894,N_31318);
nor U36081 (N_36081,N_33196,N_33262);
and U36082 (N_36082,N_33215,N_34567);
nand U36083 (N_36083,N_33567,N_33316);
nand U36084 (N_36084,N_33699,N_32564);
or U36085 (N_36085,N_33949,N_33151);
nor U36086 (N_36086,N_32900,N_33648);
xnor U36087 (N_36087,N_34971,N_33958);
nand U36088 (N_36088,N_34452,N_34620);
nor U36089 (N_36089,N_34389,N_31673);
xnor U36090 (N_36090,N_32822,N_33672);
xnor U36091 (N_36091,N_30594,N_32824);
and U36092 (N_36092,N_33799,N_30644);
nand U36093 (N_36093,N_30678,N_32593);
nand U36094 (N_36094,N_34500,N_31699);
xnor U36095 (N_36095,N_34144,N_32504);
nand U36096 (N_36096,N_31487,N_34933);
nand U36097 (N_36097,N_34715,N_30193);
xor U36098 (N_36098,N_33869,N_31479);
xnor U36099 (N_36099,N_33182,N_34401);
nor U36100 (N_36100,N_30228,N_32127);
xnor U36101 (N_36101,N_31754,N_34628);
nand U36102 (N_36102,N_33480,N_34493);
nor U36103 (N_36103,N_34949,N_32099);
or U36104 (N_36104,N_34367,N_32374);
nor U36105 (N_36105,N_32594,N_33464);
xnor U36106 (N_36106,N_30634,N_32607);
or U36107 (N_36107,N_33110,N_32294);
and U36108 (N_36108,N_30341,N_32290);
nor U36109 (N_36109,N_33093,N_32543);
or U36110 (N_36110,N_34299,N_31440);
or U36111 (N_36111,N_32141,N_31212);
nand U36112 (N_36112,N_34318,N_34584);
nor U36113 (N_36113,N_34445,N_32456);
xor U36114 (N_36114,N_32357,N_31832);
and U36115 (N_36115,N_32800,N_34044);
and U36116 (N_36116,N_30542,N_34573);
or U36117 (N_36117,N_30005,N_32390);
nand U36118 (N_36118,N_32376,N_30133);
or U36119 (N_36119,N_31697,N_31225);
or U36120 (N_36120,N_33962,N_33993);
xnor U36121 (N_36121,N_32905,N_32501);
nand U36122 (N_36122,N_34837,N_34753);
nand U36123 (N_36123,N_34416,N_30807);
nand U36124 (N_36124,N_30457,N_31934);
or U36125 (N_36125,N_32016,N_33634);
or U36126 (N_36126,N_31606,N_32134);
xor U36127 (N_36127,N_34365,N_33423);
nand U36128 (N_36128,N_30219,N_33482);
nor U36129 (N_36129,N_34854,N_30067);
and U36130 (N_36130,N_31933,N_34718);
nand U36131 (N_36131,N_33009,N_31866);
nor U36132 (N_36132,N_33348,N_31478);
nor U36133 (N_36133,N_33012,N_33927);
and U36134 (N_36134,N_32075,N_30860);
xor U36135 (N_36135,N_33826,N_33095);
or U36136 (N_36136,N_31127,N_33052);
xnor U36137 (N_36137,N_31567,N_33847);
nand U36138 (N_36138,N_33321,N_33094);
or U36139 (N_36139,N_32917,N_30601);
nand U36140 (N_36140,N_30890,N_34529);
nand U36141 (N_36141,N_31079,N_31315);
nand U36142 (N_36142,N_33339,N_30283);
or U36143 (N_36143,N_31337,N_31218);
or U36144 (N_36144,N_34442,N_30796);
or U36145 (N_36145,N_31531,N_30502);
or U36146 (N_36146,N_30985,N_33139);
or U36147 (N_36147,N_30414,N_30845);
nand U36148 (N_36148,N_34689,N_30661);
nor U36149 (N_36149,N_33232,N_34189);
xor U36150 (N_36150,N_32045,N_31282);
nor U36151 (N_36151,N_33367,N_32314);
nand U36152 (N_36152,N_30821,N_32881);
and U36153 (N_36153,N_34333,N_31100);
nor U36154 (N_36154,N_30690,N_30813);
nand U36155 (N_36155,N_33067,N_31197);
nand U36156 (N_36156,N_30703,N_32279);
nand U36157 (N_36157,N_33800,N_33056);
xor U36158 (N_36158,N_34460,N_30498);
or U36159 (N_36159,N_30677,N_34648);
and U36160 (N_36160,N_34966,N_32095);
or U36161 (N_36161,N_33785,N_33109);
xnor U36162 (N_36162,N_32588,N_33546);
xnor U36163 (N_36163,N_33345,N_32394);
nor U36164 (N_36164,N_34803,N_33585);
and U36165 (N_36165,N_30675,N_33676);
nand U36166 (N_36166,N_33400,N_33579);
nand U36167 (N_36167,N_31674,N_34553);
xnor U36168 (N_36168,N_34705,N_30706);
or U36169 (N_36169,N_34850,N_31889);
nand U36170 (N_36170,N_31277,N_30559);
nor U36171 (N_36171,N_31456,N_30589);
nor U36172 (N_36172,N_32052,N_32526);
or U36173 (N_36173,N_30880,N_32262);
xnor U36174 (N_36174,N_34035,N_33289);
xnor U36175 (N_36175,N_32228,N_34220);
nand U36176 (N_36176,N_33114,N_33838);
nor U36177 (N_36177,N_31410,N_33782);
nand U36178 (N_36178,N_30305,N_30391);
and U36179 (N_36179,N_31068,N_32203);
xor U36180 (N_36180,N_31872,N_34957);
nor U36181 (N_36181,N_30058,N_32448);
nand U36182 (N_36182,N_31969,N_32056);
and U36183 (N_36183,N_34219,N_32042);
xor U36184 (N_36184,N_32966,N_30197);
xor U36185 (N_36185,N_31826,N_31462);
xor U36186 (N_36186,N_33675,N_32316);
and U36187 (N_36187,N_30867,N_33669);
or U36188 (N_36188,N_32730,N_31394);
xor U36189 (N_36189,N_34351,N_32010);
xor U36190 (N_36190,N_34298,N_34210);
or U36191 (N_36191,N_34170,N_31664);
nor U36192 (N_36192,N_32350,N_30443);
or U36193 (N_36193,N_33132,N_33250);
nor U36194 (N_36194,N_30756,N_32759);
nand U36195 (N_36195,N_34748,N_31671);
or U36196 (N_36196,N_34494,N_31923);
nor U36197 (N_36197,N_31761,N_34845);
and U36198 (N_36198,N_30253,N_31538);
nor U36199 (N_36199,N_32411,N_33269);
nor U36200 (N_36200,N_34983,N_30646);
nand U36201 (N_36201,N_34279,N_32904);
nor U36202 (N_36202,N_30028,N_30385);
and U36203 (N_36203,N_30633,N_32269);
and U36204 (N_36204,N_31285,N_31265);
nand U36205 (N_36205,N_33282,N_33983);
nand U36206 (N_36206,N_34234,N_30106);
nand U36207 (N_36207,N_32765,N_34515);
nand U36208 (N_36208,N_31209,N_31014);
nand U36209 (N_36209,N_33494,N_32722);
or U36210 (N_36210,N_33395,N_34256);
nor U36211 (N_36211,N_32626,N_32115);
and U36212 (N_36212,N_34321,N_31666);
xor U36213 (N_36213,N_33810,N_33391);
nand U36214 (N_36214,N_30635,N_33112);
nand U36215 (N_36215,N_31314,N_33002);
xnor U36216 (N_36216,N_33408,N_34060);
nor U36217 (N_36217,N_31180,N_32793);
xnor U36218 (N_36218,N_32772,N_33552);
nor U36219 (N_36219,N_33829,N_34361);
nor U36220 (N_36220,N_34231,N_31497);
nand U36221 (N_36221,N_30755,N_32743);
xor U36222 (N_36222,N_33583,N_31355);
xnor U36223 (N_36223,N_33084,N_30048);
nor U36224 (N_36224,N_31882,N_33628);
xnor U36225 (N_36225,N_30593,N_33730);
xnor U36226 (N_36226,N_33621,N_31689);
nand U36227 (N_36227,N_31992,N_31398);
or U36228 (N_36228,N_33051,N_33864);
and U36229 (N_36229,N_30541,N_33705);
and U36230 (N_36230,N_32568,N_32328);
and U36231 (N_36231,N_33427,N_31157);
and U36232 (N_36232,N_30789,N_32365);
or U36233 (N_36233,N_33694,N_34991);
and U36234 (N_36234,N_30394,N_32417);
xnor U36235 (N_36235,N_32268,N_31119);
and U36236 (N_36236,N_30922,N_34770);
nor U36237 (N_36237,N_30962,N_32151);
xor U36238 (N_36238,N_34166,N_33609);
and U36239 (N_36239,N_30505,N_31547);
xor U36240 (N_36240,N_33314,N_32443);
nor U36241 (N_36241,N_33905,N_32061);
nand U36242 (N_36242,N_32428,N_33355);
or U36243 (N_36243,N_31756,N_30823);
or U36244 (N_36244,N_32159,N_31307);
nor U36245 (N_36245,N_34738,N_30524);
nor U36246 (N_36246,N_33478,N_30151);
or U36247 (N_36247,N_31927,N_32064);
and U36248 (N_36248,N_30345,N_30523);
or U36249 (N_36249,N_32183,N_30891);
xnor U36250 (N_36250,N_30647,N_33951);
and U36251 (N_36251,N_33878,N_32521);
and U36252 (N_36252,N_32587,N_34277);
and U36253 (N_36253,N_33881,N_32888);
xor U36254 (N_36254,N_32400,N_34691);
or U36255 (N_36255,N_34997,N_31466);
nor U36256 (N_36256,N_33522,N_31573);
and U36257 (N_36257,N_30926,N_34410);
nor U36258 (N_36258,N_32576,N_32309);
nand U36259 (N_36259,N_31102,N_34677);
and U36260 (N_36260,N_32549,N_34828);
xnor U36261 (N_36261,N_30715,N_30947);
xnor U36262 (N_36262,N_32946,N_33691);
or U36263 (N_36263,N_34816,N_31841);
and U36264 (N_36264,N_33238,N_33311);
xor U36265 (N_36265,N_33410,N_33841);
or U36266 (N_36266,N_30763,N_31519);
xnor U36267 (N_36267,N_30803,N_33746);
and U36268 (N_36268,N_31837,N_33959);
and U36269 (N_36269,N_31007,N_30227);
nand U36270 (N_36270,N_33520,N_31134);
or U36271 (N_36271,N_30486,N_32306);
xnor U36272 (N_36272,N_30149,N_32171);
and U36273 (N_36273,N_30214,N_34888);
nand U36274 (N_36274,N_33557,N_34549);
or U36275 (N_36275,N_33416,N_32044);
or U36276 (N_36276,N_30649,N_34467);
or U36277 (N_36277,N_30535,N_34977);
xor U36278 (N_36278,N_33781,N_34842);
nand U36279 (N_36279,N_33039,N_30614);
nor U36280 (N_36280,N_33071,N_32391);
xor U36281 (N_36281,N_32897,N_31338);
nor U36282 (N_36282,N_31770,N_31978);
or U36283 (N_36283,N_33101,N_34843);
nor U36284 (N_36284,N_33144,N_30851);
and U36285 (N_36285,N_32366,N_31947);
xnor U36286 (N_36286,N_31658,N_31012);
xnor U36287 (N_36287,N_31413,N_34592);
nor U36288 (N_36288,N_30940,N_34785);
and U36289 (N_36289,N_31618,N_31131);
nor U36290 (N_36290,N_33073,N_31941);
xnor U36291 (N_36291,N_30674,N_30840);
nand U36292 (N_36292,N_33278,N_30510);
xor U36293 (N_36293,N_30979,N_31428);
and U36294 (N_36294,N_30611,N_33131);
nand U36295 (N_36295,N_34505,N_34654);
and U36296 (N_36296,N_31190,N_33923);
nor U36297 (N_36297,N_31946,N_30903);
nor U36298 (N_36298,N_33967,N_32449);
and U36299 (N_36299,N_31329,N_32514);
nor U36300 (N_36300,N_34158,N_31403);
or U36301 (N_36301,N_30895,N_31187);
or U36302 (N_36302,N_34634,N_32011);
or U36303 (N_36303,N_33240,N_33431);
nor U36304 (N_36304,N_30724,N_31659);
nor U36305 (N_36305,N_31449,N_34147);
and U36306 (N_36306,N_34576,N_30412);
nor U36307 (N_36307,N_30201,N_33229);
and U36308 (N_36308,N_30299,N_34375);
nor U36309 (N_36309,N_32474,N_32485);
nor U36310 (N_36310,N_32414,N_31236);
nor U36311 (N_36311,N_32493,N_33080);
xor U36312 (N_36312,N_30846,N_31333);
xnor U36313 (N_36313,N_32711,N_31412);
xnor U36314 (N_36314,N_31584,N_30819);
xnor U36315 (N_36315,N_33802,N_30349);
or U36316 (N_36316,N_30052,N_31999);
nor U36317 (N_36317,N_33242,N_34875);
nand U36318 (N_36318,N_34898,N_34273);
xnor U36319 (N_36319,N_33398,N_30475);
nand U36320 (N_36320,N_33293,N_33372);
nand U36321 (N_36321,N_33497,N_32609);
nand U36322 (N_36322,N_33357,N_30828);
nand U36323 (N_36323,N_32574,N_30869);
xnor U36324 (N_36324,N_33243,N_31678);
and U36325 (N_36325,N_34519,N_31213);
nor U36326 (N_36326,N_32606,N_31182);
and U36327 (N_36327,N_34973,N_31493);
or U36328 (N_36328,N_32488,N_33122);
nand U36329 (N_36329,N_34055,N_32960);
or U36330 (N_36330,N_33082,N_30277);
nand U36331 (N_36331,N_32470,N_32145);
nand U36332 (N_36332,N_33738,N_31958);
nor U36333 (N_36333,N_31789,N_30950);
xnor U36334 (N_36334,N_34403,N_32377);
nand U36335 (N_36335,N_32925,N_31125);
nor U36336 (N_36336,N_33061,N_30082);
nor U36337 (N_36337,N_34794,N_31590);
and U36338 (N_36338,N_32563,N_32386);
nand U36339 (N_36339,N_31111,N_33378);
nand U36340 (N_36340,N_32860,N_30852);
nor U36341 (N_36341,N_31059,N_34690);
nand U36342 (N_36342,N_31056,N_34495);
and U36343 (N_36343,N_33313,N_30285);
xor U36344 (N_36344,N_34411,N_31776);
nor U36345 (N_36345,N_31929,N_33385);
nor U36346 (N_36346,N_34682,N_33054);
and U36347 (N_36347,N_32972,N_31054);
xor U36348 (N_36348,N_33946,N_30584);
or U36349 (N_36349,N_32807,N_31188);
and U36350 (N_36350,N_32341,N_31572);
nand U36351 (N_36351,N_33456,N_34517);
nor U36352 (N_36352,N_33463,N_30359);
or U36353 (N_36353,N_31738,N_32455);
or U36354 (N_36354,N_33004,N_30825);
nor U36355 (N_36355,N_33678,N_30458);
and U36356 (N_36356,N_30638,N_32371);
and U36357 (N_36357,N_33022,N_34280);
nor U36358 (N_36358,N_31296,N_30057);
nand U36359 (N_36359,N_34532,N_32915);
nand U36360 (N_36360,N_32545,N_34399);
nor U36361 (N_36361,N_34340,N_31383);
xnor U36362 (N_36362,N_33347,N_34757);
xor U36363 (N_36363,N_31655,N_34201);
nor U36364 (N_36364,N_30102,N_32592);
nor U36365 (N_36365,N_30892,N_30791);
and U36366 (N_36366,N_30307,N_31854);
and U36367 (N_36367,N_31956,N_32903);
and U36368 (N_36368,N_33484,N_30145);
or U36369 (N_36369,N_31748,N_30037);
or U36370 (N_36370,N_31397,N_32096);
nand U36371 (N_36371,N_33193,N_34022);
nand U36372 (N_36372,N_30602,N_31899);
and U36373 (N_36373,N_34565,N_34857);
or U36374 (N_36374,N_30220,N_33638);
or U36375 (N_36375,N_33270,N_34552);
or U36376 (N_36376,N_33509,N_31687);
and U36377 (N_36377,N_30087,N_31611);
nand U36378 (N_36378,N_33129,N_30604);
and U36379 (N_36379,N_30446,N_33908);
nand U36380 (N_36380,N_34923,N_34550);
nand U36381 (N_36381,N_32469,N_31672);
and U36382 (N_36382,N_31340,N_32799);
nand U36383 (N_36383,N_31807,N_33629);
and U36384 (N_36384,N_32595,N_34622);
or U36385 (N_36385,N_34918,N_33327);
xor U36386 (N_36386,N_32208,N_32140);
nand U36387 (N_36387,N_30156,N_34324);
nand U36388 (N_36388,N_32178,N_34477);
nand U36389 (N_36389,N_31223,N_33862);
xnor U36390 (N_36390,N_32751,N_30481);
xnor U36391 (N_36391,N_33261,N_30119);
or U36392 (N_36392,N_32332,N_34929);
nand U36393 (N_36393,N_32943,N_33111);
nand U36394 (N_36394,N_34358,N_32257);
nor U36395 (N_36395,N_33157,N_33566);
and U36396 (N_36396,N_30888,N_32081);
xor U36397 (N_36397,N_31509,N_32334);
nor U36398 (N_36398,N_32774,N_30810);
xor U36399 (N_36399,N_32031,N_31600);
nand U36400 (N_36400,N_34083,N_33769);
and U36401 (N_36401,N_34953,N_32149);
xor U36402 (N_36402,N_34729,N_32312);
or U36403 (N_36403,N_30157,N_32663);
xor U36404 (N_36404,N_32154,N_32885);
nor U36405 (N_36405,N_30045,N_32664);
nor U36406 (N_36406,N_30879,N_32542);
or U36407 (N_36407,N_30914,N_31304);
or U36408 (N_36408,N_33053,N_30320);
xnor U36409 (N_36409,N_33643,N_32858);
xor U36410 (N_36410,N_34459,N_30303);
or U36411 (N_36411,N_30173,N_32541);
nor U36412 (N_36412,N_33944,N_32846);
and U36413 (N_36413,N_34935,N_34600);
xnor U36414 (N_36414,N_30420,N_30534);
or U36415 (N_36415,N_32591,N_34804);
and U36416 (N_36416,N_31288,N_33759);
nand U36417 (N_36417,N_31810,N_33602);
or U36418 (N_36418,N_34912,N_32175);
and U36419 (N_36419,N_32551,N_32342);
nor U36420 (N_36420,N_34783,N_30777);
or U36421 (N_36421,N_33842,N_32665);
nor U36422 (N_36422,N_31772,N_31705);
xnor U36423 (N_36423,N_32094,N_30978);
nor U36424 (N_36424,N_31226,N_31434);
nand U36425 (N_36425,N_31480,N_32327);
and U36426 (N_36426,N_34486,N_32244);
or U36427 (N_36427,N_34161,N_34404);
nor U36428 (N_36428,N_30247,N_33652);
or U36429 (N_36429,N_33955,N_32779);
xor U36430 (N_36430,N_32646,N_33680);
nor U36431 (N_36431,N_33662,N_30428);
nand U36432 (N_36432,N_32650,N_31123);
nand U36433 (N_36433,N_31780,N_32492);
nor U36434 (N_36434,N_31775,N_34257);
nand U36435 (N_36435,N_34172,N_33426);
or U36436 (N_36436,N_31917,N_31011);
and U36437 (N_36437,N_34329,N_34005);
nand U36438 (N_36438,N_32875,N_31140);
and U36439 (N_36439,N_32850,N_33796);
or U36440 (N_36440,N_32420,N_30146);
and U36441 (N_36441,N_34012,N_31777);
xor U36442 (N_36442,N_30490,N_33989);
xnor U36443 (N_36443,N_33653,N_31381);
or U36444 (N_36444,N_31914,N_30624);
nand U36445 (N_36445,N_31778,N_30574);
nor U36446 (N_36446,N_30134,N_32475);
and U36447 (N_36447,N_30923,N_31001);
nor U36448 (N_36448,N_32944,N_30147);
and U36449 (N_36449,N_30866,N_33295);
or U36450 (N_36450,N_32128,N_30280);
xnor U36451 (N_36451,N_33023,N_33894);
xor U36452 (N_36452,N_33586,N_30304);
or U36453 (N_36453,N_33205,N_30897);
and U36454 (N_36454,N_30766,N_30381);
nand U36455 (N_36455,N_30255,N_32613);
nand U36456 (N_36456,N_32980,N_31471);
or U36457 (N_36457,N_31593,N_31230);
nand U36458 (N_36458,N_34522,N_30090);
and U36459 (N_36459,N_33798,N_33619);
nand U36460 (N_36460,N_32910,N_34889);
nand U36461 (N_36461,N_32319,N_31255);
or U36462 (N_36462,N_33919,N_31026);
nor U36463 (N_36463,N_31950,N_34900);
and U36464 (N_36464,N_32418,N_31161);
or U36465 (N_36465,N_33871,N_34524);
or U36466 (N_36466,N_34484,N_33911);
nor U36467 (N_36467,N_34223,N_32372);
nand U36468 (N_36468,N_31117,N_33430);
xor U36469 (N_36469,N_34400,N_32637);
nor U36470 (N_36470,N_31605,N_33030);
and U36471 (N_36471,N_32715,N_34543);
xor U36472 (N_36472,N_30570,N_33490);
nor U36473 (N_36473,N_32213,N_30127);
or U36474 (N_36474,N_32454,N_34309);
and U36475 (N_36475,N_34722,N_30822);
or U36476 (N_36476,N_33595,N_34790);
nand U36477 (N_36477,N_33340,N_33329);
xnor U36478 (N_36478,N_31076,N_33783);
nor U36479 (N_36479,N_31506,N_33630);
nand U36480 (N_36480,N_32464,N_32617);
nand U36481 (N_36481,N_31498,N_34814);
xor U36482 (N_36482,N_34425,N_31085);
nor U36483 (N_36483,N_33025,N_33170);
or U36484 (N_36484,N_31704,N_34680);
or U36485 (N_36485,N_30439,N_34937);
or U36486 (N_36486,N_32683,N_32085);
nor U36487 (N_36487,N_33338,N_33722);
nor U36488 (N_36488,N_31896,N_34751);
xor U36489 (N_36489,N_32483,N_33103);
and U36490 (N_36490,N_33599,N_34370);
or U36491 (N_36491,N_33407,N_32832);
or U36492 (N_36492,N_30569,N_30948);
or U36493 (N_36493,N_30461,N_33898);
nor U36494 (N_36494,N_32252,N_30023);
and U36495 (N_36495,N_33532,N_33640);
or U36496 (N_36496,N_32163,N_32152);
nand U36497 (N_36497,N_31864,N_33637);
or U36498 (N_36498,N_34608,N_33937);
xor U36499 (N_36499,N_32101,N_34113);
and U36500 (N_36500,N_30153,N_34423);
and U36501 (N_36501,N_30469,N_34380);
nand U36502 (N_36502,N_30812,N_32757);
or U36503 (N_36503,N_32624,N_32975);
xor U36504 (N_36504,N_31183,N_34258);
nor U36505 (N_36505,N_30360,N_30571);
or U36506 (N_36506,N_30378,N_31962);
nand U36507 (N_36507,N_32928,N_31953);
or U36508 (N_36508,N_34322,N_30464);
and U36509 (N_36509,N_30566,N_33812);
nand U36510 (N_36510,N_33354,N_30098);
or U36511 (N_36511,N_34559,N_31472);
or U36512 (N_36512,N_32479,N_30964);
or U36513 (N_36513,N_32826,N_31913);
nor U36514 (N_36514,N_31234,N_32708);
or U36515 (N_36515,N_34087,N_30358);
or U36516 (N_36516,N_30467,N_30734);
nor U36517 (N_36517,N_32569,N_34317);
xnor U36518 (N_36518,N_34053,N_32947);
nand U36519 (N_36519,N_30797,N_31613);
or U36520 (N_36520,N_32276,N_31415);
or U36521 (N_36521,N_34773,N_32053);
nor U36522 (N_36522,N_32906,N_30383);
nand U36523 (N_36523,N_31121,N_32241);
or U36524 (N_36524,N_34424,N_33779);
nand U36525 (N_36525,N_34131,N_33540);
and U36526 (N_36526,N_34047,N_34203);
nand U36527 (N_36527,N_34701,N_31737);
nand U36528 (N_36528,N_34449,N_33081);
and U36529 (N_36529,N_30418,N_31164);
nand U36530 (N_36530,N_31118,N_30489);
xor U36531 (N_36531,N_34446,N_32120);
and U36532 (N_36532,N_31513,N_33660);
nand U36533 (N_36533,N_32239,N_33390);
nand U36534 (N_36534,N_33492,N_30217);
or U36535 (N_36535,N_30877,N_33554);
xnor U36536 (N_36536,N_32956,N_32675);
nor U36537 (N_36537,N_33986,N_31221);
xor U36538 (N_36538,N_32086,N_30779);
or U36539 (N_36539,N_30913,N_34650);
or U36540 (N_36540,N_30729,N_33506);
and U36541 (N_36541,N_34325,N_34999);
and U36542 (N_36542,N_32702,N_33719);
and U36543 (N_36543,N_31719,N_33748);
or U36544 (N_36544,N_30836,N_32872);
nor U36545 (N_36545,N_34969,N_31794);
or U36546 (N_36546,N_33307,N_31634);
and U36547 (N_36547,N_34583,N_32647);
nand U36548 (N_36548,N_31753,N_31167);
or U36549 (N_36549,N_33895,N_32716);
nor U36550 (N_36550,N_33734,N_31216);
or U36551 (N_36551,N_32853,N_31215);
or U36552 (N_36552,N_33107,N_30221);
and U36553 (N_36553,N_33026,N_34603);
nand U36554 (N_36554,N_33950,N_31759);
nand U36555 (N_36555,N_30032,N_30294);
or U36556 (N_36556,N_31391,N_31752);
xnor U36557 (N_36557,N_30479,N_33104);
xnor U36558 (N_36558,N_32686,N_30751);
or U36559 (N_36559,N_31091,N_34823);
xor U36560 (N_36560,N_31375,N_31406);
and U36561 (N_36561,N_33573,N_32237);
xnor U36562 (N_36562,N_34897,N_31369);
nor U36563 (N_36563,N_34624,N_31425);
and U36564 (N_36564,N_33657,N_34276);
xnor U36565 (N_36565,N_34919,N_34697);
nor U36566 (N_36566,N_31722,N_30816);
nand U36567 (N_36567,N_34196,N_31204);
and U36568 (N_36568,N_32182,N_30754);
and U36569 (N_36569,N_31411,N_32848);
nor U36570 (N_36570,N_31444,N_32802);
and U36571 (N_36571,N_34072,N_30567);
nor U36572 (N_36572,N_34434,N_30618);
nand U36573 (N_36573,N_31247,N_34374);
and U36574 (N_36574,N_31038,N_33303);
xor U36575 (N_36575,N_30210,N_34169);
nor U36576 (N_36576,N_31208,N_34986);
nor U36577 (N_36577,N_32153,N_33974);
nand U36578 (N_36578,N_32206,N_34413);
nand U36579 (N_36579,N_32313,N_32990);
and U36580 (N_36580,N_33624,N_34050);
nand U36581 (N_36581,N_30608,N_31162);
or U36582 (N_36582,N_30415,N_31022);
nand U36583 (N_36583,N_31991,N_34067);
nand U36584 (N_36584,N_34653,N_30080);
or U36585 (N_36585,N_30683,N_33499);
nor U36586 (N_36586,N_34359,N_30551);
nand U36587 (N_36587,N_31458,N_34073);
and U36588 (N_36588,N_34018,N_33784);
or U36589 (N_36589,N_32912,N_33816);
nor U36590 (N_36590,N_31441,N_30370);
nor U36591 (N_36591,N_33574,N_34526);
xnor U36592 (N_36592,N_34346,N_33483);
nor U36593 (N_36593,N_32234,N_33189);
xor U36594 (N_36594,N_31924,N_31725);
xnor U36595 (N_36595,N_33027,N_33486);
and U36596 (N_36596,N_34934,N_34763);
xnor U36597 (N_36597,N_34659,N_30188);
xor U36598 (N_36598,N_34064,N_33368);
nand U36599 (N_36599,N_34458,N_31368);
and U36600 (N_36600,N_32066,N_32792);
nand U36601 (N_36601,N_30120,N_31104);
xnor U36602 (N_36602,N_31628,N_33283);
and U36603 (N_36603,N_32114,N_30171);
nor U36604 (N_36604,N_31818,N_33078);
xnor U36605 (N_36605,N_31844,N_30006);
and U36606 (N_36606,N_32864,N_31886);
and U36607 (N_36607,N_32434,N_31105);
or U36608 (N_36608,N_31200,N_30759);
xnor U36609 (N_36609,N_30435,N_32855);
xnor U36610 (N_36610,N_31279,N_32930);
and U36611 (N_36611,N_31957,N_32884);
nand U36612 (N_36612,N_30395,N_31343);
nand U36613 (N_36613,N_31042,N_33373);
nand U36614 (N_36614,N_31632,N_34665);
nand U36615 (N_36615,N_30261,N_33865);
and U36616 (N_36616,N_31302,N_34636);
or U36617 (N_36617,N_32347,N_31214);
or U36618 (N_36618,N_31587,N_34706);
and U36619 (N_36619,N_32408,N_30538);
xnor U36620 (N_36620,N_30971,N_33515);
nor U36621 (N_36621,N_30426,N_31828);
nor U36622 (N_36622,N_33715,N_32230);
or U36623 (N_36623,N_31549,N_31639);
xnor U36624 (N_36624,N_32090,N_34945);
and U36625 (N_36625,N_30838,N_33177);
xor U36626 (N_36626,N_31744,N_33257);
xnor U36627 (N_36627,N_30184,N_30256);
and U36628 (N_36628,N_31595,N_31955);
nor U36629 (N_36629,N_31021,N_33844);
and U36630 (N_36630,N_34678,N_30109);
nand U36631 (N_36631,N_30887,N_33322);
xor U36632 (N_36632,N_30478,N_33049);
or U36633 (N_36633,N_30970,N_30154);
and U36634 (N_36634,N_31224,N_30657);
or U36635 (N_36635,N_31202,N_30338);
and U36636 (N_36636,N_33876,N_33489);
xnor U36637 (N_36637,N_30998,N_30583);
nand U36638 (N_36638,N_31535,N_33725);
nand U36639 (N_36639,N_34448,N_31347);
and U36640 (N_36640,N_34801,N_32249);
xor U36641 (N_36641,N_34187,N_32495);
xnor U36642 (N_36642,N_33320,N_31468);
or U36643 (N_36643,N_34490,N_33823);
xor U36644 (N_36644,N_30694,N_34920);
xor U36645 (N_36645,N_33280,N_33092);
and U36646 (N_36646,N_33965,N_33005);
nor U36647 (N_36647,N_32199,N_34141);
xnor U36648 (N_36648,N_30267,N_31773);
xor U36649 (N_36649,N_30526,N_31430);
or U36650 (N_36650,N_34233,N_31594);
and U36651 (N_36651,N_30550,N_30958);
xor U36652 (N_36652,N_30605,N_33264);
nor U36653 (N_36653,N_30449,N_31229);
nor U36654 (N_36654,N_30815,N_33929);
nand U36655 (N_36655,N_34243,N_31464);
nor U36656 (N_36656,N_33389,N_31356);
or U36657 (N_36657,N_30656,N_32610);
nor U36658 (N_36658,N_33169,N_34213);
nand U36659 (N_36659,N_31069,N_34332);
and U36660 (N_36660,N_33028,N_32195);
nand U36661 (N_36661,N_31910,N_31238);
and U36662 (N_36662,N_33753,N_33707);
nand U36663 (N_36663,N_31682,N_34839);
xor U36664 (N_36664,N_30293,N_33221);
nand U36665 (N_36665,N_30356,N_33294);
nor U36666 (N_36666,N_32738,N_30996);
xnor U36667 (N_36667,N_34942,N_33659);
nand U36668 (N_36668,N_31523,N_34864);
xnor U36669 (N_36669,N_32931,N_33589);
or U36670 (N_36670,N_31082,N_32270);
or U36671 (N_36671,N_30811,N_33850);
xor U36672 (N_36672,N_32949,N_34192);
nor U36673 (N_36673,N_32471,N_31998);
nor U36674 (N_36674,N_34692,N_32006);
nand U36675 (N_36675,N_33436,N_30665);
xnor U36676 (N_36676,N_30981,N_34717);
nand U36677 (N_36677,N_30427,N_32356);
and U36678 (N_36678,N_33834,N_32658);
or U36679 (N_36679,N_30183,N_31132);
and U36680 (N_36680,N_34369,N_31501);
nor U36681 (N_36681,N_31521,N_32251);
nand U36682 (N_36682,N_33184,N_30194);
or U36683 (N_36683,N_31362,N_33807);
or U36684 (N_36684,N_33472,N_33825);
and U36685 (N_36685,N_34334,N_31588);
nor U36686 (N_36686,N_34138,N_32498);
or U36687 (N_36687,N_32844,N_32616);
and U36688 (N_36688,N_30483,N_33822);
nor U36689 (N_36689,N_33831,N_33493);
nor U36690 (N_36690,N_34941,N_32142);
and U36691 (N_36691,N_32477,N_34802);
nor U36692 (N_36692,N_33778,N_33159);
nand U36693 (N_36693,N_30942,N_30295);
xnor U36694 (N_36694,N_30238,N_33228);
or U36695 (N_36695,N_34746,N_30044);
xor U36696 (N_36696,N_30718,N_34205);
nand U36697 (N_36697,N_33945,N_32901);
or U36698 (N_36698,N_31174,N_33462);
or U36699 (N_36699,N_34341,N_33744);
nand U36700 (N_36700,N_31455,N_34248);
xnor U36701 (N_36701,N_33047,N_33757);
and U36702 (N_36702,N_33879,N_34245);
nand U36703 (N_36703,N_31984,N_33325);
and U36704 (N_36704,N_31530,N_30200);
and U36705 (N_36705,N_32381,N_32914);
xnor U36706 (N_36706,N_31565,N_32718);
nand U36707 (N_36707,N_34105,N_30577);
xnor U36708 (N_36708,N_33751,N_30402);
nor U36709 (N_36709,N_33709,N_31097);
or U36710 (N_36710,N_31080,N_34287);
xor U36711 (N_36711,N_33274,N_32821);
or U36712 (N_36712,N_33397,N_33588);
and U36713 (N_36713,N_34686,N_34760);
nand U36714 (N_36714,N_33915,N_30137);
and U36715 (N_36715,N_31949,N_34730);
or U36716 (N_36716,N_30707,N_31692);
and U36717 (N_36717,N_31145,N_32221);
or U36718 (N_36718,N_31517,N_30993);
nand U36719 (N_36719,N_32992,N_31870);
and U36720 (N_36720,N_34714,N_32709);
nor U36721 (N_36721,N_34004,N_33198);
and U36722 (N_36722,N_31308,N_31811);
or U36723 (N_36723,N_31147,N_33877);
nand U36724 (N_36724,N_34557,N_30742);
xor U36725 (N_36725,N_31482,N_31566);
or U36726 (N_36726,N_33161,N_32741);
nor U36727 (N_36727,N_34241,N_31273);
nor U36728 (N_36728,N_31260,N_30546);
or U36729 (N_36729,N_31351,N_31586);
or U36730 (N_36730,N_34396,N_31898);
nand U36731 (N_36731,N_31892,N_34909);
or U36732 (N_36732,N_30025,N_31732);
nand U36733 (N_36733,N_30160,N_32713);
nand U36734 (N_36734,N_33217,N_30337);
and U36735 (N_36735,N_33003,N_31448);
or U36736 (N_36736,N_33162,N_30316);
and U36737 (N_36737,N_32399,N_32638);
and U36738 (N_36738,N_31393,N_34594);
xnor U36739 (N_36739,N_30893,N_31736);
or U36740 (N_36740,N_30241,N_31696);
and U36741 (N_36741,N_31668,N_30158);
or U36742 (N_36742,N_32756,N_32340);
and U36743 (N_36743,N_34110,N_34457);
or U36744 (N_36744,N_33077,N_31052);
xor U36745 (N_36745,N_33452,N_32640);
nor U36746 (N_36746,N_34781,N_31074);
xor U36747 (N_36747,N_31093,N_31287);
and U36748 (N_36748,N_34616,N_30491);
xnor U36749 (N_36749,N_34640,N_34581);
and U36750 (N_36750,N_32209,N_31816);
nor U36751 (N_36751,N_34066,N_31975);
xor U36752 (N_36752,N_32058,N_30597);
nor U36753 (N_36753,N_30507,N_32007);
nor U36754 (N_36754,N_33673,N_32087);
and U36755 (N_36755,N_32760,N_32805);
nand U36756 (N_36756,N_32396,N_34304);
nand U36757 (N_36757,N_32015,N_34812);
nor U36758 (N_36758,N_31228,N_34617);
and U36759 (N_36759,N_30405,N_33488);
and U36760 (N_36760,N_31974,N_32005);
nand U36761 (N_36761,N_30509,N_34095);
or U36762 (N_36762,N_32838,N_34082);
and U36763 (N_36763,N_34776,N_30728);
nor U36764 (N_36764,N_30074,N_30753);
nand U36765 (N_36765,N_31158,N_34155);
or U36766 (N_36766,N_32633,N_33195);
nand U36767 (N_36767,N_34587,N_33063);
xor U36768 (N_36768,N_33048,N_33794);
or U36769 (N_36769,N_31965,N_30233);
xnor U36770 (N_36770,N_34076,N_34855);
xnor U36771 (N_36771,N_34930,N_34599);
xnor U36772 (N_36772,N_31396,N_34766);
nand U36773 (N_36773,N_31580,N_33620);
nand U36774 (N_36774,N_32176,N_30512);
nand U36775 (N_36775,N_30336,N_34039);
nand U36776 (N_36776,N_32890,N_33069);
nand U36777 (N_36777,N_33072,N_32733);
and U36778 (N_36778,N_34914,N_30765);
nor U36779 (N_36779,N_30321,N_34070);
xnor U36780 (N_36780,N_33568,N_33413);
nor U36781 (N_36781,N_31476,N_33175);
and U36782 (N_36782,N_32717,N_33300);
nor U36783 (N_36783,N_30918,N_31461);
nor U36784 (N_36784,N_30590,N_34198);
and U36785 (N_36785,N_30143,N_34488);
and U36786 (N_36786,N_32358,N_32935);
nand U36787 (N_36787,N_33016,N_33222);
nor U36788 (N_36788,N_34200,N_30317);
or U36789 (N_36789,N_32423,N_31758);
nor U36790 (N_36790,N_30492,N_34793);
xnor U36791 (N_36791,N_32618,N_31735);
nand U36792 (N_36792,N_33105,N_33135);
or U36793 (N_36793,N_31636,N_30049);
and U36794 (N_36794,N_31848,N_30384);
or U36795 (N_36795,N_34788,N_33563);
nor U36796 (N_36796,N_31168,N_32854);
nand U36797 (N_36797,N_32217,N_30630);
and U36798 (N_36798,N_34612,N_30182);
and U36799 (N_36799,N_33737,N_32125);
nand U36800 (N_36800,N_34308,N_33440);
nand U36801 (N_36801,N_31835,N_34151);
nor U36802 (N_36802,N_30685,N_31392);
nor U36803 (N_36803,N_30129,N_30043);
nand U36804 (N_36804,N_31357,N_34476);
and U36805 (N_36805,N_32191,N_30988);
and U36806 (N_36806,N_33447,N_34079);
nor U36807 (N_36807,N_34428,N_31793);
xnor U36808 (N_36808,N_31067,N_32642);
or U36809 (N_36809,N_30920,N_32452);
and U36810 (N_36810,N_30424,N_30757);
or U36811 (N_36811,N_30328,N_31990);
nor U36812 (N_36812,N_33632,N_31624);
nor U36813 (N_36813,N_32893,N_33288);
nand U36814 (N_36814,N_31151,N_31534);
or U36815 (N_36815,N_30536,N_33867);
nor U36816 (N_36816,N_32957,N_32436);
and U36817 (N_36817,N_31544,N_31153);
nand U36818 (N_36818,N_32788,N_31604);
xnor U36819 (N_36819,N_32049,N_30060);
nor U36820 (N_36820,N_30864,N_34127);
nor U36821 (N_36821,N_33921,N_32745);
or U36822 (N_36822,N_33631,N_32236);
and U36823 (N_36823,N_32823,N_33890);
and U36824 (N_36824,N_31563,N_34222);
or U36825 (N_36825,N_30380,N_31884);
xnor U36826 (N_36826,N_33756,N_31326);
xor U36827 (N_36827,N_32057,N_32317);
xor U36828 (N_36828,N_30413,N_31631);
or U36829 (N_36829,N_34281,N_33688);
and U36830 (N_36830,N_34885,N_33263);
xor U36831 (N_36831,N_32510,N_34921);
nor U36832 (N_36832,N_33766,N_31959);
nor U36833 (N_36833,N_31124,N_33928);
nand U36834 (N_36834,N_30610,N_32359);
or U36835 (N_36835,N_34879,N_32281);
or U36836 (N_36836,N_32131,N_31504);
xnor U36837 (N_36837,N_34685,N_33521);
and U36838 (N_36838,N_31740,N_33046);
xor U36839 (N_36839,N_32051,N_33059);
or U36840 (N_36840,N_32065,N_33086);
nor U36841 (N_36841,N_31798,N_30930);
nand U36842 (N_36842,N_30643,N_33788);
nand U36843 (N_36843,N_30083,N_33545);
xor U36844 (N_36844,N_31146,N_31175);
or U36845 (N_36845,N_33982,N_32177);
and U36846 (N_36846,N_32516,N_34026);
or U36847 (N_36847,N_34633,N_33926);
nand U36848 (N_36848,N_34731,N_33209);
or U36849 (N_36849,N_34338,N_30061);
or U36850 (N_36850,N_34606,N_32962);
xnor U36851 (N_36851,N_31823,N_34007);
xor U36852 (N_36852,N_34019,N_34427);
nand U36853 (N_36853,N_30658,N_32859);
xnor U36854 (N_36854,N_33714,N_32054);
nor U36855 (N_36855,N_33882,N_34134);
or U36856 (N_36856,N_33479,N_31116);
nor U36857 (N_36857,N_31533,N_34699);
or U36858 (N_36858,N_30949,N_32444);
or U36859 (N_36859,N_32870,N_34051);
xor U36860 (N_36860,N_31185,N_33804);
nor U36861 (N_36861,N_33663,N_32753);
nand U36862 (N_36862,N_33496,N_32614);
nor U36863 (N_36863,N_34856,N_32539);
xor U36864 (N_36864,N_32266,N_31135);
xor U36865 (N_36865,N_33827,N_32898);
nor U36866 (N_36866,N_32271,N_30631);
nand U36867 (N_36867,N_31379,N_34693);
and U36868 (N_36868,N_31179,N_30698);
and U36869 (N_36869,N_33405,N_34008);
nand U36870 (N_36870,N_34561,N_30379);
or U36871 (N_36871,N_33677,N_30995);
xnor U36872 (N_36872,N_32304,N_31799);
and U36873 (N_36873,N_33980,N_30100);
nand U36874 (N_36874,N_30239,N_30463);
nor U36875 (N_36875,N_33318,N_30107);
xnor U36876 (N_36876,N_31002,N_31240);
and U36877 (N_36877,N_31446,N_33128);
and U36878 (N_36878,N_33797,N_34646);
nand U36879 (N_36879,N_34679,N_30910);
and U36880 (N_36880,N_32465,N_33233);
xnor U36881 (N_36881,N_34395,N_32184);
xor U36882 (N_36882,N_32695,N_34858);
and U36883 (N_36883,N_33836,N_31830);
and U36884 (N_36884,N_32246,N_31802);
nor U36885 (N_36885,N_32104,N_30410);
xnor U36886 (N_36886,N_33134,N_34905);
and U36887 (N_36887,N_33889,N_31640);
xor U36888 (N_36888,N_32862,N_33044);
and U36889 (N_36889,N_31417,N_33178);
nand U36890 (N_36890,N_30355,N_31149);
xor U36891 (N_36891,N_32778,N_31982);
nor U36892 (N_36892,N_33616,N_34952);
nor U36893 (N_36893,N_31603,N_34027);
nand U36894 (N_36894,N_31801,N_33789);
xor U36895 (N_36895,N_32027,N_34964);
nor U36896 (N_36896,N_31070,N_31845);
nor U36897 (N_36897,N_34349,N_31165);
or U36898 (N_36898,N_32620,N_30902);
nor U36899 (N_36899,N_34159,N_32934);
nor U36900 (N_36900,N_32553,N_33097);
xor U36901 (N_36901,N_34392,N_32133);
or U36902 (N_36902,N_31469,N_34645);
or U36903 (N_36903,N_34782,N_32460);
or U36904 (N_36904,N_33622,N_30625);
and U36905 (N_36905,N_32674,N_33471);
or U36906 (N_36906,N_33948,N_34533);
nand U36907 (N_36907,N_30650,N_34470);
nand U36908 (N_36908,N_30244,N_31919);
xnor U36909 (N_36909,N_32940,N_30199);
nand U36910 (N_36910,N_34270,N_34353);
nor U36911 (N_36911,N_31064,N_33863);
or U36912 (N_36912,N_34742,N_34765);
and U36913 (N_36913,N_31856,N_32682);
nand U36914 (N_36914,N_34664,N_33485);
xor U36915 (N_36915,N_31781,N_34191);
and U36916 (N_36916,N_30576,N_30696);
nand U36917 (N_36917,N_30011,N_32764);
nor U36918 (N_36918,N_34618,N_30216);
and U36919 (N_36919,N_30012,N_33524);
nand U36920 (N_36920,N_31193,N_33076);
or U36921 (N_36921,N_32924,N_30667);
nor U36922 (N_36922,N_32701,N_34728);
or U36923 (N_36923,N_30501,N_34649);
nor U36924 (N_36924,N_33690,N_31852);
or U36925 (N_36925,N_32256,N_30899);
nor U36926 (N_36926,N_30203,N_32820);
or U36927 (N_36927,N_33386,N_34910);
nor U36928 (N_36928,N_32311,N_31703);
and U36929 (N_36929,N_31500,N_31876);
nand U36930 (N_36930,N_30941,N_32463);
nand U36931 (N_36931,N_33374,N_33528);
nor U36932 (N_36932,N_32834,N_33875);
and U36933 (N_36933,N_33564,N_33851);
or U36934 (N_36934,N_34379,N_34300);
or U36935 (N_36935,N_31827,N_31291);
nand U36936 (N_36936,N_34037,N_34075);
nand U36937 (N_36937,N_30513,N_31170);
or U36938 (N_36938,N_30545,N_30445);
and U36939 (N_36939,N_31727,N_33148);
nand U36940 (N_36940,N_30761,N_34221);
or U36941 (N_36941,N_33099,N_31088);
xor U36942 (N_36942,N_34809,N_33580);
nand U36943 (N_36943,N_30040,N_31568);
nor U36944 (N_36944,N_30004,N_32260);
or U36945 (N_36945,N_30161,N_31831);
nand U36946 (N_36946,N_34491,N_31349);
or U36947 (N_36947,N_30235,N_31762);
and U36948 (N_36948,N_30326,N_31649);
xnor U36949 (N_36949,N_33893,N_30873);
xor U36950 (N_36950,N_30997,N_31176);
xor U36951 (N_36951,N_34666,N_30163);
xor U36952 (N_36952,N_31423,N_31971);
and U36953 (N_36953,N_30786,N_31358);
xnor U36954 (N_36954,N_32457,N_33272);
nor U36955 (N_36955,N_32719,N_33860);
or U36956 (N_36956,N_30245,N_33171);
xor U36957 (N_36957,N_32137,N_32361);
and U36958 (N_36958,N_30839,N_30883);
or U36959 (N_36959,N_31620,N_31401);
or U36960 (N_36960,N_31195,N_31646);
nand U36961 (N_36961,N_34890,N_34314);
xnor U36962 (N_36962,N_32710,N_33938);
and U36963 (N_36963,N_32993,N_33777);
nor U36964 (N_36964,N_34224,N_34808);
xnor U36965 (N_36965,N_31241,N_32679);
nor U36966 (N_36966,N_30743,N_32794);
nor U36967 (N_36967,N_34563,N_34904);
and U36968 (N_36968,N_34081,N_33041);
xor U36969 (N_36969,N_34344,N_33913);
or U36970 (N_36970,N_33750,N_30270);
nor U36971 (N_36971,N_30854,N_32560);
and U36972 (N_36972,N_30243,N_31908);
xnor U36973 (N_36973,N_33333,N_31250);
or U36974 (N_36974,N_34244,N_34078);
nor U36975 (N_36975,N_30560,N_32345);
nand U36976 (N_36976,N_31376,N_34468);
nand U36977 (N_36977,N_30833,N_31877);
xor U36978 (N_36978,N_34058,N_34695);
or U36979 (N_36979,N_31850,N_32468);
or U36980 (N_36980,N_32547,N_32522);
nand U36981 (N_36981,N_34884,N_30390);
nor U36982 (N_36982,N_30327,N_33910);
xor U36983 (N_36983,N_31597,N_31378);
and U36984 (N_36984,N_34128,N_32438);
nand U36985 (N_36985,N_31101,N_32584);
xor U36986 (N_36986,N_30456,N_30954);
xnor U36987 (N_36987,N_33213,N_34768);
xnor U36988 (N_36988,N_34140,N_32336);
nand U36989 (N_36989,N_30374,N_32952);
nand U36990 (N_36990,N_30676,N_30782);
nand U36991 (N_36991,N_32107,N_30367);
nor U36992 (N_36992,N_34102,N_33465);
xor U36993 (N_36993,N_33330,N_30956);
nor U36994 (N_36994,N_33932,N_34548);
nand U36995 (N_36995,N_34284,N_33754);
or U36996 (N_36996,N_34727,N_30462);
and U36997 (N_36997,N_32373,N_33543);
nor U36998 (N_36998,N_31645,N_30070);
nand U36999 (N_36999,N_34635,N_30671);
or U37000 (N_37000,N_31928,N_34840);
nand U37001 (N_37001,N_33469,N_34381);
xor U37002 (N_37002,N_30874,N_34377);
nand U37003 (N_37003,N_31868,N_34146);
xor U37004 (N_37004,N_31486,N_30079);
xnor U37005 (N_37005,N_31730,N_32060);
or U37006 (N_37006,N_33070,N_30177);
or U37007 (N_37007,N_33032,N_33726);
nor U37008 (N_37008,N_30774,N_32727);
nand U37009 (N_37009,N_31460,N_32117);
and U37010 (N_37010,N_32118,N_31483);
or U37011 (N_37011,N_30081,N_33849);
and U37012 (N_37012,N_34384,N_30176);
nor U37013 (N_37013,N_34260,N_32486);
or U37014 (N_37014,N_32397,N_31994);
or U37015 (N_37015,N_34197,N_32354);
nor U37016 (N_37016,N_32652,N_33625);
nor U37017 (N_37017,N_33596,N_32729);
xnor U37018 (N_37018,N_30272,N_31973);
xnor U37019 (N_37019,N_33376,N_33455);
nor U37020 (N_37020,N_33896,N_34895);
nand U37021 (N_37021,N_33835,N_31602);
xor U37022 (N_37022,N_34259,N_30516);
nand U37023 (N_37023,N_33265,N_33897);
nand U37024 (N_37024,N_32288,N_31731);
xnor U37025 (N_37025,N_31427,N_32653);
nand U37026 (N_37026,N_30579,N_32921);
and U37027 (N_37027,N_30783,N_32157);
or U37028 (N_37028,N_34710,N_33349);
and U37029 (N_37029,N_34463,N_34740);
nand U37030 (N_37030,N_30555,N_33006);
nor U37031 (N_37031,N_32689,N_32441);
nand U37032 (N_37032,N_34849,N_34696);
or U37033 (N_37033,N_32723,N_32506);
and U37034 (N_37034,N_31019,N_33468);
and U37035 (N_37035,N_30549,N_31693);
or U37036 (N_37036,N_32791,N_30078);
or U37037 (N_37037,N_31887,N_33342);
nor U37038 (N_37038,N_33008,N_30529);
or U37039 (N_37039,N_32955,N_31360);
nand U37040 (N_37040,N_32478,N_32530);
or U37041 (N_37041,N_34246,N_31363);
xnor U37042 (N_37042,N_30036,N_33604);
nand U37043 (N_37043,N_34630,N_30682);
or U37044 (N_37044,N_30312,N_32333);
and U37045 (N_37045,N_31660,N_32272);
nand U37046 (N_37046,N_31231,N_30108);
nor U37047 (N_37047,N_34651,N_33384);
or U37048 (N_37048,N_34350,N_34331);
or U37049 (N_37049,N_31173,N_34663);
nand U37050 (N_37050,N_31717,N_33998);
and U37051 (N_37051,N_33858,N_33326);
xor U37052 (N_37052,N_34595,N_33820);
xnor U37053 (N_37053,N_31635,N_30393);
and U37054 (N_37054,N_31252,N_33767);
and U37055 (N_37055,N_32958,N_34826);
nand U37056 (N_37056,N_34112,N_34882);
nor U37057 (N_37057,N_33382,N_30168);
xnor U37058 (N_37058,N_34759,N_32193);
nand U37059 (N_37059,N_32989,N_30155);
nor U37060 (N_37060,N_34421,N_32325);
or U37061 (N_37061,N_32909,N_30376);
or U37062 (N_37062,N_31888,N_30875);
nand U37063 (N_37063,N_30820,N_31685);
nor U37064 (N_37064,N_34703,N_33977);
and U37065 (N_37065,N_32214,N_31642);
xnor U37066 (N_37066,N_30350,N_31878);
xor U37067 (N_37067,N_30343,N_30533);
xnor U37068 (N_37068,N_32938,N_31422);
or U37069 (N_37069,N_32427,N_30919);
nand U37070 (N_37070,N_33527,N_31833);
xor U37071 (N_37071,N_32245,N_30453);
xor U37072 (N_37072,N_34800,N_31081);
nor U37073 (N_37073,N_31325,N_30396);
nor U37074 (N_37074,N_30092,N_34173);
or U37075 (N_37075,N_30975,N_31129);
nor U37076 (N_37076,N_34975,N_34045);
or U37077 (N_37077,N_33286,N_32451);
and U37078 (N_37078,N_30056,N_30539);
nand U37079 (N_37079,N_34625,N_31575);
and U37080 (N_37080,N_34720,N_31253);
xor U37081 (N_37081,N_30333,N_32896);
nor U37082 (N_37082,N_34043,N_33559);
and U37083 (N_37083,N_34873,N_34707);
and U37084 (N_37084,N_32558,N_33613);
nand U37085 (N_37085,N_30863,N_30963);
nor U37086 (N_37086,N_31543,N_34586);
and U37087 (N_37087,N_30609,N_30804);
nand U37088 (N_37088,N_30152,N_32409);
or U37089 (N_37089,N_30857,N_34364);
nand U37090 (N_37090,N_30240,N_30351);
nor U37091 (N_37091,N_30144,N_32050);
or U37092 (N_37092,N_32511,N_32602);
and U37093 (N_37093,N_34667,N_31301);
xor U37094 (N_37094,N_31154,N_33275);
nor U37095 (N_37095,N_31305,N_34755);
and U37096 (N_37096,N_32138,N_30659);
and U37097 (N_37097,N_31843,N_31885);
nor U37098 (N_37098,N_34537,N_30440);
and U37099 (N_37099,N_30065,N_33201);
xnor U37100 (N_37100,N_34186,N_33441);
nand U37101 (N_37101,N_34336,N_32619);
nand U37102 (N_37102,N_31122,N_33323);
xor U37103 (N_37103,N_34001,N_33704);
and U37104 (N_37104,N_33793,N_33231);
xnor U37105 (N_37105,N_34226,N_30407);
or U37106 (N_37106,N_31246,N_33308);
xor U37107 (N_37107,N_30748,N_31505);
and U37108 (N_37108,N_32981,N_30540);
xor U37109 (N_37109,N_34613,N_32787);
xor U37110 (N_37110,N_33058,N_30617);
nor U37111 (N_37111,N_34772,N_31790);
xor U37112 (N_37112,N_32113,N_33582);
xor U37113 (N_37113,N_32220,N_32254);
nand U37114 (N_37114,N_30983,N_34621);
and U37115 (N_37115,N_34756,N_30064);
xnor U37116 (N_37116,N_32920,N_33203);
nor U37117 (N_37117,N_30162,N_30497);
or U37118 (N_37118,N_32668,N_33125);
or U37119 (N_37119,N_33773,N_31617);
and U37120 (N_37120,N_33106,N_33801);
nand U37121 (N_37121,N_34218,N_34604);
nand U37122 (N_37122,N_32235,N_33821);
nor U37123 (N_37123,N_30347,N_34156);
or U37124 (N_37124,N_32939,N_32069);
nand U37125 (N_37125,N_32895,N_32517);
or U37126 (N_37126,N_31842,N_31331);
nor U37127 (N_37127,N_30896,N_32255);
or U37128 (N_37128,N_31142,N_34683);
and U37129 (N_37129,N_31621,N_32899);
nor U37130 (N_37130,N_33207,N_34996);
xor U37131 (N_37131,N_30842,N_30126);
and U37132 (N_37132,N_34525,N_31609);
and U37133 (N_37133,N_31749,N_32310);
and U37134 (N_37134,N_34805,N_34511);
or U37135 (N_37135,N_32412,N_30672);
nor U37136 (N_37136,N_34779,N_34499);
nor U37137 (N_37137,N_31066,N_31033);
xnor U37138 (N_37138,N_31548,N_31083);
or U37139 (N_37139,N_32724,N_32538);
nand U37140 (N_37140,N_31073,N_33762);
and U37141 (N_37141,N_34405,N_31663);
and U37142 (N_37142,N_32977,N_30072);
nor U37143 (N_37143,N_32459,N_32080);
xor U37144 (N_37144,N_34866,N_30557);
nand U37145 (N_37145,N_30992,N_31980);
or U37146 (N_37146,N_33815,N_32527);
or U37147 (N_37147,N_31137,N_33534);
nor U37148 (N_37148,N_33147,N_30713);
nor U37149 (N_37149,N_33284,N_33979);
nand U37150 (N_37150,N_33931,N_32301);
or U37151 (N_37151,N_31233,N_32352);
or U37152 (N_37152,N_34639,N_34061);
nand U37153 (N_37153,N_33732,N_30369);
nor U37154 (N_37154,N_32508,N_34822);
nand U37155 (N_37155,N_30764,N_31495);
nor U37156 (N_37156,N_33684,N_32083);
nand U37157 (N_37157,N_33626,N_34249);
nor U37158 (N_37158,N_33001,N_31784);
or U37159 (N_37159,N_32440,N_31729);
or U37160 (N_37160,N_34306,N_33210);
nor U37161 (N_37161,N_32942,N_34579);
and U37162 (N_37162,N_32216,N_30990);
xnor U37163 (N_37163,N_33745,N_32437);
nor U37164 (N_37164,N_34305,N_34641);
and U37165 (N_37165,N_34676,N_30027);
nand U37166 (N_37166,N_32552,N_30711);
nor U37167 (N_37167,N_32871,N_31902);
nand U37168 (N_37168,N_34713,N_30433);
nand U37169 (N_37169,N_31883,N_32926);
and U37170 (N_37170,N_30858,N_30438);
nor U37171 (N_37171,N_32961,N_34397);
xnor U37172 (N_37172,N_34282,N_30448);
nor U37173 (N_37173,N_30585,N_32818);
xnor U37174 (N_37174,N_33154,N_32923);
nor U37175 (N_37175,N_31138,N_30727);
xnor U37176 (N_37176,N_30640,N_31499);
and U37177 (N_37177,N_30834,N_33749);
and U37178 (N_37178,N_33852,N_33832);
xor U37179 (N_37179,N_33687,N_33062);
or U37180 (N_37180,N_32223,N_30375);
or U37181 (N_37181,N_30572,N_32337);
xor U37182 (N_37182,N_33790,N_34657);
and U37183 (N_37183,N_30330,N_34209);
xnor U37184 (N_37184,N_34239,N_30503);
xnor U37185 (N_37185,N_33350,N_34531);
nor U37186 (N_37186,N_31194,N_30496);
or U37187 (N_37187,N_30939,N_34859);
nand U37188 (N_37188,N_31993,N_32546);
or U37189 (N_37189,N_31242,N_34509);
or U37190 (N_37190,N_34501,N_31078);
nor U37191 (N_37191,N_33487,N_33547);
nor U37192 (N_37192,N_31865,N_33689);
nor U37193 (N_37193,N_34893,N_32491);
nand U37194 (N_37194,N_30055,N_30726);
nand U37195 (N_37195,N_33886,N_34437);
or U37196 (N_37196,N_30606,N_30898);
or U37197 (N_37197,N_31006,N_30029);
nor U37198 (N_37198,N_33934,N_30131);
or U37199 (N_37199,N_32300,N_31244);
and U37200 (N_37200,N_32194,N_30297);
nor U37201 (N_37201,N_34386,N_34250);
and U37202 (N_37202,N_34372,N_31271);
nand U37203 (N_37203,N_33317,N_33593);
xor U37204 (N_37204,N_34632,N_32362);
or U37205 (N_37205,N_30289,N_30932);
or U37206 (N_37206,N_33994,N_33113);
nand U37207 (N_37207,N_32430,N_30148);
nor U37208 (N_37208,N_30257,N_34289);
xnor U37209 (N_37209,N_31438,N_31656);
nor U37210 (N_37210,N_33996,N_34441);
nand U37211 (N_37211,N_33214,N_31036);
and U37212 (N_37212,N_31952,N_33140);
nor U37213 (N_37213,N_33736,N_33667);
and U37214 (N_37214,N_33218,N_34175);
or U37215 (N_37215,N_34153,N_31622);
nor U37216 (N_37216,N_33246,N_32442);
xor U37217 (N_37217,N_34655,N_33819);
nand U37218 (N_37218,N_34815,N_34461);
xor U37219 (N_37219,N_31742,N_31545);
or U37220 (N_37220,N_30989,N_31536);
xor U37221 (N_37221,N_34431,N_33943);
or U37222 (N_37222,N_31964,N_32029);
nor U37223 (N_37223,N_33253,N_30762);
or U37224 (N_37224,N_33646,N_33273);
and U37225 (N_37225,N_31630,N_32815);
nor U37226 (N_37226,N_32916,N_33010);
nand U37227 (N_37227,N_34094,N_31477);
and U37228 (N_37228,N_32507,N_30929);
or U37229 (N_37229,N_31245,N_30103);
xor U37230 (N_37230,N_34984,N_32648);
or U37231 (N_37231,N_33548,N_33553);
or U37232 (N_37232,N_33608,N_31029);
nand U37233 (N_37233,N_31096,N_30886);
or U37234 (N_37234,N_32435,N_33434);
nor U37235 (N_37235,N_31904,N_32615);
or U37236 (N_37236,N_34148,N_32143);
nor U37237 (N_37237,N_34262,N_30053);
nand U37238 (N_37238,N_31385,N_30016);
xor U37239 (N_37239,N_32579,N_32707);
nor U37240 (N_37240,N_34556,N_30191);
nor U37241 (N_37241,N_33771,N_34868);
xnor U37242 (N_37242,N_30262,N_30994);
nand U37243 (N_37243,N_33365,N_30265);
and U37244 (N_37244,N_32782,N_34883);
or U37245 (N_37245,N_30278,N_34601);
xor U37246 (N_37246,N_33085,N_31075);
and U37247 (N_37247,N_34870,N_31524);
or U37248 (N_37248,N_31824,N_30026);
nand U37249 (N_37249,N_31972,N_33237);
xor U37250 (N_37250,N_31808,N_32523);
or U37251 (N_37251,N_31490,N_32840);
xor U37252 (N_37252,N_33142,N_34558);
and U37253 (N_37253,N_31510,N_32003);
and U37254 (N_37254,N_32130,N_34704);
nand U37255 (N_37255,N_34264,N_31025);
xor U37256 (N_37256,N_30018,N_30101);
nand U37257 (N_37257,N_32432,N_33127);
nand U37258 (N_37258,N_32537,N_31782);
or U37259 (N_37259,N_34555,N_32305);
or U37260 (N_37260,N_32817,N_32315);
xnor U37261 (N_37261,N_33234,N_32556);
nor U37262 (N_37262,N_30518,N_34433);
nor U37263 (N_37263,N_30159,N_32562);
or U37264 (N_37264,N_30788,N_33123);
nor U37265 (N_37265,N_31055,N_32932);
or U37266 (N_37266,N_31577,N_34228);
and U37267 (N_37267,N_30946,N_31647);
nand U37268 (N_37268,N_30202,N_34171);
nor U37269 (N_37269,N_30603,N_33542);
nor U37270 (N_37270,N_30365,N_32673);
nand U37271 (N_37271,N_31724,N_30844);
xnor U37272 (N_37272,N_34605,N_34464);
xor U37273 (N_37273,N_33244,N_30530);
xnor U37274 (N_37274,N_32258,N_30830);
nor U37275 (N_37275,N_32326,N_31317);
xnor U37276 (N_37276,N_31512,N_31948);
xnor U37277 (N_37277,N_32520,N_34577);
or U37278 (N_37278,N_30423,N_31836);
nand U37279 (N_37279,N_34825,N_33259);
xor U37280 (N_37280,N_32611,N_31723);
xnor U37281 (N_37281,N_30805,N_34926);
xor U37282 (N_37282,N_34130,N_30514);
nor U37283 (N_37283,N_32098,N_30259);
nand U37284 (N_37284,N_34780,N_33298);
nand U37285 (N_37285,N_32267,N_33467);
nand U37286 (N_37286,N_31788,N_31177);
xor U37287 (N_37287,N_33961,N_32139);
xor U37288 (N_37288,N_34227,N_32997);
nor U37289 (N_37289,N_30344,N_34021);
or U37290 (N_37290,N_30544,N_31897);
xnor U37291 (N_37291,N_34502,N_31935);
or U37292 (N_37292,N_33446,N_34959);
nand U37293 (N_37293,N_31771,N_32385);
and U37294 (N_37294,N_34098,N_31496);
nand U37295 (N_37295,N_30528,N_34743);
nor U37296 (N_37296,N_30470,N_34752);
xnor U37297 (N_37297,N_34907,N_34090);
or U37298 (N_37298,N_31861,N_30944);
xor U37299 (N_37299,N_32887,N_32344);
xor U37300 (N_37300,N_30781,N_33843);
nand U37301 (N_37301,N_33304,N_33306);
and U37302 (N_37302,N_32169,N_32559);
nor U37303 (N_37303,N_34754,N_33141);
nand U37304 (N_37304,N_33268,N_33891);
or U37305 (N_37305,N_31909,N_32205);
nor U37306 (N_37306,N_31743,N_34737);
or U37307 (N_37307,N_33448,N_32762);
or U37308 (N_37308,N_31936,N_31053);
xor U37309 (N_37309,N_31834,N_32403);
nor U37310 (N_37310,N_31792,N_32712);
or U37311 (N_37311,N_30042,N_30758);
xor U37312 (N_37312,N_31270,N_33824);
or U37313 (N_37313,N_32073,N_34482);
and U37314 (N_37314,N_31891,N_32575);
nor U37315 (N_37315,N_32282,N_30352);
xor U37316 (N_37316,N_33696,N_30292);
and U37317 (N_37317,N_31484,N_34301);
nor U37318 (N_37318,N_34056,N_31418);
nor U37319 (N_37319,N_32012,N_32110);
or U37320 (N_37320,N_34758,N_30318);
nand U37321 (N_37321,N_34041,N_33451);
or U37322 (N_37322,N_33670,N_31686);
and U37323 (N_37323,N_30965,N_32404);
or U37324 (N_37324,N_31747,N_32911);
and U37325 (N_37325,N_33212,N_30258);
and U37326 (N_37326,N_32531,N_31402);
or U37327 (N_37327,N_34865,N_31341);
xor U37328 (N_37328,N_30051,N_32000);
or U37329 (N_37329,N_33226,N_30167);
or U37330 (N_37330,N_32102,N_31541);
nor U37331 (N_37331,N_33695,N_33650);
and U37332 (N_37332,N_31387,N_30925);
nor U37333 (N_37333,N_30911,N_30170);
nor U37334 (N_37334,N_32092,N_33190);
nor U37335 (N_37335,N_31372,N_30790);
nor U37336 (N_37336,N_34444,N_33633);
nand U37337 (N_37337,N_30387,N_31714);
and U37338 (N_37338,N_32019,N_33997);
nand U37339 (N_37339,N_32813,N_31720);
nand U37340 (N_37340,N_31551,N_32803);
nand U37341 (N_37341,N_31698,N_30826);
nand U37342 (N_37342,N_34313,N_31661);
nand U37343 (N_37343,N_34207,N_31525);
nand U37344 (N_37344,N_32389,N_33976);
nand U37345 (N_37345,N_34523,N_34994);
and U37346 (N_37346,N_31353,N_33541);
nand U37347 (N_37347,N_32929,N_30735);
xnor U37348 (N_37348,N_32204,N_31172);
and U37349 (N_37349,N_33665,N_30651);
xor U37350 (N_37350,N_31733,N_34124);
and U37351 (N_37351,N_31840,N_30824);
nand U37352 (N_37352,N_33731,N_31023);
or U37353 (N_37353,N_34412,N_30508);
nor U37354 (N_37354,N_33936,N_30334);
nand U37355 (N_37355,N_31791,N_30652);
xnor U37356 (N_37356,N_32387,N_31035);
nor U37357 (N_37357,N_33187,N_34157);
nor U37358 (N_37358,N_34944,N_33953);
nand U37359 (N_37359,N_33438,N_33156);
nand U37360 (N_37360,N_34407,N_34165);
nor U37361 (N_37361,N_30943,N_32825);
xor U37362 (N_37362,N_34660,N_33517);
nor U37363 (N_37363,N_31249,N_33102);
xor U37364 (N_37364,N_34029,N_32622);
and U37365 (N_37365,N_34031,N_31324);
or U37366 (N_37366,N_33830,N_32192);
or U37367 (N_37367,N_34059,N_30115);
nand U37368 (N_37368,N_32843,N_31783);
nand U37369 (N_37369,N_33334,N_30451);
or U37370 (N_37370,N_31937,N_34570);
xor U37371 (N_37371,N_33975,N_32259);
and U37372 (N_37372,N_30230,N_30264);
or U37373 (N_37373,N_32662,N_31821);
nand U37374 (N_37374,N_31986,N_30882);
xor U37375 (N_37375,N_32461,N_31445);
or U37376 (N_37376,N_32028,N_30733);
or U37377 (N_37377,N_31330,N_31062);
nand U37378 (N_37378,N_31746,N_34254);
nor U37379 (N_37379,N_33248,N_30499);
or U37380 (N_37380,N_34472,N_30655);
nor U37381 (N_37381,N_32040,N_31276);
and U37382 (N_37382,N_33839,N_30666);
nand U37383 (N_37383,N_30187,N_34512);
xnor U37384 (N_37384,N_32009,N_33752);
and U37385 (N_37385,N_30003,N_31619);
nor U37386 (N_37386,N_33765,N_34807);
and U37387 (N_37387,N_32540,N_31895);
xnor U37388 (N_37388,N_33741,N_34958);
and U37389 (N_37389,N_31680,N_34028);
or U37390 (N_37390,N_33458,N_34065);
nor U37391 (N_37391,N_33383,N_31280);
nand U37392 (N_37392,N_32623,N_34819);
or U37393 (N_37393,N_33206,N_33504);
nor U37394 (N_37394,N_32331,N_33138);
nor U37395 (N_37395,N_31065,N_30399);
and U37396 (N_37396,N_31616,N_32218);
or U37397 (N_37397,N_30494,N_34422);
and U37398 (N_37398,N_34435,N_32806);
nand U37399 (N_37399,N_30362,N_34835);
nor U37400 (N_37400,N_33584,N_31893);
nand U37401 (N_37401,N_32446,N_32022);
xor U37402 (N_37402,N_34345,N_34438);
xor U37403 (N_37403,N_32502,N_31989);
nor U37404 (N_37404,N_34057,N_33137);
and U37405 (N_37405,N_32982,N_33309);
xor U37406 (N_37406,N_32039,N_33302);
nand U37407 (N_37407,N_30030,N_30377);
nor U37408 (N_37408,N_34995,N_31849);
nor U37409 (N_37409,N_32597,N_31681);
nand U37410 (N_37410,N_30342,N_32857);
and U37411 (N_37411,N_32963,N_30578);
and U37412 (N_37412,N_31443,N_33476);
or U37413 (N_37413,N_30853,N_31159);
and U37414 (N_37414,N_31106,N_32557);
nand U37415 (N_37415,N_33021,N_33336);
nand U37416 (N_37416,N_34010,N_30190);
nand U37417 (N_37417,N_30688,N_30164);
and U37418 (N_37418,N_32959,N_33969);
xnor U37419 (N_37419,N_32671,N_30031);
nor U37420 (N_37420,N_30687,N_32555);
and U37421 (N_37421,N_33614,N_31181);
nor U37422 (N_37422,N_33393,N_32967);
or U37423 (N_37423,N_30961,N_31292);
and U37424 (N_37424,N_34899,N_34627);
nor U37425 (N_37425,N_32651,N_34774);
nand U37426 (N_37426,N_31334,N_31863);
nor U37427 (N_37427,N_31155,N_34719);
nor U37428 (N_37428,N_30429,N_34518);
or U37429 (N_37429,N_30668,N_32746);
and U37430 (N_37430,N_30124,N_33192);
xnor U37431 (N_37431,N_31554,N_31262);
and U37432 (N_37432,N_30827,N_34042);
or U37433 (N_37433,N_30769,N_33686);
nor U37434 (N_37434,N_31641,N_30150);
or U37435 (N_37435,N_33164,N_32100);
xor U37436 (N_37436,N_34932,N_30945);
nand U37437 (N_37437,N_33133,N_34275);
nand U37438 (N_37438,N_32740,N_30422);
and U37439 (N_37439,N_32533,N_33902);
nand U37440 (N_37440,N_33220,N_33271);
nor U37441 (N_37441,N_32672,N_30069);
xor U37442 (N_37442,N_32135,N_31684);
nor U37443 (N_37443,N_34292,N_30767);
xor U37444 (N_37444,N_32865,N_30166);
or U37445 (N_37445,N_33429,N_30710);
xor U37446 (N_37446,N_32108,N_32248);
nor U37447 (N_37447,N_32293,N_32109);
nand U37448 (N_37448,N_34596,N_32168);
xor U37449 (N_37449,N_32030,N_34496);
or U37450 (N_37450,N_30309,N_30686);
xor U37451 (N_37451,N_33200,N_30673);
nand U37452 (N_37452,N_33635,N_33947);
and U37453 (N_37453,N_31322,N_32466);
nand U37454 (N_37454,N_30476,N_33319);
or U37455 (N_37455,N_31653,N_34360);
nor U37456 (N_37456,N_32680,N_32777);
nand U37457 (N_37457,N_34020,N_34886);
xnor U37458 (N_37458,N_34955,N_30849);
xnor U37459 (N_37459,N_34462,N_32035);
xnor U37460 (N_37460,N_34821,N_30010);
or U37461 (N_37461,N_33442,N_32242);
nor U37462 (N_37462,N_33991,N_31475);
and U37463 (N_37463,N_32422,N_34342);
and U37464 (N_37464,N_33538,N_34475);
or U37465 (N_37465,N_34732,N_32880);
nand U37466 (N_37466,N_30681,N_30224);
and U37467 (N_37467,N_34480,N_33555);
nor U37468 (N_37468,N_32628,N_32842);
or U37469 (N_37469,N_32696,N_34261);
nand U37470 (N_37470,N_31970,N_33700);
and U37471 (N_37471,N_30664,N_34419);
nand U37472 (N_37472,N_30770,N_30250);
and U37473 (N_37473,N_32698,N_31706);
nor U37474 (N_37474,N_32450,N_30452);
xor U37475 (N_37475,N_30928,N_31967);
nand U37476 (N_37476,N_31034,N_34033);
nor U37477 (N_37477,N_34724,N_32433);
xnor U37478 (N_37478,N_32725,N_34327);
nor U37479 (N_37479,N_31298,N_32126);
xnor U37480 (N_37480,N_30130,N_34744);
or U37481 (N_37481,N_33724,N_32699);
nand U37482 (N_37482,N_34852,N_30504);
and U37483 (N_37483,N_32830,N_33615);
nand U37484 (N_37484,N_31297,N_33343);
nand U37485 (N_37485,N_32692,N_34976);
xnor U37486 (N_37486,N_31365,N_30722);
nand U37487 (N_37487,N_30859,N_33859);
and U37488 (N_37488,N_30730,N_34180);
nand U37489 (N_37489,N_32694,N_33043);
or U37490 (N_37490,N_30286,N_32046);
and U37491 (N_37491,N_34126,N_32999);
xor U37492 (N_37492,N_30977,N_31359);
nand U37493 (N_37493,N_33245,N_33352);
xor U37494 (N_37494,N_33606,N_32320);
and U37495 (N_37495,N_33775,N_31086);
or U37496 (N_37496,N_31694,N_30296);
or U37497 (N_37497,N_32122,N_31352);
and U37498 (N_37498,N_32749,N_31871);
xnor U37499 (N_37499,N_33868,N_32048);
nor U37500 (N_37500,N_34398,N_34134);
or U37501 (N_37501,N_33334,N_32590);
nand U37502 (N_37502,N_31339,N_30650);
nor U37503 (N_37503,N_30372,N_32394);
or U37504 (N_37504,N_31600,N_31387);
and U37505 (N_37505,N_33578,N_34758);
or U37506 (N_37506,N_31615,N_30799);
nor U37507 (N_37507,N_32583,N_32832);
nand U37508 (N_37508,N_31856,N_31388);
nand U37509 (N_37509,N_33138,N_33126);
nand U37510 (N_37510,N_33234,N_33416);
and U37511 (N_37511,N_33637,N_31701);
nand U37512 (N_37512,N_31791,N_31437);
or U37513 (N_37513,N_32193,N_32255);
and U37514 (N_37514,N_31020,N_30026);
and U37515 (N_37515,N_30236,N_34433);
nor U37516 (N_37516,N_32658,N_34893);
or U37517 (N_37517,N_34120,N_31678);
xnor U37518 (N_37518,N_30057,N_33135);
nand U37519 (N_37519,N_30782,N_34058);
xnor U37520 (N_37520,N_30396,N_32868);
and U37521 (N_37521,N_33864,N_31231);
nand U37522 (N_37522,N_31238,N_30693);
xnor U37523 (N_37523,N_33619,N_31271);
or U37524 (N_37524,N_34310,N_30422);
and U37525 (N_37525,N_30176,N_30763);
and U37526 (N_37526,N_30008,N_33491);
xnor U37527 (N_37527,N_31572,N_30586);
and U37528 (N_37528,N_31189,N_31483);
or U37529 (N_37529,N_33487,N_32224);
xor U37530 (N_37530,N_30468,N_32224);
nand U37531 (N_37531,N_33786,N_32369);
nand U37532 (N_37532,N_30594,N_31090);
nor U37533 (N_37533,N_34528,N_30036);
or U37534 (N_37534,N_32775,N_34739);
or U37535 (N_37535,N_32939,N_34894);
xor U37536 (N_37536,N_33718,N_33725);
and U37537 (N_37537,N_34563,N_33563);
xor U37538 (N_37538,N_32574,N_33886);
nand U37539 (N_37539,N_31536,N_34423);
or U37540 (N_37540,N_32556,N_31887);
xnor U37541 (N_37541,N_34718,N_30993);
or U37542 (N_37542,N_32878,N_34796);
nand U37543 (N_37543,N_32242,N_30119);
nor U37544 (N_37544,N_30426,N_30519);
nor U37545 (N_37545,N_32044,N_34354);
nor U37546 (N_37546,N_33962,N_33001);
or U37547 (N_37547,N_34054,N_30761);
xnor U37548 (N_37548,N_33663,N_32163);
xnor U37549 (N_37549,N_32504,N_30215);
xor U37550 (N_37550,N_32146,N_33824);
xor U37551 (N_37551,N_32763,N_34609);
nor U37552 (N_37552,N_33992,N_33658);
xnor U37553 (N_37553,N_33256,N_31473);
nand U37554 (N_37554,N_31210,N_33123);
or U37555 (N_37555,N_34847,N_32232);
and U37556 (N_37556,N_34029,N_34221);
and U37557 (N_37557,N_33982,N_32666);
nand U37558 (N_37558,N_30166,N_32366);
nor U37559 (N_37559,N_30601,N_30511);
xnor U37560 (N_37560,N_33711,N_34676);
and U37561 (N_37561,N_30423,N_30894);
xor U37562 (N_37562,N_30239,N_31911);
xnor U37563 (N_37563,N_32363,N_31014);
nand U37564 (N_37564,N_33419,N_31439);
or U37565 (N_37565,N_34953,N_31825);
xor U37566 (N_37566,N_33148,N_34009);
and U37567 (N_37567,N_32805,N_30341);
xor U37568 (N_37568,N_31300,N_34984);
nand U37569 (N_37569,N_31315,N_34709);
nand U37570 (N_37570,N_32810,N_30538);
xnor U37571 (N_37571,N_33021,N_34037);
nand U37572 (N_37572,N_32079,N_33348);
nor U37573 (N_37573,N_32807,N_33334);
or U37574 (N_37574,N_30868,N_30315);
and U37575 (N_37575,N_31838,N_34472);
or U37576 (N_37576,N_31552,N_30821);
or U37577 (N_37577,N_31099,N_31945);
xor U37578 (N_37578,N_30276,N_30448);
nand U37579 (N_37579,N_32834,N_31522);
and U37580 (N_37580,N_33808,N_34765);
nor U37581 (N_37581,N_34712,N_32126);
nand U37582 (N_37582,N_31577,N_34983);
and U37583 (N_37583,N_34450,N_34273);
and U37584 (N_37584,N_33480,N_33401);
or U37585 (N_37585,N_31751,N_30629);
and U37586 (N_37586,N_33182,N_33990);
xor U37587 (N_37587,N_34437,N_33189);
or U37588 (N_37588,N_32311,N_31496);
or U37589 (N_37589,N_30128,N_33026);
or U37590 (N_37590,N_33826,N_34774);
nor U37591 (N_37591,N_31757,N_32869);
and U37592 (N_37592,N_34081,N_30526);
nand U37593 (N_37593,N_33022,N_31683);
nor U37594 (N_37594,N_33747,N_30885);
nor U37595 (N_37595,N_33379,N_34639);
nand U37596 (N_37596,N_33142,N_31214);
and U37597 (N_37597,N_31943,N_32032);
nand U37598 (N_37598,N_32075,N_33266);
or U37599 (N_37599,N_33703,N_31616);
nor U37600 (N_37600,N_33408,N_31335);
nand U37601 (N_37601,N_31208,N_30132);
nand U37602 (N_37602,N_32127,N_32913);
or U37603 (N_37603,N_31421,N_34716);
or U37604 (N_37604,N_33200,N_33169);
nor U37605 (N_37605,N_30142,N_31001);
nor U37606 (N_37606,N_33415,N_32740);
or U37607 (N_37607,N_32910,N_31153);
and U37608 (N_37608,N_31863,N_33334);
and U37609 (N_37609,N_34905,N_32850);
nand U37610 (N_37610,N_34019,N_31477);
or U37611 (N_37611,N_32434,N_34415);
nand U37612 (N_37612,N_31689,N_32977);
nor U37613 (N_37613,N_30941,N_31557);
nand U37614 (N_37614,N_34392,N_31882);
nor U37615 (N_37615,N_33448,N_31386);
xnor U37616 (N_37616,N_32997,N_30020);
and U37617 (N_37617,N_30568,N_30481);
or U37618 (N_37618,N_34170,N_32367);
and U37619 (N_37619,N_34658,N_32806);
nand U37620 (N_37620,N_32968,N_31643);
or U37621 (N_37621,N_32027,N_32717);
or U37622 (N_37622,N_33977,N_30078);
nand U37623 (N_37623,N_31513,N_30693);
xor U37624 (N_37624,N_30998,N_32334);
or U37625 (N_37625,N_31046,N_32982);
nand U37626 (N_37626,N_33069,N_33757);
nand U37627 (N_37627,N_34440,N_31776);
and U37628 (N_37628,N_34580,N_30358);
nor U37629 (N_37629,N_32521,N_31882);
nor U37630 (N_37630,N_31943,N_30098);
nor U37631 (N_37631,N_31963,N_34763);
nor U37632 (N_37632,N_31623,N_30085);
nor U37633 (N_37633,N_32302,N_33439);
xor U37634 (N_37634,N_32293,N_31595);
and U37635 (N_37635,N_34693,N_33548);
and U37636 (N_37636,N_32577,N_32618);
xor U37637 (N_37637,N_31676,N_34010);
nand U37638 (N_37638,N_34444,N_32072);
or U37639 (N_37639,N_34110,N_30808);
nand U37640 (N_37640,N_30421,N_31722);
xor U37641 (N_37641,N_33789,N_34085);
nor U37642 (N_37642,N_32261,N_32098);
and U37643 (N_37643,N_32957,N_32109);
and U37644 (N_37644,N_34733,N_31586);
and U37645 (N_37645,N_34925,N_30945);
or U37646 (N_37646,N_31442,N_32556);
nor U37647 (N_37647,N_31604,N_33349);
nor U37648 (N_37648,N_33128,N_34473);
nor U37649 (N_37649,N_33232,N_34511);
nor U37650 (N_37650,N_34047,N_34138);
nor U37651 (N_37651,N_31966,N_33486);
xnor U37652 (N_37652,N_30915,N_33237);
xnor U37653 (N_37653,N_32938,N_32832);
or U37654 (N_37654,N_31961,N_33904);
or U37655 (N_37655,N_32823,N_31589);
xor U37656 (N_37656,N_34565,N_34956);
nand U37657 (N_37657,N_34077,N_30186);
nand U37658 (N_37658,N_31267,N_30571);
nor U37659 (N_37659,N_33766,N_30835);
nor U37660 (N_37660,N_34985,N_30515);
and U37661 (N_37661,N_32091,N_33857);
or U37662 (N_37662,N_34399,N_34581);
nand U37663 (N_37663,N_30307,N_31643);
and U37664 (N_37664,N_30109,N_31727);
nand U37665 (N_37665,N_32277,N_33928);
xnor U37666 (N_37666,N_31058,N_34727);
xnor U37667 (N_37667,N_33647,N_30567);
and U37668 (N_37668,N_33473,N_30271);
or U37669 (N_37669,N_33582,N_30273);
and U37670 (N_37670,N_34509,N_33400);
and U37671 (N_37671,N_31488,N_34006);
or U37672 (N_37672,N_33031,N_34870);
or U37673 (N_37673,N_34274,N_33086);
xor U37674 (N_37674,N_31045,N_32613);
xnor U37675 (N_37675,N_30741,N_31727);
xor U37676 (N_37676,N_32322,N_32894);
xnor U37677 (N_37677,N_33506,N_32558);
and U37678 (N_37678,N_33597,N_33864);
nand U37679 (N_37679,N_32850,N_30111);
nand U37680 (N_37680,N_34543,N_32018);
nand U37681 (N_37681,N_33919,N_33899);
and U37682 (N_37682,N_34818,N_30373);
or U37683 (N_37683,N_31255,N_34505);
nor U37684 (N_37684,N_31783,N_34778);
xnor U37685 (N_37685,N_34705,N_32706);
or U37686 (N_37686,N_30606,N_31709);
or U37687 (N_37687,N_31731,N_34157);
or U37688 (N_37688,N_30832,N_30974);
xnor U37689 (N_37689,N_31255,N_32571);
or U37690 (N_37690,N_33916,N_31146);
nor U37691 (N_37691,N_34957,N_32444);
nor U37692 (N_37692,N_34062,N_33643);
nand U37693 (N_37693,N_34902,N_33786);
xnor U37694 (N_37694,N_30648,N_30839);
xnor U37695 (N_37695,N_34949,N_31163);
nand U37696 (N_37696,N_33947,N_34845);
nand U37697 (N_37697,N_31028,N_30580);
and U37698 (N_37698,N_34896,N_31103);
or U37699 (N_37699,N_31604,N_31205);
xnor U37700 (N_37700,N_34345,N_34985);
and U37701 (N_37701,N_32093,N_31021);
nor U37702 (N_37702,N_33679,N_30364);
nor U37703 (N_37703,N_31142,N_33563);
nor U37704 (N_37704,N_31890,N_30300);
xor U37705 (N_37705,N_33401,N_32249);
and U37706 (N_37706,N_32007,N_31282);
nand U37707 (N_37707,N_31152,N_31102);
or U37708 (N_37708,N_33683,N_33285);
nor U37709 (N_37709,N_33562,N_33940);
or U37710 (N_37710,N_33760,N_31980);
nor U37711 (N_37711,N_30799,N_32563);
and U37712 (N_37712,N_32132,N_32643);
and U37713 (N_37713,N_33272,N_31336);
nand U37714 (N_37714,N_31620,N_30897);
xor U37715 (N_37715,N_31793,N_33588);
nor U37716 (N_37716,N_32047,N_32694);
xor U37717 (N_37717,N_31847,N_33322);
nand U37718 (N_37718,N_32937,N_34984);
and U37719 (N_37719,N_30389,N_30462);
or U37720 (N_37720,N_34792,N_32933);
nand U37721 (N_37721,N_32914,N_33928);
xor U37722 (N_37722,N_34408,N_34043);
xnor U37723 (N_37723,N_34756,N_34886);
or U37724 (N_37724,N_33111,N_30473);
nor U37725 (N_37725,N_31915,N_34101);
nor U37726 (N_37726,N_33595,N_34584);
nand U37727 (N_37727,N_33387,N_33658);
and U37728 (N_37728,N_30382,N_31791);
and U37729 (N_37729,N_30359,N_33906);
nor U37730 (N_37730,N_32903,N_31693);
and U37731 (N_37731,N_33782,N_32984);
nor U37732 (N_37732,N_31814,N_30491);
or U37733 (N_37733,N_31007,N_33443);
nand U37734 (N_37734,N_31167,N_34065);
nor U37735 (N_37735,N_31753,N_33816);
or U37736 (N_37736,N_33375,N_30287);
and U37737 (N_37737,N_31977,N_30614);
and U37738 (N_37738,N_30140,N_34531);
xnor U37739 (N_37739,N_31526,N_30473);
nor U37740 (N_37740,N_30240,N_31189);
nor U37741 (N_37741,N_33880,N_33405);
and U37742 (N_37742,N_34102,N_31678);
or U37743 (N_37743,N_30348,N_31339);
nor U37744 (N_37744,N_30673,N_30628);
nand U37745 (N_37745,N_33825,N_34766);
nor U37746 (N_37746,N_33807,N_32584);
and U37747 (N_37747,N_30311,N_31418);
xnor U37748 (N_37748,N_33545,N_33040);
or U37749 (N_37749,N_31945,N_33007);
nor U37750 (N_37750,N_31696,N_30048);
nor U37751 (N_37751,N_31368,N_32265);
or U37752 (N_37752,N_34948,N_30271);
nand U37753 (N_37753,N_30915,N_30211);
nand U37754 (N_37754,N_33308,N_32298);
and U37755 (N_37755,N_32341,N_34290);
xnor U37756 (N_37756,N_33632,N_33362);
nand U37757 (N_37757,N_32729,N_34199);
nor U37758 (N_37758,N_30400,N_31576);
nand U37759 (N_37759,N_34713,N_32074);
nand U37760 (N_37760,N_31275,N_30509);
or U37761 (N_37761,N_30638,N_33157);
xor U37762 (N_37762,N_32443,N_30275);
and U37763 (N_37763,N_34034,N_33692);
or U37764 (N_37764,N_30211,N_34212);
xor U37765 (N_37765,N_31400,N_33119);
xor U37766 (N_37766,N_34109,N_32528);
nor U37767 (N_37767,N_32898,N_30905);
nand U37768 (N_37768,N_33705,N_31906);
or U37769 (N_37769,N_34261,N_34580);
nor U37770 (N_37770,N_34059,N_33992);
nor U37771 (N_37771,N_30554,N_31725);
or U37772 (N_37772,N_32603,N_31681);
xor U37773 (N_37773,N_33975,N_30648);
xnor U37774 (N_37774,N_32821,N_30589);
or U37775 (N_37775,N_30551,N_32432);
nand U37776 (N_37776,N_32740,N_32634);
nand U37777 (N_37777,N_31693,N_32720);
nand U37778 (N_37778,N_31261,N_31662);
nand U37779 (N_37779,N_30201,N_34788);
and U37780 (N_37780,N_33834,N_32400);
nor U37781 (N_37781,N_34293,N_32617);
or U37782 (N_37782,N_33003,N_31407);
and U37783 (N_37783,N_33659,N_30466);
or U37784 (N_37784,N_30868,N_34830);
nor U37785 (N_37785,N_30690,N_30952);
xnor U37786 (N_37786,N_33758,N_30581);
xnor U37787 (N_37787,N_33864,N_33951);
nand U37788 (N_37788,N_34052,N_31502);
or U37789 (N_37789,N_30238,N_32399);
nand U37790 (N_37790,N_33620,N_32764);
nand U37791 (N_37791,N_33181,N_34153);
and U37792 (N_37792,N_30027,N_31419);
nand U37793 (N_37793,N_32928,N_31446);
nand U37794 (N_37794,N_30956,N_33255);
nand U37795 (N_37795,N_33386,N_33261);
and U37796 (N_37796,N_32942,N_33060);
xnor U37797 (N_37797,N_30181,N_34176);
nor U37798 (N_37798,N_34841,N_32424);
and U37799 (N_37799,N_34336,N_34543);
and U37800 (N_37800,N_32707,N_34904);
and U37801 (N_37801,N_32087,N_32671);
nor U37802 (N_37802,N_31064,N_34489);
or U37803 (N_37803,N_32561,N_30768);
nand U37804 (N_37804,N_33439,N_31034);
or U37805 (N_37805,N_31826,N_34364);
xnor U37806 (N_37806,N_32778,N_31163);
and U37807 (N_37807,N_32085,N_31194);
and U37808 (N_37808,N_31264,N_30454);
nor U37809 (N_37809,N_32214,N_32792);
nand U37810 (N_37810,N_34249,N_31943);
and U37811 (N_37811,N_31690,N_33601);
and U37812 (N_37812,N_30076,N_34176);
nor U37813 (N_37813,N_34281,N_30970);
nand U37814 (N_37814,N_32086,N_33697);
nand U37815 (N_37815,N_30797,N_30988);
xor U37816 (N_37816,N_34882,N_33890);
xor U37817 (N_37817,N_34943,N_32480);
and U37818 (N_37818,N_34901,N_31257);
or U37819 (N_37819,N_33579,N_31776);
and U37820 (N_37820,N_30667,N_34601);
and U37821 (N_37821,N_33337,N_31186);
nor U37822 (N_37822,N_31019,N_30037);
nor U37823 (N_37823,N_32794,N_31372);
nor U37824 (N_37824,N_32229,N_32878);
or U37825 (N_37825,N_30398,N_33902);
and U37826 (N_37826,N_30761,N_30154);
nand U37827 (N_37827,N_31493,N_33640);
or U37828 (N_37828,N_34511,N_33750);
nor U37829 (N_37829,N_33306,N_31476);
nand U37830 (N_37830,N_34210,N_33697);
nor U37831 (N_37831,N_30432,N_32251);
nor U37832 (N_37832,N_34182,N_32116);
xnor U37833 (N_37833,N_32481,N_34009);
or U37834 (N_37834,N_34526,N_30168);
nor U37835 (N_37835,N_33640,N_31470);
nand U37836 (N_37836,N_34219,N_32585);
xor U37837 (N_37837,N_33454,N_31698);
or U37838 (N_37838,N_31311,N_34206);
nand U37839 (N_37839,N_34314,N_34233);
xor U37840 (N_37840,N_31229,N_33343);
and U37841 (N_37841,N_33775,N_32594);
or U37842 (N_37842,N_30784,N_32101);
and U37843 (N_37843,N_31687,N_34525);
and U37844 (N_37844,N_33587,N_33038);
and U37845 (N_37845,N_30701,N_31708);
nand U37846 (N_37846,N_30943,N_34720);
nand U37847 (N_37847,N_34196,N_31590);
or U37848 (N_37848,N_33355,N_33038);
nand U37849 (N_37849,N_33391,N_32706);
or U37850 (N_37850,N_33755,N_33058);
or U37851 (N_37851,N_31477,N_31969);
nor U37852 (N_37852,N_30395,N_32362);
and U37853 (N_37853,N_30752,N_33190);
or U37854 (N_37854,N_31643,N_34172);
nor U37855 (N_37855,N_30425,N_33987);
nor U37856 (N_37856,N_33026,N_30142);
or U37857 (N_37857,N_31194,N_34212);
nor U37858 (N_37858,N_32336,N_32384);
or U37859 (N_37859,N_30133,N_32078);
xor U37860 (N_37860,N_30005,N_32992);
and U37861 (N_37861,N_31326,N_33999);
xnor U37862 (N_37862,N_32154,N_34881);
nor U37863 (N_37863,N_32826,N_33648);
xnor U37864 (N_37864,N_31556,N_31021);
nand U37865 (N_37865,N_30037,N_34142);
xnor U37866 (N_37866,N_33878,N_31581);
and U37867 (N_37867,N_34599,N_32845);
and U37868 (N_37868,N_31784,N_31182);
and U37869 (N_37869,N_31423,N_30475);
or U37870 (N_37870,N_30838,N_31829);
nand U37871 (N_37871,N_34484,N_32728);
nand U37872 (N_37872,N_34987,N_32526);
nor U37873 (N_37873,N_33546,N_32357);
or U37874 (N_37874,N_32373,N_30628);
nor U37875 (N_37875,N_34240,N_33047);
and U37876 (N_37876,N_32375,N_30245);
nor U37877 (N_37877,N_33162,N_33953);
and U37878 (N_37878,N_34431,N_31379);
or U37879 (N_37879,N_34143,N_34777);
xor U37880 (N_37880,N_33868,N_31572);
nor U37881 (N_37881,N_32705,N_30292);
and U37882 (N_37882,N_33522,N_31671);
or U37883 (N_37883,N_32107,N_34171);
nand U37884 (N_37884,N_34492,N_32890);
and U37885 (N_37885,N_30787,N_33446);
and U37886 (N_37886,N_33306,N_32461);
nor U37887 (N_37887,N_33589,N_34388);
or U37888 (N_37888,N_34700,N_34577);
or U37889 (N_37889,N_31405,N_31868);
or U37890 (N_37890,N_33949,N_33270);
and U37891 (N_37891,N_33986,N_30941);
nor U37892 (N_37892,N_32436,N_33598);
nand U37893 (N_37893,N_30249,N_31431);
and U37894 (N_37894,N_34524,N_33728);
nand U37895 (N_37895,N_33636,N_30950);
and U37896 (N_37896,N_31832,N_33517);
nor U37897 (N_37897,N_32819,N_32397);
xnor U37898 (N_37898,N_34927,N_32920);
or U37899 (N_37899,N_30030,N_34115);
or U37900 (N_37900,N_30545,N_32703);
nand U37901 (N_37901,N_30152,N_30514);
nor U37902 (N_37902,N_33762,N_34443);
and U37903 (N_37903,N_34525,N_33753);
nor U37904 (N_37904,N_33153,N_30035);
xor U37905 (N_37905,N_32879,N_33379);
xor U37906 (N_37906,N_30081,N_31918);
nand U37907 (N_37907,N_34904,N_30912);
nand U37908 (N_37908,N_33327,N_30514);
nor U37909 (N_37909,N_30887,N_32028);
and U37910 (N_37910,N_34335,N_33233);
or U37911 (N_37911,N_32028,N_32730);
or U37912 (N_37912,N_30127,N_34252);
or U37913 (N_37913,N_33505,N_32379);
or U37914 (N_37914,N_31605,N_30484);
or U37915 (N_37915,N_33874,N_34447);
xor U37916 (N_37916,N_33541,N_34468);
or U37917 (N_37917,N_34362,N_31020);
xor U37918 (N_37918,N_33618,N_32328);
xnor U37919 (N_37919,N_31123,N_34417);
nor U37920 (N_37920,N_31944,N_31662);
nand U37921 (N_37921,N_30433,N_31575);
xnor U37922 (N_37922,N_33021,N_32015);
and U37923 (N_37923,N_34243,N_34270);
nor U37924 (N_37924,N_31959,N_30842);
nand U37925 (N_37925,N_31371,N_31409);
nor U37926 (N_37926,N_30902,N_30018);
and U37927 (N_37927,N_31975,N_34817);
or U37928 (N_37928,N_32644,N_33881);
and U37929 (N_37929,N_34103,N_32480);
nand U37930 (N_37930,N_34049,N_30331);
and U37931 (N_37931,N_30743,N_32494);
nand U37932 (N_37932,N_33195,N_30579);
and U37933 (N_37933,N_34848,N_31772);
xor U37934 (N_37934,N_34827,N_30004);
nand U37935 (N_37935,N_34913,N_34785);
nor U37936 (N_37936,N_31472,N_33517);
nor U37937 (N_37937,N_30335,N_34610);
nand U37938 (N_37938,N_33278,N_31472);
xnor U37939 (N_37939,N_32253,N_32723);
nor U37940 (N_37940,N_31008,N_31232);
and U37941 (N_37941,N_32278,N_31166);
and U37942 (N_37942,N_31563,N_33184);
xor U37943 (N_37943,N_34844,N_30133);
xnor U37944 (N_37944,N_33938,N_31279);
xnor U37945 (N_37945,N_32708,N_32459);
or U37946 (N_37946,N_33280,N_31125);
xor U37947 (N_37947,N_31987,N_32044);
or U37948 (N_37948,N_31345,N_30518);
nor U37949 (N_37949,N_31322,N_34763);
or U37950 (N_37950,N_31681,N_33625);
or U37951 (N_37951,N_31047,N_30666);
xnor U37952 (N_37952,N_32245,N_32666);
nor U37953 (N_37953,N_30535,N_34671);
and U37954 (N_37954,N_32996,N_33752);
and U37955 (N_37955,N_33147,N_33971);
xor U37956 (N_37956,N_30604,N_33033);
or U37957 (N_37957,N_33375,N_33961);
xnor U37958 (N_37958,N_30021,N_30314);
xnor U37959 (N_37959,N_31956,N_32429);
or U37960 (N_37960,N_30297,N_32567);
and U37961 (N_37961,N_31807,N_31059);
xor U37962 (N_37962,N_30799,N_32074);
nand U37963 (N_37963,N_33946,N_34798);
or U37964 (N_37964,N_33185,N_34093);
nand U37965 (N_37965,N_33067,N_30522);
and U37966 (N_37966,N_30553,N_33855);
and U37967 (N_37967,N_34103,N_34903);
and U37968 (N_37968,N_32804,N_32680);
nor U37969 (N_37969,N_34986,N_30934);
and U37970 (N_37970,N_32327,N_32814);
nand U37971 (N_37971,N_32397,N_30666);
nand U37972 (N_37972,N_30546,N_33969);
nand U37973 (N_37973,N_33304,N_31138);
xor U37974 (N_37974,N_32725,N_33228);
and U37975 (N_37975,N_31378,N_33388);
and U37976 (N_37976,N_32773,N_34245);
nand U37977 (N_37977,N_32233,N_30891);
nand U37978 (N_37978,N_33933,N_34264);
or U37979 (N_37979,N_33873,N_33453);
and U37980 (N_37980,N_31300,N_33415);
xor U37981 (N_37981,N_30346,N_30527);
nand U37982 (N_37982,N_34548,N_34137);
xor U37983 (N_37983,N_33419,N_31377);
nor U37984 (N_37984,N_30374,N_32333);
or U37985 (N_37985,N_32131,N_33972);
or U37986 (N_37986,N_34833,N_33271);
xnor U37987 (N_37987,N_31987,N_33404);
and U37988 (N_37988,N_34330,N_34780);
or U37989 (N_37989,N_31057,N_33180);
xnor U37990 (N_37990,N_32410,N_30606);
nor U37991 (N_37991,N_30089,N_31542);
xnor U37992 (N_37992,N_33296,N_30575);
or U37993 (N_37993,N_31008,N_32948);
and U37994 (N_37994,N_33737,N_34747);
or U37995 (N_37995,N_31738,N_30254);
xnor U37996 (N_37996,N_31728,N_34630);
nand U37997 (N_37997,N_33498,N_34527);
or U37998 (N_37998,N_34003,N_31214);
and U37999 (N_37999,N_32819,N_32419);
nand U38000 (N_38000,N_33824,N_33496);
and U38001 (N_38001,N_31866,N_32974);
nor U38002 (N_38002,N_31334,N_30223);
nor U38003 (N_38003,N_34367,N_31660);
or U38004 (N_38004,N_32418,N_31236);
nand U38005 (N_38005,N_34775,N_30249);
or U38006 (N_38006,N_33521,N_32278);
nor U38007 (N_38007,N_32672,N_31624);
xor U38008 (N_38008,N_33622,N_32744);
nor U38009 (N_38009,N_32783,N_32933);
nor U38010 (N_38010,N_32802,N_31862);
and U38011 (N_38011,N_34800,N_30964);
or U38012 (N_38012,N_34515,N_32447);
nor U38013 (N_38013,N_32014,N_33794);
nand U38014 (N_38014,N_31938,N_34361);
or U38015 (N_38015,N_30566,N_32294);
nor U38016 (N_38016,N_31020,N_30352);
xor U38017 (N_38017,N_31254,N_31190);
nor U38018 (N_38018,N_30722,N_32102);
or U38019 (N_38019,N_31412,N_32296);
and U38020 (N_38020,N_33617,N_34200);
nor U38021 (N_38021,N_34123,N_31976);
xnor U38022 (N_38022,N_34005,N_34877);
and U38023 (N_38023,N_34861,N_33597);
xor U38024 (N_38024,N_31197,N_34450);
nand U38025 (N_38025,N_31202,N_32731);
nand U38026 (N_38026,N_33999,N_31126);
and U38027 (N_38027,N_34520,N_31436);
and U38028 (N_38028,N_32299,N_30180);
xor U38029 (N_38029,N_30310,N_30978);
nand U38030 (N_38030,N_32097,N_34347);
nor U38031 (N_38031,N_30859,N_31309);
xor U38032 (N_38032,N_33948,N_30266);
xor U38033 (N_38033,N_31733,N_34839);
xor U38034 (N_38034,N_30083,N_31486);
xnor U38035 (N_38035,N_30564,N_31079);
nor U38036 (N_38036,N_34607,N_34308);
xnor U38037 (N_38037,N_32233,N_31300);
xnor U38038 (N_38038,N_30120,N_31963);
nor U38039 (N_38039,N_33927,N_32367);
and U38040 (N_38040,N_34006,N_33885);
and U38041 (N_38041,N_30175,N_34057);
nor U38042 (N_38042,N_30395,N_34621);
xor U38043 (N_38043,N_31497,N_31069);
and U38044 (N_38044,N_34806,N_30557);
or U38045 (N_38045,N_31378,N_30477);
and U38046 (N_38046,N_30636,N_31077);
xnor U38047 (N_38047,N_31714,N_31448);
nand U38048 (N_38048,N_32767,N_33537);
nand U38049 (N_38049,N_34524,N_31447);
nand U38050 (N_38050,N_34914,N_30223);
and U38051 (N_38051,N_34855,N_31949);
xnor U38052 (N_38052,N_34369,N_34786);
xor U38053 (N_38053,N_34508,N_31533);
nand U38054 (N_38054,N_30385,N_31756);
nor U38055 (N_38055,N_30010,N_31231);
xor U38056 (N_38056,N_34685,N_31860);
nand U38057 (N_38057,N_34478,N_33633);
nor U38058 (N_38058,N_30542,N_32209);
nor U38059 (N_38059,N_30618,N_32957);
nor U38060 (N_38060,N_30131,N_32424);
xor U38061 (N_38061,N_33485,N_30439);
nor U38062 (N_38062,N_33244,N_33618);
xor U38063 (N_38063,N_31322,N_30981);
or U38064 (N_38064,N_31409,N_34973);
nand U38065 (N_38065,N_33083,N_33944);
nand U38066 (N_38066,N_31929,N_34800);
nand U38067 (N_38067,N_32483,N_34655);
nor U38068 (N_38068,N_33499,N_34690);
or U38069 (N_38069,N_34655,N_34441);
or U38070 (N_38070,N_34525,N_33097);
xnor U38071 (N_38071,N_30329,N_34590);
nand U38072 (N_38072,N_30862,N_31957);
and U38073 (N_38073,N_33221,N_31721);
xor U38074 (N_38074,N_34555,N_34799);
nand U38075 (N_38075,N_32546,N_30897);
xnor U38076 (N_38076,N_31774,N_32853);
xor U38077 (N_38077,N_31269,N_34152);
and U38078 (N_38078,N_30082,N_31693);
and U38079 (N_38079,N_34562,N_32933);
or U38080 (N_38080,N_33938,N_32011);
nand U38081 (N_38081,N_32966,N_34695);
xor U38082 (N_38082,N_31402,N_30377);
or U38083 (N_38083,N_34667,N_32467);
nor U38084 (N_38084,N_30595,N_31513);
nand U38085 (N_38085,N_33230,N_30849);
nand U38086 (N_38086,N_32803,N_30303);
nand U38087 (N_38087,N_30110,N_31094);
and U38088 (N_38088,N_33741,N_32303);
nand U38089 (N_38089,N_31102,N_30129);
or U38090 (N_38090,N_34165,N_31150);
or U38091 (N_38091,N_34421,N_31245);
or U38092 (N_38092,N_30867,N_33316);
or U38093 (N_38093,N_30975,N_34172);
or U38094 (N_38094,N_30191,N_30002);
nor U38095 (N_38095,N_32993,N_33226);
or U38096 (N_38096,N_32617,N_31516);
nand U38097 (N_38097,N_32936,N_32585);
nand U38098 (N_38098,N_33044,N_34947);
or U38099 (N_38099,N_31642,N_33416);
xnor U38100 (N_38100,N_30437,N_32640);
nor U38101 (N_38101,N_30070,N_30736);
and U38102 (N_38102,N_30765,N_34382);
nand U38103 (N_38103,N_33401,N_32618);
xor U38104 (N_38104,N_32395,N_33914);
nor U38105 (N_38105,N_34276,N_32603);
nand U38106 (N_38106,N_33321,N_30152);
and U38107 (N_38107,N_34211,N_30822);
nor U38108 (N_38108,N_33488,N_32432);
nor U38109 (N_38109,N_32390,N_31075);
or U38110 (N_38110,N_32422,N_34081);
or U38111 (N_38111,N_32105,N_33122);
nor U38112 (N_38112,N_33078,N_32940);
nand U38113 (N_38113,N_30168,N_31736);
xor U38114 (N_38114,N_31947,N_32607);
nor U38115 (N_38115,N_30707,N_33325);
or U38116 (N_38116,N_34102,N_34535);
nand U38117 (N_38117,N_34521,N_32511);
nand U38118 (N_38118,N_34179,N_34909);
xnor U38119 (N_38119,N_30294,N_33317);
nor U38120 (N_38120,N_31058,N_33459);
nand U38121 (N_38121,N_34960,N_34947);
xor U38122 (N_38122,N_34481,N_30897);
nor U38123 (N_38123,N_34699,N_30132);
and U38124 (N_38124,N_33443,N_34618);
or U38125 (N_38125,N_33732,N_30558);
and U38126 (N_38126,N_34526,N_32754);
or U38127 (N_38127,N_33210,N_32704);
or U38128 (N_38128,N_33323,N_32768);
or U38129 (N_38129,N_34830,N_31884);
nand U38130 (N_38130,N_32949,N_33390);
or U38131 (N_38131,N_31604,N_34439);
or U38132 (N_38132,N_31822,N_33178);
and U38133 (N_38133,N_34517,N_34939);
xor U38134 (N_38134,N_33679,N_30645);
xnor U38135 (N_38135,N_31106,N_33409);
or U38136 (N_38136,N_31636,N_32000);
xnor U38137 (N_38137,N_34060,N_32437);
nor U38138 (N_38138,N_33806,N_31349);
or U38139 (N_38139,N_32163,N_33964);
and U38140 (N_38140,N_34639,N_31599);
and U38141 (N_38141,N_31680,N_33084);
or U38142 (N_38142,N_30564,N_30252);
xnor U38143 (N_38143,N_30273,N_33650);
and U38144 (N_38144,N_31729,N_32805);
xnor U38145 (N_38145,N_30752,N_31604);
nand U38146 (N_38146,N_33866,N_32740);
nand U38147 (N_38147,N_34938,N_31657);
nand U38148 (N_38148,N_32227,N_34572);
nand U38149 (N_38149,N_34744,N_33888);
nor U38150 (N_38150,N_31508,N_32267);
and U38151 (N_38151,N_33480,N_30956);
xor U38152 (N_38152,N_30183,N_31902);
nand U38153 (N_38153,N_34424,N_31125);
nor U38154 (N_38154,N_32260,N_33929);
nor U38155 (N_38155,N_32693,N_34266);
nand U38156 (N_38156,N_32475,N_32935);
nand U38157 (N_38157,N_30570,N_34032);
or U38158 (N_38158,N_32120,N_32298);
xor U38159 (N_38159,N_30892,N_30834);
nand U38160 (N_38160,N_31692,N_32793);
or U38161 (N_38161,N_32141,N_34290);
or U38162 (N_38162,N_32031,N_34968);
and U38163 (N_38163,N_32085,N_30013);
xor U38164 (N_38164,N_34659,N_31854);
or U38165 (N_38165,N_34160,N_30647);
xnor U38166 (N_38166,N_31794,N_34038);
xnor U38167 (N_38167,N_33729,N_30236);
nor U38168 (N_38168,N_33437,N_34559);
or U38169 (N_38169,N_32634,N_34598);
nor U38170 (N_38170,N_31121,N_30536);
nand U38171 (N_38171,N_33784,N_32371);
xnor U38172 (N_38172,N_31004,N_34046);
and U38173 (N_38173,N_32862,N_32475);
nor U38174 (N_38174,N_32069,N_33323);
nor U38175 (N_38175,N_33071,N_33153);
nor U38176 (N_38176,N_33636,N_34789);
and U38177 (N_38177,N_31479,N_31622);
or U38178 (N_38178,N_33456,N_32582);
or U38179 (N_38179,N_32012,N_32157);
nor U38180 (N_38180,N_32744,N_32038);
or U38181 (N_38181,N_32538,N_34328);
nand U38182 (N_38182,N_34884,N_30938);
xnor U38183 (N_38183,N_32694,N_34655);
xor U38184 (N_38184,N_32096,N_33575);
and U38185 (N_38185,N_34942,N_33937);
or U38186 (N_38186,N_34584,N_33936);
and U38187 (N_38187,N_31284,N_32057);
xor U38188 (N_38188,N_30316,N_34157);
nor U38189 (N_38189,N_30587,N_31729);
nor U38190 (N_38190,N_34213,N_32331);
and U38191 (N_38191,N_32389,N_31930);
nand U38192 (N_38192,N_34464,N_33172);
and U38193 (N_38193,N_30786,N_33570);
and U38194 (N_38194,N_31877,N_32124);
nor U38195 (N_38195,N_33457,N_34471);
or U38196 (N_38196,N_31327,N_34984);
xor U38197 (N_38197,N_33536,N_33848);
xnor U38198 (N_38198,N_32318,N_33362);
nor U38199 (N_38199,N_31197,N_30921);
nand U38200 (N_38200,N_34315,N_31356);
and U38201 (N_38201,N_32865,N_31768);
or U38202 (N_38202,N_31562,N_33566);
or U38203 (N_38203,N_32474,N_30756);
or U38204 (N_38204,N_34444,N_31648);
nor U38205 (N_38205,N_34006,N_30184);
nand U38206 (N_38206,N_31699,N_31500);
nand U38207 (N_38207,N_30177,N_33691);
xnor U38208 (N_38208,N_33294,N_33377);
or U38209 (N_38209,N_32018,N_30555);
and U38210 (N_38210,N_33709,N_32233);
nand U38211 (N_38211,N_31602,N_32572);
and U38212 (N_38212,N_31040,N_30584);
or U38213 (N_38213,N_32131,N_31869);
or U38214 (N_38214,N_34319,N_33907);
nor U38215 (N_38215,N_31920,N_31627);
nand U38216 (N_38216,N_32745,N_31708);
xnor U38217 (N_38217,N_33572,N_33224);
nand U38218 (N_38218,N_34465,N_31890);
nor U38219 (N_38219,N_33667,N_31702);
nand U38220 (N_38220,N_31972,N_33849);
or U38221 (N_38221,N_33583,N_30453);
and U38222 (N_38222,N_30454,N_31597);
nor U38223 (N_38223,N_30822,N_32000);
or U38224 (N_38224,N_32661,N_33700);
nand U38225 (N_38225,N_33347,N_32296);
xnor U38226 (N_38226,N_31146,N_33833);
or U38227 (N_38227,N_30674,N_34342);
nor U38228 (N_38228,N_31302,N_33790);
or U38229 (N_38229,N_33409,N_30419);
or U38230 (N_38230,N_34846,N_34134);
nor U38231 (N_38231,N_30482,N_33090);
xor U38232 (N_38232,N_31015,N_32382);
nand U38233 (N_38233,N_31713,N_30639);
nand U38234 (N_38234,N_34034,N_30132);
and U38235 (N_38235,N_30637,N_30968);
or U38236 (N_38236,N_34334,N_33985);
nor U38237 (N_38237,N_34205,N_31132);
and U38238 (N_38238,N_30950,N_31082);
nand U38239 (N_38239,N_34934,N_31888);
and U38240 (N_38240,N_34312,N_32715);
or U38241 (N_38241,N_32293,N_30196);
xor U38242 (N_38242,N_30534,N_32587);
nor U38243 (N_38243,N_30550,N_30222);
or U38244 (N_38244,N_33587,N_33325);
xor U38245 (N_38245,N_33628,N_33151);
nor U38246 (N_38246,N_31157,N_33094);
and U38247 (N_38247,N_34824,N_30138);
nor U38248 (N_38248,N_31824,N_32454);
or U38249 (N_38249,N_31148,N_31020);
and U38250 (N_38250,N_32223,N_33922);
or U38251 (N_38251,N_30368,N_33017);
nand U38252 (N_38252,N_30589,N_31446);
or U38253 (N_38253,N_33141,N_30668);
nor U38254 (N_38254,N_31131,N_32886);
nor U38255 (N_38255,N_30171,N_30744);
and U38256 (N_38256,N_33393,N_30440);
nor U38257 (N_38257,N_30509,N_32852);
or U38258 (N_38258,N_34574,N_33672);
nand U38259 (N_38259,N_32666,N_33957);
xor U38260 (N_38260,N_31528,N_33808);
and U38261 (N_38261,N_30366,N_31464);
xnor U38262 (N_38262,N_34798,N_32996);
xor U38263 (N_38263,N_30315,N_33847);
or U38264 (N_38264,N_33204,N_33812);
or U38265 (N_38265,N_34892,N_33681);
nand U38266 (N_38266,N_31085,N_31991);
nand U38267 (N_38267,N_31784,N_32015);
nand U38268 (N_38268,N_31648,N_33130);
xor U38269 (N_38269,N_30777,N_33393);
nand U38270 (N_38270,N_34422,N_30596);
nor U38271 (N_38271,N_34162,N_30851);
or U38272 (N_38272,N_34132,N_32728);
nor U38273 (N_38273,N_33967,N_30331);
nand U38274 (N_38274,N_34731,N_34501);
nand U38275 (N_38275,N_34443,N_33599);
or U38276 (N_38276,N_32188,N_32073);
nor U38277 (N_38277,N_34477,N_31295);
xor U38278 (N_38278,N_30608,N_33742);
and U38279 (N_38279,N_33606,N_31372);
and U38280 (N_38280,N_30456,N_31564);
nor U38281 (N_38281,N_30021,N_30232);
and U38282 (N_38282,N_32237,N_33521);
nand U38283 (N_38283,N_30852,N_32767);
nand U38284 (N_38284,N_33774,N_33219);
nor U38285 (N_38285,N_31833,N_30057);
nand U38286 (N_38286,N_30170,N_33049);
nand U38287 (N_38287,N_31299,N_34468);
or U38288 (N_38288,N_31094,N_34062);
nor U38289 (N_38289,N_31712,N_34822);
or U38290 (N_38290,N_34476,N_31033);
nor U38291 (N_38291,N_32443,N_32173);
and U38292 (N_38292,N_32242,N_30345);
nor U38293 (N_38293,N_33106,N_32617);
or U38294 (N_38294,N_33883,N_30933);
or U38295 (N_38295,N_31743,N_31855);
and U38296 (N_38296,N_31618,N_32702);
or U38297 (N_38297,N_32305,N_31682);
and U38298 (N_38298,N_32199,N_30661);
and U38299 (N_38299,N_31381,N_33891);
xor U38300 (N_38300,N_32887,N_32846);
xnor U38301 (N_38301,N_31492,N_32246);
and U38302 (N_38302,N_30501,N_34788);
nand U38303 (N_38303,N_33519,N_34005);
and U38304 (N_38304,N_33172,N_31259);
or U38305 (N_38305,N_34652,N_30504);
nor U38306 (N_38306,N_33224,N_31036);
and U38307 (N_38307,N_31515,N_34653);
or U38308 (N_38308,N_30642,N_34873);
or U38309 (N_38309,N_34112,N_33797);
nor U38310 (N_38310,N_33590,N_31017);
nor U38311 (N_38311,N_30961,N_31799);
xnor U38312 (N_38312,N_32494,N_30551);
xnor U38313 (N_38313,N_33062,N_30411);
and U38314 (N_38314,N_32864,N_30623);
nand U38315 (N_38315,N_31824,N_34255);
xnor U38316 (N_38316,N_31021,N_34427);
or U38317 (N_38317,N_31519,N_31593);
nor U38318 (N_38318,N_32464,N_34551);
nor U38319 (N_38319,N_34347,N_34255);
nand U38320 (N_38320,N_34825,N_31787);
nor U38321 (N_38321,N_30884,N_33513);
nor U38322 (N_38322,N_34144,N_31634);
nor U38323 (N_38323,N_32125,N_34650);
and U38324 (N_38324,N_31869,N_33992);
nand U38325 (N_38325,N_34947,N_31332);
xor U38326 (N_38326,N_33229,N_33193);
and U38327 (N_38327,N_32548,N_30885);
xor U38328 (N_38328,N_33373,N_33641);
nor U38329 (N_38329,N_32004,N_31896);
nand U38330 (N_38330,N_31046,N_32731);
and U38331 (N_38331,N_32959,N_32850);
nor U38332 (N_38332,N_30161,N_33946);
or U38333 (N_38333,N_34098,N_31256);
or U38334 (N_38334,N_33036,N_32745);
nand U38335 (N_38335,N_31043,N_31182);
and U38336 (N_38336,N_31039,N_32867);
xnor U38337 (N_38337,N_32557,N_30626);
nor U38338 (N_38338,N_31214,N_31444);
nand U38339 (N_38339,N_34712,N_33352);
xnor U38340 (N_38340,N_31879,N_30504);
nand U38341 (N_38341,N_31308,N_30344);
nand U38342 (N_38342,N_31400,N_31052);
or U38343 (N_38343,N_30101,N_33110);
nand U38344 (N_38344,N_31376,N_30807);
nor U38345 (N_38345,N_31746,N_31404);
and U38346 (N_38346,N_32913,N_31875);
nor U38347 (N_38347,N_33233,N_33604);
and U38348 (N_38348,N_30480,N_34985);
nand U38349 (N_38349,N_33592,N_34644);
nand U38350 (N_38350,N_33888,N_32746);
and U38351 (N_38351,N_32784,N_33746);
xor U38352 (N_38352,N_30986,N_32215);
nand U38353 (N_38353,N_34173,N_34110);
xor U38354 (N_38354,N_34080,N_33994);
and U38355 (N_38355,N_30725,N_33643);
nor U38356 (N_38356,N_34038,N_31224);
or U38357 (N_38357,N_30356,N_30855);
nand U38358 (N_38358,N_31789,N_31920);
nand U38359 (N_38359,N_32513,N_30414);
nand U38360 (N_38360,N_31454,N_30222);
nor U38361 (N_38361,N_32599,N_34133);
and U38362 (N_38362,N_34765,N_30538);
xor U38363 (N_38363,N_30742,N_32639);
or U38364 (N_38364,N_33175,N_34121);
xor U38365 (N_38365,N_33178,N_34896);
nor U38366 (N_38366,N_34889,N_34706);
nor U38367 (N_38367,N_33358,N_32952);
and U38368 (N_38368,N_30812,N_31987);
and U38369 (N_38369,N_32925,N_34772);
nor U38370 (N_38370,N_34275,N_33704);
and U38371 (N_38371,N_30449,N_30450);
xor U38372 (N_38372,N_31510,N_33063);
nand U38373 (N_38373,N_30793,N_30042);
nor U38374 (N_38374,N_31169,N_30446);
and U38375 (N_38375,N_30256,N_31581);
xnor U38376 (N_38376,N_34666,N_31171);
nor U38377 (N_38377,N_30927,N_34439);
nand U38378 (N_38378,N_31890,N_33847);
or U38379 (N_38379,N_32195,N_32697);
xor U38380 (N_38380,N_32455,N_32521);
xnor U38381 (N_38381,N_33189,N_31823);
nor U38382 (N_38382,N_30209,N_31389);
nand U38383 (N_38383,N_30351,N_32622);
and U38384 (N_38384,N_33385,N_34898);
xor U38385 (N_38385,N_32888,N_33872);
and U38386 (N_38386,N_32158,N_34560);
nand U38387 (N_38387,N_34671,N_31634);
nand U38388 (N_38388,N_30864,N_32020);
xnor U38389 (N_38389,N_30400,N_30265);
and U38390 (N_38390,N_31007,N_33123);
and U38391 (N_38391,N_30195,N_34081);
or U38392 (N_38392,N_33623,N_31681);
and U38393 (N_38393,N_33726,N_30438);
or U38394 (N_38394,N_31516,N_34087);
nor U38395 (N_38395,N_32598,N_33131);
nor U38396 (N_38396,N_31496,N_30263);
nand U38397 (N_38397,N_34875,N_34985);
nand U38398 (N_38398,N_31087,N_32317);
nor U38399 (N_38399,N_31457,N_30365);
nor U38400 (N_38400,N_30260,N_30719);
nand U38401 (N_38401,N_31117,N_31531);
nand U38402 (N_38402,N_32430,N_31247);
and U38403 (N_38403,N_30171,N_34630);
nor U38404 (N_38404,N_33100,N_34406);
nand U38405 (N_38405,N_32342,N_32065);
nor U38406 (N_38406,N_31631,N_30054);
nand U38407 (N_38407,N_34917,N_30045);
or U38408 (N_38408,N_30915,N_31684);
xnor U38409 (N_38409,N_31241,N_32428);
xnor U38410 (N_38410,N_33467,N_33257);
or U38411 (N_38411,N_34415,N_33369);
xor U38412 (N_38412,N_31421,N_33901);
xor U38413 (N_38413,N_34379,N_30102);
or U38414 (N_38414,N_30840,N_31437);
nor U38415 (N_38415,N_31998,N_31340);
and U38416 (N_38416,N_32689,N_30883);
nor U38417 (N_38417,N_30929,N_34342);
and U38418 (N_38418,N_32030,N_30913);
and U38419 (N_38419,N_32655,N_31629);
nand U38420 (N_38420,N_30670,N_32001);
or U38421 (N_38421,N_32994,N_33389);
xor U38422 (N_38422,N_30192,N_30828);
nand U38423 (N_38423,N_34004,N_34199);
xor U38424 (N_38424,N_30855,N_32426);
nand U38425 (N_38425,N_32346,N_33815);
or U38426 (N_38426,N_30286,N_34899);
nand U38427 (N_38427,N_33588,N_31994);
nor U38428 (N_38428,N_31418,N_30477);
xnor U38429 (N_38429,N_31644,N_31198);
and U38430 (N_38430,N_34029,N_34166);
nand U38431 (N_38431,N_34114,N_34574);
and U38432 (N_38432,N_30170,N_33028);
nand U38433 (N_38433,N_33142,N_33370);
nor U38434 (N_38434,N_31465,N_34821);
or U38435 (N_38435,N_31688,N_33355);
xnor U38436 (N_38436,N_30477,N_33779);
or U38437 (N_38437,N_30127,N_31322);
nand U38438 (N_38438,N_30409,N_31202);
nand U38439 (N_38439,N_31007,N_34107);
or U38440 (N_38440,N_33382,N_34519);
or U38441 (N_38441,N_33992,N_32052);
nand U38442 (N_38442,N_32375,N_32445);
xnor U38443 (N_38443,N_31076,N_33784);
and U38444 (N_38444,N_32240,N_31477);
and U38445 (N_38445,N_30881,N_34207);
xnor U38446 (N_38446,N_34672,N_32945);
xor U38447 (N_38447,N_30495,N_34756);
or U38448 (N_38448,N_32400,N_34626);
nor U38449 (N_38449,N_33525,N_33989);
and U38450 (N_38450,N_32032,N_34731);
nand U38451 (N_38451,N_34543,N_34362);
nor U38452 (N_38452,N_33124,N_34351);
nor U38453 (N_38453,N_30241,N_33715);
or U38454 (N_38454,N_32964,N_31044);
xor U38455 (N_38455,N_31695,N_33624);
nand U38456 (N_38456,N_32898,N_31799);
nand U38457 (N_38457,N_30269,N_31174);
xor U38458 (N_38458,N_32184,N_34875);
nor U38459 (N_38459,N_30139,N_33889);
and U38460 (N_38460,N_34678,N_33257);
xor U38461 (N_38461,N_31332,N_30147);
or U38462 (N_38462,N_30671,N_33125);
and U38463 (N_38463,N_31975,N_31908);
xor U38464 (N_38464,N_34624,N_32164);
xnor U38465 (N_38465,N_32333,N_32484);
nor U38466 (N_38466,N_32555,N_30288);
or U38467 (N_38467,N_31719,N_30349);
nor U38468 (N_38468,N_34883,N_32300);
nand U38469 (N_38469,N_30113,N_33804);
and U38470 (N_38470,N_32943,N_32717);
nand U38471 (N_38471,N_30836,N_31298);
nand U38472 (N_38472,N_34081,N_31430);
nand U38473 (N_38473,N_33182,N_30379);
or U38474 (N_38474,N_32236,N_33381);
xor U38475 (N_38475,N_34586,N_32925);
xnor U38476 (N_38476,N_32239,N_32506);
nor U38477 (N_38477,N_30998,N_34879);
nand U38478 (N_38478,N_30066,N_30840);
xor U38479 (N_38479,N_30888,N_34340);
xor U38480 (N_38480,N_34794,N_32972);
nor U38481 (N_38481,N_33555,N_32115);
nand U38482 (N_38482,N_34456,N_32571);
nand U38483 (N_38483,N_32601,N_30860);
and U38484 (N_38484,N_33241,N_32185);
nor U38485 (N_38485,N_30274,N_34260);
xor U38486 (N_38486,N_32302,N_31764);
or U38487 (N_38487,N_30052,N_32325);
or U38488 (N_38488,N_33847,N_34748);
nand U38489 (N_38489,N_32317,N_30583);
and U38490 (N_38490,N_34110,N_33843);
and U38491 (N_38491,N_31766,N_33765);
and U38492 (N_38492,N_34689,N_34398);
nor U38493 (N_38493,N_30661,N_30755);
nand U38494 (N_38494,N_32386,N_31881);
or U38495 (N_38495,N_34988,N_30242);
xor U38496 (N_38496,N_33083,N_32779);
or U38497 (N_38497,N_30059,N_33194);
or U38498 (N_38498,N_33396,N_34969);
xor U38499 (N_38499,N_34971,N_32135);
and U38500 (N_38500,N_34129,N_34090);
or U38501 (N_38501,N_33852,N_34723);
or U38502 (N_38502,N_34745,N_32510);
nand U38503 (N_38503,N_31721,N_33683);
or U38504 (N_38504,N_32082,N_30659);
and U38505 (N_38505,N_32062,N_31857);
and U38506 (N_38506,N_32399,N_33759);
nand U38507 (N_38507,N_30123,N_33261);
or U38508 (N_38508,N_34326,N_31238);
nor U38509 (N_38509,N_31925,N_32162);
nor U38510 (N_38510,N_34983,N_30266);
nor U38511 (N_38511,N_31340,N_31650);
nand U38512 (N_38512,N_33018,N_30797);
xnor U38513 (N_38513,N_31493,N_34711);
nor U38514 (N_38514,N_32704,N_32359);
nand U38515 (N_38515,N_34258,N_32714);
and U38516 (N_38516,N_30182,N_30712);
or U38517 (N_38517,N_31344,N_30596);
nand U38518 (N_38518,N_30288,N_33418);
nor U38519 (N_38519,N_31676,N_34352);
nand U38520 (N_38520,N_33260,N_32521);
nand U38521 (N_38521,N_33244,N_34222);
nand U38522 (N_38522,N_31249,N_31214);
nor U38523 (N_38523,N_30015,N_32923);
and U38524 (N_38524,N_34565,N_33292);
xor U38525 (N_38525,N_31652,N_30064);
nor U38526 (N_38526,N_30039,N_32267);
nand U38527 (N_38527,N_31944,N_32117);
nor U38528 (N_38528,N_33318,N_34009);
nor U38529 (N_38529,N_30917,N_34811);
nand U38530 (N_38530,N_32091,N_31074);
or U38531 (N_38531,N_32199,N_34397);
or U38532 (N_38532,N_31726,N_30872);
and U38533 (N_38533,N_34673,N_34248);
or U38534 (N_38534,N_32486,N_33936);
nor U38535 (N_38535,N_32871,N_30616);
nand U38536 (N_38536,N_32338,N_34581);
and U38537 (N_38537,N_33580,N_32602);
or U38538 (N_38538,N_30638,N_33207);
nor U38539 (N_38539,N_30606,N_31330);
xor U38540 (N_38540,N_33166,N_33178);
nor U38541 (N_38541,N_30372,N_31755);
or U38542 (N_38542,N_30907,N_32298);
nor U38543 (N_38543,N_30160,N_32249);
nor U38544 (N_38544,N_34548,N_30202);
nor U38545 (N_38545,N_33325,N_31378);
nor U38546 (N_38546,N_30239,N_34309);
and U38547 (N_38547,N_32970,N_31157);
nor U38548 (N_38548,N_33146,N_34091);
nor U38549 (N_38549,N_32411,N_31345);
xnor U38550 (N_38550,N_34012,N_33357);
nand U38551 (N_38551,N_33533,N_30108);
or U38552 (N_38552,N_31117,N_30688);
or U38553 (N_38553,N_33614,N_34605);
nor U38554 (N_38554,N_32062,N_32209);
nor U38555 (N_38555,N_34929,N_32749);
nor U38556 (N_38556,N_30622,N_31224);
xor U38557 (N_38557,N_30417,N_31588);
xor U38558 (N_38558,N_31575,N_31813);
nand U38559 (N_38559,N_33151,N_30714);
and U38560 (N_38560,N_31539,N_34498);
and U38561 (N_38561,N_32104,N_31188);
and U38562 (N_38562,N_31598,N_33188);
nor U38563 (N_38563,N_34931,N_34669);
and U38564 (N_38564,N_31019,N_34413);
xnor U38565 (N_38565,N_32903,N_31143);
xnor U38566 (N_38566,N_30392,N_30896);
or U38567 (N_38567,N_30119,N_32646);
nand U38568 (N_38568,N_34103,N_30901);
or U38569 (N_38569,N_33386,N_33441);
nand U38570 (N_38570,N_34900,N_34106);
or U38571 (N_38571,N_33907,N_33865);
nand U38572 (N_38572,N_33936,N_30088);
or U38573 (N_38573,N_33499,N_34565);
and U38574 (N_38574,N_31502,N_30324);
nor U38575 (N_38575,N_34131,N_34958);
or U38576 (N_38576,N_31432,N_30601);
or U38577 (N_38577,N_34516,N_34361);
xnor U38578 (N_38578,N_30755,N_30460);
nand U38579 (N_38579,N_33325,N_31136);
nor U38580 (N_38580,N_30381,N_33218);
or U38581 (N_38581,N_31946,N_33318);
xnor U38582 (N_38582,N_31121,N_32223);
nand U38583 (N_38583,N_34303,N_31183);
xor U38584 (N_38584,N_31864,N_31815);
nand U38585 (N_38585,N_33194,N_34525);
or U38586 (N_38586,N_33824,N_31398);
nor U38587 (N_38587,N_30598,N_31104);
or U38588 (N_38588,N_30113,N_33348);
nand U38589 (N_38589,N_33173,N_31819);
xor U38590 (N_38590,N_31883,N_32130);
nand U38591 (N_38591,N_32029,N_32590);
xnor U38592 (N_38592,N_33519,N_32608);
nand U38593 (N_38593,N_30808,N_32679);
or U38594 (N_38594,N_33040,N_30659);
nor U38595 (N_38595,N_31118,N_33457);
xnor U38596 (N_38596,N_30432,N_34044);
nor U38597 (N_38597,N_32933,N_32371);
xnor U38598 (N_38598,N_33048,N_33949);
xor U38599 (N_38599,N_34183,N_31418);
and U38600 (N_38600,N_33822,N_34915);
and U38601 (N_38601,N_32182,N_33845);
or U38602 (N_38602,N_33419,N_34002);
or U38603 (N_38603,N_31060,N_32611);
and U38604 (N_38604,N_32022,N_32624);
nand U38605 (N_38605,N_30850,N_30758);
nor U38606 (N_38606,N_32454,N_30299);
nand U38607 (N_38607,N_33668,N_32067);
nor U38608 (N_38608,N_30232,N_34892);
xnor U38609 (N_38609,N_33702,N_32317);
xnor U38610 (N_38610,N_32609,N_30499);
and U38611 (N_38611,N_32494,N_34571);
and U38612 (N_38612,N_33530,N_31116);
nor U38613 (N_38613,N_31991,N_32265);
or U38614 (N_38614,N_30860,N_31307);
nor U38615 (N_38615,N_30837,N_33806);
nor U38616 (N_38616,N_33036,N_33072);
xnor U38617 (N_38617,N_31093,N_31387);
nor U38618 (N_38618,N_32901,N_33132);
nor U38619 (N_38619,N_32609,N_30912);
or U38620 (N_38620,N_33918,N_34986);
xor U38621 (N_38621,N_32995,N_31720);
nand U38622 (N_38622,N_34835,N_34250);
nor U38623 (N_38623,N_31367,N_34069);
nand U38624 (N_38624,N_33039,N_33691);
nand U38625 (N_38625,N_33372,N_31679);
xor U38626 (N_38626,N_31967,N_32370);
or U38627 (N_38627,N_32443,N_32184);
nor U38628 (N_38628,N_32978,N_34884);
and U38629 (N_38629,N_34741,N_30541);
nor U38630 (N_38630,N_30810,N_33474);
or U38631 (N_38631,N_32306,N_33808);
and U38632 (N_38632,N_31941,N_30173);
and U38633 (N_38633,N_33169,N_33292);
nor U38634 (N_38634,N_34814,N_33091);
or U38635 (N_38635,N_31887,N_30086);
nor U38636 (N_38636,N_32124,N_32403);
xor U38637 (N_38637,N_30805,N_34818);
and U38638 (N_38638,N_32847,N_34919);
xor U38639 (N_38639,N_30336,N_33785);
nor U38640 (N_38640,N_33398,N_34348);
nor U38641 (N_38641,N_30964,N_30416);
nor U38642 (N_38642,N_31461,N_33589);
nor U38643 (N_38643,N_32309,N_31789);
nor U38644 (N_38644,N_31062,N_30399);
nand U38645 (N_38645,N_33140,N_30035);
nor U38646 (N_38646,N_30665,N_33598);
and U38647 (N_38647,N_34823,N_34870);
nor U38648 (N_38648,N_34512,N_30453);
or U38649 (N_38649,N_33504,N_31242);
xor U38650 (N_38650,N_30368,N_33245);
xor U38651 (N_38651,N_34867,N_32574);
and U38652 (N_38652,N_31039,N_33440);
nor U38653 (N_38653,N_34224,N_30880);
nor U38654 (N_38654,N_34361,N_30430);
nor U38655 (N_38655,N_30470,N_31372);
or U38656 (N_38656,N_31236,N_32094);
nor U38657 (N_38657,N_32640,N_32751);
or U38658 (N_38658,N_30202,N_30968);
or U38659 (N_38659,N_33794,N_30683);
or U38660 (N_38660,N_32366,N_33696);
xnor U38661 (N_38661,N_31971,N_31560);
nor U38662 (N_38662,N_30476,N_34680);
nand U38663 (N_38663,N_33019,N_34963);
nand U38664 (N_38664,N_31523,N_34758);
and U38665 (N_38665,N_32080,N_30876);
or U38666 (N_38666,N_33656,N_32662);
nand U38667 (N_38667,N_30799,N_30168);
nor U38668 (N_38668,N_33107,N_33975);
nand U38669 (N_38669,N_34553,N_32343);
or U38670 (N_38670,N_34726,N_32342);
xnor U38671 (N_38671,N_34523,N_33344);
or U38672 (N_38672,N_34862,N_33649);
and U38673 (N_38673,N_32756,N_30624);
or U38674 (N_38674,N_31291,N_33781);
nand U38675 (N_38675,N_30943,N_31912);
nor U38676 (N_38676,N_30586,N_30116);
nor U38677 (N_38677,N_34922,N_30147);
or U38678 (N_38678,N_31128,N_34125);
nand U38679 (N_38679,N_31030,N_34025);
xnor U38680 (N_38680,N_32234,N_32100);
or U38681 (N_38681,N_32176,N_30434);
nor U38682 (N_38682,N_34486,N_31303);
xor U38683 (N_38683,N_30672,N_30479);
xnor U38684 (N_38684,N_31852,N_32708);
nand U38685 (N_38685,N_33449,N_32326);
xor U38686 (N_38686,N_31852,N_34205);
and U38687 (N_38687,N_34067,N_30835);
nand U38688 (N_38688,N_32027,N_31794);
and U38689 (N_38689,N_32592,N_34251);
or U38690 (N_38690,N_33865,N_34502);
nor U38691 (N_38691,N_34310,N_34153);
nor U38692 (N_38692,N_33784,N_31459);
nor U38693 (N_38693,N_34475,N_30366);
xnor U38694 (N_38694,N_33114,N_33893);
or U38695 (N_38695,N_34526,N_30427);
nand U38696 (N_38696,N_32611,N_31226);
nand U38697 (N_38697,N_31573,N_30956);
nand U38698 (N_38698,N_34251,N_30450);
and U38699 (N_38699,N_33023,N_32271);
xor U38700 (N_38700,N_34033,N_30737);
xnor U38701 (N_38701,N_33965,N_31614);
xor U38702 (N_38702,N_31732,N_30851);
or U38703 (N_38703,N_30968,N_32527);
and U38704 (N_38704,N_33516,N_32674);
or U38705 (N_38705,N_32731,N_31029);
and U38706 (N_38706,N_30010,N_33209);
xor U38707 (N_38707,N_34311,N_34890);
nand U38708 (N_38708,N_34394,N_30546);
nor U38709 (N_38709,N_32072,N_33130);
nand U38710 (N_38710,N_34402,N_34185);
nor U38711 (N_38711,N_34030,N_32879);
nor U38712 (N_38712,N_30927,N_30529);
xor U38713 (N_38713,N_34244,N_30431);
and U38714 (N_38714,N_32925,N_34271);
or U38715 (N_38715,N_32564,N_33667);
and U38716 (N_38716,N_30172,N_30647);
or U38717 (N_38717,N_32919,N_32204);
xor U38718 (N_38718,N_32263,N_34909);
xnor U38719 (N_38719,N_33743,N_30030);
nor U38720 (N_38720,N_30057,N_31230);
nand U38721 (N_38721,N_34451,N_30900);
xnor U38722 (N_38722,N_32887,N_31582);
and U38723 (N_38723,N_34579,N_31639);
nor U38724 (N_38724,N_31850,N_34995);
nor U38725 (N_38725,N_33945,N_34391);
nand U38726 (N_38726,N_30766,N_34183);
xnor U38727 (N_38727,N_33896,N_32757);
xor U38728 (N_38728,N_30132,N_34303);
xnor U38729 (N_38729,N_32783,N_32505);
nand U38730 (N_38730,N_34900,N_30633);
nand U38731 (N_38731,N_32151,N_34939);
xnor U38732 (N_38732,N_34877,N_30389);
nand U38733 (N_38733,N_32653,N_31787);
nand U38734 (N_38734,N_31769,N_32846);
nand U38735 (N_38735,N_34801,N_31579);
or U38736 (N_38736,N_32918,N_30619);
and U38737 (N_38737,N_30955,N_33757);
or U38738 (N_38738,N_33227,N_30664);
and U38739 (N_38739,N_33289,N_32024);
xnor U38740 (N_38740,N_34419,N_30805);
nand U38741 (N_38741,N_33612,N_30958);
nand U38742 (N_38742,N_34406,N_31178);
or U38743 (N_38743,N_31606,N_32268);
and U38744 (N_38744,N_32191,N_31656);
and U38745 (N_38745,N_33202,N_33838);
nor U38746 (N_38746,N_32226,N_33770);
and U38747 (N_38747,N_31557,N_33865);
nand U38748 (N_38748,N_30016,N_30616);
nand U38749 (N_38749,N_33767,N_30049);
xnor U38750 (N_38750,N_32991,N_32343);
or U38751 (N_38751,N_30015,N_31500);
nand U38752 (N_38752,N_32328,N_31845);
and U38753 (N_38753,N_33177,N_31891);
nand U38754 (N_38754,N_33709,N_33562);
and U38755 (N_38755,N_32998,N_31544);
or U38756 (N_38756,N_32305,N_32573);
and U38757 (N_38757,N_31537,N_34394);
xnor U38758 (N_38758,N_31422,N_31940);
or U38759 (N_38759,N_33053,N_30730);
and U38760 (N_38760,N_34930,N_31491);
and U38761 (N_38761,N_30709,N_30594);
xnor U38762 (N_38762,N_34558,N_31578);
or U38763 (N_38763,N_33385,N_31046);
or U38764 (N_38764,N_32298,N_30964);
or U38765 (N_38765,N_34242,N_33551);
nor U38766 (N_38766,N_30104,N_34998);
and U38767 (N_38767,N_33457,N_30429);
nor U38768 (N_38768,N_31836,N_34007);
or U38769 (N_38769,N_34672,N_32909);
nor U38770 (N_38770,N_31709,N_34156);
and U38771 (N_38771,N_30215,N_32843);
or U38772 (N_38772,N_33677,N_32759);
nand U38773 (N_38773,N_30343,N_34208);
xor U38774 (N_38774,N_31940,N_33409);
xor U38775 (N_38775,N_33365,N_34131);
nand U38776 (N_38776,N_30095,N_33806);
nand U38777 (N_38777,N_32713,N_34649);
nand U38778 (N_38778,N_34112,N_31556);
xor U38779 (N_38779,N_32992,N_33917);
nor U38780 (N_38780,N_34660,N_34461);
or U38781 (N_38781,N_30177,N_30316);
nor U38782 (N_38782,N_34343,N_34349);
nand U38783 (N_38783,N_33930,N_34255);
or U38784 (N_38784,N_33456,N_34384);
or U38785 (N_38785,N_33696,N_32715);
nor U38786 (N_38786,N_30337,N_30013);
nor U38787 (N_38787,N_31195,N_32936);
nor U38788 (N_38788,N_30542,N_31044);
nor U38789 (N_38789,N_33431,N_33360);
nand U38790 (N_38790,N_31774,N_30452);
xor U38791 (N_38791,N_34845,N_31303);
xor U38792 (N_38792,N_33115,N_33275);
or U38793 (N_38793,N_30652,N_33061);
xnor U38794 (N_38794,N_33909,N_30937);
or U38795 (N_38795,N_34720,N_32663);
and U38796 (N_38796,N_30280,N_34231);
and U38797 (N_38797,N_31139,N_30825);
or U38798 (N_38798,N_30300,N_33260);
nand U38799 (N_38799,N_34519,N_30977);
xnor U38800 (N_38800,N_30373,N_32979);
nor U38801 (N_38801,N_33628,N_34382);
nand U38802 (N_38802,N_34673,N_31263);
or U38803 (N_38803,N_34545,N_30820);
xnor U38804 (N_38804,N_34055,N_30442);
or U38805 (N_38805,N_34316,N_34591);
and U38806 (N_38806,N_30004,N_30469);
and U38807 (N_38807,N_34692,N_34690);
and U38808 (N_38808,N_31017,N_34982);
and U38809 (N_38809,N_34015,N_31650);
nand U38810 (N_38810,N_30455,N_32152);
and U38811 (N_38811,N_33038,N_31902);
nor U38812 (N_38812,N_34380,N_34029);
nand U38813 (N_38813,N_33640,N_30880);
and U38814 (N_38814,N_33089,N_32946);
nand U38815 (N_38815,N_32552,N_30781);
and U38816 (N_38816,N_31755,N_31847);
xor U38817 (N_38817,N_32403,N_33918);
nor U38818 (N_38818,N_31813,N_30656);
xor U38819 (N_38819,N_33240,N_30559);
nand U38820 (N_38820,N_31437,N_34384);
nor U38821 (N_38821,N_31248,N_32027);
nor U38822 (N_38822,N_34017,N_34376);
nor U38823 (N_38823,N_34044,N_31956);
xor U38824 (N_38824,N_34091,N_34923);
and U38825 (N_38825,N_32260,N_33545);
xor U38826 (N_38826,N_34399,N_30076);
nand U38827 (N_38827,N_30508,N_32295);
or U38828 (N_38828,N_31899,N_33308);
xor U38829 (N_38829,N_32365,N_33577);
nor U38830 (N_38830,N_32407,N_34137);
or U38831 (N_38831,N_31802,N_33713);
nand U38832 (N_38832,N_33121,N_33176);
or U38833 (N_38833,N_31527,N_33523);
xnor U38834 (N_38834,N_30919,N_30509);
nor U38835 (N_38835,N_34857,N_33683);
xor U38836 (N_38836,N_34914,N_30334);
nand U38837 (N_38837,N_34092,N_32174);
xor U38838 (N_38838,N_33388,N_33779);
nand U38839 (N_38839,N_30282,N_32637);
or U38840 (N_38840,N_31814,N_34978);
xor U38841 (N_38841,N_33345,N_34953);
or U38842 (N_38842,N_30431,N_30287);
nor U38843 (N_38843,N_31884,N_30455);
nand U38844 (N_38844,N_32568,N_31949);
or U38845 (N_38845,N_34370,N_30082);
xor U38846 (N_38846,N_33735,N_33812);
nor U38847 (N_38847,N_34066,N_31484);
nor U38848 (N_38848,N_31242,N_31365);
nand U38849 (N_38849,N_30899,N_33854);
and U38850 (N_38850,N_30194,N_30875);
and U38851 (N_38851,N_32903,N_33848);
xnor U38852 (N_38852,N_34626,N_33177);
xor U38853 (N_38853,N_34439,N_33062);
xnor U38854 (N_38854,N_34200,N_32712);
xor U38855 (N_38855,N_34838,N_32108);
nand U38856 (N_38856,N_34924,N_30329);
or U38857 (N_38857,N_33314,N_34090);
nand U38858 (N_38858,N_33446,N_30838);
xor U38859 (N_38859,N_30043,N_33357);
xnor U38860 (N_38860,N_33752,N_31983);
xor U38861 (N_38861,N_33792,N_34370);
xor U38862 (N_38862,N_33232,N_31007);
nor U38863 (N_38863,N_33533,N_34670);
and U38864 (N_38864,N_32724,N_32025);
xor U38865 (N_38865,N_32916,N_33707);
xor U38866 (N_38866,N_32563,N_30478);
xnor U38867 (N_38867,N_31894,N_31743);
xnor U38868 (N_38868,N_34629,N_33416);
xor U38869 (N_38869,N_34257,N_31249);
xor U38870 (N_38870,N_31614,N_32613);
and U38871 (N_38871,N_34518,N_32674);
nor U38872 (N_38872,N_34628,N_30179);
or U38873 (N_38873,N_30631,N_30229);
and U38874 (N_38874,N_30559,N_30533);
nor U38875 (N_38875,N_30301,N_33876);
or U38876 (N_38876,N_31078,N_32799);
xor U38877 (N_38877,N_30069,N_33481);
nor U38878 (N_38878,N_34844,N_32147);
and U38879 (N_38879,N_34494,N_31905);
or U38880 (N_38880,N_30374,N_31748);
xor U38881 (N_38881,N_31994,N_31641);
nand U38882 (N_38882,N_30584,N_30021);
xnor U38883 (N_38883,N_32535,N_31135);
xor U38884 (N_38884,N_33324,N_34565);
and U38885 (N_38885,N_34790,N_30698);
nand U38886 (N_38886,N_31298,N_32470);
xnor U38887 (N_38887,N_33124,N_34883);
nor U38888 (N_38888,N_34347,N_33906);
and U38889 (N_38889,N_34472,N_30064);
nand U38890 (N_38890,N_32530,N_33173);
or U38891 (N_38891,N_32828,N_32462);
or U38892 (N_38892,N_32668,N_34125);
nor U38893 (N_38893,N_33653,N_31873);
or U38894 (N_38894,N_34607,N_33928);
and U38895 (N_38895,N_32198,N_30818);
and U38896 (N_38896,N_32166,N_31926);
or U38897 (N_38897,N_34062,N_34006);
or U38898 (N_38898,N_30047,N_33185);
and U38899 (N_38899,N_34087,N_34490);
and U38900 (N_38900,N_30705,N_31042);
and U38901 (N_38901,N_31111,N_30197);
nor U38902 (N_38902,N_32377,N_32881);
or U38903 (N_38903,N_33347,N_32875);
nor U38904 (N_38904,N_33850,N_31189);
and U38905 (N_38905,N_32370,N_31433);
nor U38906 (N_38906,N_34010,N_31571);
xor U38907 (N_38907,N_32799,N_31456);
xnor U38908 (N_38908,N_32447,N_32295);
nor U38909 (N_38909,N_33611,N_33794);
nand U38910 (N_38910,N_30576,N_33031);
or U38911 (N_38911,N_32056,N_30557);
or U38912 (N_38912,N_32112,N_33140);
nor U38913 (N_38913,N_33954,N_34970);
nor U38914 (N_38914,N_31170,N_34768);
nor U38915 (N_38915,N_31062,N_30078);
and U38916 (N_38916,N_34668,N_32777);
or U38917 (N_38917,N_30422,N_32964);
nand U38918 (N_38918,N_33520,N_31641);
nand U38919 (N_38919,N_34701,N_31989);
nand U38920 (N_38920,N_34751,N_34454);
xor U38921 (N_38921,N_32156,N_30433);
nand U38922 (N_38922,N_34269,N_34520);
nand U38923 (N_38923,N_30685,N_31583);
or U38924 (N_38924,N_33241,N_33011);
and U38925 (N_38925,N_31115,N_34801);
xor U38926 (N_38926,N_30771,N_32590);
xor U38927 (N_38927,N_32057,N_30209);
nand U38928 (N_38928,N_34241,N_31163);
and U38929 (N_38929,N_32907,N_34506);
nand U38930 (N_38930,N_30712,N_33614);
nand U38931 (N_38931,N_33914,N_34824);
xnor U38932 (N_38932,N_30106,N_32510);
xor U38933 (N_38933,N_32012,N_34273);
nor U38934 (N_38934,N_31160,N_30111);
xor U38935 (N_38935,N_30027,N_33388);
xor U38936 (N_38936,N_31489,N_34922);
and U38937 (N_38937,N_31050,N_30039);
nand U38938 (N_38938,N_33747,N_30122);
nand U38939 (N_38939,N_30261,N_34026);
xor U38940 (N_38940,N_32240,N_30439);
and U38941 (N_38941,N_33109,N_34230);
nand U38942 (N_38942,N_32527,N_34126);
xor U38943 (N_38943,N_33640,N_33634);
and U38944 (N_38944,N_34233,N_31232);
nor U38945 (N_38945,N_32293,N_34534);
nor U38946 (N_38946,N_34325,N_32565);
or U38947 (N_38947,N_32079,N_33923);
xnor U38948 (N_38948,N_31342,N_31644);
xor U38949 (N_38949,N_31288,N_31652);
and U38950 (N_38950,N_34438,N_34012);
nor U38951 (N_38951,N_32193,N_33806);
or U38952 (N_38952,N_32527,N_34117);
nor U38953 (N_38953,N_31183,N_31717);
or U38954 (N_38954,N_32194,N_33731);
or U38955 (N_38955,N_33694,N_34516);
xnor U38956 (N_38956,N_33598,N_33314);
and U38957 (N_38957,N_30242,N_31456);
xor U38958 (N_38958,N_33660,N_32517);
xnor U38959 (N_38959,N_32859,N_30950);
nand U38960 (N_38960,N_30426,N_33410);
xor U38961 (N_38961,N_30478,N_33011);
or U38962 (N_38962,N_30035,N_33175);
and U38963 (N_38963,N_30736,N_30632);
or U38964 (N_38964,N_33895,N_31834);
xnor U38965 (N_38965,N_33175,N_31915);
or U38966 (N_38966,N_32747,N_33028);
or U38967 (N_38967,N_31405,N_30154);
or U38968 (N_38968,N_33183,N_31867);
nand U38969 (N_38969,N_32099,N_31720);
nand U38970 (N_38970,N_33363,N_33864);
and U38971 (N_38971,N_31387,N_34498);
nand U38972 (N_38972,N_33024,N_31709);
xnor U38973 (N_38973,N_32824,N_33909);
nand U38974 (N_38974,N_31181,N_31517);
nor U38975 (N_38975,N_31067,N_31313);
and U38976 (N_38976,N_32714,N_33018);
nand U38977 (N_38977,N_32188,N_30870);
xnor U38978 (N_38978,N_33073,N_30657);
xor U38979 (N_38979,N_32549,N_31020);
nor U38980 (N_38980,N_30918,N_30347);
nand U38981 (N_38981,N_33484,N_33724);
nor U38982 (N_38982,N_34332,N_30334);
nor U38983 (N_38983,N_31940,N_34105);
nand U38984 (N_38984,N_34237,N_31806);
nand U38985 (N_38985,N_31258,N_32539);
and U38986 (N_38986,N_30016,N_32186);
and U38987 (N_38987,N_32897,N_31635);
or U38988 (N_38988,N_34717,N_33473);
or U38989 (N_38989,N_31048,N_32529);
or U38990 (N_38990,N_33531,N_30518);
xnor U38991 (N_38991,N_33916,N_31284);
or U38992 (N_38992,N_33337,N_31434);
or U38993 (N_38993,N_31236,N_33465);
nor U38994 (N_38994,N_32083,N_32015);
nand U38995 (N_38995,N_33757,N_31235);
or U38996 (N_38996,N_30671,N_32411);
or U38997 (N_38997,N_30731,N_32769);
and U38998 (N_38998,N_30277,N_32763);
and U38999 (N_38999,N_31134,N_31067);
nand U39000 (N_39000,N_31395,N_33899);
nand U39001 (N_39001,N_30263,N_32319);
xnor U39002 (N_39002,N_33641,N_30484);
and U39003 (N_39003,N_32816,N_34790);
xnor U39004 (N_39004,N_33471,N_31870);
nor U39005 (N_39005,N_30264,N_33137);
nor U39006 (N_39006,N_32427,N_31871);
xnor U39007 (N_39007,N_31125,N_32436);
nor U39008 (N_39008,N_32821,N_30361);
and U39009 (N_39009,N_34664,N_33341);
and U39010 (N_39010,N_30139,N_32230);
nor U39011 (N_39011,N_33555,N_32660);
xor U39012 (N_39012,N_32597,N_31611);
nor U39013 (N_39013,N_32334,N_33703);
nand U39014 (N_39014,N_31089,N_33791);
or U39015 (N_39015,N_31183,N_30124);
xor U39016 (N_39016,N_31161,N_31093);
xor U39017 (N_39017,N_32391,N_30223);
xnor U39018 (N_39018,N_31119,N_34470);
nor U39019 (N_39019,N_34352,N_30023);
nand U39020 (N_39020,N_31719,N_31656);
nor U39021 (N_39021,N_30032,N_34039);
nand U39022 (N_39022,N_34942,N_31348);
nor U39023 (N_39023,N_32418,N_33432);
nand U39024 (N_39024,N_31350,N_33355);
nand U39025 (N_39025,N_34983,N_33275);
and U39026 (N_39026,N_31197,N_34232);
nand U39027 (N_39027,N_34790,N_30116);
or U39028 (N_39028,N_32025,N_31621);
or U39029 (N_39029,N_33810,N_33320);
nand U39030 (N_39030,N_33689,N_34139);
nor U39031 (N_39031,N_30698,N_32738);
or U39032 (N_39032,N_31467,N_33725);
nor U39033 (N_39033,N_33574,N_33887);
nand U39034 (N_39034,N_34273,N_33697);
nor U39035 (N_39035,N_31715,N_32192);
or U39036 (N_39036,N_33572,N_30062);
nor U39037 (N_39037,N_34953,N_31617);
nand U39038 (N_39038,N_33021,N_30815);
and U39039 (N_39039,N_34084,N_30958);
xor U39040 (N_39040,N_31168,N_32162);
nor U39041 (N_39041,N_31919,N_31566);
xnor U39042 (N_39042,N_34408,N_34992);
or U39043 (N_39043,N_32339,N_31631);
nand U39044 (N_39044,N_31304,N_33412);
or U39045 (N_39045,N_31789,N_34506);
nand U39046 (N_39046,N_34720,N_32369);
xor U39047 (N_39047,N_34863,N_34307);
nand U39048 (N_39048,N_30133,N_31863);
nand U39049 (N_39049,N_30570,N_33275);
nand U39050 (N_39050,N_34869,N_32308);
or U39051 (N_39051,N_30399,N_31500);
xor U39052 (N_39052,N_34364,N_33513);
nor U39053 (N_39053,N_31294,N_33122);
nor U39054 (N_39054,N_32161,N_31757);
xnor U39055 (N_39055,N_33360,N_32614);
xnor U39056 (N_39056,N_31267,N_32366);
nor U39057 (N_39057,N_33632,N_32596);
xor U39058 (N_39058,N_34763,N_31350);
nand U39059 (N_39059,N_31721,N_34623);
or U39060 (N_39060,N_31187,N_31203);
nand U39061 (N_39061,N_32110,N_31671);
and U39062 (N_39062,N_32682,N_30784);
nor U39063 (N_39063,N_34376,N_31065);
nand U39064 (N_39064,N_34618,N_30581);
nand U39065 (N_39065,N_33034,N_30205);
nand U39066 (N_39066,N_34075,N_33843);
or U39067 (N_39067,N_30155,N_31797);
and U39068 (N_39068,N_33459,N_33583);
xnor U39069 (N_39069,N_34393,N_30945);
and U39070 (N_39070,N_32077,N_31096);
and U39071 (N_39071,N_30704,N_32326);
nor U39072 (N_39072,N_34121,N_33994);
or U39073 (N_39073,N_31321,N_31429);
nand U39074 (N_39074,N_31081,N_30077);
nand U39075 (N_39075,N_32396,N_31286);
nor U39076 (N_39076,N_30957,N_31414);
nor U39077 (N_39077,N_32695,N_31669);
nor U39078 (N_39078,N_33008,N_32091);
nand U39079 (N_39079,N_30075,N_33447);
xnor U39080 (N_39080,N_34980,N_34259);
xor U39081 (N_39081,N_30141,N_33062);
and U39082 (N_39082,N_31608,N_31866);
nand U39083 (N_39083,N_30488,N_30862);
xor U39084 (N_39084,N_32962,N_32086);
xnor U39085 (N_39085,N_34522,N_30731);
or U39086 (N_39086,N_31996,N_30937);
and U39087 (N_39087,N_33477,N_34885);
nor U39088 (N_39088,N_31089,N_33085);
or U39089 (N_39089,N_34527,N_30152);
xor U39090 (N_39090,N_31799,N_32735);
and U39091 (N_39091,N_32441,N_34790);
nor U39092 (N_39092,N_34152,N_33373);
or U39093 (N_39093,N_32628,N_32469);
xnor U39094 (N_39094,N_34938,N_34160);
nor U39095 (N_39095,N_30947,N_34643);
nand U39096 (N_39096,N_30809,N_33647);
nor U39097 (N_39097,N_34890,N_34940);
nor U39098 (N_39098,N_31478,N_32902);
and U39099 (N_39099,N_33232,N_30443);
and U39100 (N_39100,N_34319,N_33283);
nor U39101 (N_39101,N_34770,N_30373);
xnor U39102 (N_39102,N_34907,N_31905);
nand U39103 (N_39103,N_34848,N_31137);
nor U39104 (N_39104,N_32360,N_30157);
or U39105 (N_39105,N_30507,N_34878);
nand U39106 (N_39106,N_34661,N_34945);
xnor U39107 (N_39107,N_31098,N_34978);
nand U39108 (N_39108,N_31363,N_33764);
nor U39109 (N_39109,N_32857,N_34344);
nand U39110 (N_39110,N_33650,N_34807);
or U39111 (N_39111,N_31398,N_32472);
xor U39112 (N_39112,N_30205,N_32985);
nor U39113 (N_39113,N_31773,N_31384);
and U39114 (N_39114,N_31427,N_31769);
or U39115 (N_39115,N_32199,N_30785);
xor U39116 (N_39116,N_30577,N_33049);
xnor U39117 (N_39117,N_34678,N_34959);
nand U39118 (N_39118,N_31829,N_30656);
or U39119 (N_39119,N_32996,N_32082);
and U39120 (N_39120,N_32557,N_32609);
nand U39121 (N_39121,N_34096,N_33660);
nor U39122 (N_39122,N_34118,N_30681);
nand U39123 (N_39123,N_33723,N_32447);
nand U39124 (N_39124,N_30056,N_33200);
xnor U39125 (N_39125,N_32940,N_31789);
and U39126 (N_39126,N_34809,N_32755);
nor U39127 (N_39127,N_30234,N_31311);
xor U39128 (N_39128,N_33671,N_34355);
nand U39129 (N_39129,N_33527,N_31084);
xnor U39130 (N_39130,N_32088,N_30469);
xnor U39131 (N_39131,N_30093,N_30920);
or U39132 (N_39132,N_31457,N_30650);
nand U39133 (N_39133,N_33530,N_30793);
nand U39134 (N_39134,N_30985,N_30010);
and U39135 (N_39135,N_34860,N_31148);
nand U39136 (N_39136,N_34327,N_34959);
nand U39137 (N_39137,N_34909,N_31793);
xnor U39138 (N_39138,N_34504,N_31991);
nor U39139 (N_39139,N_32976,N_30177);
nand U39140 (N_39140,N_30783,N_31379);
nor U39141 (N_39141,N_34065,N_33482);
xnor U39142 (N_39142,N_30802,N_32889);
and U39143 (N_39143,N_30269,N_32696);
or U39144 (N_39144,N_32600,N_31360);
nand U39145 (N_39145,N_33447,N_33935);
nor U39146 (N_39146,N_31489,N_33012);
xnor U39147 (N_39147,N_32368,N_31491);
xor U39148 (N_39148,N_34505,N_32963);
and U39149 (N_39149,N_30136,N_31150);
or U39150 (N_39150,N_30050,N_33881);
or U39151 (N_39151,N_34057,N_33916);
nor U39152 (N_39152,N_34320,N_33104);
nand U39153 (N_39153,N_33215,N_34308);
nor U39154 (N_39154,N_34655,N_33381);
nor U39155 (N_39155,N_31694,N_31184);
nand U39156 (N_39156,N_32321,N_33560);
nor U39157 (N_39157,N_32907,N_31371);
nor U39158 (N_39158,N_32544,N_31464);
or U39159 (N_39159,N_30871,N_30728);
or U39160 (N_39160,N_32407,N_32674);
or U39161 (N_39161,N_30758,N_32097);
or U39162 (N_39162,N_33063,N_31464);
xnor U39163 (N_39163,N_33596,N_32614);
xnor U39164 (N_39164,N_32418,N_32334);
nor U39165 (N_39165,N_34332,N_32763);
xnor U39166 (N_39166,N_30163,N_33975);
and U39167 (N_39167,N_32855,N_30487);
and U39168 (N_39168,N_34220,N_30861);
xor U39169 (N_39169,N_31204,N_32471);
and U39170 (N_39170,N_34972,N_31048);
xor U39171 (N_39171,N_34430,N_32576);
xor U39172 (N_39172,N_30804,N_30530);
and U39173 (N_39173,N_32507,N_31498);
and U39174 (N_39174,N_30301,N_30081);
and U39175 (N_39175,N_30604,N_31963);
nand U39176 (N_39176,N_34008,N_31633);
nand U39177 (N_39177,N_30374,N_33835);
nand U39178 (N_39178,N_33948,N_34597);
nand U39179 (N_39179,N_30269,N_32167);
or U39180 (N_39180,N_33020,N_30135);
and U39181 (N_39181,N_30713,N_31545);
nand U39182 (N_39182,N_31669,N_33879);
nor U39183 (N_39183,N_34820,N_34320);
nand U39184 (N_39184,N_33374,N_33014);
and U39185 (N_39185,N_33479,N_30689);
and U39186 (N_39186,N_31944,N_34857);
nand U39187 (N_39187,N_30900,N_32284);
xor U39188 (N_39188,N_31526,N_33131);
xnor U39189 (N_39189,N_34469,N_31770);
and U39190 (N_39190,N_32465,N_34943);
and U39191 (N_39191,N_32777,N_33660);
nor U39192 (N_39192,N_30153,N_34545);
nor U39193 (N_39193,N_32314,N_31904);
xor U39194 (N_39194,N_34631,N_34633);
and U39195 (N_39195,N_30046,N_30467);
or U39196 (N_39196,N_32633,N_32732);
and U39197 (N_39197,N_34063,N_31459);
nand U39198 (N_39198,N_33771,N_33927);
xor U39199 (N_39199,N_34059,N_31026);
and U39200 (N_39200,N_33816,N_33999);
nand U39201 (N_39201,N_31404,N_31587);
and U39202 (N_39202,N_34496,N_30838);
and U39203 (N_39203,N_34764,N_30402);
nor U39204 (N_39204,N_32517,N_30976);
and U39205 (N_39205,N_32818,N_32007);
and U39206 (N_39206,N_31044,N_30871);
and U39207 (N_39207,N_33105,N_33132);
xnor U39208 (N_39208,N_31038,N_33895);
xnor U39209 (N_39209,N_34125,N_31949);
nand U39210 (N_39210,N_32788,N_34120);
nand U39211 (N_39211,N_31258,N_34454);
or U39212 (N_39212,N_30258,N_34189);
or U39213 (N_39213,N_30818,N_31422);
nand U39214 (N_39214,N_30691,N_33003);
nor U39215 (N_39215,N_33899,N_34086);
or U39216 (N_39216,N_32067,N_30424);
and U39217 (N_39217,N_33347,N_33171);
xor U39218 (N_39218,N_33862,N_33327);
nor U39219 (N_39219,N_30820,N_34992);
xnor U39220 (N_39220,N_33806,N_30960);
xor U39221 (N_39221,N_34748,N_31388);
nand U39222 (N_39222,N_34295,N_31120);
and U39223 (N_39223,N_31684,N_30587);
and U39224 (N_39224,N_31441,N_30751);
and U39225 (N_39225,N_33183,N_34115);
or U39226 (N_39226,N_30012,N_32812);
nor U39227 (N_39227,N_32790,N_34929);
nor U39228 (N_39228,N_31023,N_34858);
nand U39229 (N_39229,N_34274,N_30891);
and U39230 (N_39230,N_34869,N_31759);
xor U39231 (N_39231,N_33873,N_32542);
nand U39232 (N_39232,N_34931,N_33688);
nand U39233 (N_39233,N_33145,N_34998);
nor U39234 (N_39234,N_34209,N_31854);
xor U39235 (N_39235,N_31025,N_34190);
nor U39236 (N_39236,N_30556,N_34281);
nand U39237 (N_39237,N_34507,N_34607);
xnor U39238 (N_39238,N_33681,N_32510);
and U39239 (N_39239,N_34852,N_30253);
nand U39240 (N_39240,N_33946,N_34951);
xor U39241 (N_39241,N_34934,N_31984);
xor U39242 (N_39242,N_32598,N_30085);
and U39243 (N_39243,N_31318,N_32232);
nand U39244 (N_39244,N_32412,N_30913);
and U39245 (N_39245,N_33242,N_31730);
or U39246 (N_39246,N_30661,N_33936);
nor U39247 (N_39247,N_30022,N_30378);
and U39248 (N_39248,N_34494,N_34029);
nand U39249 (N_39249,N_33831,N_33846);
nand U39250 (N_39250,N_31894,N_33101);
nor U39251 (N_39251,N_30400,N_30411);
nand U39252 (N_39252,N_32582,N_32583);
and U39253 (N_39253,N_34245,N_34689);
and U39254 (N_39254,N_32151,N_30104);
and U39255 (N_39255,N_31983,N_34864);
and U39256 (N_39256,N_32839,N_31720);
nand U39257 (N_39257,N_30428,N_31496);
and U39258 (N_39258,N_30737,N_32128);
nand U39259 (N_39259,N_30250,N_34697);
nand U39260 (N_39260,N_30225,N_33377);
xor U39261 (N_39261,N_33971,N_33239);
or U39262 (N_39262,N_30377,N_30484);
or U39263 (N_39263,N_31669,N_32279);
nand U39264 (N_39264,N_34569,N_32577);
and U39265 (N_39265,N_31898,N_30316);
or U39266 (N_39266,N_32575,N_34551);
or U39267 (N_39267,N_32299,N_33716);
nand U39268 (N_39268,N_32273,N_30388);
nand U39269 (N_39269,N_30365,N_30221);
or U39270 (N_39270,N_30696,N_30934);
or U39271 (N_39271,N_34185,N_30135);
or U39272 (N_39272,N_30431,N_33123);
nor U39273 (N_39273,N_33108,N_34013);
or U39274 (N_39274,N_32323,N_30064);
xnor U39275 (N_39275,N_33826,N_31046);
nand U39276 (N_39276,N_30175,N_33612);
or U39277 (N_39277,N_33514,N_33348);
or U39278 (N_39278,N_32177,N_32313);
xor U39279 (N_39279,N_32283,N_31622);
nor U39280 (N_39280,N_31863,N_33317);
or U39281 (N_39281,N_34699,N_34416);
and U39282 (N_39282,N_30020,N_32097);
nor U39283 (N_39283,N_34977,N_33838);
xnor U39284 (N_39284,N_34999,N_33609);
or U39285 (N_39285,N_32794,N_32447);
xnor U39286 (N_39286,N_31126,N_32914);
or U39287 (N_39287,N_31711,N_32354);
and U39288 (N_39288,N_30890,N_31708);
or U39289 (N_39289,N_32422,N_34837);
and U39290 (N_39290,N_34116,N_30724);
nor U39291 (N_39291,N_32493,N_31825);
xor U39292 (N_39292,N_31925,N_32451);
and U39293 (N_39293,N_34819,N_34738);
and U39294 (N_39294,N_31536,N_34026);
xnor U39295 (N_39295,N_32108,N_32833);
and U39296 (N_39296,N_31525,N_33646);
and U39297 (N_39297,N_30466,N_33233);
or U39298 (N_39298,N_32094,N_32549);
xor U39299 (N_39299,N_34380,N_30467);
or U39300 (N_39300,N_33713,N_32963);
and U39301 (N_39301,N_34479,N_31328);
nor U39302 (N_39302,N_31930,N_31090);
nand U39303 (N_39303,N_30227,N_33374);
and U39304 (N_39304,N_34446,N_33711);
nand U39305 (N_39305,N_30667,N_34610);
or U39306 (N_39306,N_30520,N_30090);
and U39307 (N_39307,N_30805,N_32968);
nor U39308 (N_39308,N_30857,N_31884);
and U39309 (N_39309,N_33445,N_30310);
nor U39310 (N_39310,N_30232,N_32798);
or U39311 (N_39311,N_34835,N_30203);
xor U39312 (N_39312,N_31055,N_33632);
nand U39313 (N_39313,N_32622,N_34779);
or U39314 (N_39314,N_31603,N_34749);
xnor U39315 (N_39315,N_31518,N_32888);
nor U39316 (N_39316,N_34405,N_33832);
nand U39317 (N_39317,N_31122,N_31965);
or U39318 (N_39318,N_34127,N_30516);
xnor U39319 (N_39319,N_34491,N_34180);
nor U39320 (N_39320,N_30329,N_31666);
nand U39321 (N_39321,N_32564,N_31002);
and U39322 (N_39322,N_30264,N_33334);
nand U39323 (N_39323,N_31249,N_32185);
nor U39324 (N_39324,N_32068,N_32559);
nor U39325 (N_39325,N_32636,N_31109);
nand U39326 (N_39326,N_34474,N_30504);
nor U39327 (N_39327,N_30897,N_32557);
xor U39328 (N_39328,N_30519,N_32417);
or U39329 (N_39329,N_33094,N_31501);
or U39330 (N_39330,N_34121,N_30651);
and U39331 (N_39331,N_32014,N_34977);
nor U39332 (N_39332,N_33308,N_30031);
nor U39333 (N_39333,N_30151,N_33377);
nand U39334 (N_39334,N_30881,N_32402);
nand U39335 (N_39335,N_31447,N_34223);
or U39336 (N_39336,N_34670,N_33861);
or U39337 (N_39337,N_32076,N_30102);
or U39338 (N_39338,N_33658,N_33462);
nand U39339 (N_39339,N_33599,N_33411);
nand U39340 (N_39340,N_34862,N_33796);
nand U39341 (N_39341,N_33221,N_33709);
nor U39342 (N_39342,N_33926,N_31064);
nor U39343 (N_39343,N_33934,N_30867);
nand U39344 (N_39344,N_32753,N_34959);
nand U39345 (N_39345,N_34357,N_33558);
and U39346 (N_39346,N_32311,N_33135);
or U39347 (N_39347,N_30105,N_31162);
and U39348 (N_39348,N_31348,N_33425);
nor U39349 (N_39349,N_31880,N_33886);
and U39350 (N_39350,N_30809,N_30512);
and U39351 (N_39351,N_33922,N_34747);
xor U39352 (N_39352,N_31536,N_33709);
nor U39353 (N_39353,N_30887,N_34679);
or U39354 (N_39354,N_30836,N_32184);
nand U39355 (N_39355,N_30639,N_34367);
xor U39356 (N_39356,N_34168,N_31093);
nand U39357 (N_39357,N_33151,N_31542);
and U39358 (N_39358,N_32251,N_34553);
and U39359 (N_39359,N_33150,N_31359);
nor U39360 (N_39360,N_33104,N_34034);
or U39361 (N_39361,N_31538,N_31314);
or U39362 (N_39362,N_30715,N_33140);
or U39363 (N_39363,N_33623,N_30068);
and U39364 (N_39364,N_31798,N_32408);
xor U39365 (N_39365,N_31107,N_31072);
nor U39366 (N_39366,N_32818,N_34051);
nor U39367 (N_39367,N_34624,N_31632);
and U39368 (N_39368,N_34380,N_32957);
xor U39369 (N_39369,N_32217,N_30838);
or U39370 (N_39370,N_34855,N_33610);
xnor U39371 (N_39371,N_30665,N_33350);
xnor U39372 (N_39372,N_31448,N_30685);
xor U39373 (N_39373,N_30851,N_34403);
or U39374 (N_39374,N_30361,N_31858);
xnor U39375 (N_39375,N_30350,N_32250);
and U39376 (N_39376,N_34022,N_32390);
nand U39377 (N_39377,N_32306,N_31747);
nor U39378 (N_39378,N_32733,N_33128);
nor U39379 (N_39379,N_33906,N_32739);
or U39380 (N_39380,N_33615,N_33956);
nor U39381 (N_39381,N_33475,N_32059);
or U39382 (N_39382,N_34108,N_31469);
and U39383 (N_39383,N_34853,N_32654);
nor U39384 (N_39384,N_30403,N_33449);
xnor U39385 (N_39385,N_33863,N_31844);
nor U39386 (N_39386,N_33101,N_31208);
xnor U39387 (N_39387,N_34388,N_30442);
or U39388 (N_39388,N_30092,N_32704);
nand U39389 (N_39389,N_31998,N_34352);
or U39390 (N_39390,N_30072,N_34282);
or U39391 (N_39391,N_32402,N_31608);
nand U39392 (N_39392,N_30362,N_32249);
and U39393 (N_39393,N_31763,N_32330);
nor U39394 (N_39394,N_33794,N_33751);
and U39395 (N_39395,N_33252,N_33727);
or U39396 (N_39396,N_31180,N_31103);
nor U39397 (N_39397,N_30106,N_30097);
nor U39398 (N_39398,N_31641,N_34280);
nand U39399 (N_39399,N_32400,N_34928);
or U39400 (N_39400,N_33830,N_34207);
xnor U39401 (N_39401,N_31760,N_30153);
or U39402 (N_39402,N_32245,N_34998);
nand U39403 (N_39403,N_33783,N_33637);
or U39404 (N_39404,N_32477,N_34879);
xnor U39405 (N_39405,N_30975,N_31158);
xor U39406 (N_39406,N_34062,N_32373);
or U39407 (N_39407,N_32844,N_32809);
and U39408 (N_39408,N_31355,N_33219);
and U39409 (N_39409,N_32517,N_32326);
and U39410 (N_39410,N_33617,N_33871);
nand U39411 (N_39411,N_31903,N_30174);
xnor U39412 (N_39412,N_32946,N_33898);
nand U39413 (N_39413,N_30927,N_33394);
and U39414 (N_39414,N_30212,N_30061);
or U39415 (N_39415,N_34612,N_31072);
or U39416 (N_39416,N_33594,N_30993);
xnor U39417 (N_39417,N_33298,N_31858);
nand U39418 (N_39418,N_31420,N_33660);
and U39419 (N_39419,N_32787,N_31074);
nor U39420 (N_39420,N_33043,N_30446);
or U39421 (N_39421,N_33728,N_32701);
nor U39422 (N_39422,N_33996,N_31701);
xnor U39423 (N_39423,N_31491,N_32866);
and U39424 (N_39424,N_30480,N_32163);
nand U39425 (N_39425,N_34011,N_30376);
nor U39426 (N_39426,N_33557,N_33219);
xor U39427 (N_39427,N_34657,N_30484);
or U39428 (N_39428,N_30067,N_32622);
nand U39429 (N_39429,N_30542,N_30615);
or U39430 (N_39430,N_32595,N_32837);
nor U39431 (N_39431,N_31647,N_34024);
xnor U39432 (N_39432,N_33849,N_30387);
xnor U39433 (N_39433,N_34629,N_33300);
nor U39434 (N_39434,N_32224,N_34227);
xnor U39435 (N_39435,N_30434,N_30389);
nand U39436 (N_39436,N_31251,N_30466);
or U39437 (N_39437,N_31305,N_34610);
xor U39438 (N_39438,N_33288,N_31821);
nand U39439 (N_39439,N_31981,N_32440);
and U39440 (N_39440,N_30154,N_34176);
nand U39441 (N_39441,N_34864,N_31007);
and U39442 (N_39442,N_31779,N_32882);
nor U39443 (N_39443,N_33189,N_34334);
nor U39444 (N_39444,N_31256,N_30169);
xnor U39445 (N_39445,N_31047,N_34706);
or U39446 (N_39446,N_33064,N_34949);
and U39447 (N_39447,N_34539,N_34158);
or U39448 (N_39448,N_33352,N_34091);
or U39449 (N_39449,N_34753,N_31059);
or U39450 (N_39450,N_31583,N_30441);
xnor U39451 (N_39451,N_31353,N_34444);
or U39452 (N_39452,N_32285,N_34415);
nor U39453 (N_39453,N_32179,N_33515);
xnor U39454 (N_39454,N_30743,N_33817);
and U39455 (N_39455,N_33348,N_32966);
and U39456 (N_39456,N_31094,N_33900);
xnor U39457 (N_39457,N_34971,N_33281);
xnor U39458 (N_39458,N_31362,N_31782);
nor U39459 (N_39459,N_33553,N_30327);
nand U39460 (N_39460,N_30932,N_31297);
nand U39461 (N_39461,N_31539,N_33927);
or U39462 (N_39462,N_30236,N_34057);
nor U39463 (N_39463,N_30158,N_30186);
xnor U39464 (N_39464,N_34173,N_32702);
xnor U39465 (N_39465,N_33089,N_33874);
nand U39466 (N_39466,N_34928,N_32140);
or U39467 (N_39467,N_31153,N_34343);
nor U39468 (N_39468,N_33221,N_32291);
or U39469 (N_39469,N_31447,N_34955);
nand U39470 (N_39470,N_31002,N_33515);
and U39471 (N_39471,N_32572,N_33568);
nor U39472 (N_39472,N_34260,N_33480);
or U39473 (N_39473,N_32007,N_33124);
or U39474 (N_39474,N_30125,N_33625);
xor U39475 (N_39475,N_31476,N_32272);
xnor U39476 (N_39476,N_30075,N_33020);
and U39477 (N_39477,N_32885,N_34901);
xor U39478 (N_39478,N_31014,N_32234);
nand U39479 (N_39479,N_32893,N_34510);
nor U39480 (N_39480,N_31468,N_32385);
nor U39481 (N_39481,N_32065,N_30919);
or U39482 (N_39482,N_32683,N_32862);
xor U39483 (N_39483,N_32449,N_31540);
nand U39484 (N_39484,N_31125,N_32311);
nor U39485 (N_39485,N_31020,N_32245);
nor U39486 (N_39486,N_33978,N_33942);
or U39487 (N_39487,N_31606,N_31926);
xnor U39488 (N_39488,N_34079,N_34407);
nand U39489 (N_39489,N_33748,N_33412);
xor U39490 (N_39490,N_34814,N_33113);
xnor U39491 (N_39491,N_30080,N_34430);
nand U39492 (N_39492,N_33851,N_32044);
and U39493 (N_39493,N_31866,N_30833);
and U39494 (N_39494,N_32975,N_30606);
nor U39495 (N_39495,N_34006,N_32772);
and U39496 (N_39496,N_33107,N_32212);
nand U39497 (N_39497,N_34841,N_32855);
and U39498 (N_39498,N_34661,N_32386);
and U39499 (N_39499,N_34517,N_30797);
and U39500 (N_39500,N_31124,N_31798);
or U39501 (N_39501,N_33959,N_34304);
nand U39502 (N_39502,N_31528,N_34417);
nand U39503 (N_39503,N_34327,N_33510);
or U39504 (N_39504,N_30806,N_33702);
and U39505 (N_39505,N_32837,N_32491);
nand U39506 (N_39506,N_32773,N_31247);
and U39507 (N_39507,N_31375,N_31249);
and U39508 (N_39508,N_32917,N_32337);
nand U39509 (N_39509,N_33398,N_31978);
or U39510 (N_39510,N_33807,N_31258);
xnor U39511 (N_39511,N_30329,N_31830);
or U39512 (N_39512,N_34716,N_34051);
nand U39513 (N_39513,N_33147,N_33833);
nand U39514 (N_39514,N_31369,N_34746);
nand U39515 (N_39515,N_32309,N_30382);
nor U39516 (N_39516,N_34886,N_31426);
xor U39517 (N_39517,N_30808,N_33759);
xnor U39518 (N_39518,N_30624,N_32944);
nor U39519 (N_39519,N_31530,N_34625);
nor U39520 (N_39520,N_33175,N_32923);
or U39521 (N_39521,N_32313,N_34754);
or U39522 (N_39522,N_31075,N_31795);
or U39523 (N_39523,N_30850,N_31217);
nor U39524 (N_39524,N_33487,N_34340);
and U39525 (N_39525,N_32146,N_30413);
xor U39526 (N_39526,N_34061,N_33196);
nor U39527 (N_39527,N_33033,N_31719);
or U39528 (N_39528,N_34133,N_32743);
nor U39529 (N_39529,N_34459,N_32337);
or U39530 (N_39530,N_33097,N_34888);
and U39531 (N_39531,N_32475,N_34278);
nand U39532 (N_39532,N_33747,N_34580);
and U39533 (N_39533,N_34149,N_34721);
or U39534 (N_39534,N_32679,N_34508);
and U39535 (N_39535,N_34230,N_31752);
or U39536 (N_39536,N_31264,N_30581);
nand U39537 (N_39537,N_34396,N_30045);
nand U39538 (N_39538,N_34415,N_34376);
xnor U39539 (N_39539,N_33300,N_32878);
xnor U39540 (N_39540,N_33300,N_34860);
and U39541 (N_39541,N_31616,N_31435);
xor U39542 (N_39542,N_31934,N_34096);
xor U39543 (N_39543,N_30904,N_30926);
or U39544 (N_39544,N_30636,N_34365);
and U39545 (N_39545,N_32356,N_33236);
nor U39546 (N_39546,N_30296,N_32507);
xnor U39547 (N_39547,N_33043,N_32851);
nand U39548 (N_39548,N_30087,N_32361);
nand U39549 (N_39549,N_33299,N_31815);
nor U39550 (N_39550,N_32795,N_32492);
nand U39551 (N_39551,N_33383,N_30524);
and U39552 (N_39552,N_34233,N_33904);
xor U39553 (N_39553,N_33499,N_32449);
nor U39554 (N_39554,N_32808,N_34637);
or U39555 (N_39555,N_34109,N_32680);
or U39556 (N_39556,N_34158,N_33221);
nor U39557 (N_39557,N_31929,N_31555);
and U39558 (N_39558,N_31851,N_30069);
nor U39559 (N_39559,N_30763,N_31828);
and U39560 (N_39560,N_30116,N_34455);
and U39561 (N_39561,N_34121,N_31001);
nand U39562 (N_39562,N_33876,N_33945);
nor U39563 (N_39563,N_30031,N_32773);
and U39564 (N_39564,N_31334,N_31427);
nor U39565 (N_39565,N_32867,N_34530);
nand U39566 (N_39566,N_33357,N_33096);
nor U39567 (N_39567,N_34848,N_30969);
and U39568 (N_39568,N_33253,N_31496);
or U39569 (N_39569,N_30298,N_30619);
nor U39570 (N_39570,N_34737,N_30290);
or U39571 (N_39571,N_32536,N_31060);
nor U39572 (N_39572,N_30701,N_32452);
xor U39573 (N_39573,N_30756,N_30804);
xnor U39574 (N_39574,N_31341,N_30342);
or U39575 (N_39575,N_30894,N_33963);
or U39576 (N_39576,N_30516,N_31420);
xor U39577 (N_39577,N_34155,N_33497);
nand U39578 (N_39578,N_32384,N_33699);
or U39579 (N_39579,N_32585,N_31811);
or U39580 (N_39580,N_30272,N_32124);
and U39581 (N_39581,N_32829,N_30664);
and U39582 (N_39582,N_34459,N_30250);
and U39583 (N_39583,N_32647,N_30298);
nand U39584 (N_39584,N_33656,N_33771);
nand U39585 (N_39585,N_32216,N_31960);
and U39586 (N_39586,N_33703,N_33463);
xnor U39587 (N_39587,N_31236,N_32492);
or U39588 (N_39588,N_32025,N_34727);
and U39589 (N_39589,N_32623,N_34697);
and U39590 (N_39590,N_30810,N_31045);
xor U39591 (N_39591,N_33882,N_31676);
xor U39592 (N_39592,N_33817,N_33039);
nand U39593 (N_39593,N_30422,N_33813);
xnor U39594 (N_39594,N_31817,N_34718);
or U39595 (N_39595,N_33415,N_30398);
and U39596 (N_39596,N_32187,N_33344);
nand U39597 (N_39597,N_34802,N_32796);
nand U39598 (N_39598,N_30241,N_33495);
nor U39599 (N_39599,N_32797,N_32484);
nor U39600 (N_39600,N_30056,N_31312);
nand U39601 (N_39601,N_33161,N_30820);
or U39602 (N_39602,N_30355,N_30232);
or U39603 (N_39603,N_32266,N_32534);
and U39604 (N_39604,N_30873,N_30218);
or U39605 (N_39605,N_32966,N_32984);
xnor U39606 (N_39606,N_33250,N_32001);
or U39607 (N_39607,N_33732,N_31554);
and U39608 (N_39608,N_32534,N_34968);
and U39609 (N_39609,N_33039,N_32613);
nor U39610 (N_39610,N_32300,N_31697);
nand U39611 (N_39611,N_31475,N_34325);
nor U39612 (N_39612,N_31718,N_33383);
and U39613 (N_39613,N_30985,N_34836);
xnor U39614 (N_39614,N_33374,N_30745);
xnor U39615 (N_39615,N_33214,N_30312);
or U39616 (N_39616,N_31870,N_30139);
or U39617 (N_39617,N_30083,N_33788);
nand U39618 (N_39618,N_32092,N_34278);
and U39619 (N_39619,N_31625,N_31277);
or U39620 (N_39620,N_31097,N_31192);
or U39621 (N_39621,N_31430,N_34734);
xor U39622 (N_39622,N_30145,N_34651);
or U39623 (N_39623,N_31747,N_33017);
xor U39624 (N_39624,N_33886,N_32782);
nor U39625 (N_39625,N_33529,N_31411);
or U39626 (N_39626,N_32618,N_34674);
xor U39627 (N_39627,N_31508,N_33160);
nand U39628 (N_39628,N_32952,N_32865);
nand U39629 (N_39629,N_32932,N_34722);
and U39630 (N_39630,N_32364,N_32231);
and U39631 (N_39631,N_34186,N_33070);
nand U39632 (N_39632,N_33983,N_31320);
or U39633 (N_39633,N_32990,N_33384);
or U39634 (N_39634,N_34642,N_32797);
xnor U39635 (N_39635,N_32258,N_30073);
xnor U39636 (N_39636,N_30267,N_33044);
nand U39637 (N_39637,N_34943,N_31095);
nor U39638 (N_39638,N_32593,N_32438);
and U39639 (N_39639,N_33870,N_31810);
nand U39640 (N_39640,N_30288,N_31500);
and U39641 (N_39641,N_34969,N_33834);
nor U39642 (N_39642,N_31174,N_30297);
xnor U39643 (N_39643,N_33993,N_34759);
and U39644 (N_39644,N_33023,N_30416);
nand U39645 (N_39645,N_34205,N_32203);
nor U39646 (N_39646,N_31207,N_30458);
nor U39647 (N_39647,N_31421,N_31128);
nand U39648 (N_39648,N_34873,N_31034);
nor U39649 (N_39649,N_34196,N_33043);
or U39650 (N_39650,N_30759,N_31485);
nor U39651 (N_39651,N_32852,N_34855);
or U39652 (N_39652,N_34840,N_32012);
xor U39653 (N_39653,N_32797,N_31260);
xor U39654 (N_39654,N_30222,N_33088);
xnor U39655 (N_39655,N_34490,N_30759);
and U39656 (N_39656,N_34867,N_30666);
or U39657 (N_39657,N_34325,N_34597);
nand U39658 (N_39658,N_32112,N_30002);
nand U39659 (N_39659,N_32775,N_31405);
nand U39660 (N_39660,N_34461,N_34602);
nor U39661 (N_39661,N_30701,N_32837);
nand U39662 (N_39662,N_33027,N_30725);
nand U39663 (N_39663,N_34238,N_34717);
and U39664 (N_39664,N_34622,N_34598);
nor U39665 (N_39665,N_33056,N_31281);
or U39666 (N_39666,N_31780,N_31488);
or U39667 (N_39667,N_32668,N_32390);
xnor U39668 (N_39668,N_30640,N_31233);
and U39669 (N_39669,N_30354,N_30605);
xnor U39670 (N_39670,N_31839,N_34256);
and U39671 (N_39671,N_31125,N_30811);
nor U39672 (N_39672,N_30358,N_30070);
or U39673 (N_39673,N_31774,N_30974);
nand U39674 (N_39674,N_33085,N_30205);
nor U39675 (N_39675,N_30334,N_31703);
nor U39676 (N_39676,N_33910,N_30880);
or U39677 (N_39677,N_33784,N_34346);
and U39678 (N_39678,N_33114,N_31985);
or U39679 (N_39679,N_31901,N_31294);
nand U39680 (N_39680,N_32117,N_30673);
nor U39681 (N_39681,N_34874,N_31767);
nand U39682 (N_39682,N_30091,N_34422);
or U39683 (N_39683,N_33141,N_34755);
nor U39684 (N_39684,N_31045,N_33566);
and U39685 (N_39685,N_30803,N_33576);
nand U39686 (N_39686,N_30640,N_31131);
xor U39687 (N_39687,N_30232,N_30943);
or U39688 (N_39688,N_30948,N_33707);
and U39689 (N_39689,N_34378,N_34463);
or U39690 (N_39690,N_33290,N_34368);
or U39691 (N_39691,N_31934,N_34272);
nor U39692 (N_39692,N_33714,N_34234);
xor U39693 (N_39693,N_33486,N_30788);
or U39694 (N_39694,N_31518,N_34705);
nand U39695 (N_39695,N_31656,N_31280);
xor U39696 (N_39696,N_34546,N_34586);
nor U39697 (N_39697,N_34929,N_30449);
nand U39698 (N_39698,N_34023,N_31407);
or U39699 (N_39699,N_34608,N_30751);
nand U39700 (N_39700,N_32339,N_34264);
nand U39701 (N_39701,N_33959,N_32226);
nor U39702 (N_39702,N_33040,N_31849);
nand U39703 (N_39703,N_31752,N_31864);
and U39704 (N_39704,N_31461,N_31463);
nand U39705 (N_39705,N_34598,N_31952);
xor U39706 (N_39706,N_33876,N_32536);
xnor U39707 (N_39707,N_31804,N_32425);
nand U39708 (N_39708,N_34235,N_34497);
xor U39709 (N_39709,N_31825,N_30826);
nand U39710 (N_39710,N_32758,N_30202);
nand U39711 (N_39711,N_30535,N_32848);
nand U39712 (N_39712,N_33333,N_31452);
nand U39713 (N_39713,N_31074,N_33480);
nand U39714 (N_39714,N_30846,N_32309);
xnor U39715 (N_39715,N_31352,N_33099);
nand U39716 (N_39716,N_30962,N_32129);
nor U39717 (N_39717,N_31394,N_33671);
nor U39718 (N_39718,N_32599,N_30078);
nor U39719 (N_39719,N_34728,N_34522);
and U39720 (N_39720,N_33730,N_32381);
nor U39721 (N_39721,N_30241,N_30721);
nor U39722 (N_39722,N_33556,N_30526);
nand U39723 (N_39723,N_31347,N_33642);
nand U39724 (N_39724,N_32891,N_34532);
nand U39725 (N_39725,N_33965,N_31409);
nand U39726 (N_39726,N_30246,N_30822);
xnor U39727 (N_39727,N_33965,N_32074);
xnor U39728 (N_39728,N_30850,N_33529);
and U39729 (N_39729,N_31225,N_31297);
nand U39730 (N_39730,N_34365,N_34453);
and U39731 (N_39731,N_32336,N_34114);
nor U39732 (N_39732,N_31668,N_34708);
and U39733 (N_39733,N_33212,N_30715);
nor U39734 (N_39734,N_30356,N_32595);
and U39735 (N_39735,N_32135,N_33179);
xnor U39736 (N_39736,N_30347,N_30018);
and U39737 (N_39737,N_31949,N_33423);
and U39738 (N_39738,N_33936,N_33663);
nand U39739 (N_39739,N_33117,N_33440);
xnor U39740 (N_39740,N_30191,N_30462);
nand U39741 (N_39741,N_30321,N_30413);
nand U39742 (N_39742,N_31551,N_33927);
and U39743 (N_39743,N_33195,N_33478);
nand U39744 (N_39744,N_32809,N_30799);
and U39745 (N_39745,N_33590,N_30851);
nand U39746 (N_39746,N_33118,N_30607);
and U39747 (N_39747,N_33122,N_31679);
and U39748 (N_39748,N_32042,N_32008);
and U39749 (N_39749,N_31668,N_31765);
nor U39750 (N_39750,N_34137,N_31291);
nor U39751 (N_39751,N_31861,N_30851);
or U39752 (N_39752,N_32964,N_33903);
xor U39753 (N_39753,N_31818,N_33808);
nor U39754 (N_39754,N_33904,N_30051);
nor U39755 (N_39755,N_31739,N_31354);
nand U39756 (N_39756,N_30022,N_31657);
nor U39757 (N_39757,N_32049,N_33719);
xnor U39758 (N_39758,N_34915,N_33429);
or U39759 (N_39759,N_32514,N_31128);
nor U39760 (N_39760,N_31797,N_33448);
nand U39761 (N_39761,N_34827,N_30472);
and U39762 (N_39762,N_31584,N_31183);
xor U39763 (N_39763,N_34644,N_32018);
or U39764 (N_39764,N_34506,N_33316);
and U39765 (N_39765,N_30653,N_33799);
nor U39766 (N_39766,N_34418,N_31196);
xnor U39767 (N_39767,N_32610,N_31092);
nor U39768 (N_39768,N_31533,N_33660);
or U39769 (N_39769,N_31661,N_31875);
or U39770 (N_39770,N_31488,N_32629);
or U39771 (N_39771,N_34827,N_33581);
and U39772 (N_39772,N_34270,N_31907);
nor U39773 (N_39773,N_32900,N_33514);
xnor U39774 (N_39774,N_33936,N_30924);
xnor U39775 (N_39775,N_34705,N_32004);
and U39776 (N_39776,N_32195,N_32023);
and U39777 (N_39777,N_34812,N_34111);
xnor U39778 (N_39778,N_31188,N_31685);
xnor U39779 (N_39779,N_32698,N_30152);
or U39780 (N_39780,N_32356,N_31551);
and U39781 (N_39781,N_34038,N_33643);
and U39782 (N_39782,N_34313,N_34429);
nor U39783 (N_39783,N_34281,N_32807);
nand U39784 (N_39784,N_32827,N_30452);
or U39785 (N_39785,N_33549,N_33381);
xor U39786 (N_39786,N_33892,N_31712);
or U39787 (N_39787,N_34215,N_33247);
nor U39788 (N_39788,N_33413,N_31092);
or U39789 (N_39789,N_33803,N_34329);
and U39790 (N_39790,N_33783,N_34998);
nor U39791 (N_39791,N_30648,N_30314);
and U39792 (N_39792,N_34939,N_33264);
nand U39793 (N_39793,N_32981,N_34971);
or U39794 (N_39794,N_34968,N_33794);
or U39795 (N_39795,N_31322,N_34676);
nand U39796 (N_39796,N_31126,N_33956);
nor U39797 (N_39797,N_33378,N_31641);
xor U39798 (N_39798,N_32260,N_33040);
nor U39799 (N_39799,N_31453,N_30226);
nand U39800 (N_39800,N_31859,N_32813);
xor U39801 (N_39801,N_31947,N_30910);
and U39802 (N_39802,N_33125,N_32910);
xor U39803 (N_39803,N_34277,N_34451);
or U39804 (N_39804,N_33368,N_34405);
and U39805 (N_39805,N_34918,N_31719);
xor U39806 (N_39806,N_32440,N_32874);
or U39807 (N_39807,N_32460,N_31673);
or U39808 (N_39808,N_34525,N_30031);
nor U39809 (N_39809,N_33169,N_33063);
or U39810 (N_39810,N_34543,N_33445);
and U39811 (N_39811,N_30627,N_34821);
nor U39812 (N_39812,N_30839,N_31318);
xnor U39813 (N_39813,N_31628,N_33230);
nor U39814 (N_39814,N_31809,N_34032);
nor U39815 (N_39815,N_31399,N_31542);
and U39816 (N_39816,N_31658,N_31902);
nor U39817 (N_39817,N_31552,N_30926);
and U39818 (N_39818,N_33563,N_34392);
xnor U39819 (N_39819,N_32507,N_32427);
xor U39820 (N_39820,N_34278,N_30771);
nor U39821 (N_39821,N_30877,N_32187);
nor U39822 (N_39822,N_31850,N_33127);
or U39823 (N_39823,N_32282,N_33700);
or U39824 (N_39824,N_31078,N_30234);
xnor U39825 (N_39825,N_34518,N_31772);
and U39826 (N_39826,N_34861,N_31247);
nand U39827 (N_39827,N_33897,N_33132);
nand U39828 (N_39828,N_33895,N_33234);
and U39829 (N_39829,N_30887,N_30546);
nor U39830 (N_39830,N_32836,N_33661);
and U39831 (N_39831,N_32223,N_34018);
and U39832 (N_39832,N_32298,N_34126);
xor U39833 (N_39833,N_32666,N_34590);
or U39834 (N_39834,N_32149,N_33044);
and U39835 (N_39835,N_30170,N_34389);
nor U39836 (N_39836,N_33492,N_31031);
nand U39837 (N_39837,N_32064,N_34150);
xnor U39838 (N_39838,N_34804,N_34328);
or U39839 (N_39839,N_33156,N_30580);
or U39840 (N_39840,N_30401,N_31926);
and U39841 (N_39841,N_30587,N_33524);
nor U39842 (N_39842,N_31602,N_31419);
and U39843 (N_39843,N_32998,N_30017);
or U39844 (N_39844,N_34997,N_32101);
nor U39845 (N_39845,N_31400,N_30958);
or U39846 (N_39846,N_31116,N_31702);
nand U39847 (N_39847,N_33066,N_30211);
xnor U39848 (N_39848,N_31673,N_30375);
nand U39849 (N_39849,N_33169,N_31708);
or U39850 (N_39850,N_34962,N_30159);
xnor U39851 (N_39851,N_34838,N_33717);
or U39852 (N_39852,N_32572,N_33641);
xor U39853 (N_39853,N_31735,N_33576);
and U39854 (N_39854,N_32681,N_31408);
nand U39855 (N_39855,N_32678,N_32219);
nand U39856 (N_39856,N_31702,N_30177);
nand U39857 (N_39857,N_33969,N_33130);
xor U39858 (N_39858,N_31796,N_34614);
xor U39859 (N_39859,N_33029,N_31545);
and U39860 (N_39860,N_31189,N_32734);
or U39861 (N_39861,N_30389,N_30501);
nor U39862 (N_39862,N_30359,N_31911);
and U39863 (N_39863,N_30119,N_33243);
nor U39864 (N_39864,N_32393,N_34686);
and U39865 (N_39865,N_31514,N_31427);
nor U39866 (N_39866,N_33651,N_32394);
xor U39867 (N_39867,N_31865,N_33629);
nor U39868 (N_39868,N_34116,N_32421);
nand U39869 (N_39869,N_33554,N_33656);
and U39870 (N_39870,N_32054,N_31987);
nor U39871 (N_39871,N_33768,N_32100);
or U39872 (N_39872,N_33456,N_33980);
and U39873 (N_39873,N_34722,N_30663);
and U39874 (N_39874,N_31699,N_31803);
or U39875 (N_39875,N_34100,N_34093);
xor U39876 (N_39876,N_32999,N_34948);
xnor U39877 (N_39877,N_33545,N_33260);
nand U39878 (N_39878,N_34331,N_31117);
and U39879 (N_39879,N_31698,N_34990);
xnor U39880 (N_39880,N_32041,N_32443);
nor U39881 (N_39881,N_32084,N_30355);
or U39882 (N_39882,N_33522,N_31846);
nor U39883 (N_39883,N_30665,N_31263);
or U39884 (N_39884,N_33676,N_30453);
nand U39885 (N_39885,N_32325,N_31642);
nand U39886 (N_39886,N_30902,N_30042);
xor U39887 (N_39887,N_32139,N_32282);
nand U39888 (N_39888,N_34825,N_34719);
or U39889 (N_39889,N_32446,N_33077);
nor U39890 (N_39890,N_33106,N_34291);
nand U39891 (N_39891,N_31413,N_32263);
and U39892 (N_39892,N_33568,N_32100);
xor U39893 (N_39893,N_31901,N_33458);
xnor U39894 (N_39894,N_33455,N_31037);
xor U39895 (N_39895,N_32287,N_33224);
nor U39896 (N_39896,N_32384,N_30578);
xnor U39897 (N_39897,N_31942,N_31034);
xor U39898 (N_39898,N_34921,N_33552);
nor U39899 (N_39899,N_33305,N_32784);
nor U39900 (N_39900,N_32381,N_31251);
or U39901 (N_39901,N_33647,N_30338);
and U39902 (N_39902,N_30247,N_32347);
or U39903 (N_39903,N_30918,N_32133);
nand U39904 (N_39904,N_33896,N_31602);
nand U39905 (N_39905,N_33157,N_34031);
or U39906 (N_39906,N_34438,N_33988);
and U39907 (N_39907,N_32846,N_30325);
and U39908 (N_39908,N_34518,N_30330);
or U39909 (N_39909,N_34004,N_33873);
nand U39910 (N_39910,N_34725,N_31777);
nor U39911 (N_39911,N_34491,N_30911);
nand U39912 (N_39912,N_32847,N_33023);
or U39913 (N_39913,N_33609,N_31314);
xnor U39914 (N_39914,N_31924,N_30563);
xnor U39915 (N_39915,N_34979,N_31531);
nand U39916 (N_39916,N_30119,N_33960);
nor U39917 (N_39917,N_33525,N_33955);
or U39918 (N_39918,N_33148,N_30884);
nor U39919 (N_39919,N_33898,N_34342);
xnor U39920 (N_39920,N_32976,N_32309);
nor U39921 (N_39921,N_33955,N_33201);
or U39922 (N_39922,N_31578,N_33007);
xnor U39923 (N_39923,N_31846,N_34651);
nor U39924 (N_39924,N_33611,N_32898);
or U39925 (N_39925,N_33703,N_33808);
or U39926 (N_39926,N_34796,N_31737);
and U39927 (N_39927,N_33547,N_30417);
and U39928 (N_39928,N_32775,N_30895);
or U39929 (N_39929,N_33351,N_30951);
nor U39930 (N_39930,N_34860,N_34108);
or U39931 (N_39931,N_32890,N_33166);
xnor U39932 (N_39932,N_30963,N_31838);
nor U39933 (N_39933,N_33941,N_33861);
nor U39934 (N_39934,N_34360,N_31678);
nand U39935 (N_39935,N_32021,N_30509);
nand U39936 (N_39936,N_33359,N_30038);
nand U39937 (N_39937,N_32007,N_31104);
nand U39938 (N_39938,N_32558,N_32513);
and U39939 (N_39939,N_34734,N_30727);
xor U39940 (N_39940,N_32909,N_32902);
and U39941 (N_39941,N_34032,N_34421);
nand U39942 (N_39942,N_31606,N_34322);
xnor U39943 (N_39943,N_33915,N_34762);
xnor U39944 (N_39944,N_32755,N_30581);
and U39945 (N_39945,N_33333,N_34194);
xor U39946 (N_39946,N_34605,N_33385);
or U39947 (N_39947,N_34043,N_31522);
or U39948 (N_39948,N_34077,N_31811);
or U39949 (N_39949,N_32018,N_34166);
and U39950 (N_39950,N_34996,N_33735);
or U39951 (N_39951,N_31690,N_31615);
xor U39952 (N_39952,N_32328,N_31554);
nand U39953 (N_39953,N_30162,N_32560);
or U39954 (N_39954,N_34372,N_32135);
and U39955 (N_39955,N_32021,N_30152);
xor U39956 (N_39956,N_30136,N_31366);
nand U39957 (N_39957,N_31760,N_33920);
nand U39958 (N_39958,N_33929,N_30419);
or U39959 (N_39959,N_33713,N_32024);
nor U39960 (N_39960,N_32183,N_31227);
nand U39961 (N_39961,N_34333,N_34438);
or U39962 (N_39962,N_34725,N_34667);
nor U39963 (N_39963,N_33201,N_33971);
or U39964 (N_39964,N_34282,N_31085);
nand U39965 (N_39965,N_33467,N_30818);
nor U39966 (N_39966,N_34085,N_33919);
nand U39967 (N_39967,N_30812,N_34752);
or U39968 (N_39968,N_31482,N_30274);
nand U39969 (N_39969,N_30108,N_31335);
nand U39970 (N_39970,N_34282,N_30597);
xnor U39971 (N_39971,N_34045,N_32628);
xor U39972 (N_39972,N_32441,N_32139);
and U39973 (N_39973,N_33847,N_31841);
xnor U39974 (N_39974,N_31635,N_30574);
or U39975 (N_39975,N_32737,N_34813);
nor U39976 (N_39976,N_34903,N_34615);
xnor U39977 (N_39977,N_32419,N_33598);
or U39978 (N_39978,N_32789,N_30471);
or U39979 (N_39979,N_33163,N_31403);
nand U39980 (N_39980,N_34219,N_34426);
and U39981 (N_39981,N_34059,N_31739);
or U39982 (N_39982,N_32056,N_33417);
and U39983 (N_39983,N_33943,N_34191);
and U39984 (N_39984,N_31086,N_34534);
and U39985 (N_39985,N_34414,N_31739);
nand U39986 (N_39986,N_33689,N_31525);
and U39987 (N_39987,N_32626,N_34364);
nand U39988 (N_39988,N_34915,N_32258);
nand U39989 (N_39989,N_31264,N_30873);
xor U39990 (N_39990,N_33737,N_30379);
nor U39991 (N_39991,N_30628,N_30907);
xnor U39992 (N_39992,N_31727,N_32074);
xor U39993 (N_39993,N_34573,N_33775);
nand U39994 (N_39994,N_34315,N_30363);
nand U39995 (N_39995,N_31911,N_30622);
and U39996 (N_39996,N_32527,N_33140);
nand U39997 (N_39997,N_32472,N_30615);
xor U39998 (N_39998,N_30593,N_33499);
nand U39999 (N_39999,N_32305,N_34045);
and U40000 (N_40000,N_38595,N_38553);
and U40001 (N_40001,N_35823,N_39705);
or U40002 (N_40002,N_38646,N_36311);
nand U40003 (N_40003,N_37954,N_38739);
nand U40004 (N_40004,N_36065,N_36153);
nand U40005 (N_40005,N_37735,N_38070);
xnor U40006 (N_40006,N_35730,N_36725);
nor U40007 (N_40007,N_39198,N_38356);
nor U40008 (N_40008,N_39357,N_39296);
nor U40009 (N_40009,N_39416,N_36588);
and U40010 (N_40010,N_37652,N_35598);
nand U40011 (N_40011,N_35695,N_35046);
and U40012 (N_40012,N_38610,N_39900);
nand U40013 (N_40013,N_38150,N_39631);
and U40014 (N_40014,N_37071,N_38639);
and U40015 (N_40015,N_39129,N_38557);
and U40016 (N_40016,N_35120,N_35790);
nor U40017 (N_40017,N_35160,N_37092);
and U40018 (N_40018,N_39204,N_35729);
nand U40019 (N_40019,N_36705,N_39516);
xor U40020 (N_40020,N_37523,N_38538);
xor U40021 (N_40021,N_38265,N_38143);
nand U40022 (N_40022,N_37074,N_38080);
nor U40023 (N_40023,N_38619,N_36056);
nor U40024 (N_40024,N_37687,N_37266);
nand U40025 (N_40025,N_38941,N_38732);
nand U40026 (N_40026,N_38787,N_39911);
nor U40027 (N_40027,N_38936,N_39724);
nand U40028 (N_40028,N_39811,N_38602);
or U40029 (N_40029,N_37208,N_38370);
and U40030 (N_40030,N_36748,N_37199);
xnor U40031 (N_40031,N_36080,N_39322);
and U40032 (N_40032,N_35216,N_35306);
or U40033 (N_40033,N_39594,N_37632);
nand U40034 (N_40034,N_36148,N_39879);
xnor U40035 (N_40035,N_37673,N_37176);
or U40036 (N_40036,N_39781,N_38653);
and U40037 (N_40037,N_35409,N_39346);
nand U40038 (N_40038,N_36838,N_38103);
or U40039 (N_40039,N_35118,N_37766);
and U40040 (N_40040,N_37893,N_38854);
nand U40041 (N_40041,N_39604,N_37636);
and U40042 (N_40042,N_39959,N_39017);
nor U40043 (N_40043,N_38466,N_39327);
or U40044 (N_40044,N_37680,N_37471);
and U40045 (N_40045,N_35948,N_36602);
nor U40046 (N_40046,N_35491,N_35609);
nand U40047 (N_40047,N_35067,N_38226);
nor U40048 (N_40048,N_38870,N_39754);
nand U40049 (N_40049,N_35566,N_36836);
xnor U40050 (N_40050,N_37103,N_39250);
nand U40051 (N_40051,N_38428,N_37884);
or U40052 (N_40052,N_39392,N_35440);
nor U40053 (N_40053,N_39007,N_37098);
or U40054 (N_40054,N_39200,N_38841);
nand U40055 (N_40055,N_36009,N_38568);
xor U40056 (N_40056,N_38254,N_38305);
nor U40057 (N_40057,N_38352,N_35559);
xor U40058 (N_40058,N_37007,N_39192);
xnor U40059 (N_40059,N_36561,N_38076);
nor U40060 (N_40060,N_37291,N_38307);
nor U40061 (N_40061,N_36414,N_36547);
nand U40062 (N_40062,N_38430,N_38863);
xor U40063 (N_40063,N_39929,N_35548);
nor U40064 (N_40064,N_39430,N_35125);
nand U40065 (N_40065,N_38446,N_39630);
nor U40066 (N_40066,N_38228,N_35465);
nor U40067 (N_40067,N_36323,N_35346);
or U40068 (N_40068,N_39719,N_35466);
nor U40069 (N_40069,N_36223,N_38661);
or U40070 (N_40070,N_39009,N_36644);
and U40071 (N_40071,N_38484,N_37231);
xnor U40072 (N_40072,N_35378,N_35229);
and U40073 (N_40073,N_37530,N_36142);
nor U40074 (N_40074,N_35347,N_36304);
nand U40075 (N_40075,N_37234,N_38346);
and U40076 (N_40076,N_36957,N_39972);
and U40077 (N_40077,N_36136,N_37505);
and U40078 (N_40078,N_36699,N_39442);
nand U40079 (N_40079,N_39868,N_35807);
xnor U40080 (N_40080,N_39949,N_36097);
and U40081 (N_40081,N_39272,N_37567);
nor U40082 (N_40082,N_36190,N_38458);
nor U40083 (N_40083,N_35716,N_37209);
xor U40084 (N_40084,N_38810,N_37412);
or U40085 (N_40085,N_39539,N_39030);
xnor U40086 (N_40086,N_36746,N_39497);
nand U40087 (N_40087,N_35536,N_39559);
nor U40088 (N_40088,N_36295,N_38620);
xnor U40089 (N_40089,N_39544,N_36900);
xnor U40090 (N_40090,N_35742,N_36254);
nor U40091 (N_40091,N_38770,N_38894);
and U40092 (N_40092,N_38139,N_39358);
xnor U40093 (N_40093,N_36884,N_37923);
nand U40094 (N_40094,N_38337,N_36260);
and U40095 (N_40095,N_37001,N_39141);
or U40096 (N_40096,N_35177,N_37562);
nand U40097 (N_40097,N_36268,N_37977);
and U40098 (N_40098,N_38581,N_37821);
or U40099 (N_40099,N_35145,N_38858);
or U40100 (N_40100,N_38644,N_39688);
or U40101 (N_40101,N_38845,N_36166);
nand U40102 (N_40102,N_39634,N_38249);
and U40103 (N_40103,N_35723,N_38611);
or U40104 (N_40104,N_37386,N_35843);
nor U40105 (N_40105,N_36848,N_38410);
xor U40106 (N_40106,N_39000,N_35093);
or U40107 (N_40107,N_39156,N_36845);
and U40108 (N_40108,N_39143,N_36904);
xor U40109 (N_40109,N_38758,N_35001);
xor U40110 (N_40110,N_39954,N_38270);
xnor U40111 (N_40111,N_37552,N_38792);
nand U40112 (N_40112,N_36639,N_36060);
xor U40113 (N_40113,N_36971,N_39838);
nand U40114 (N_40114,N_36182,N_39469);
or U40115 (N_40115,N_36025,N_37722);
or U40116 (N_40116,N_36513,N_37214);
or U40117 (N_40117,N_39494,N_38688);
or U40118 (N_40118,N_37450,N_35954);
or U40119 (N_40119,N_35249,N_38118);
nand U40120 (N_40120,N_38395,N_35579);
or U40121 (N_40121,N_35848,N_35867);
or U40122 (N_40122,N_37716,N_35567);
and U40123 (N_40123,N_38622,N_36171);
or U40124 (N_40124,N_38773,N_35753);
and U40125 (N_40125,N_36730,N_39027);
nor U40126 (N_40126,N_37187,N_39314);
nand U40127 (N_40127,N_39668,N_38185);
and U40128 (N_40128,N_37331,N_36791);
nor U40129 (N_40129,N_37065,N_35167);
and U40130 (N_40130,N_36839,N_39656);
or U40131 (N_40131,N_36282,N_35601);
nand U40132 (N_40132,N_35617,N_35087);
or U40133 (N_40133,N_36234,N_35907);
and U40134 (N_40134,N_38401,N_38396);
or U40135 (N_40135,N_39955,N_37759);
or U40136 (N_40136,N_36527,N_37825);
nand U40137 (N_40137,N_38426,N_37992);
or U40138 (N_40138,N_38393,N_35822);
nand U40139 (N_40139,N_39591,N_38585);
nand U40140 (N_40140,N_39093,N_37747);
nand U40141 (N_40141,N_38807,N_36494);
nor U40142 (N_40142,N_35999,N_36595);
nor U40143 (N_40143,N_35366,N_38981);
nor U40144 (N_40144,N_35205,N_36897);
and U40145 (N_40145,N_38781,N_36071);
nand U40146 (N_40146,N_39203,N_35824);
or U40147 (N_40147,N_36818,N_38210);
nor U40148 (N_40148,N_39536,N_37792);
nor U40149 (N_40149,N_38464,N_35626);
xnor U40150 (N_40150,N_37134,N_39409);
nand U40151 (N_40151,N_36445,N_38286);
nor U40152 (N_40152,N_36164,N_35804);
nand U40153 (N_40153,N_38282,N_39892);
and U40154 (N_40154,N_37996,N_35071);
xor U40155 (N_40155,N_37645,N_36870);
nor U40156 (N_40156,N_36624,N_39390);
nor U40157 (N_40157,N_39659,N_37487);
and U40158 (N_40158,N_39175,N_38264);
nor U40159 (N_40159,N_38711,N_37712);
nor U40160 (N_40160,N_37382,N_35452);
nand U40161 (N_40161,N_35628,N_35284);
or U40162 (N_40162,N_36331,N_39152);
nand U40163 (N_40163,N_35873,N_39712);
nor U40164 (N_40164,N_36714,N_38048);
or U40165 (N_40165,N_39827,N_39128);
xnor U40166 (N_40166,N_38895,N_39682);
nor U40167 (N_40167,N_39511,N_37162);
and U40168 (N_40168,N_37519,N_35812);
nor U40169 (N_40169,N_36069,N_37697);
nor U40170 (N_40170,N_39655,N_39839);
or U40171 (N_40171,N_36867,N_38178);
nand U40172 (N_40172,N_38660,N_38405);
nor U40173 (N_40173,N_36849,N_39064);
and U40174 (N_40174,N_39297,N_37038);
or U40175 (N_40175,N_37196,N_37940);
or U40176 (N_40176,N_35307,N_37273);
nor U40177 (N_40177,N_38234,N_38705);
nand U40178 (N_40178,N_39582,N_36517);
and U40179 (N_40179,N_36612,N_39319);
or U40180 (N_40180,N_35554,N_38427);
or U40181 (N_40181,N_39862,N_38368);
and U40182 (N_40182,N_35434,N_37077);
or U40183 (N_40183,N_38258,N_36021);
or U40184 (N_40184,N_38508,N_38175);
nor U40185 (N_40185,N_35015,N_38983);
xnor U40186 (N_40186,N_37922,N_36643);
or U40187 (N_40187,N_37517,N_35778);
nor U40188 (N_40188,N_36537,N_36873);
nand U40189 (N_40189,N_37477,N_36091);
and U40190 (N_40190,N_37538,N_39541);
nand U40191 (N_40191,N_39915,N_39350);
nor U40192 (N_40192,N_37686,N_37484);
nand U40193 (N_40193,N_39550,N_36912);
and U40194 (N_40194,N_38062,N_39347);
and U40195 (N_40195,N_36421,N_38822);
xor U40196 (N_40196,N_38495,N_38703);
and U40197 (N_40197,N_39041,N_36729);
nor U40198 (N_40198,N_38716,N_39340);
xor U40199 (N_40199,N_36023,N_35429);
and U40200 (N_40200,N_39570,N_39167);
or U40201 (N_40201,N_37627,N_36147);
xor U40202 (N_40202,N_37107,N_38003);
nand U40203 (N_40203,N_39254,N_38663);
or U40204 (N_40204,N_36563,N_35750);
and U40205 (N_40205,N_36666,N_37679);
and U40206 (N_40206,N_38712,N_36188);
nor U40207 (N_40207,N_38556,N_37560);
nand U40208 (N_40208,N_37163,N_36478);
and U40209 (N_40209,N_38179,N_37495);
xor U40210 (N_40210,N_37808,N_36345);
xor U40211 (N_40211,N_36129,N_37643);
xor U40212 (N_40212,N_39553,N_39320);
and U40213 (N_40213,N_38349,N_39509);
or U40214 (N_40214,N_35304,N_38676);
and U40215 (N_40215,N_36964,N_35510);
nand U40216 (N_40216,N_39366,N_38919);
nor U40217 (N_40217,N_36703,N_35870);
xnor U40218 (N_40218,N_37934,N_35631);
and U40219 (N_40219,N_36459,N_39782);
and U40220 (N_40220,N_38054,N_37730);
nand U40221 (N_40221,N_39482,N_35326);
nand U40222 (N_40222,N_35321,N_38574);
or U40223 (N_40223,N_36278,N_39211);
nand U40224 (N_40224,N_36031,N_39563);
and U40225 (N_40225,N_38387,N_37292);
or U40226 (N_40226,N_36231,N_37666);
or U40227 (N_40227,N_37483,N_39775);
xnor U40228 (N_40228,N_38905,N_36274);
or U40229 (N_40229,N_39164,N_36436);
xnor U40230 (N_40230,N_38443,N_36767);
nand U40231 (N_40231,N_36698,N_36202);
nor U40232 (N_40232,N_36638,N_38641);
nor U40233 (N_40233,N_36859,N_39987);
and U40234 (N_40234,N_36128,N_36280);
or U40235 (N_40235,N_38238,N_39794);
nand U40236 (N_40236,N_39124,N_37013);
and U40237 (N_40237,N_39413,N_39969);
xor U40238 (N_40238,N_39081,N_39617);
xor U40239 (N_40239,N_37704,N_35996);
nand U40240 (N_40240,N_37955,N_38885);
nand U40241 (N_40241,N_35426,N_37403);
nand U40242 (N_40242,N_36045,N_36843);
xor U40243 (N_40243,N_35511,N_35128);
nor U40244 (N_40244,N_36238,N_39807);
nor U40245 (N_40245,N_37556,N_35481);
or U40246 (N_40246,N_36435,N_36815);
and U40247 (N_40247,N_39339,N_37784);
and U40248 (N_40248,N_37375,N_35264);
xor U40249 (N_40249,N_35076,N_37201);
or U40250 (N_40250,N_38692,N_39680);
xor U40251 (N_40251,N_37698,N_36036);
xor U40252 (N_40252,N_36251,N_39005);
nand U40253 (N_40253,N_39336,N_35386);
nor U40254 (N_40254,N_38526,N_37540);
xor U40255 (N_40255,N_39377,N_38964);
or U40256 (N_40256,N_39761,N_35581);
or U40257 (N_40257,N_37016,N_39556);
nand U40258 (N_40258,N_37788,N_39595);
xnor U40259 (N_40259,N_35575,N_37758);
or U40260 (N_40260,N_39088,N_39084);
or U40261 (N_40261,N_38698,N_38880);
or U40262 (N_40262,N_35171,N_37387);
nand U40263 (N_40263,N_35668,N_37886);
nor U40264 (N_40264,N_36403,N_37147);
nor U40265 (N_40265,N_39345,N_35974);
or U40266 (N_40266,N_39528,N_39957);
xor U40267 (N_40267,N_37379,N_39445);
or U40268 (N_40268,N_38035,N_35134);
nand U40269 (N_40269,N_36784,N_38389);
nand U40270 (N_40270,N_35315,N_39933);
or U40271 (N_40271,N_38169,N_39732);
nand U40272 (N_40272,N_35914,N_39543);
xnor U40273 (N_40273,N_39993,N_35780);
and U40274 (N_40274,N_38051,N_38294);
nand U40275 (N_40275,N_35660,N_36505);
or U40276 (N_40276,N_37975,N_36812);
and U40277 (N_40277,N_35501,N_36012);
or U40278 (N_40278,N_38903,N_39814);
and U40279 (N_40279,N_35802,N_35963);
and U40280 (N_40280,N_35888,N_37101);
or U40281 (N_40281,N_36568,N_36918);
nand U40282 (N_40282,N_35016,N_36138);
or U40283 (N_40283,N_39845,N_39755);
and U40284 (N_40284,N_37261,N_35402);
xor U40285 (N_40285,N_35913,N_38757);
xor U40286 (N_40286,N_39239,N_35296);
and U40287 (N_40287,N_36498,N_38655);
and U40288 (N_40288,N_39676,N_35417);
and U40289 (N_40289,N_37568,N_39245);
nand U40290 (N_40290,N_36562,N_35681);
and U40291 (N_40291,N_37002,N_37858);
or U40292 (N_40292,N_37141,N_39852);
and U40293 (N_40293,N_38984,N_39998);
nor U40294 (N_40294,N_35165,N_39836);
nand U40295 (N_40295,N_36616,N_35130);
xnor U40296 (N_40296,N_37528,N_35073);
xor U40297 (N_40297,N_37145,N_37883);
and U40298 (N_40298,N_37976,N_37376);
and U40299 (N_40299,N_39766,N_37937);
and U40300 (N_40300,N_37900,N_39519);
nor U40301 (N_40301,N_39734,N_39759);
nor U40302 (N_40302,N_38291,N_37939);
nand U40303 (N_40303,N_39560,N_35184);
or U40304 (N_40304,N_39770,N_35140);
and U40305 (N_40305,N_36384,N_38252);
xor U40306 (N_40306,N_38884,N_38564);
or U40307 (N_40307,N_37212,N_37917);
nand U40308 (N_40308,N_35545,N_35217);
and U40309 (N_40309,N_36766,N_36104);
or U40310 (N_40310,N_36163,N_37526);
nand U40311 (N_40311,N_38119,N_38081);
or U40312 (N_40312,N_37449,N_39613);
or U40313 (N_40313,N_37596,N_39090);
or U40314 (N_40314,N_38956,N_35223);
nand U40315 (N_40315,N_35114,N_38162);
nor U40316 (N_40316,N_36370,N_37437);
or U40317 (N_40317,N_37272,N_37641);
xor U40318 (N_40318,N_36089,N_37262);
nand U40319 (N_40319,N_38590,N_36346);
and U40320 (N_40320,N_39155,N_37109);
and U40321 (N_40321,N_35613,N_37081);
nor U40322 (N_40322,N_36885,N_35933);
or U40323 (N_40323,N_38338,N_39580);
and U40324 (N_40324,N_39908,N_39707);
nand U40325 (N_40325,N_38631,N_37941);
or U40326 (N_40326,N_39873,N_37317);
and U40327 (N_40327,N_38753,N_39665);
or U40328 (N_40328,N_39384,N_36078);
and U40329 (N_40329,N_38125,N_38324);
nand U40330 (N_40330,N_39213,N_36875);
nand U40331 (N_40331,N_36948,N_37819);
or U40332 (N_40332,N_37935,N_37621);
xor U40333 (N_40333,N_37997,N_36755);
nand U40334 (N_40334,N_38690,N_35708);
nor U40335 (N_40335,N_36126,N_35692);
nor U40336 (N_40336,N_35270,N_35398);
and U40337 (N_40337,N_38820,N_39793);
or U40338 (N_40338,N_39332,N_35624);
xor U40339 (N_40339,N_35667,N_36158);
nor U40340 (N_40340,N_39660,N_36470);
nor U40341 (N_40341,N_39710,N_39795);
nor U40342 (N_40342,N_37860,N_37294);
nor U40343 (N_40343,N_39279,N_38422);
and U40344 (N_40344,N_36004,N_36541);
and U40345 (N_40345,N_38402,N_39367);
nor U40346 (N_40346,N_38207,N_36701);
nor U40347 (N_40347,N_35836,N_35285);
nand U40348 (N_40348,N_37415,N_36864);
or U40349 (N_40349,N_37994,N_35657);
xor U40350 (N_40350,N_38419,N_35693);
or U40351 (N_40351,N_39714,N_35754);
or U40352 (N_40352,N_35241,N_36749);
and U40353 (N_40353,N_36728,N_37658);
nand U40354 (N_40354,N_36143,N_36246);
or U40355 (N_40355,N_38134,N_38713);
or U40356 (N_40356,N_38367,N_35132);
nor U40357 (N_40357,N_35748,N_37775);
or U40358 (N_40358,N_38722,N_37773);
nand U40359 (N_40359,N_36259,N_38550);
and U40360 (N_40360,N_37910,N_38257);
xor U40361 (N_40361,N_36565,N_35320);
nand U40362 (N_40362,N_38491,N_39087);
xnor U40363 (N_40363,N_39293,N_38177);
nand U40364 (N_40364,N_36711,N_37255);
xnor U40365 (N_40365,N_35190,N_37420);
nand U40366 (N_40366,N_39153,N_37338);
and U40367 (N_40367,N_36642,N_39488);
or U40368 (N_40368,N_36908,N_35866);
nand U40369 (N_40369,N_38489,N_37473);
or U40370 (N_40370,N_37979,N_39312);
nand U40371 (N_40371,N_37578,N_35627);
xor U40372 (N_40372,N_37408,N_35206);
nand U40373 (N_40373,N_35871,N_35961);
and U40374 (N_40374,N_39257,N_36649);
nand U40375 (N_40375,N_36230,N_35047);
nand U40376 (N_40376,N_37793,N_38844);
nor U40377 (N_40377,N_38159,N_39028);
nand U40378 (N_40378,N_35053,N_37618);
nor U40379 (N_40379,N_36216,N_36671);
and U40380 (N_40380,N_35074,N_37323);
and U40381 (N_40381,N_36248,N_36019);
or U40382 (N_40382,N_37158,N_36217);
nor U40383 (N_40383,N_35162,N_36687);
nand U40384 (N_40384,N_36872,N_36115);
and U40385 (N_40385,N_39006,N_35300);
nand U40386 (N_40386,N_37781,N_39383);
and U40387 (N_40387,N_36033,N_36584);
nand U40388 (N_40388,N_37510,N_38677);
nor U40389 (N_40389,N_35019,N_37206);
and U40390 (N_40390,N_37080,N_38866);
nand U40391 (N_40391,N_38771,N_39378);
nor U40392 (N_40392,N_39227,N_35865);
or U40393 (N_40393,N_38651,N_36531);
and U40394 (N_40394,N_35457,N_35944);
nor U40395 (N_40395,N_35064,N_39032);
xnor U40396 (N_40396,N_36708,N_39179);
nor U40397 (N_40397,N_37901,N_38607);
or U40398 (N_40398,N_36330,N_37813);
and U40399 (N_40399,N_36844,N_35146);
nand U40400 (N_40400,N_37490,N_38369);
nand U40401 (N_40401,N_39258,N_38436);
nor U40402 (N_40402,N_38358,N_38227);
nand U40403 (N_40403,N_38671,N_35738);
xor U40404 (N_40404,N_39532,N_36183);
and U40405 (N_40405,N_37009,N_37529);
or U40406 (N_40406,N_38214,N_37429);
and U40407 (N_40407,N_36360,N_39120);
or U40408 (N_40408,N_36830,N_38482);
nand U40409 (N_40409,N_37502,N_35213);
or U40410 (N_40410,N_37282,N_38633);
nor U40411 (N_40411,N_35376,N_39496);
nor U40412 (N_40412,N_36938,N_38961);
or U40413 (N_40413,N_35007,N_35168);
nand U40414 (N_40414,N_39628,N_36466);
nand U40415 (N_40415,N_38323,N_36795);
xor U40416 (N_40416,N_38089,N_36737);
nor U40417 (N_40417,N_36363,N_35825);
nor U40418 (N_40418,N_38120,N_39489);
and U40419 (N_40419,N_38907,N_39746);
nor U40420 (N_40420,N_39909,N_37524);
or U40421 (N_40421,N_38988,N_39566);
xor U40422 (N_40422,N_35385,N_36450);
and U40423 (N_40423,N_37458,N_35401);
xor U40424 (N_40424,N_35864,N_36385);
xor U40425 (N_40425,N_35048,N_38780);
or U40426 (N_40426,N_36763,N_39468);
nor U40427 (N_40427,N_38206,N_37648);
nor U40428 (N_40428,N_39871,N_35311);
and U40429 (N_40429,N_35027,N_35930);
nand U40430 (N_40430,N_37689,N_37832);
xnor U40431 (N_40431,N_36674,N_38709);
nand U40432 (N_40432,N_38283,N_39804);
nor U40433 (N_40433,N_37126,N_37435);
nor U40434 (N_40434,N_37764,N_39423);
and U40435 (N_40435,N_35516,N_36215);
and U40436 (N_40436,N_35230,N_35680);
xnor U40437 (N_40437,N_37918,N_39303);
nor U40438 (N_40438,N_36018,N_38440);
xnor U40439 (N_40439,N_39289,N_36189);
or U40440 (N_40440,N_37761,N_37797);
xor U40441 (N_40441,N_35594,N_38437);
xor U40442 (N_40442,N_35449,N_38355);
or U40443 (N_40443,N_39122,N_38719);
nor U40444 (N_40444,N_36598,N_38522);
or U40445 (N_40445,N_38582,N_38546);
xor U40446 (N_40446,N_37824,N_37247);
or U40447 (N_40447,N_37851,N_37978);
and U40448 (N_40448,N_37018,N_37224);
nor U40449 (N_40449,N_35964,N_38030);
and U40450 (N_40450,N_36244,N_39669);
xnor U40451 (N_40451,N_35088,N_39237);
nor U40452 (N_40452,N_37252,N_38480);
and U40453 (N_40453,N_36847,N_36118);
nand U40454 (N_40454,N_38790,N_37363);
nand U40455 (N_40455,N_38906,N_39898);
or U40456 (N_40456,N_37566,N_37607);
and U40457 (N_40457,N_38542,N_39251);
xor U40458 (N_40458,N_38106,N_39177);
or U40459 (N_40459,N_37059,N_37827);
xor U40460 (N_40460,N_39777,N_35322);
xnor U40461 (N_40461,N_35069,N_37343);
or U40462 (N_40462,N_37816,N_39529);
and U40463 (N_40463,N_37659,N_35600);
nor U40464 (N_40464,N_36342,N_37242);
nand U40465 (N_40465,N_37414,N_37493);
or U40466 (N_40466,N_39583,N_37057);
nor U40467 (N_40467,N_39542,N_36076);
nor U40468 (N_40468,N_38104,N_39751);
nor U40469 (N_40469,N_38832,N_37744);
xnor U40470 (N_40470,N_36310,N_39049);
nor U40471 (N_40471,N_36754,N_38225);
xor U40472 (N_40472,N_35797,N_36857);
or U40473 (N_40473,N_37877,N_35784);
xnor U40474 (N_40474,N_36712,N_36267);
xor U40475 (N_40475,N_37307,N_36374);
xnor U40476 (N_40476,N_39050,N_35794);
and U40477 (N_40477,N_36756,N_39452);
or U40478 (N_40478,N_35878,N_35147);
nor U40479 (N_40479,N_39620,N_35595);
or U40480 (N_40480,N_39222,N_38621);
nand U40481 (N_40481,N_39882,N_38414);
and U40482 (N_40482,N_38833,N_39031);
nand U40483 (N_40483,N_39510,N_37019);
or U40484 (N_40484,N_39965,N_37078);
or U40485 (N_40485,N_37482,N_37908);
nor U40486 (N_40486,N_35161,N_39412);
and U40487 (N_40487,N_36130,N_36566);
and U40488 (N_40488,N_38558,N_39762);
or U40489 (N_40489,N_39411,N_38317);
and U40490 (N_40490,N_38505,N_38730);
nand U40491 (N_40491,N_35525,N_39044);
nand U40492 (N_40492,N_39568,N_39826);
nor U40493 (N_40493,N_35887,N_39420);
and U40494 (N_40494,N_36357,N_35091);
nor U40495 (N_40495,N_37801,N_37283);
or U40496 (N_40496,N_39561,N_37963);
or U40497 (N_40497,N_38220,N_38392);
nand U40498 (N_40498,N_35782,N_37846);
nor U40499 (N_40499,N_37512,N_39348);
xnor U40500 (N_40500,N_38696,N_38005);
nand U40501 (N_40501,N_35834,N_36831);
and U40502 (N_40502,N_39992,N_35446);
or U40503 (N_40503,N_37037,N_38969);
xor U40504 (N_40504,N_38973,N_38312);
and U40505 (N_40505,N_38597,N_37417);
or U40506 (N_40506,N_38586,N_36124);
nor U40507 (N_40507,N_38132,N_36232);
nand U40508 (N_40508,N_35547,N_38019);
and U40509 (N_40509,N_39525,N_36770);
or U40510 (N_40510,N_36905,N_35353);
nor U40511 (N_40511,N_38737,N_35638);
nor U40512 (N_40512,N_38359,N_39663);
and U40513 (N_40513,N_35406,N_37656);
xor U40514 (N_40514,N_39947,N_35092);
nor U40515 (N_40515,N_37913,N_36178);
xnor U40516 (N_40516,N_39076,N_39308);
and U40517 (N_40517,N_38612,N_35399);
or U40518 (N_40518,N_38399,N_36528);
nand U40519 (N_40519,N_36937,N_35099);
or U40520 (N_40520,N_35095,N_36395);
nor U40521 (N_40521,N_37944,N_35275);
and U40522 (N_40522,N_39521,N_37527);
or U40523 (N_40523,N_36418,N_36054);
xor U40524 (N_40524,N_38604,N_37005);
and U40525 (N_40525,N_38088,N_38231);
nand U40526 (N_40526,N_37866,N_35442);
nor U40527 (N_40527,N_36522,N_38090);
and U40528 (N_40528,N_38348,N_39870);
and U40529 (N_40529,N_35766,N_38767);
nor U40530 (N_40530,N_35454,N_39256);
xnor U40531 (N_40531,N_37384,N_36404);
and U40532 (N_40532,N_39573,N_37066);
or U40533 (N_40533,N_35191,N_37842);
nand U40534 (N_40534,N_37820,N_36529);
and U40535 (N_40535,N_36002,N_35798);
nor U40536 (N_40536,N_35393,N_38735);
or U40537 (N_40537,N_38540,N_39290);
nand U40538 (N_40538,N_39033,N_39535);
and U40539 (N_40539,N_38935,N_37151);
nand U40540 (N_40540,N_38998,N_37806);
or U40541 (N_40541,N_36073,N_38007);
nor U40542 (N_40542,N_36362,N_39443);
nand U40543 (N_40543,N_39618,N_35131);
and U40544 (N_40544,N_36287,N_39381);
xor U40545 (N_40545,N_38112,N_37287);
and U40546 (N_40546,N_38253,N_37156);
or U40547 (N_40547,N_39495,N_35492);
nand U40548 (N_40548,N_39847,N_38235);
nor U40549 (N_40549,N_38157,N_35653);
or U40550 (N_40550,N_39438,N_35892);
nand U40551 (N_40551,N_36865,N_36526);
nor U40552 (N_40552,N_36402,N_39531);
xnor U40553 (N_40553,N_36695,N_39456);
nand U40554 (N_40554,N_36798,N_39522);
nand U40555 (N_40555,N_37555,N_35493);
nor U40556 (N_40556,N_37579,N_36100);
xor U40557 (N_40557,N_37198,N_38403);
and U40558 (N_40558,N_39785,N_36633);
nor U40559 (N_40559,N_35316,N_37146);
xor U40560 (N_40560,N_36944,N_36366);
xnor U40561 (N_40561,N_36999,N_37559);
xnor U40562 (N_40562,N_35447,N_35546);
and U40563 (N_40563,N_39765,N_37776);
xnor U40564 (N_40564,N_37237,N_38587);
nand U40565 (N_40565,N_35665,N_38830);
or U40566 (N_40566,N_36394,N_36736);
and U40567 (N_40567,N_39238,N_36449);
nand U40568 (N_40568,N_38778,N_38171);
xor U40569 (N_40569,N_36303,N_39074);
or U40570 (N_40570,N_38271,N_39702);
and U40571 (N_40571,N_37116,N_36778);
and U40572 (N_40572,N_35137,N_38433);
nand U40573 (N_40573,N_35207,N_38775);
or U40574 (N_40574,N_37903,N_38567);
nor U40575 (N_40575,N_35862,N_39963);
or U40576 (N_40576,N_38533,N_35332);
nand U40577 (N_40577,N_39173,N_36973);
xnor U40578 (N_40578,N_38860,N_37181);
nor U40579 (N_40579,N_35931,N_36894);
or U40580 (N_40580,N_36866,N_38615);
and U40581 (N_40581,N_37448,N_36167);
or U40582 (N_40582,N_37028,N_36924);
nor U40583 (N_40583,N_35461,N_37542);
nor U40584 (N_40584,N_37678,N_35257);
xnor U40585 (N_40585,N_37577,N_37909);
xnor U40586 (N_40586,N_38476,N_36208);
and U40587 (N_40587,N_37251,N_38275);
and U40588 (N_40588,N_37289,N_37128);
xnor U40589 (N_40589,N_38927,N_38878);
and U40590 (N_40590,N_37389,N_35576);
and U40591 (N_40591,N_38212,N_38708);
xor U40592 (N_40592,N_37393,N_36535);
nand U40593 (N_40593,N_35816,N_39371);
and U40594 (N_40594,N_38733,N_36213);
xnor U40595 (N_40595,N_39638,N_35482);
nand U40596 (N_40596,N_37603,N_38955);
or U40597 (N_40597,N_39763,N_38451);
or U40598 (N_40598,N_39099,N_36490);
xor U40599 (N_40599,N_37699,N_36192);
nand U40600 (N_40600,N_39422,N_38219);
nor U40601 (N_40601,N_36651,N_38189);
and U40602 (N_40602,N_35395,N_37324);
xnor U40603 (N_40603,N_39723,N_35829);
xnor U40604 (N_40604,N_39230,N_35083);
nor U40605 (N_40605,N_39788,N_36631);
and U40606 (N_40606,N_39140,N_35676);
nand U40607 (N_40607,N_37902,N_36028);
nor U40608 (N_40608,N_35713,N_38700);
nor U40609 (N_40609,N_38751,N_38520);
or U40610 (N_40610,N_38325,N_36281);
and U40611 (N_40611,N_36053,N_38811);
or U40612 (N_40612,N_35992,N_35502);
nor U40613 (N_40613,N_38001,N_38952);
or U40614 (N_40614,N_35345,N_39548);
and U40615 (N_40615,N_38881,N_39917);
xnor U40616 (N_40616,N_35475,N_38456);
xnor U40617 (N_40617,N_36485,N_37352);
nand U40618 (N_40618,N_39154,N_37779);
nor U40619 (N_40619,N_36840,N_36442);
and U40620 (N_40620,N_37157,N_35818);
xor U40621 (N_40621,N_37867,N_39113);
and U40622 (N_40622,N_37485,N_36391);
xnor U40623 (N_40623,N_36794,N_37588);
nor U40624 (N_40624,N_38181,N_38506);
and U40625 (N_40625,N_36181,N_38366);
nor U40626 (N_40626,N_37783,N_39061);
and U40627 (N_40627,N_37366,N_38626);
and U40628 (N_40628,N_38105,N_37682);
or U40629 (N_40629,N_37563,N_39872);
or U40630 (N_40630,N_39641,N_38184);
xnor U40631 (N_40631,N_36623,N_38327);
and U40632 (N_40632,N_35384,N_37166);
and U40633 (N_40633,N_36017,N_35698);
and U40634 (N_40634,N_36797,N_36606);
xor U40635 (N_40635,N_38930,N_38503);
and U40636 (N_40636,N_38536,N_36684);
and U40637 (N_40637,N_36235,N_39267);
nor U40638 (N_40638,N_37494,N_36051);
xnor U40639 (N_40639,N_35211,N_39160);
and U40640 (N_40640,N_35874,N_35276);
nor U40641 (N_40641,N_35622,N_39803);
nand U40642 (N_40642,N_39739,N_36064);
and U40643 (N_40643,N_35247,N_35443);
xnor U40644 (N_40644,N_39855,N_38345);
nand U40645 (N_40645,N_37210,N_38752);
xnor U40646 (N_40646,N_35799,N_39191);
or U40647 (N_40647,N_35476,N_39119);
xor U40648 (N_40648,N_36947,N_39060);
nor U40649 (N_40649,N_38384,N_36473);
nand U40650 (N_40650,N_38371,N_35605);
nor U40651 (N_40651,N_38233,N_35833);
nor U40652 (N_40652,N_38123,N_39945);
or U40653 (N_40653,N_38823,N_36863);
or U40654 (N_40654,N_39818,N_35543);
xor U40655 (N_40655,N_36276,N_39171);
or U40656 (N_40656,N_36397,N_38873);
xnor U40657 (N_40657,N_36656,N_36087);
or U40658 (N_40658,N_36874,N_35341);
or U40659 (N_40659,N_36889,N_38269);
nor U40660 (N_40660,N_37186,N_35634);
xor U40661 (N_40661,N_38316,N_37180);
and U40662 (N_40662,N_35339,N_38848);
and U40663 (N_40663,N_37791,N_39999);
nand U40664 (N_40664,N_35540,N_36453);
and U40665 (N_40665,N_38710,N_37489);
or U40666 (N_40666,N_36162,N_36159);
and U40667 (N_40667,N_36586,N_39436);
xor U40668 (N_40668,N_37890,N_39833);
nand U40669 (N_40669,N_36061,N_35237);
or U40670 (N_40670,N_37207,N_35768);
xor U40671 (N_40671,N_38102,N_39013);
xor U40672 (N_40672,N_38056,N_38499);
xnor U40673 (N_40673,N_36461,N_38658);
xnor U40674 (N_40674,N_35648,N_37161);
nand U40675 (N_40675,N_35846,N_36882);
nor U40676 (N_40676,N_37912,N_36271);
nor U40677 (N_40677,N_37812,N_36039);
nor U40678 (N_40678,N_36931,N_37507);
or U40679 (N_40679,N_36092,N_38545);
nand U40680 (N_40680,N_39019,N_37506);
xnor U40681 (N_40681,N_38295,N_39625);
nand U40682 (N_40682,N_37177,N_38268);
and U40683 (N_40683,N_37639,N_39695);
nor U40684 (N_40684,N_36354,N_35392);
xor U40685 (N_40685,N_39502,N_37117);
and U40686 (N_40686,N_39484,N_37068);
or U40687 (N_40687,N_37665,N_37476);
or U40688 (N_40688,N_36608,N_35185);
or U40689 (N_40689,N_36558,N_35283);
or U40690 (N_40690,N_35608,N_35119);
xnor U40691 (N_40691,N_39431,N_39182);
xnor U40692 (N_40692,N_39515,N_36454);
xor U40693 (N_40693,N_37119,N_38024);
and U40694 (N_40694,N_37582,N_36827);
or U40695 (N_40695,N_38498,N_37122);
xnor U40696 (N_40696,N_39454,N_37543);
nand U40697 (N_40697,N_35483,N_37660);
xor U40698 (N_40698,N_36997,N_37149);
nand U40699 (N_40699,N_38576,N_38783);
xnor U40700 (N_40700,N_38638,N_38819);
and U40701 (N_40701,N_35941,N_36249);
and U40702 (N_40702,N_35448,N_35329);
or U40703 (N_40703,N_37246,N_37723);
and U40704 (N_40704,N_37432,N_37953);
and U40705 (N_40705,N_39414,N_39572);
or U40706 (N_40706,N_36321,N_36349);
nor U40707 (N_40707,N_38261,N_36329);
and U40708 (N_40708,N_37202,N_35050);
xor U40709 (N_40709,N_36438,N_36811);
or U40710 (N_40710,N_39147,N_38762);
and U40711 (N_40711,N_39942,N_36383);
or U40712 (N_40712,N_39517,N_36343);
nor U40713 (N_40713,N_36982,N_38085);
or U40714 (N_40714,N_36479,N_36146);
and U40715 (N_40715,N_35330,N_36518);
nor U40716 (N_40716,N_36851,N_38086);
or U40717 (N_40717,N_39220,N_35494);
or U40718 (N_40718,N_38304,N_39385);
and U40719 (N_40719,N_38846,N_35984);
nand U40720 (N_40720,N_35861,N_38388);
or U40721 (N_40721,N_38281,N_35066);
or U40722 (N_40722,N_36822,N_38068);
nand U40723 (N_40723,N_35830,N_39178);
nor U40724 (N_40724,N_37411,N_39218);
xnor U40725 (N_40725,N_38192,N_35682);
and U40726 (N_40726,N_37143,N_37782);
nor U40727 (N_40727,N_38298,N_38251);
and U40728 (N_40728,N_39287,N_38624);
and U40729 (N_40729,N_37032,N_37848);
or U40730 (N_40730,N_38869,N_36488);
xor U40731 (N_40731,N_38318,N_37347);
nand U40732 (N_40732,N_36483,N_35801);
or U40733 (N_40733,N_37349,N_38018);
and U40734 (N_40734,N_39810,N_35102);
nor U40735 (N_40735,N_38850,N_35254);
nor U40736 (N_40736,N_39860,N_36946);
nand U40737 (N_40737,N_37222,N_35173);
nand U40738 (N_40738,N_37693,N_39577);
nand U40739 (N_40739,N_38948,N_36401);
xor U40740 (N_40740,N_37991,N_38645);
nand U40741 (N_40741,N_39207,N_37628);
xor U40742 (N_40742,N_38072,N_38311);
or U40743 (N_40743,N_35416,N_39605);
nor U40744 (N_40744,N_36992,N_39235);
or U40745 (N_40745,N_39886,N_36621);
or U40746 (N_40746,N_38113,N_39086);
nor U40747 (N_40747,N_36144,N_37974);
nand U40748 (N_40748,N_39897,N_38578);
and U40749 (N_40749,N_35686,N_38297);
nor U40750 (N_40750,N_38029,N_35827);
or U40751 (N_40751,N_38040,N_35891);
and U40752 (N_40752,N_38217,N_38246);
nor U40753 (N_40753,N_37045,N_35868);
xnor U40754 (N_40754,N_37063,N_38652);
or U40755 (N_40755,N_35263,N_36081);
and U40756 (N_40756,N_38902,N_37481);
xnor U40757 (N_40757,N_36266,N_35923);
nor U40758 (N_40758,N_35497,N_39878);
xnor U40759 (N_40759,N_35025,N_39453);
or U40760 (N_40760,N_36057,N_35256);
and U40761 (N_40761,N_39215,N_37929);
and U40762 (N_40762,N_38041,N_38372);
or U40763 (N_40763,N_38452,N_36151);
or U40764 (N_40764,N_36952,N_35412);
xnor U40765 (N_40765,N_39666,N_39552);
and U40766 (N_40766,N_35077,N_38909);
and U40767 (N_40767,N_39075,N_36145);
nor U40768 (N_40768,N_37219,N_37035);
xnor U40769 (N_40769,N_37139,N_38648);
nand U40770 (N_40770,N_36302,N_35070);
xor U40771 (N_40771,N_38055,N_35135);
xnor U40772 (N_40772,N_39151,N_39784);
and U40773 (N_40773,N_36691,N_37558);
nor U40774 (N_40774,N_36876,N_37710);
and U40775 (N_40775,N_39474,N_35116);
xnor U40776 (N_40776,N_35977,N_38643);
and U40777 (N_40777,N_39701,N_35924);
nand U40778 (N_40778,N_37599,N_38434);
nand U40779 (N_40779,N_37030,N_36492);
or U40780 (N_40780,N_35539,N_39355);
or U40781 (N_40781,N_38827,N_39252);
nor U40782 (N_40782,N_35572,N_35551);
or U40783 (N_40783,N_37966,N_36696);
nor U40784 (N_40784,N_35603,N_38997);
or U40785 (N_40785,N_37600,N_37445);
and U40786 (N_40786,N_39768,N_37280);
or U40787 (N_40787,N_35040,N_38014);
nand U40788 (N_40788,N_39421,N_36921);
and U40789 (N_40789,N_37985,N_35879);
nor U40790 (N_40790,N_38695,N_35728);
and U40791 (N_40791,N_38890,N_37661);
and U40792 (N_40792,N_35022,N_36983);
xnor U40793 (N_40793,N_37551,N_38552);
and U40794 (N_40794,N_38279,N_39816);
xnor U40795 (N_40795,N_36389,N_35265);
or U40796 (N_40796,N_36368,N_36682);
xnor U40797 (N_40797,N_39645,N_37350);
or U40798 (N_40798,N_38413,N_38013);
or U40799 (N_40799,N_35441,N_39458);
xnor U40800 (N_40800,N_35560,N_39596);
nand U40801 (N_40801,N_37085,N_37229);
nand U40802 (N_40802,N_35940,N_37051);
or U40803 (N_40803,N_37742,N_37232);
nand U40804 (N_40804,N_35732,N_38842);
nor U40805 (N_40805,N_37719,N_36622);
nand U40806 (N_40806,N_39072,N_37919);
nor U40807 (N_40807,N_35394,N_38789);
or U40808 (N_40808,N_35342,N_36241);
and U40809 (N_40809,N_35200,N_37967);
xor U40810 (N_40810,N_35552,N_39864);
or U40811 (N_40811,N_39386,N_36585);
xnor U40812 (N_40812,N_37946,N_37034);
or U40813 (N_40813,N_36673,N_35375);
nor U40814 (N_40814,N_38874,N_39311);
xnor U40815 (N_40815,N_35419,N_37048);
nor U40816 (N_40816,N_38687,N_36253);
and U40817 (N_40817,N_39111,N_39792);
nor U40818 (N_40818,N_38673,N_36290);
nor U40819 (N_40819,N_36429,N_36419);
nor U40820 (N_40820,N_37740,N_39144);
xor U40821 (N_40821,N_39123,N_36125);
and U40822 (N_40822,N_37036,N_36913);
nand U40823 (N_40823,N_38933,N_38320);
or U40824 (N_40824,N_38263,N_39372);
xnor U40825 (N_40825,N_38101,N_35463);
xnor U40826 (N_40826,N_38728,N_37316);
or U40827 (N_40827,N_35352,N_36035);
nand U40828 (N_40828,N_37855,N_36113);
xnor U40829 (N_40829,N_35437,N_35100);
nand U40830 (N_40830,N_38559,N_38944);
and U40831 (N_40831,N_39313,N_35520);
and U40832 (N_40832,N_39744,N_35509);
and U40833 (N_40833,N_35507,N_36678);
and U40834 (N_40834,N_39936,N_35541);
nor U40835 (N_40835,N_39967,N_38524);
nand U40836 (N_40836,N_35273,N_39194);
nor U40837 (N_40837,N_38036,N_35029);
or U40838 (N_40838,N_37584,N_38668);
xor U40839 (N_40839,N_35431,N_37278);
xor U40840 (N_40840,N_39685,N_38078);
nor U40841 (N_40841,N_35989,N_39592);
nand U40842 (N_40842,N_38158,N_37340);
or U40843 (N_40843,N_39874,N_35718);
and U40844 (N_40844,N_39268,N_35472);
nor U40845 (N_40845,N_39696,N_38764);
and U40846 (N_40846,N_37619,N_39709);
or U40847 (N_40847,N_38802,N_36298);
and U40848 (N_40848,N_36236,N_36532);
or U40849 (N_40849,N_37205,N_35488);
nor U40850 (N_40850,N_37521,N_39642);
and U40851 (N_40851,N_38156,N_36133);
and U40852 (N_40852,N_35272,N_36779);
nand U40853 (N_40853,N_39341,N_38815);
xnor U40854 (N_40854,N_36353,N_39354);
or U40855 (N_40855,N_39973,N_35959);
nor U40856 (N_40856,N_35260,N_39170);
and U40857 (N_40857,N_36487,N_38202);
and U40858 (N_40858,N_35410,N_36068);
or U40859 (N_40859,N_39426,N_38501);
and U40860 (N_40860,N_36853,N_37859);
xnor U40861 (N_40861,N_35997,N_35647);
nand U40862 (N_40862,N_37572,N_36074);
and U40863 (N_40863,N_37311,N_35152);
or U40864 (N_40864,N_37642,N_36976);
or U40865 (N_40865,N_38531,N_39736);
nand U40866 (N_40866,N_37253,N_37936);
and U40867 (N_40867,N_38583,N_35635);
and U40868 (N_40868,N_39733,N_37112);
nand U40869 (N_40869,N_38682,N_37168);
nand U40870 (N_40870,N_39083,N_39769);
or U40871 (N_40871,N_35039,N_39865);
nor U40872 (N_40872,N_38743,N_36361);
or U40873 (N_40873,N_38630,N_39174);
or U40874 (N_40874,N_35208,N_37322);
or U40875 (N_40875,N_35783,N_36059);
or U40876 (N_40876,N_38809,N_35240);
xor U40877 (N_40877,N_35683,N_35972);
and U40878 (N_40878,N_36603,N_37227);
xnor U40879 (N_40879,N_39646,N_39619);
and U40880 (N_40880,N_37681,N_37011);
nand U40881 (N_40881,N_38847,N_35532);
and U40882 (N_40882,N_36933,N_36037);
or U40883 (N_40883,N_39741,N_37200);
nor U40884 (N_40884,N_37787,N_35242);
or U40885 (N_40885,N_39637,N_38377);
or U40886 (N_40886,N_38879,N_36709);
nor U40887 (N_40887,N_37594,N_37442);
xnor U40888 (N_40888,N_37353,N_35370);
xor U40889 (N_40889,N_38195,N_36317);
nor U40890 (N_40890,N_37213,N_35904);
nor U40891 (N_40891,N_37277,N_39370);
nand U40892 (N_40892,N_37014,N_38731);
or U40893 (N_40893,N_36817,N_37614);
xnor U40894 (N_40894,N_38341,N_38444);
xor U40895 (N_40895,N_35504,N_39229);
nor U40896 (N_40896,N_35480,N_36917);
and U40897 (N_40897,N_35607,N_37131);
or U40898 (N_40898,N_39518,N_38798);
nand U40899 (N_40899,N_36925,N_38592);
nand U40900 (N_40900,N_35435,N_37020);
or U40901 (N_40901,N_39407,N_35633);
nor U40902 (N_40902,N_37197,N_38130);
and U40903 (N_40903,N_35623,N_39970);
nand U40904 (N_40904,N_35710,N_36781);
xor U40905 (N_40905,N_39305,N_38114);
nand U40906 (N_40906,N_37999,N_35354);
nor U40907 (N_40907,N_39562,N_38589);
nand U40908 (N_40908,N_36325,N_36338);
or U40909 (N_40909,N_38813,N_38313);
nor U40910 (N_40910,N_39224,N_38834);
nand U40911 (N_40911,N_36657,N_37836);
and U40912 (N_40912,N_39939,N_37367);
xnor U40913 (N_40913,N_38435,N_38934);
xnor U40914 (N_40914,N_36273,N_35599);
or U40915 (N_40915,N_36637,N_35305);
nor U40916 (N_40916,N_39840,N_36523);
and U40917 (N_40917,N_39233,N_35045);
nor U40918 (N_40918,N_38861,N_35156);
and U40919 (N_40919,N_38603,N_37441);
xor U40920 (N_40920,N_39545,N_37630);
nor U40921 (N_40921,N_36681,N_39584);
xnor U40922 (N_40922,N_37416,N_38987);
nor U40923 (N_40923,N_35231,N_35117);
and U40924 (N_40924,N_36358,N_39404);
xor U40925 (N_40925,N_39771,N_36837);
and U40926 (N_40926,N_39697,N_35267);
xnor U40927 (N_40927,N_37123,N_39767);
xor U40928 (N_40928,N_37633,N_38203);
xnor U40929 (N_40929,N_36519,N_35893);
xor U40930 (N_40930,N_37286,N_39106);
nor U40931 (N_40931,N_36318,N_35003);
and U40932 (N_40932,N_38618,N_35644);
and U40933 (N_40933,N_36545,N_36356);
xnor U40934 (N_40934,N_37142,N_36502);
and U40935 (N_40935,N_38840,N_36510);
and U40936 (N_40936,N_39921,N_36557);
or U40937 (N_40937,N_38438,N_38459);
xor U40938 (N_40938,N_35697,N_37337);
nor U40939 (N_40939,N_39121,N_36289);
nand U40940 (N_40940,N_37907,N_38598);
or U40941 (N_40941,N_35072,N_38685);
nand U40942 (N_40942,N_38996,N_39589);
nand U40943 (N_40943,N_37986,N_38563);
nor U40944 (N_40944,N_36350,N_39169);
and U40945 (N_40945,N_37585,N_36579);
xor U40946 (N_40946,N_35826,N_38774);
or U40947 (N_40947,N_37690,N_38950);
xnor U40948 (N_40948,N_38074,N_37136);
and U40949 (N_40949,N_36137,N_36620);
nand U40950 (N_40950,N_37427,N_36420);
or U40951 (N_40951,N_35970,N_36928);
or U40952 (N_40952,N_39806,N_35872);
xnor U40953 (N_40953,N_35912,N_36883);
or U40954 (N_40954,N_36850,N_37118);
or U40955 (N_40955,N_39098,N_37105);
or U40956 (N_40956,N_37932,N_37882);
nor U40957 (N_40957,N_38493,N_37586);
nor U40958 (N_40958,N_39928,N_35456);
nand U40959 (N_40959,N_38839,N_37410);
or U40960 (N_40960,N_38502,N_39925);
and U40961 (N_40961,N_37576,N_37916);
nand U40962 (N_40962,N_36277,N_38469);
xnor U40963 (N_40963,N_37407,N_39112);
nand U40964 (N_40964,N_35121,N_35439);
nor U40965 (N_40965,N_38519,N_36826);
nand U40966 (N_40966,N_35980,N_39018);
or U40967 (N_40967,N_37221,N_36929);
nor U40968 (N_40968,N_39884,N_35719);
and U40969 (N_40969,N_36959,N_35123);
nor U40970 (N_40970,N_39546,N_36203);
nand U40971 (N_40971,N_39394,N_36871);
nor U40972 (N_40972,N_39116,N_39479);
nand U40973 (N_40973,N_39219,N_37115);
or U40974 (N_40974,N_38859,N_36854);
nor U40975 (N_40975,N_39990,N_35564);
or U40976 (N_40976,N_38315,N_36626);
or U40977 (N_40977,N_36632,N_38960);
and U40978 (N_40978,N_38262,N_39001);
xnor U40979 (N_40979,N_37664,N_39760);
nor U40980 (N_40980,N_36969,N_37310);
xor U40981 (N_40981,N_37024,N_35373);
and U40982 (N_40982,N_39232,N_35453);
or U40983 (N_40983,N_39787,N_39388);
or U40984 (N_40984,N_37754,N_35744);
and U40985 (N_40985,N_38115,N_38966);
or U40986 (N_40986,N_36556,N_38882);
nor U40987 (N_40987,N_35244,N_39540);
and U40988 (N_40988,N_35832,N_37325);
and U40989 (N_40989,N_37258,N_36263);
nand U40990 (N_40990,N_38071,N_37400);
and U40991 (N_40991,N_38479,N_37082);
nor U40992 (N_40992,N_36109,N_39166);
or U40993 (N_40993,N_38154,N_35655);
nor U40994 (N_40994,N_38486,N_38801);
and U40995 (N_40995,N_37137,N_37515);
and U40996 (N_40996,N_38198,N_36710);
nand U40997 (N_40997,N_37508,N_39581);
xor U40998 (N_40998,N_36010,N_38145);
xnor U40999 (N_40999,N_39318,N_37313);
or U41000 (N_41000,N_37269,N_35023);
or U41001 (N_41001,N_39491,N_37823);
xnor U41002 (N_41002,N_39636,N_39379);
nand U41003 (N_41003,N_37150,N_36141);
and U41004 (N_41004,N_37841,N_38032);
and U41005 (N_41005,N_35885,N_36769);
nand U41006 (N_41006,N_39687,N_39226);
nand U41007 (N_41007,N_36740,N_38701);
xor U41008 (N_41008,N_36825,N_39593);
or U41009 (N_41009,N_39070,N_39052);
nand U41010 (N_41010,N_35301,N_39960);
nand U41011 (N_41011,N_38180,N_37184);
xor U41012 (N_41012,N_35288,N_35772);
nand U41013 (N_41013,N_39325,N_38704);
and U41014 (N_41014,N_38373,N_38849);
or U41015 (N_41015,N_35712,N_36706);
nor U41016 (N_41016,N_39731,N_35994);
and U41017 (N_41017,N_39603,N_35170);
xor U41018 (N_41018,N_38947,N_35142);
and U41019 (N_41019,N_35884,N_36806);
and U41020 (N_41020,N_39449,N_36194);
or U41021 (N_41021,N_35172,N_36347);
or U41022 (N_41022,N_36083,N_35245);
nand U41023 (N_41023,N_36199,N_38922);
nand U41024 (N_41024,N_38678,N_36352);
xnor U41025 (N_41025,N_37795,N_37488);
and U41026 (N_41026,N_37993,N_36291);
and U41027 (N_41027,N_35182,N_38570);
nor U41028 (N_41028,N_38339,N_36998);
and U41029 (N_41029,N_35335,N_36834);
or U41030 (N_41030,N_39146,N_37694);
or U41031 (N_41031,N_38962,N_36451);
and U41032 (N_41032,N_35451,N_39208);
nand U41033 (N_41033,N_38245,N_37569);
nor U41034 (N_41034,N_36893,N_35280);
nand U41035 (N_41035,N_35236,N_35255);
or U41036 (N_41036,N_39248,N_38957);
xor U41037 (N_41037,N_38867,N_38928);
nand U41038 (N_41038,N_39398,N_36247);
nand U41039 (N_41039,N_37728,N_37091);
nand U41040 (N_41040,N_36177,N_36675);
xor U41041 (N_41041,N_36890,N_38699);
xnor U41042 (N_41042,N_37676,N_37739);
or U41043 (N_41043,N_39048,N_35512);
xor U41044 (N_41044,N_36371,N_36856);
or U41045 (N_41045,N_36772,N_38361);
and U41046 (N_41046,N_35960,N_39894);
and U41047 (N_41047,N_37734,N_36262);
nor U41048 (N_41048,N_38303,N_38300);
nand U41049 (N_41049,N_37054,N_37818);
and U41050 (N_41050,N_37342,N_39148);
xor U41051 (N_41051,N_38424,N_38656);
nand U41052 (N_41052,N_35596,N_38975);
xor U41053 (N_41053,N_38293,N_35759);
nor U41054 (N_41054,N_35858,N_35291);
nand U41055 (N_41055,N_39353,N_36962);
or U41056 (N_41056,N_36284,N_36264);
and U41057 (N_41057,N_35059,N_36668);
nor U41058 (N_41058,N_39481,N_35390);
nor U41059 (N_41059,N_37657,N_35684);
and U41060 (N_41060,N_39281,N_39869);
nor U41061 (N_41061,N_38407,N_38067);
or U41062 (N_41062,N_37086,N_38060);
or U41063 (N_41063,N_36040,N_36738);
nor U41064 (N_41064,N_36950,N_37840);
and U41065 (N_41065,N_38855,N_39437);
xor U41066 (N_41066,N_37465,N_37460);
nor U41067 (N_41067,N_37732,N_37079);
nand U41068 (N_41068,N_36095,N_36088);
and U41069 (N_41069,N_38513,N_35938);
nor U41070 (N_41070,N_39202,N_35979);
or U41071 (N_41071,N_35942,N_38487);
xnor U41072 (N_41072,N_38200,N_38548);
nor U41073 (N_41073,N_36994,N_37768);
nand U41074 (N_41074,N_39743,N_39077);
and U41075 (N_41075,N_38929,N_36240);
nor U41076 (N_41076,N_36210,N_37617);
xor U41077 (N_41077,N_37817,N_37319);
or U41078 (N_41078,N_35703,N_39190);
xor U41079 (N_41079,N_36662,N_39590);
and U41080 (N_41080,N_35901,N_35282);
xnor U41081 (N_41081,N_36760,N_37022);
nand U41082 (N_41082,N_36717,N_38971);
nor U41083 (N_41083,N_39924,N_37951);
nor U41084 (N_41084,N_38416,N_36465);
and U41085 (N_41085,N_39020,N_36359);
and U41086 (N_41086,N_38970,N_39285);
nand U41087 (N_41087,N_35990,N_39351);
xor U41088 (N_41088,N_38223,N_36140);
nor U41089 (N_41089,N_39460,N_35246);
nand U41090 (N_41090,N_37872,N_35344);
nor U41091 (N_41091,N_36942,N_39406);
xor U41092 (N_41092,N_36887,N_37956);
and U41093 (N_41093,N_38992,N_37511);
nor U41094 (N_41094,N_36934,N_36433);
and U41095 (N_41095,N_39387,N_38278);
nor U41096 (N_41096,N_38593,N_35467);
or U41097 (N_41097,N_35646,N_35898);
nor U41098 (N_41098,N_35736,N_39040);
nor U41099 (N_41099,N_37298,N_38609);
nand U41100 (N_41100,N_37204,N_38693);
nor U41101 (N_41101,N_35847,N_38379);
xnor U41102 (N_41102,N_39653,N_35936);
nor U41103 (N_41103,N_35031,N_36458);
and U41104 (N_41104,N_37497,N_35407);
nor U41105 (N_41105,N_36984,N_39415);
nand U41106 (N_41106,N_37401,N_36550);
nor U41107 (N_41107,N_36765,N_35965);
nand U41108 (N_41108,N_36776,N_37729);
nor U41109 (N_41109,N_35030,N_37326);
and U41110 (N_41110,N_39791,N_39996);
nand U41111 (N_41111,N_38729,N_37861);
nand U41112 (N_41112,N_39704,N_39264);
xor U41113 (N_41113,N_35400,N_39131);
or U41114 (N_41114,N_38423,N_37058);
and U41115 (N_41115,N_37561,N_37854);
nor U41116 (N_41116,N_37748,N_35700);
or U41117 (N_41117,N_35808,N_37043);
xnor U41118 (N_41118,N_37171,N_38033);
nand U41119 (N_41119,N_38167,N_39633);
xnor U41120 (N_41120,N_36107,N_37275);
nor U41121 (N_41121,N_37905,N_35925);
xor U41122 (N_41122,N_38176,N_36452);
nand U41123 (N_41123,N_36174,N_36334);
xor U41124 (N_41124,N_35583,N_39158);
or U41125 (N_41125,N_38577,N_35139);
or U41126 (N_41126,N_37042,N_37605);
and U41127 (N_41127,N_39772,N_39700);
nand U41128 (N_41128,N_38448,N_36858);
nor U41129 (N_41129,N_36583,N_39014);
nand U41130 (N_41130,N_38073,N_38190);
nor U41131 (N_41131,N_35702,N_38864);
or U41132 (N_41132,N_39051,N_36988);
nor U41133 (N_41133,N_37031,N_36257);
nand U41134 (N_41134,N_36560,N_38547);
and U41135 (N_41135,N_36604,N_39114);
nand U41136 (N_41136,N_35886,N_39692);
xor U41137 (N_41137,N_38429,N_39376);
nand U41138 (N_41138,N_36879,N_35020);
xor U41139 (N_41139,N_38628,N_39997);
nor U41140 (N_41140,N_39199,N_36160);
xor U41141 (N_41141,N_36409,N_39780);
nor U41142 (N_41142,N_39664,N_37492);
nor U41143 (N_41143,N_36689,N_35591);
xor U41144 (N_41144,N_39823,N_35962);
or U41145 (N_41145,N_39773,N_38406);
xnor U41146 (N_41146,N_39841,N_37973);
xor U41147 (N_41147,N_35460,N_38449);
and U41148 (N_41148,N_39615,N_39565);
nand U41149 (N_41149,N_36659,N_35334);
nor U41150 (N_41150,N_35228,N_37865);
or U41151 (N_41151,N_35889,N_37547);
or U41152 (N_41152,N_35365,N_36543);
nand U41153 (N_41153,N_38008,N_38383);
nor U41154 (N_41154,N_36680,N_39508);
nor U41155 (N_41155,N_39201,N_39306);
nand U41156 (N_41156,N_38138,N_39362);
or U41157 (N_41157,N_37622,N_38344);
nor U41158 (N_41158,N_39717,N_36486);
xnor U41159 (N_41159,N_35849,N_38121);
or U41160 (N_41160,N_39330,N_35553);
and U41161 (N_41161,N_35707,N_36569);
nand U41162 (N_41162,N_36250,N_38496);
nand U41163 (N_41163,N_37701,N_38910);
and U41164 (N_41164,N_35549,N_39461);
nor U41165 (N_41165,N_39966,N_35174);
or U41166 (N_41166,N_39338,N_36226);
or U41167 (N_41167,N_36610,N_39466);
xor U41168 (N_41168,N_39885,N_38172);
xor U41169 (N_41169,N_36020,N_39524);
xor U41170 (N_41170,N_37378,N_38099);
nand U41171 (N_41171,N_39586,N_39564);
nand U41172 (N_41172,N_36105,N_39247);
or U41173 (N_41173,N_38893,N_37076);
and U41174 (N_41174,N_39490,N_39323);
nand U41175 (N_41175,N_37265,N_39132);
nand U41176 (N_41176,N_35639,N_36048);
nor U41177 (N_41177,N_36546,N_36764);
nor U41178 (N_41178,N_39690,N_35340);
nand U41179 (N_41179,N_36808,N_38852);
nand U41180 (N_41180,N_38376,N_37446);
nand U41181 (N_41181,N_35157,N_37933);
nand U41182 (N_41182,N_37033,N_35528);
nor U41183 (N_41183,N_36860,N_38812);
and U41184 (N_41184,N_37464,N_37862);
nor U41185 (N_41185,N_35508,N_39798);
nand U41186 (N_41186,N_37751,N_35379);
xnor U41187 (N_41187,N_39910,N_39240);
xnor U41188 (N_41188,N_39657,N_36955);
xnor U41189 (N_41189,N_38900,N_37583);
nand U41190 (N_41190,N_35597,N_35489);
or U41191 (N_41191,N_38336,N_36055);
and U41192 (N_41192,N_39599,N_35771);
nor U41193 (N_41193,N_35922,N_39002);
nor U41194 (N_41194,N_35002,N_35524);
nor U41195 (N_41195,N_35214,N_36496);
nand U41196 (N_41196,N_37155,N_35042);
nand U41197 (N_41197,N_35221,N_39317);
or U41198 (N_41198,N_35756,N_39432);
nand U41199 (N_41199,N_36434,N_38092);
and U41200 (N_41200,N_39417,N_36499);
xnor U41201 (N_41201,N_36732,N_38724);
xnor U41202 (N_41202,N_38290,N_38897);
nand U41203 (N_41203,N_35527,N_37925);
xnor U41204 (N_41204,N_37952,N_35436);
nand U41205 (N_41205,N_37777,N_39789);
and U41206 (N_41206,N_36497,N_38201);
nor U41207 (N_41207,N_35327,N_35422);
nand U41208 (N_41208,N_39316,N_35317);
and U41209 (N_41209,N_37803,N_38015);
and U41210 (N_41210,N_37010,N_37140);
xor U41211 (N_41211,N_38329,N_39530);
xnor U41212 (N_41212,N_39790,N_35966);
xnor U41213 (N_41213,N_38721,N_38098);
and U41214 (N_41214,N_36255,N_36376);
nor U41215 (N_41215,N_35659,N_38474);
or U41216 (N_41216,N_39678,N_36075);
nor U41217 (N_41217,N_37948,N_39089);
nand U41218 (N_41218,N_36965,N_35619);
nor U41219 (N_41219,N_39858,N_37467);
nand U41220 (N_41220,N_39036,N_35478);
and U41221 (N_41221,N_37845,N_37240);
xor U41222 (N_41222,N_36549,N_36669);
and U41223 (N_41223,N_37926,N_35302);
nand U41224 (N_41224,N_36503,N_38267);
nor U41225 (N_41225,N_37731,N_36411);
nand U41226 (N_41226,N_36949,N_35943);
nor U41227 (N_41227,N_35474,N_38779);
xor U41228 (N_41228,N_37360,N_37609);
xor U41229 (N_41229,N_38052,N_38967);
xnor U41230 (N_41230,N_35987,N_37029);
and U41231 (N_41231,N_37879,N_35760);
or U41232 (N_41232,N_37553,N_36219);
nand U41233 (N_41233,N_38004,N_35580);
xnor U41234 (N_41234,N_35556,N_35201);
or U41235 (N_41235,N_36653,N_38963);
nor U41236 (N_41236,N_37371,N_37746);
xnor U41237 (N_41237,N_38170,N_35793);
nand U41238 (N_41238,N_37479,N_37892);
xnor U41239 (N_41239,N_38974,N_35324);
nor U41240 (N_41240,N_38173,N_37914);
and U41241 (N_41241,N_38537,N_38445);
nand U41242 (N_41242,N_38675,N_39253);
and U41243 (N_41243,N_35731,N_39932);
nor U41244 (N_41244,N_36062,N_37046);
xor U41245 (N_41245,N_38127,N_37876);
nor U41246 (N_41246,N_38862,N_36700);
xor U41247 (N_41247,N_36613,N_36443);
nor U41248 (N_41248,N_36072,N_35126);
and U41249 (N_41249,N_35821,N_38391);
nor U41250 (N_41250,N_35309,N_35252);
nor U41251 (N_41251,N_35852,N_36533);
xor U41252 (N_41252,N_39485,N_39024);
and U41253 (N_41253,N_36685,N_35640);
xor U41254 (N_41254,N_37301,N_35318);
xor U41255 (N_41255,N_37546,N_37364);
and U41256 (N_41256,N_36576,N_36707);
xnor U41257 (N_41257,N_39434,N_36180);
or U41258 (N_41258,N_36316,N_39859);
nand U41259 (N_41259,N_39943,N_37459);
and U41260 (N_41260,N_37921,N_35049);
and U41261 (N_41261,N_35903,N_37550);
and U41262 (N_41262,N_38521,N_37708);
nor U41263 (N_41263,N_37988,N_36297);
or U41264 (N_41264,N_36423,N_39360);
xnor U41265 (N_41265,N_35266,N_35767);
and U41266 (N_41266,N_38494,N_35909);
or U41267 (N_41267,N_35953,N_36022);
and U41268 (N_41268,N_35333,N_35918);
and U41269 (N_41269,N_37629,N_39995);
and U41270 (N_41270,N_38744,N_39214);
nand U41271 (N_41271,N_35204,N_37341);
xor U41272 (N_41272,N_35741,N_37785);
xnor U41273 (N_41273,N_36204,N_36406);
or U41274 (N_41274,N_36816,N_35189);
nor U41275 (N_41275,N_37423,N_37499);
nor U41276 (N_41276,N_35408,N_37822);
or U41277 (N_41277,N_36196,N_39056);
nand U41278 (N_41278,N_36390,N_35606);
nor U41279 (N_41279,N_37496,N_39661);
or U41280 (N_41280,N_35991,N_37541);
nor U41281 (N_41281,N_37800,N_39506);
nand U41282 (N_41282,N_35998,N_36265);
and U41283 (N_41283,N_38321,N_35985);
nand U41284 (N_41284,N_36759,N_35498);
and U41285 (N_41285,N_39241,N_36577);
nand U41286 (N_41286,N_39301,N_39889);
nand U41287 (N_41287,N_38302,N_39711);
nand U41288 (N_41288,N_37513,N_38310);
and U41289 (N_41289,N_37475,N_36050);
nand U41290 (N_41290,N_38871,N_35391);
and U41291 (N_41291,N_36986,N_36618);
xor U41292 (N_41292,N_37762,N_35198);
xnor U41293 (N_41293,N_35735,N_35538);
nor U41294 (N_41294,N_38000,N_36553);
or U41295 (N_41295,N_37612,N_36991);
nand U41296 (N_41296,N_35986,N_35013);
nand U41297 (N_41297,N_35179,N_38566);
nand U41298 (N_41298,N_39209,N_38818);
xor U41299 (N_41299,N_36220,N_35261);
xor U41300 (N_41300,N_35258,N_36393);
or U41301 (N_41301,N_37203,N_38284);
nand U41302 (N_41302,N_35051,N_39650);
xor U41303 (N_41303,N_39185,N_39365);
or U41304 (N_41304,N_37830,N_37095);
xnor U41305 (N_41305,N_36516,N_39186);
nor U41306 (N_41306,N_39729,N_36437);
or U41307 (N_41307,N_36096,N_39335);
nor U41308 (N_41308,N_36380,N_37597);
and U41309 (N_41309,N_36197,N_37491);
and U41310 (N_41310,N_35085,N_36936);
xor U41311 (N_41311,N_36507,N_37881);
and U41312 (N_41312,N_35381,N_36961);
nor U41313 (N_41313,N_36744,N_36762);
nand U41314 (N_41314,N_35537,N_39815);
xor U41315 (N_41315,N_36337,N_38133);
nand U41316 (N_41316,N_37470,N_38017);
nor U41317 (N_41317,N_38985,N_38804);
nand U41318 (N_41318,N_39748,N_39899);
xnor U41319 (N_41319,N_35629,N_36683);
and U41320 (N_41320,N_35164,N_35094);
and U41321 (N_41321,N_39159,N_39919);
xnor U41322 (N_41322,N_35835,N_39809);
or U41323 (N_41323,N_35129,N_36333);
and U41324 (N_41324,N_38471,N_36801);
nand U41325 (N_41325,N_38877,N_39986);
or U41326 (N_41326,N_37587,N_39295);
and U41327 (N_41327,N_37635,N_39977);
nor U41328 (N_41328,N_36407,N_35424);
xor U41329 (N_41329,N_35210,N_39549);
or U41330 (N_41330,N_39627,N_39021);
nor U41331 (N_41331,N_38255,N_38642);
xor U41332 (N_41332,N_36919,N_35098);
xnor U41333 (N_41333,N_35691,N_38972);
xnor U41334 (N_41334,N_35041,N_39459);
xor U41335 (N_41335,N_37904,N_37276);
nor U41336 (N_41336,N_38912,N_38853);
nor U41337 (N_41337,N_35983,N_35969);
nand U41338 (N_41338,N_39464,N_37368);
or U41339 (N_41339,N_38650,N_36886);
nor U41340 (N_41340,N_35149,N_36605);
nand U41341 (N_41341,N_36116,N_36686);
or U41342 (N_41342,N_37455,N_37864);
or U41343 (N_41343,N_39008,N_36590);
nand U41344 (N_41344,N_36630,N_35722);
nor U41345 (N_41345,N_38924,N_35144);
nand U41346 (N_41346,N_35584,N_36891);
xnor U41347 (N_41347,N_35238,N_37314);
and U41348 (N_41348,N_35054,N_39391);
nand U41349 (N_41349,N_39276,N_37573);
nor U41350 (N_41350,N_38151,N_35374);
and U41351 (N_41351,N_36652,N_36377);
and U41352 (N_41352,N_38555,N_37179);
and U41353 (N_41353,N_35534,N_37070);
nand U41354 (N_41354,N_37688,N_37486);
xor U41355 (N_41355,N_37789,N_38065);
xnor U41356 (N_41356,N_38527,N_37950);
nand U41357 (N_41357,N_36293,N_38084);
and U41358 (N_41358,N_39930,N_35194);
xor U41359 (N_41359,N_38124,N_35084);
and U41360 (N_41360,N_37896,N_38551);
and U41361 (N_41361,N_38991,N_36269);
and U41362 (N_41362,N_36512,N_37615);
and U41363 (N_41363,N_35956,N_36641);
nor U41364 (N_41364,N_37684,N_38009);
xor U41365 (N_41365,N_35544,N_37654);
or U41366 (N_41366,N_39065,N_37320);
and U41367 (N_41367,N_36294,N_37653);
xor U41368 (N_41368,N_39103,N_39961);
and U41369 (N_41369,N_37395,N_37545);
xnor U41370 (N_41370,N_38805,N_39265);
xor U41371 (N_41371,N_38034,N_35387);
nor U41372 (N_41372,N_35112,N_39284);
and U41373 (N_41373,N_37703,N_36152);
nand U41374 (N_41374,N_38136,N_37170);
and U41375 (N_41375,N_38534,N_38083);
or U41376 (N_41376,N_37254,N_36580);
and U41377 (N_41377,N_35670,N_37500);
nand U41378 (N_41378,N_38571,N_36932);
and U41379 (N_41379,N_38357,N_38632);
nor U41380 (N_41380,N_35733,N_39150);
nor U41381 (N_41381,N_35034,N_38500);
and U41382 (N_41382,N_37195,N_38797);
nand U41383 (N_41383,N_39609,N_37835);
nand U41384 (N_41384,N_38408,N_35268);
nand U41385 (N_41385,N_36344,N_38049);
xor U41386 (N_41386,N_36899,N_37906);
nand U41387 (N_41387,N_38461,N_38213);
or U41388 (N_41388,N_38525,N_39983);
nand U41389 (N_41389,N_35672,N_35615);
nor U41390 (N_41390,N_39608,N_36910);
nand U41391 (N_41391,N_36106,N_36833);
and U41392 (N_41392,N_37924,N_35065);
nand U41393 (N_41393,N_39402,N_35004);
and U41394 (N_41394,N_36066,N_36430);
nand U41395 (N_41395,N_36821,N_37837);
nor U41396 (N_41396,N_39092,N_38285);
nand U41397 (N_41397,N_35469,N_38876);
nand U41398 (N_41398,N_37315,N_35000);
or U41399 (N_41399,N_35503,N_39480);
nand U41400 (N_41400,N_35427,N_36862);
or U41401 (N_41401,N_36322,N_38335);
xnor U41402 (N_41402,N_39667,N_35745);
or U41403 (N_41403,N_35180,N_36408);
xor U41404 (N_41404,N_39361,N_37096);
nor U41405 (N_41405,N_36306,N_35971);
nand U41406 (N_41406,N_37241,N_37190);
nor U41407 (N_41407,N_35968,N_35773);
nand U41408 (N_41408,N_37099,N_37575);
nor U41409 (N_41409,N_35569,N_35762);
nand U41410 (N_41410,N_38800,N_38875);
and U41411 (N_41411,N_37392,N_37279);
or U41412 (N_41412,N_37958,N_36058);
nor U41413 (N_41413,N_38353,N_38528);
or U41414 (N_41414,N_37284,N_36941);
nor U41415 (N_41415,N_35900,N_37646);
nor U41416 (N_41416,N_35786,N_37638);
or U41417 (N_41417,N_39863,N_36536);
nor U41418 (N_41418,N_37718,N_39368);
and U41419 (N_41419,N_39010,N_37072);
or U41420 (N_41420,N_39333,N_38940);
nand U41421 (N_41421,N_39629,N_36615);
nor U41422 (N_41422,N_37192,N_35805);
nand U41423 (N_41423,N_39828,N_37549);
nor U41424 (N_41424,N_38478,N_36386);
nand U41425 (N_41425,N_39139,N_38796);
nand U41426 (N_41426,N_39439,N_35505);
nand U41427 (N_41427,N_39797,N_39016);
and U41428 (N_41428,N_38194,N_38938);
nor U41429 (N_41429,N_39938,N_38794);
and U41430 (N_41430,N_36581,N_36351);
or U41431 (N_41431,N_36582,N_36191);
nor U41432 (N_41432,N_36024,N_39419);
nand U41433 (N_41433,N_39162,N_38736);
and U41434 (N_41434,N_38250,N_39393);
nor U41435 (N_41435,N_38274,N_39585);
and U41436 (N_41436,N_37705,N_39117);
xnor U41437 (N_41437,N_39331,N_38431);
or U41438 (N_41438,N_37911,N_38750);
or U41439 (N_41439,N_36179,N_35251);
or U41440 (N_41440,N_37452,N_37332);
or U41441 (N_41441,N_35810,N_37102);
xor U41442 (N_41442,N_38468,N_39025);
nand U41443 (N_41443,N_39866,N_38976);
and U41444 (N_41444,N_37268,N_37047);
nand U41445 (N_41445,N_37050,N_36723);
or U41446 (N_41446,N_36364,N_38636);
nor U41447 (N_41447,N_39115,N_39538);
or U41448 (N_41448,N_39428,N_37539);
and U41449 (N_41449,N_39321,N_37397);
xor U41450 (N_41450,N_38765,N_39952);
xor U41451 (N_41451,N_38467,N_35929);
xor U41452 (N_41452,N_39901,N_37327);
xor U41453 (N_41453,N_36648,N_39135);
and U41454 (N_41454,N_35286,N_37433);
or U41455 (N_41455,N_37501,N_37357);
nand U41456 (N_41456,N_37772,N_37970);
and U41457 (N_41457,N_38043,N_39985);
or U41458 (N_41458,N_39300,N_36319);
nor U41459 (N_41459,N_35701,N_37888);
or U41460 (N_41460,N_35079,N_36654);
xnor U41461 (N_41461,N_35561,N_36491);
nand U41462 (N_41462,N_37960,N_36966);
or U41463 (N_41463,N_35674,N_36034);
nor U41464 (N_41464,N_36457,N_37839);
nor U41465 (N_41465,N_38155,N_39926);
nor U41466 (N_41466,N_35568,N_39465);
or U41467 (N_41467,N_35506,N_39738);
xnor U41468 (N_41468,N_35438,N_35917);
nand U41469 (N_41469,N_39217,N_35806);
xor U41470 (N_41470,N_35517,N_35565);
nor U41471 (N_41471,N_38937,N_38470);
nand U41472 (N_41472,N_35060,N_38747);
and U41473 (N_41473,N_35651,N_38738);
nand U41474 (N_41474,N_35058,N_37391);
and U41475 (N_41475,N_37602,N_38949);
xor U41476 (N_41476,N_38606,N_37649);
nor U41477 (N_41477,N_37853,N_37104);
nor U41478 (N_41478,N_35592,N_35222);
nand U41479 (N_41479,N_36201,N_37702);
and U41480 (N_41480,N_38483,N_36332);
and U41481 (N_41481,N_36482,N_38886);
or U41482 (N_41482,N_38069,N_39275);
nor U41483 (N_41483,N_38772,N_36627);
nand U41484 (N_41484,N_39118,N_39903);
or U41485 (N_41485,N_38164,N_35796);
xnor U41486 (N_41486,N_36412,N_39486);
xnor U41487 (N_41487,N_38094,N_37083);
or U41488 (N_41488,N_37581,N_38280);
xor U41489 (N_41489,N_35380,N_37114);
xnor U41490 (N_41490,N_37193,N_36609);
nor U41491 (N_41491,N_37295,N_36206);
nand U41492 (N_41492,N_35678,N_35586);
nand U41493 (N_41493,N_36127,N_39259);
or U41494 (N_41494,N_37256,N_39686);
and U41495 (N_41495,N_38193,N_39534);
nand U41496 (N_41496,N_37843,N_38965);
nand U41497 (N_41497,N_38958,N_36530);
or U41498 (N_41498,N_37434,N_36935);
xnor U41499 (N_41499,N_35574,N_39424);
nor U41500 (N_41500,N_37004,N_35018);
nor U41501 (N_41501,N_35696,N_35278);
or U41502 (N_41502,N_35838,N_39216);
nand U41503 (N_41503,N_38580,N_38450);
nor U41504 (N_41504,N_36225,N_39451);
or U41505 (N_41505,N_36099,N_38364);
nand U41506 (N_41506,N_39328,N_35178);
and U41507 (N_41507,N_38454,N_39343);
and U41508 (N_41508,N_35277,N_36474);
nand U41509 (N_41509,N_35981,N_39273);
or U41510 (N_41510,N_38788,N_37466);
xnor U41511 (N_41511,N_37440,N_37438);
and U41512 (N_41512,N_36861,N_35611);
and U41513 (N_41513,N_36800,N_36587);
and U41514 (N_41514,N_38488,N_38740);
or U41515 (N_41515,N_35235,N_39105);
and U41516 (N_41516,N_38755,N_39579);
nand U41517 (N_41517,N_39071,N_35988);
or U41518 (N_41518,N_36441,N_38857);
or U41519 (N_41519,N_38053,N_35078);
nor U41520 (N_41520,N_38904,N_36165);
or U41521 (N_41521,N_37534,N_36741);
xor U41522 (N_41522,N_35289,N_39487);
xor U41523 (N_41523,N_36154,N_37133);
nor U41524 (N_41524,N_36646,N_37405);
and U41525 (N_41525,N_37067,N_35795);
and U41526 (N_41526,N_38702,N_37874);
xnor U41527 (N_41527,N_36665,N_39652);
xor U41528 (N_41528,N_37023,N_38562);
nor U41529 (N_41529,N_39893,N_35645);
nand U41530 (N_41530,N_36424,N_37182);
xnor U41531 (N_41531,N_36275,N_39649);
xor U41532 (N_41532,N_37040,N_37844);
or U41533 (N_41533,N_39448,N_37873);
nand U41534 (N_41534,N_38306,N_38946);
nor U41535 (N_41535,N_37249,N_38786);
xnor U41536 (N_41536,N_35014,N_39622);
and U41537 (N_41537,N_37672,N_36573);
nor U41538 (N_41538,N_36221,N_38541);
xnor U41539 (N_41539,N_39752,N_39612);
xnor U41540 (N_41540,N_39462,N_36731);
nor U41541 (N_41541,N_35169,N_37598);
xnor U41542 (N_41542,N_39493,N_39263);
xnor U41543 (N_41543,N_39621,N_36974);
and U41544 (N_41544,N_39805,N_36774);
nand U41545 (N_41545,N_36824,N_36979);
nor U41546 (N_41546,N_39369,N_35958);
or U41547 (N_41547,N_38147,N_37947);
nor U41548 (N_41548,N_39635,N_39473);
and U41549 (N_41549,N_35749,N_36987);
nand U41550 (N_41550,N_35578,N_38803);
xnor U41551 (N_41551,N_39713,N_37296);
nand U41552 (N_41552,N_39547,N_35202);
xnor U41553 (N_41553,N_39703,N_36693);
and U41554 (N_41554,N_35432,N_36702);
xor U41555 (N_41555,N_35331,N_36739);
nor U41556 (N_41556,N_38390,N_35920);
and U41557 (N_41557,N_38759,N_36464);
nor U41558 (N_41558,N_35690,N_37106);
xor U41559 (N_41559,N_35839,N_38979);
nand U41560 (N_41560,N_38326,N_35035);
xor U41561 (N_41561,N_38714,N_38037);
nand U41562 (N_41562,N_35915,N_36670);
xor U41563 (N_41563,N_38793,N_39127);
nor U41564 (N_41564,N_39137,N_36378);
and U41565 (N_41565,N_35110,N_39425);
xor U41566 (N_41566,N_38543,N_36209);
nand U41567 (N_41567,N_37194,N_37898);
nor U41568 (N_41568,N_37239,N_37398);
nand U41569 (N_41569,N_38050,N_37931);
and U41570 (N_41570,N_37755,N_36820);
and U41571 (N_41571,N_35444,N_35462);
nand U41572 (N_41572,N_39708,N_36077);
nor U41573 (N_41573,N_38107,N_37998);
and U41574 (N_41574,N_35314,N_38925);
and U41575 (N_41575,N_37591,N_36079);
xnor U41576 (N_41576,N_36103,N_36381);
nand U41577 (N_41577,N_37738,N_38397);
or U41578 (N_41578,N_37880,N_36098);
nor U41579 (N_41579,N_38137,N_37154);
nand U41580 (N_41580,N_39356,N_35017);
nand U41581 (N_41581,N_38616,N_36951);
or U41582 (N_41582,N_35883,N_36829);
nand U41583 (N_41583,N_35518,N_37299);
nor U41584 (N_41584,N_37663,N_36954);
or U41585 (N_41585,N_35514,N_36398);
or U41586 (N_41586,N_35485,N_35150);
nor U41587 (N_41587,N_37733,N_35143);
nor U41588 (N_41588,N_35043,N_38485);
nand U41589 (N_41589,N_37724,N_35471);
or U41590 (N_41590,N_36943,N_37365);
or U41591 (N_41591,N_39101,N_36501);
nand U41592 (N_41592,N_37089,N_35009);
or U41593 (N_41593,N_36256,N_37164);
nor U41594 (N_41594,N_38328,N_35899);
nand U41595 (N_41595,N_35299,N_39844);
xor U41596 (N_41596,N_37152,N_38340);
nor U41597 (N_41597,N_38322,N_36327);
and U41598 (N_41598,N_38095,N_35845);
and U41599 (N_41599,N_35687,N_36985);
or U41600 (N_41600,N_36572,N_35227);
nand U41601 (N_41601,N_38681,N_36773);
nor U41602 (N_41602,N_36123,N_36243);
or U41603 (N_41603,N_35368,N_39606);
nand U41604 (N_41604,N_39906,N_39244);
xor U41605 (N_41605,N_38354,N_38144);
nor U41606 (N_41606,N_36484,N_39974);
xor U41607 (N_41607,N_37426,N_35303);
nor U41608 (N_41608,N_38913,N_37260);
nand U41609 (N_41609,N_39195,N_37518);
nand U41610 (N_41610,N_38166,N_35496);
xor U41611 (N_41611,N_38259,N_37113);
nand U41612 (N_41612,N_38745,N_39134);
and U41613 (N_41613,N_36907,N_35075);
nand U41614 (N_41614,N_37604,N_38657);
xnor U41615 (N_41615,N_38455,N_39504);
or U41616 (N_41616,N_36117,N_36041);
and U41617 (N_41617,N_37765,N_35593);
xor U41618 (N_41618,N_38381,N_38659);
xor U41619 (N_41619,N_35388,N_39455);
and U41620 (N_41620,N_39389,N_35588);
nor U41621 (N_41621,N_36745,N_36301);
and U41622 (N_41622,N_39429,N_37554);
nor U41623 (N_41623,N_38920,N_38865);
nor U41624 (N_41624,N_36619,N_35815);
xor U41625 (N_41625,N_39796,N_37380);
nor U41626 (N_41626,N_35187,N_36186);
or U41627 (N_41627,N_39951,N_39382);
xor U41628 (N_41628,N_35181,N_39096);
nand U41629 (N_41629,N_38896,N_39758);
nand U41630 (N_41630,N_39047,N_39600);
nor U41631 (N_41631,N_37570,N_35661);
or U41632 (N_41632,N_39978,N_37794);
nand U41633 (N_41633,N_38640,N_38059);
or U41634 (N_41634,N_38579,N_36600);
or U41635 (N_41635,N_39557,N_35726);
and U41636 (N_41636,N_37969,N_37418);
nor U41637 (N_41637,N_35310,N_38763);
nand U41638 (N_41638,N_36493,N_39359);
or U41639 (N_41639,N_36005,N_36313);
nand U41640 (N_41640,N_36601,N_36743);
nand U41641 (N_41641,N_36614,N_39610);
nand U41642 (N_41642,N_37061,N_38669);
nor U41643 (N_41643,N_39799,N_37692);
xor U41644 (N_41644,N_38463,N_38561);
nand U41645 (N_41645,N_39991,N_38412);
and U41646 (N_41646,N_38776,N_39533);
and U41647 (N_41647,N_35470,N_37799);
or U41648 (N_41648,N_35932,N_36679);
or U41649 (N_41649,N_37451,N_35677);
nor U41650 (N_41650,N_35563,N_35005);
or U41651 (N_41651,N_36481,N_38816);
or U41652 (N_41652,N_39037,N_39395);
and U41653 (N_41653,N_39206,N_39982);
and U41654 (N_41654,N_35109,N_39640);
or U41655 (N_41655,N_36469,N_38472);
xnor U41656 (N_41656,N_37090,N_39699);
and U41657 (N_41657,N_38761,N_36742);
or U41658 (N_41658,N_36539,N_35290);
nand U41659 (N_41659,N_35006,N_36156);
or U41660 (N_41660,N_39720,N_38047);
nand U41661 (N_41661,N_38199,N_35689);
and U41662 (N_41662,N_38492,N_36299);
nor U41663 (N_41663,N_35935,N_38573);
nor U41664 (N_41664,N_37421,N_37536);
nor U41665 (N_41665,N_39157,N_35484);
and U41666 (N_41666,N_37235,N_37430);
and U41667 (N_41667,N_35350,N_37404);
or U41668 (N_41668,N_37949,N_35248);
nor U41669 (N_41669,N_38330,N_36977);
nor U41670 (N_41670,N_38504,N_38243);
nor U41671 (N_41671,N_37402,N_36155);
and U41672 (N_41672,N_38943,N_39483);
nand U41673 (N_41673,N_37616,N_36046);
nor U41674 (N_41674,N_39817,N_37174);
nor U41675 (N_41675,N_35911,N_36233);
and U41676 (N_41676,N_36660,N_37183);
and U41677 (N_41677,N_36697,N_35542);
xor U41678 (N_41678,N_36926,N_36694);
xor U41679 (N_41679,N_38292,N_35720);
nand U41680 (N_41680,N_35106,N_36307);
xnor U41681 (N_41681,N_39611,N_39597);
or U41682 (N_41682,N_39410,N_35209);
nor U41683 (N_41683,N_39944,N_37691);
nand U41684 (N_41684,N_35840,N_39043);
or U41685 (N_41685,N_35850,N_35377);
and U41686 (N_41686,N_38152,N_35195);
nor U41687 (N_41687,N_37942,N_37637);
xnor U41688 (N_41688,N_37778,N_36172);
xnor U41689 (N_41689,N_37930,N_36953);
and U41690 (N_41690,N_35515,N_38308);
or U41691 (N_41691,N_38400,N_38160);
or U41692 (N_41692,N_36462,N_37743);
nor U41693 (N_41693,N_36597,N_36455);
or U41694 (N_41694,N_39324,N_37601);
and U41695 (N_41695,N_35011,N_39102);
and U41696 (N_41696,N_37121,N_38002);
and U41697 (N_41697,N_37760,N_35967);
xor U41698 (N_41698,N_35364,N_37717);
xor U41699 (N_41699,N_37055,N_39015);
nand U41700 (N_41700,N_35727,N_38599);
nor U41701 (N_41701,N_36788,N_39374);
or U41702 (N_41702,N_37695,N_39956);
nor U41703 (N_41703,N_39513,N_38824);
nor U41704 (N_41704,N_36783,N_39172);
and U41705 (N_41705,N_38140,N_37303);
nand U41706 (N_41706,N_35602,N_37564);
xnor U41707 (N_41707,N_35312,N_39887);
and U41708 (N_41708,N_38260,N_37685);
or U41709 (N_41709,N_38723,N_37228);
or U41710 (N_41710,N_39003,N_36920);
nand U41711 (N_41711,N_37700,N_37667);
nand U41712 (N_41712,N_39914,N_35637);
and U41713 (N_41713,N_35910,N_37381);
xnor U41714 (N_41714,N_38507,N_38091);
nor U41715 (N_41715,N_35033,N_35225);
nor U41716 (N_41716,N_38888,N_35636);
xor U41717 (N_41717,N_36288,N_39950);
xnor U41718 (N_41718,N_36320,N_37498);
and U41719 (N_41719,N_36629,N_38301);
or U41720 (N_41720,N_37191,N_37424);
nor U41721 (N_41721,N_37060,N_39674);
xor U41722 (N_41722,N_35789,N_37983);
or U41723 (N_41723,N_38128,N_35706);
nand U41724 (N_41724,N_38497,N_39980);
nand U41725 (N_41725,N_36328,N_36252);
nor U41726 (N_41726,N_35679,N_38182);
xnor U41727 (N_41727,N_36688,N_39831);
nand U41728 (N_41728,N_39912,N_38923);
nor U41729 (N_41729,N_35947,N_37725);
xor U41730 (N_41730,N_37345,N_38057);
xnor U41731 (N_41731,N_39693,N_35945);
or U41732 (N_41732,N_38994,N_39681);
nand U41733 (N_41733,N_37189,N_36480);
xnor U41734 (N_41734,N_38462,N_35423);
and U41735 (N_41735,N_35671,N_37592);
and U41736 (N_41736,N_36567,N_39689);
and U41737 (N_41737,N_39740,N_38208);
and U41738 (N_41738,N_36432,N_39691);
nand U41739 (N_41739,N_36477,N_38891);
xnor U41740 (N_41740,N_38679,N_37737);
and U41741 (N_41741,N_39672,N_38196);
nor U41742 (N_41742,N_37075,N_39624);
or U41743 (N_41743,N_36898,N_38791);
or U41744 (N_41744,N_35809,N_38473);
nor U41745 (N_41745,N_38915,N_38453);
xor U41746 (N_41746,N_35298,N_36339);
nor U41747 (N_41747,N_39891,N_36664);
or U41748 (N_41748,N_35372,N_39309);
nor U41749 (N_41749,N_36869,N_35175);
and U41750 (N_41750,N_38523,N_38016);
xor U41751 (N_41751,N_39125,N_35367);
xnor U41752 (N_41752,N_37611,N_38826);
xnor U41753 (N_41753,N_36832,N_38510);
and U41754 (N_41754,N_36111,N_39880);
nor U41755 (N_41755,N_35928,N_38649);
nand U41756 (N_41756,N_36218,N_39427);
nand U41757 (N_41757,N_37431,N_35604);
nand U41758 (N_41758,N_38432,N_38836);
nor U41759 (N_41759,N_36283,N_37574);
and U41760 (N_41760,N_39843,N_37608);
or U41761 (N_41761,N_35975,N_37409);
xnor U41762 (N_41762,N_38662,N_37419);
and U41763 (N_41763,N_38109,N_38795);
nor U41764 (N_41764,N_36995,N_37590);
xor U41765 (N_41765,N_38707,N_35115);
nand U41766 (N_41766,N_37243,N_36495);
nor U41767 (N_41767,N_39059,N_38331);
and U41768 (N_41768,N_39138,N_37175);
xor U41769 (N_41769,N_35253,N_35791);
nor U41770 (N_41770,N_38664,N_35415);
xor U41771 (N_41771,N_39079,N_38116);
or U41772 (N_41772,N_39575,N_39742);
nor U41773 (N_41773,N_35881,N_38058);
nor U41774 (N_41774,N_39401,N_38222);
nor U41775 (N_41775,N_38012,N_39503);
and U41776 (N_41776,N_36511,N_38817);
nand U41777 (N_41777,N_37786,N_35530);
nand U41778 (N_41778,N_38942,N_39142);
nand U41779 (N_41779,N_36413,N_35590);
nand U41780 (N_41780,N_39614,N_36027);
xor U41781 (N_41781,N_35855,N_39026);
or U41782 (N_41782,N_37757,N_37462);
nor U41783 (N_41783,N_37571,N_35127);
and U41784 (N_41784,N_37211,N_35587);
nor U41785 (N_41785,N_38221,N_39363);
xnor U41786 (N_41786,N_38978,N_35711);
and U41787 (N_41787,N_39149,N_38569);
xnor U41788 (N_41788,N_35151,N_36102);
xor U41789 (N_41789,N_38342,N_36721);
or U41790 (N_41790,N_35413,N_39042);
and U41791 (N_41791,N_39189,N_39571);
nand U41792 (N_41792,N_35220,N_37153);
nor U41793 (N_41793,N_36747,N_36132);
nor U41794 (N_41794,N_36084,N_37727);
or U41795 (N_41795,N_39989,N_38777);
xor U41796 (N_41796,N_38061,N_37094);
or U41797 (N_41797,N_36070,N_35995);
or U41798 (N_41798,N_38077,N_39246);
nor U41799 (N_41799,N_36785,N_39307);
nand U41800 (N_41800,N_38204,N_39034);
xnor U41801 (N_41801,N_35008,N_37478);
and U41802 (N_41802,N_39262,N_35396);
and U41803 (N_41803,N_37270,N_35688);
nor U41804 (N_41804,N_36915,N_36200);
nand U41805 (N_41805,N_39876,N_38333);
nand U41806 (N_41806,N_36515,N_37248);
nor U41807 (N_41807,N_35652,N_37713);
and U41808 (N_41808,N_36324,N_38319);
nand U41809 (N_41809,N_35215,N_35658);
nand U41810 (N_41810,N_39813,N_39774);
and U41811 (N_41811,N_39108,N_38415);
and U41812 (N_41812,N_37084,N_39801);
and U41813 (N_41813,N_35705,N_39569);
nor U41814 (N_41814,N_37100,N_36647);
nand U41815 (N_41815,N_36422,N_37520);
nand U41816 (N_41816,N_35650,N_39881);
and U41817 (N_41817,N_35949,N_35363);
and U41818 (N_41818,N_36052,N_36504);
nor U41819 (N_41819,N_37463,N_35664);
nor U41820 (N_41820,N_37927,N_37982);
nor U41821 (N_41821,N_35281,N_39722);
xor U41822 (N_41822,N_36903,N_39514);
nor U41823 (N_41823,N_37336,N_37720);
or U41824 (N_41824,N_38010,N_38554);
nand U41825 (N_41825,N_39271,N_36110);
or U41826 (N_41826,N_39067,N_39819);
nand U41827 (N_41827,N_38908,N_35876);
or U41828 (N_41828,N_35978,N_35669);
nand U41829 (N_41829,N_37468,N_37312);
nand U41830 (N_41830,N_37027,N_37377);
xnor U41831 (N_41831,N_37346,N_38411);
nor U41832 (N_41832,N_39011,N_35360);
nand U41833 (N_41833,N_37711,N_38215);
or U41834 (N_41834,N_37297,N_39288);
and U41835 (N_41835,N_39922,N_35828);
nand U41836 (N_41836,N_39778,N_36270);
nor U41837 (N_41837,N_37062,N_39725);
xnor U41838 (N_41838,N_39299,N_36574);
and U41839 (N_41839,N_35952,N_38126);
nand U41840 (N_41840,N_37300,N_36846);
xnor U41841 (N_41841,N_37962,N_37088);
nand U41842 (N_41842,N_38694,N_39269);
and U41843 (N_41843,N_37428,N_37756);
and U41844 (N_41844,N_39188,N_37339);
nor U41845 (N_41845,N_37236,N_38951);
or U41846 (N_41846,N_37443,N_38457);
or U41847 (N_41847,N_36157,N_35445);
nor U41848 (N_41848,N_35269,N_39326);
xnor U41849 (N_41849,N_38398,N_36131);
xnor U41850 (N_41850,N_38544,N_37780);
xnor U41851 (N_41851,N_39243,N_38205);
xor U41852 (N_41852,N_35853,N_36168);
nor U41853 (N_41853,N_38725,N_36285);
nor U41854 (N_41854,N_35529,N_35356);
xor U41855 (N_41855,N_38635,N_36596);
xnor U41856 (N_41856,N_37714,N_35063);
or U41857 (N_41857,N_36032,N_39904);
xor U41858 (N_41858,N_35250,N_36786);
nor U41859 (N_41859,N_36551,N_37769);
or U41860 (N_41860,N_39976,N_37671);
nor U41861 (N_41861,N_37041,N_36538);
nor U41862 (N_41862,N_38945,N_37388);
and U41863 (N_41863,N_39107,N_36771);
nor U41864 (N_41864,N_35717,N_39104);
nand U41865 (N_41865,N_36211,N_35418);
nor U41866 (N_41866,N_39329,N_37220);
xnor U41867 (N_41867,N_35082,N_35389);
nor U41868 (N_41868,N_37039,N_39835);
xor U41869 (N_41869,N_36355,N_35699);
and U41870 (N_41870,N_37233,N_35662);
nand U41871 (N_41871,N_35487,N_35061);
xnor U41872 (N_41872,N_37257,N_39883);
xnor U41873 (N_41873,N_35199,N_38314);
and U41874 (N_41874,N_36506,N_36038);
xnor U41875 (N_41875,N_35239,N_36227);
nor U41876 (N_41876,N_36388,N_38549);
nand U41877 (N_41877,N_38382,N_39842);
xor U41878 (N_41878,N_39278,N_36400);
and U41879 (N_41879,N_37285,N_38637);
nand U41880 (N_41880,N_36724,N_38237);
or U41881 (N_41881,N_35026,N_38363);
nand U41882 (N_41882,N_35362,N_39405);
nor U41883 (N_41883,N_35788,N_39941);
and U41884 (N_41884,N_39670,N_35800);
xor U41885 (N_41885,N_39907,N_38914);
nand U41886 (N_41886,N_38837,N_39337);
nor U41887 (N_41887,N_36309,N_35420);
and U41888 (N_41888,N_39078,N_35081);
nor U41889 (N_41889,N_37589,N_35856);
or U41890 (N_41890,N_39058,N_37610);
xor U41891 (N_41891,N_38667,N_37828);
or U41892 (N_41892,N_36525,N_36326);
and U41893 (N_41893,N_38038,N_37516);
nor U41894 (N_41894,N_38530,N_37533);
or U41895 (N_41895,N_36471,N_39953);
nor U41896 (N_41896,N_38244,N_39315);
nor U41897 (N_41897,N_36169,N_37439);
nand U41898 (N_41898,N_37741,N_39598);
and U41899 (N_41899,N_36286,N_36690);
and U41900 (N_41900,N_36135,N_37159);
xor U41901 (N_41901,N_35787,N_39747);
and U41902 (N_41902,N_35232,N_39334);
or U41903 (N_41903,N_38288,N_37522);
and U41904 (N_41904,N_36426,N_38647);
xor U41905 (N_41905,N_39012,N_36335);
and U41906 (N_41906,N_37456,N_36634);
nor U41907 (N_41907,N_38596,N_38066);
and U41908 (N_41908,N_39073,N_35522);
nand U41909 (N_41909,N_38784,N_39282);
nand U41910 (N_41910,N_39984,N_36676);
and U41911 (N_41911,N_37897,N_37006);
and U41912 (N_41912,N_38749,N_35224);
and U41913 (N_41913,N_38509,N_37453);
nor U41914 (N_41914,N_37238,N_35279);
or U41915 (N_41915,N_39786,N_37288);
and U41916 (N_41916,N_38247,N_39856);
nand U41917 (N_41917,N_38990,N_38808);
or U41918 (N_41918,N_35663,N_37838);
and U41919 (N_41919,N_39261,N_35763);
and U41920 (N_41920,N_39082,N_38921);
xor U41921 (N_41921,N_37390,N_35052);
and U41922 (N_41922,N_36752,N_39472);
nand U41923 (N_41923,N_39850,N_37120);
and U41924 (N_41924,N_39602,N_39913);
xor U41925 (N_41925,N_39935,N_37957);
nor U41926 (N_41926,N_38380,N_38901);
nand U41927 (N_41927,N_38715,N_36405);
nand U41928 (N_41928,N_36980,N_39004);
or U41929 (N_41929,N_39444,N_38148);
xnor U41930 (N_41930,N_37334,N_39902);
or U41931 (N_41931,N_39964,N_37165);
xnor U41932 (N_41932,N_36636,N_37980);
nand U41933 (N_41933,N_35875,N_35133);
nor U41934 (N_41934,N_36119,N_38986);
and U41935 (N_41935,N_38096,N_37625);
nor U41936 (N_41936,N_36868,N_38417);
xnor U41937 (N_41937,N_35521,N_35486);
or U41938 (N_41938,N_36042,N_38165);
or U41939 (N_41939,N_37012,N_37267);
nor U41940 (N_41940,N_37971,N_38230);
or U41941 (N_41941,N_39375,N_39937);
nor U41942 (N_41942,N_39344,N_36757);
xor U41943 (N_41943,N_36001,N_38959);
nor U41944 (N_41944,N_36396,N_38517);
and U41945 (N_41945,N_36108,N_39820);
and U41946 (N_41946,N_35894,N_35976);
xnor U41947 (N_41947,N_35183,N_38829);
or U41948 (N_41948,N_36542,N_35411);
or U41949 (N_41949,N_38277,N_37525);
or U41950 (N_41950,N_36751,N_35571);
or U41951 (N_41951,N_39145,N_35776);
nand U41952 (N_41952,N_39446,N_35616);
nor U41953 (N_41953,N_37815,N_37829);
xor U41954 (N_41954,N_37810,N_39673);
nor U41955 (N_41955,N_36237,N_39053);
and U41956 (N_41956,N_37959,N_38760);
nand U41957 (N_41957,N_35649,N_36888);
nand U41958 (N_41958,N_36975,N_38720);
or U41959 (N_41959,N_38591,N_39662);
and U41960 (N_41960,N_38011,N_37767);
nor U41961 (N_41961,N_35383,N_36272);
xor U41962 (N_41962,N_36768,N_39824);
and U41963 (N_41963,N_37021,N_38365);
nand U41964 (N_41964,N_38027,N_37826);
or U41965 (N_41965,N_36410,N_39588);
and U41966 (N_41966,N_38022,N_37125);
nand U41967 (N_41967,N_36758,N_39923);
nand U41968 (N_41968,N_39554,N_38334);
or U41969 (N_41969,N_39716,N_35758);
nand U41970 (N_41970,N_37354,N_35573);
or U41971 (N_41971,N_36978,N_37372);
and U41972 (N_41972,N_36150,N_37290);
and U41973 (N_41973,N_38939,N_37548);
nor U41974 (N_41974,N_38512,N_37752);
xor U41975 (N_41975,N_35761,N_36672);
nand U41976 (N_41976,N_36799,N_37677);
and U41977 (N_41977,N_39094,N_36956);
nand U41978 (N_41978,N_36667,N_36805);
nand U41979 (N_41979,N_37351,N_38031);
and U41980 (N_41980,N_39971,N_36914);
nand U41981 (N_41981,N_37850,N_37373);
and U41982 (N_41982,N_36713,N_35358);
nor U41983 (N_41983,N_35557,N_39779);
nor U41984 (N_41984,N_38425,N_36939);
xor U41985 (N_41985,N_36575,N_39867);
or U41986 (N_41986,N_39753,N_35950);
xnor U41987 (N_41987,N_38995,N_36015);
nand U41988 (N_41988,N_39578,N_39916);
and U41989 (N_41989,N_37348,N_39764);
nand U41990 (N_41990,N_36967,N_36564);
or U41991 (N_41991,N_36855,N_36828);
nor U41992 (N_41992,N_39776,N_37899);
nand U41993 (N_41993,N_35262,N_38982);
and U41994 (N_41994,N_37833,N_38898);
xor U41995 (N_41995,N_37964,N_37715);
and U41996 (N_41996,N_37318,N_39644);
xor U41997 (N_41997,N_35919,N_35337);
and U41998 (N_41998,N_38672,N_35271);
nand U41999 (N_41999,N_37650,N_37025);
xnor U42000 (N_42000,N_36540,N_35153);
nor U42001 (N_42001,N_38475,N_37623);
nor U42002 (N_42002,N_35155,N_37965);
nor U42003 (N_42003,N_36187,N_39399);
or U42004 (N_42004,N_38575,N_36902);
xnor U42005 (N_42005,N_39975,N_38146);
and U42006 (N_42006,N_37606,N_38042);
nand U42007 (N_42007,N_36901,N_39821);
xor U42008 (N_42008,N_37436,N_38768);
and U42009 (N_42009,N_36534,N_35951);
nand U42010 (N_42010,N_38421,N_37721);
and U42011 (N_42011,N_35021,N_37683);
or U42012 (N_42012,N_38831,N_39054);
or U42013 (N_42013,N_39249,N_35523);
nand U42014 (N_42014,N_35176,N_39829);
and U42015 (N_42015,N_39100,N_39475);
or U42016 (N_42016,N_35851,N_37108);
nor U42017 (N_42017,N_36677,N_37811);
and U42018 (N_42018,N_38718,N_36086);
xor U42019 (N_42019,N_39623,N_37557);
nand U42020 (N_42020,N_39683,N_39298);
xnor U42021 (N_42021,N_35860,N_35819);
xnor U42022 (N_42022,N_36802,N_37640);
xor U42023 (N_42023,N_39500,N_35877);
and U42024 (N_42024,N_37736,N_38168);
and U42025 (N_42025,N_38360,N_36049);
and U42026 (N_42026,N_35770,N_35355);
and U42027 (N_42027,N_36911,N_38683);
nand U42028 (N_42028,N_39193,N_35757);
and U42029 (N_42029,N_36789,N_39857);
or U42030 (N_42030,N_37770,N_36945);
xnor U42031 (N_42031,N_38766,N_39715);
and U42032 (N_42032,N_36296,N_36063);
and U42033 (N_42033,N_37595,N_39310);
nand U42034 (N_42034,N_38851,N_35405);
and U42035 (N_42035,N_35831,N_39958);
nand U42036 (N_42036,N_39694,N_39735);
nor U42037 (N_42037,N_38028,N_36521);
nor U42038 (N_42038,N_38748,N_37130);
and U42039 (N_42039,N_36008,N_35038);
or U42040 (N_42040,N_36916,N_38025);
or U42041 (N_42041,N_38872,N_35902);
nand U42042 (N_42042,N_35643,N_38216);
or U42043 (N_42043,N_39274,N_39197);
and U42044 (N_42044,N_36416,N_37044);
nand U42045 (N_42045,N_36593,N_35057);
xor U42046 (N_42046,N_38856,N_39994);
or U42047 (N_42047,N_35103,N_38968);
nand U42048 (N_42048,N_35896,N_39626);
xor U42049 (N_42049,N_39205,N_35630);
or U42050 (N_42050,N_37889,N_37774);
or U42051 (N_42051,N_38666,N_39045);
nor U42052 (N_42052,N_36981,N_35743);
xnor U42053 (N_42053,N_36082,N_38931);
nand U42054 (N_42054,N_38535,N_39418);
nor U42055 (N_42055,N_35068,N_36895);
xnor U42056 (N_42056,N_36803,N_36993);
nor U42057 (N_42057,N_36719,N_35535);
or U42058 (N_42058,N_36121,N_35937);
and U42059 (N_42059,N_39196,N_37358);
nor U42060 (N_42060,N_35714,N_39447);
nand U42061 (N_42061,N_37593,N_37852);
nor U42062 (N_42062,N_38601,N_39830);
and U42063 (N_42063,N_35159,N_35775);
or U42064 (N_42064,N_38006,N_36176);
nand U42065 (N_42065,N_37264,N_37304);
and U42066 (N_42066,N_38980,N_38209);
and U42067 (N_42067,N_39342,N_35880);
nand U42068 (N_42068,N_36594,N_37129);
nand U42069 (N_42069,N_39463,N_37406);
nand U42070 (N_42070,N_38111,N_38256);
or U42071 (N_42071,N_37369,N_37798);
nand U42072 (N_42072,N_35811,N_37328);
nand U42073 (N_42073,N_35468,N_36514);
xnor U42074 (N_42074,N_37857,N_35863);
xor U42075 (N_42075,N_35122,N_38289);
nand U42076 (N_42076,N_35641,N_35632);
and U42077 (N_42077,N_38746,N_36793);
xor U42078 (N_42078,N_35233,N_37537);
xor U42079 (N_42079,N_37394,N_39523);
nor U42080 (N_42080,N_35765,N_37834);
nor U42081 (N_42081,N_35028,N_39110);
nor U42082 (N_42082,N_39181,N_37895);
xor U42083 (N_42083,N_36878,N_36645);
and U42084 (N_42084,N_39022,N_37362);
nor U42085 (N_42085,N_35916,N_38691);
or U42086 (N_42086,N_38515,N_36047);
nand U42087 (N_42087,N_36735,N_38374);
nand U42088 (N_42088,N_39783,N_35854);
xnor U42089 (N_42089,N_38565,N_36628);
nand U42090 (N_42090,N_37474,N_38977);
and U42091 (N_42091,N_38932,N_35656);
xnor U42092 (N_42092,N_36835,N_36940);
nand U42093 (N_42093,N_38239,N_39397);
and U42094 (N_42094,N_38916,N_39706);
or U42095 (N_42095,N_39403,N_37981);
xnor U42096 (N_42096,N_38351,N_37675);
or U42097 (N_42097,N_39698,N_37749);
nand U42098 (N_42098,N_37444,N_39846);
nand U42099 (N_42099,N_38272,N_35921);
nor U42100 (N_42100,N_37532,N_39851);
or U42101 (N_42101,N_36242,N_37620);
or U42102 (N_42102,N_37631,N_38623);
nor U42103 (N_42103,N_38110,N_36733);
xnor U42104 (N_42104,N_35562,N_38490);
nor U42105 (N_42105,N_35188,N_37696);
or U42106 (N_42106,N_36578,N_35101);
xor U42107 (N_42107,N_35328,N_38629);
nor U42108 (N_42108,N_38756,N_37709);
xor U42109 (N_42109,N_35897,N_38917);
or U42110 (N_42110,N_39408,N_37281);
nand U42111 (N_42111,N_36704,N_35056);
nor U42112 (N_42112,N_39130,N_39745);
or U42113 (N_42113,N_36279,N_36382);
xnor U42114 (N_42114,N_36841,N_37753);
nand U42115 (N_42115,N_37230,N_38296);
nor U42116 (N_42116,N_35089,N_35274);
nand U42117 (N_42117,N_37052,N_39567);
or U42118 (N_42118,N_35490,N_38838);
nand U42119 (N_42119,N_35425,N_35428);
nand U42120 (N_42120,N_36599,N_38654);
nand U42121 (N_42121,N_39176,N_38362);
and U42122 (N_42122,N_35397,N_36509);
nand U42123 (N_42123,N_38727,N_36880);
xor U42124 (N_42124,N_36369,N_35585);
xnor U42125 (N_42125,N_35751,N_38142);
nor U42126 (N_42126,N_37356,N_36224);
nand U42127 (N_42127,N_36205,N_36044);
nand U42128 (N_42128,N_37802,N_36011);
nand U42129 (N_42129,N_39512,N_36635);
xnor U42130 (N_42130,N_37132,N_36134);
nor U42131 (N_42131,N_35513,N_37454);
or U42132 (N_42132,N_38634,N_37875);
nor U42133 (N_42133,N_36761,N_38686);
nor U42134 (N_42134,N_36090,N_36440);
nor U42135 (N_42135,N_35219,N_37135);
or U42136 (N_42136,N_36790,N_37185);
nand U42137 (N_42137,N_39727,N_39223);
nor U42138 (N_42138,N_36807,N_39837);
nand U42139 (N_42139,N_36026,N_36448);
nand U42140 (N_42140,N_37245,N_36212);
or U42141 (N_42141,N_36782,N_39895);
nand U42142 (N_42142,N_39527,N_38608);
xor U42143 (N_42143,N_38020,N_37863);
xor U42144 (N_42144,N_36029,N_37706);
or U42145 (N_42145,N_35973,N_37928);
nand U42146 (N_42146,N_37370,N_39035);
and U42147 (N_42147,N_36372,N_38674);
nor U42148 (N_42148,N_36456,N_39520);
nand U42149 (N_42149,N_36544,N_37790);
xor U42150 (N_42150,N_35357,N_35499);
or U42151 (N_42151,N_35519,N_38248);
nor U42152 (N_42152,N_35148,N_37504);
and U42153 (N_42153,N_36607,N_36810);
nor U42154 (N_42154,N_36308,N_39616);
nand U42155 (N_42155,N_38093,N_37670);
or U42156 (N_42156,N_37565,N_35946);
nor U42157 (N_42157,N_38266,N_36261);
or U42158 (N_42158,N_35163,N_37223);
or U42159 (N_42159,N_39537,N_37509);
xnor U42160 (N_42160,N_35479,N_38063);
xnor U42161 (N_42161,N_35926,N_38131);
nand U42162 (N_42162,N_36415,N_37968);
xor U42163 (N_42163,N_35715,N_38868);
nor U42164 (N_42164,N_36399,N_39601);
or U42165 (N_42165,N_38386,N_37226);
nor U42166 (N_42166,N_36305,N_38665);
xnor U42167 (N_42167,N_38477,N_35837);
nand U42168 (N_42168,N_35032,N_39587);
and U42169 (N_42169,N_36427,N_38347);
or U42170 (N_42170,N_35781,N_36881);
nor U42171 (N_42171,N_38046,N_38287);
or U42172 (N_42172,N_38892,N_38843);
nand U42173 (N_42173,N_35734,N_37218);
and U42174 (N_42174,N_36804,N_35610);
or U42175 (N_42175,N_36417,N_35621);
or U42176 (N_42176,N_37017,N_37422);
nor U42177 (N_42177,N_38242,N_35414);
xor U42178 (N_42178,N_36655,N_37814);
nand U42179 (N_42179,N_37144,N_36819);
xor U42180 (N_42180,N_36094,N_37008);
nand U42181 (N_42181,N_35769,N_39210);
and U42182 (N_42182,N_35779,N_35096);
xor U42183 (N_42183,N_38100,N_39242);
or U42184 (N_42184,N_39808,N_35721);
nor U42185 (N_42185,N_37856,N_39286);
or U42186 (N_42186,N_36003,N_37127);
and U42187 (N_42187,N_37064,N_36500);
or U42188 (N_42188,N_36524,N_36852);
nor U42189 (N_42189,N_37938,N_38439);
nand U42190 (N_42190,N_39643,N_39126);
nand U42191 (N_42191,N_36006,N_35136);
nand U42192 (N_42192,N_39607,N_35725);
or U42193 (N_42193,N_35450,N_36173);
nor U42194 (N_42194,N_35292,N_36229);
nor U42195 (N_42195,N_36016,N_35037);
and U42196 (N_42196,N_35642,N_37330);
or U42197 (N_42197,N_36312,N_38465);
nor U42198 (N_42198,N_38511,N_38309);
and U42199 (N_42199,N_39576,N_36960);
or U42200 (N_42200,N_37891,N_37943);
nand U42201 (N_42201,N_35090,N_38799);
and U42202 (N_42202,N_38378,N_37138);
and U42203 (N_42203,N_37644,N_35097);
or U42204 (N_42204,N_39492,N_39470);
nand U42205 (N_42205,N_38149,N_37894);
and U42206 (N_42206,N_38560,N_37110);
and U42207 (N_42207,N_39046,N_35993);
nor U42208 (N_42208,N_39968,N_37984);
nor U42209 (N_42209,N_39062,N_36722);
nor U42210 (N_42210,N_36085,N_39834);
nand U42211 (N_42211,N_37167,N_35589);
nor U42212 (N_42212,N_36718,N_38299);
nand U42213 (N_42213,N_38276,N_37990);
nor U42214 (N_42214,N_36650,N_36617);
xnor U42215 (N_42215,N_36692,N_35293);
nor U42216 (N_42216,N_37472,N_39380);
or U42217 (N_42217,N_35403,N_35193);
nor U42218 (N_42218,N_38684,N_38122);
xor U42219 (N_42219,N_35141,N_35905);
and U42220 (N_42220,N_38785,N_37215);
and U42221 (N_42221,N_36387,N_35319);
nand U42222 (N_42222,N_36726,N_39812);
nand U42223 (N_42223,N_38627,N_38188);
xor U42224 (N_42224,N_38588,N_35803);
and U42225 (N_42225,N_37651,N_36175);
nor U42226 (N_42226,N_39648,N_39136);
nand U42227 (N_42227,N_39981,N_35841);
xor U42228 (N_42228,N_35382,N_38385);
or U42229 (N_42229,N_39212,N_36508);
and U42230 (N_42230,N_38617,N_36367);
nor U42231 (N_42231,N_35458,N_36475);
and U42232 (N_42232,N_39364,N_37887);
xnor U42233 (N_42233,N_38918,N_38224);
or U42234 (N_42234,N_37274,N_39163);
and U42235 (N_42235,N_38064,N_37961);
xor U42236 (N_42236,N_39373,N_39896);
and U42237 (N_42237,N_35012,N_37217);
xor U42238 (N_42238,N_39023,N_37244);
nor U42239 (N_42239,N_38532,N_39854);
and U42240 (N_42240,N_36161,N_36611);
xnor U42241 (N_42241,N_39931,N_36120);
nor U42242 (N_42242,N_38481,N_36139);
nor U42243 (N_42243,N_36972,N_35558);
nand U42244 (N_42244,N_37374,N_36014);
or U42245 (N_42245,N_38883,N_36663);
xnor U42246 (N_42246,N_37329,N_36896);
nor U42247 (N_42247,N_39757,N_36927);
xor U42248 (N_42248,N_37745,N_35348);
and U42249 (N_42249,N_35226,N_36989);
or U42250 (N_42250,N_39940,N_35654);
nand U42251 (N_42251,N_38782,N_36431);
and U42252 (N_42252,N_36787,N_37771);
or U42253 (N_42253,N_35234,N_35044);
xnor U42254 (N_42254,N_36112,N_39651);
or U42255 (N_42255,N_39639,N_38741);
xor U42256 (N_42256,N_36463,N_35570);
nand U42257 (N_42257,N_35196,N_39180);
and U42258 (N_42258,N_37188,N_37613);
or U42259 (N_42259,N_38117,N_37634);
or U42260 (N_42260,N_39097,N_36468);
and U42261 (N_42261,N_39849,N_38420);
nor U42262 (N_42262,N_36185,N_38899);
nor U42263 (N_42263,N_39988,N_36559);
xnor U42264 (N_42264,N_38186,N_35746);
and U42265 (N_42265,N_35055,N_35433);
xor U42266 (N_42266,N_35313,N_36439);
or U42267 (N_42267,N_37535,N_37053);
and U42268 (N_42268,N_39038,N_36013);
and U42269 (N_42269,N_39270,N_37259);
or U42270 (N_42270,N_37293,N_35666);
nand U42271 (N_42271,N_38697,N_35495);
and U42272 (N_42272,N_39800,N_36906);
xor U42273 (N_42273,N_38625,N_37355);
nand U42274 (N_42274,N_35105,N_38135);
nand U42275 (N_42275,N_36373,N_36170);
xor U42276 (N_42276,N_38828,N_35859);
nand U42277 (N_42277,N_35336,N_39260);
nor U42278 (N_42278,N_38442,N_37216);
nand U42279 (N_42279,N_35166,N_36122);
or U42280 (N_42280,N_39091,N_39352);
and U42281 (N_42281,N_36970,N_39918);
nor U42282 (N_42282,N_36348,N_38814);
and U42283 (N_42283,N_39433,N_35430);
or U42284 (N_42284,N_38953,N_36548);
xnor U42285 (N_42285,N_36043,N_35533);
nand U42286 (N_42286,N_38039,N_38516);
or U42287 (N_42287,N_37674,N_35882);
xor U42288 (N_42288,N_37148,N_37849);
and U42289 (N_42289,N_39277,N_38825);
nand U42290 (N_42290,N_38045,N_35939);
nor U42291 (N_42291,N_36661,N_35820);
and U42292 (N_42292,N_37271,N_37668);
nand U42293 (N_42293,N_38742,N_38021);
or U42294 (N_42294,N_35982,N_35526);
nand U42295 (N_42295,N_38680,N_37624);
nor U42296 (N_42296,N_39875,N_37945);
and U42297 (N_42297,N_36476,N_35817);
or U42298 (N_42298,N_37647,N_36777);
nand U42299 (N_42299,N_36922,N_36447);
nor U42300 (N_42300,N_39730,N_35620);
xnor U42301 (N_42301,N_37480,N_39853);
or U42302 (N_42302,N_39109,N_36570);
nand U42303 (N_42303,N_38572,N_36340);
or U42304 (N_42304,N_36930,N_36842);
or U42305 (N_42305,N_38689,N_36007);
nor U42306 (N_42306,N_38350,N_37263);
nand U42307 (N_42307,N_35550,N_36228);
or U42308 (N_42308,N_36715,N_38926);
or U42309 (N_42309,N_35359,N_35186);
nor U42310 (N_42310,N_35455,N_35212);
nand U42311 (N_42311,N_38183,N_37073);
xor U42312 (N_42312,N_35154,N_36392);
xnor U42313 (N_42313,N_39080,N_37995);
nor U42314 (N_42314,N_39822,N_35192);
xor U42315 (N_42315,N_39221,N_38082);
and U42316 (N_42316,N_36258,N_37868);
and U42317 (N_42317,N_39574,N_35138);
xor U42318 (N_42318,N_35582,N_39920);
nand U42319 (N_42319,N_38887,N_37831);
nand U42320 (N_42320,N_39677,N_37457);
and U42321 (N_42321,N_37049,N_37333);
nor U42322 (N_42322,N_39962,N_39477);
xor U42323 (N_42323,N_35343,N_36809);
or U42324 (N_42324,N_35308,N_37111);
xnor U42325 (N_42325,N_36720,N_39396);
and U42326 (N_42326,N_39684,N_39471);
nand U42327 (N_42327,N_35124,N_36990);
and U42328 (N_42328,N_37026,N_38594);
nor U42329 (N_42329,N_38087,N_36909);
xor U42330 (N_42330,N_37385,N_35500);
or U42331 (N_42331,N_37399,N_38460);
and U42332 (N_42332,N_36571,N_37915);
nor U42333 (N_42333,N_37087,N_39675);
xor U42334 (N_42334,N_36750,N_37173);
and U42335 (N_42335,N_36300,N_36552);
or U42336 (N_42336,N_38600,N_38769);
and U42337 (N_42337,N_37669,N_38418);
or U42338 (N_42338,N_38447,N_36555);
xor U42339 (N_42339,N_38539,N_38734);
or U42340 (N_42340,N_35351,N_39187);
nor U42341 (N_42341,N_37306,N_39658);
nor U42342 (N_42342,N_37626,N_37308);
nand U42343 (N_42343,N_39551,N_35813);
nor U42344 (N_42344,N_38614,N_38613);
nor U42345 (N_42345,N_36792,N_35421);
and U42346 (N_42346,N_35325,N_39291);
nor U42347 (N_42347,N_35890,N_35724);
xor U42348 (N_42348,N_36428,N_37531);
and U42349 (N_42349,N_35294,N_37383);
nand U42350 (N_42350,N_38806,N_35338);
or U42351 (N_42351,N_37809,N_39228);
nand U42352 (N_42352,N_35361,N_39231);
or U42353 (N_42353,N_39756,N_38211);
or U42354 (N_42354,N_35297,N_35111);
and U42355 (N_42355,N_35477,N_38605);
nand U42356 (N_42356,N_35024,N_36780);
xnor U42357 (N_42357,N_38889,N_35774);
nand U42358 (N_42358,N_38197,N_35062);
and U42359 (N_42359,N_38129,N_39055);
and U42360 (N_42360,N_37124,N_39069);
nand U42361 (N_42361,N_35086,N_37870);
or U42362 (N_42362,N_35792,N_39161);
and U42363 (N_42363,N_39304,N_38191);
or U42364 (N_42364,N_37413,N_37305);
or U42365 (N_42365,N_39294,N_36375);
and U42366 (N_42366,N_37000,N_35218);
nor U42367 (N_42367,N_39234,N_39632);
or U42368 (N_42368,N_38026,N_39255);
and U42369 (N_42369,N_39165,N_36193);
xor U42370 (N_42370,N_35740,N_36184);
xor U42371 (N_42371,N_39948,N_38232);
nor U42372 (N_42372,N_39168,N_35243);
nor U42373 (N_42373,N_36716,N_36796);
or U42374 (N_42374,N_37805,N_37056);
xnor U42375 (N_42375,N_39266,N_37396);
nor U42376 (N_42376,N_39737,N_37750);
nor U42377 (N_42377,N_37172,N_37885);
nand U42378 (N_42378,N_36379,N_36222);
xor U42379 (N_42379,N_38989,N_37804);
nand U42380 (N_42380,N_38409,N_39979);
nand U42381 (N_42381,N_36753,N_35906);
xor U42382 (N_42382,N_36968,N_37425);
nand U42383 (N_42383,N_38993,N_35473);
and U42384 (N_42384,N_37469,N_36923);
xnor U42385 (N_42385,N_38518,N_39749);
or U42386 (N_42386,N_37796,N_39457);
xnor U42387 (N_42387,N_39728,N_36214);
nor U42388 (N_42388,N_39718,N_35737);
and U42389 (N_42389,N_36775,N_36425);
or U42390 (N_42390,N_35777,N_35857);
nand U42391 (N_42391,N_37662,N_36114);
xor U42392 (N_42392,N_35955,N_35614);
nor U42393 (N_42393,N_35785,N_35287);
or U42394 (N_42394,N_38141,N_39499);
and U42395 (N_42395,N_37726,N_39726);
nor U42396 (N_42396,N_35349,N_36446);
or U42397 (N_42397,N_39507,N_39441);
nand U42398 (N_42398,N_35158,N_39133);
nor U42399 (N_42399,N_36658,N_39802);
xor U42400 (N_42400,N_38717,N_38236);
and U42401 (N_42401,N_38273,N_38079);
and U42402 (N_42402,N_35957,N_37447);
nor U42403 (N_42403,N_35927,N_39068);
nor U42404 (N_42404,N_39888,N_37250);
xor U42405 (N_42405,N_36239,N_36292);
xor U42406 (N_42406,N_38240,N_36892);
nand U42407 (N_42407,N_39476,N_35869);
xnor U42408 (N_42408,N_39526,N_36996);
nand U42409 (N_42409,N_35577,N_35323);
xor U42410 (N_42410,N_37580,N_37003);
or U42411 (N_42411,N_36067,N_38174);
nor U42412 (N_42412,N_36823,N_39861);
nor U42413 (N_42413,N_35464,N_39467);
xnor U42414 (N_42414,N_39085,N_37987);
nor U42415 (N_42415,N_38584,N_35908);
xor U42416 (N_42416,N_38108,N_37160);
and U42417 (N_42417,N_39654,N_36814);
and U42418 (N_42418,N_35104,N_38097);
and U42419 (N_42419,N_35259,N_36365);
nand U42420 (N_42420,N_35814,N_39066);
or U42421 (N_42421,N_36314,N_39184);
nor U42422 (N_42422,N_39292,N_35459);
nand U42423 (N_42423,N_36198,N_35036);
or U42424 (N_42424,N_38954,N_36149);
and U42425 (N_42425,N_35369,N_37920);
nor U42426 (N_42426,N_38163,N_36958);
or U42427 (N_42427,N_38332,N_37302);
nand U42428 (N_42428,N_37655,N_39825);
and U42429 (N_42429,N_37015,N_35764);
and U42430 (N_42430,N_35747,N_38529);
xor U42431 (N_42431,N_37807,N_38404);
and U42432 (N_42432,N_36093,N_38394);
nor U42433 (N_42433,N_39647,N_38670);
or U42434 (N_42434,N_38911,N_37361);
or U42435 (N_42435,N_37871,N_35295);
xor U42436 (N_42436,N_35739,N_35010);
and U42437 (N_42437,N_35555,N_35113);
or U42438 (N_42438,N_36813,N_35704);
nor U42439 (N_42439,N_39183,N_38514);
or U42440 (N_42440,N_35625,N_39236);
or U42441 (N_42441,N_39555,N_36554);
xor U42442 (N_42442,N_39501,N_39039);
nand U42443 (N_42443,N_35404,N_35203);
nand U42444 (N_42444,N_38999,N_37847);
xor U42445 (N_42445,N_37878,N_39349);
and U42446 (N_42446,N_35531,N_39750);
xor U42447 (N_42447,N_37503,N_39505);
or U42448 (N_42448,N_37972,N_36640);
or U42449 (N_42449,N_39890,N_35842);
nor U42450 (N_42450,N_36625,N_37093);
and U42451 (N_42451,N_35080,N_39832);
or U42452 (N_42452,N_38075,N_38375);
nor U42453 (N_42453,N_36315,N_39280);
or U42454 (N_42454,N_37763,N_35694);
nor U42455 (N_42455,N_39848,N_35673);
nand U42456 (N_42456,N_36030,N_38821);
xnor U42457 (N_42457,N_38706,N_35618);
and U42458 (N_42458,N_38044,N_37544);
nand U42459 (N_42459,N_39435,N_38241);
or U42460 (N_42460,N_37989,N_38726);
nor U42461 (N_42461,N_39905,N_36592);
xor U42462 (N_42462,N_38754,N_39057);
or U42463 (N_42463,N_39063,N_36472);
nor U42464 (N_42464,N_35197,N_35685);
or U42465 (N_42465,N_37344,N_38343);
or U42466 (N_42466,N_35895,N_39440);
or U42467 (N_42467,N_39671,N_36101);
and U42468 (N_42468,N_36207,N_38229);
nand U42469 (N_42469,N_39877,N_36727);
and U42470 (N_42470,N_37069,N_35108);
xnor U42471 (N_42471,N_37309,N_39498);
nand U42472 (N_42472,N_37461,N_39927);
xor U42473 (N_42473,N_37169,N_38023);
xor U42474 (N_42474,N_37097,N_36341);
or U42475 (N_42475,N_39302,N_39095);
nor U42476 (N_42476,N_36460,N_36589);
and U42477 (N_42477,N_36734,N_37514);
and U42478 (N_42478,N_36444,N_35934);
and U42479 (N_42479,N_38835,N_38153);
nand U42480 (N_42480,N_37869,N_39283);
nor U42481 (N_42481,N_35752,N_36963);
and U42482 (N_42482,N_37225,N_39478);
nand U42483 (N_42483,N_38161,N_35709);
nor U42484 (N_42484,N_39558,N_39946);
and U42485 (N_42485,N_39400,N_36489);
xor U42486 (N_42486,N_39679,N_35844);
xnor U42487 (N_42487,N_38441,N_36520);
nand U42488 (N_42488,N_36336,N_35612);
nand U42489 (N_42489,N_36467,N_36000);
and U42490 (N_42490,N_37359,N_37178);
or U42491 (N_42491,N_37707,N_36877);
or U42492 (N_42492,N_38187,N_36245);
or U42493 (N_42493,N_37335,N_35755);
nand U42494 (N_42494,N_36195,N_39225);
nor U42495 (N_42495,N_35107,N_38218);
and U42496 (N_42496,N_39934,N_37321);
and U42497 (N_42497,N_39721,N_39029);
xnor U42498 (N_42498,N_39450,N_35675);
and U42499 (N_42499,N_36591,N_35371);
nand U42500 (N_42500,N_38512,N_39987);
and U42501 (N_42501,N_39278,N_39577);
nor U42502 (N_42502,N_38670,N_38892);
nor U42503 (N_42503,N_36401,N_35256);
nor U42504 (N_42504,N_35356,N_37635);
or U42505 (N_42505,N_37362,N_35555);
and U42506 (N_42506,N_35178,N_37790);
nand U42507 (N_42507,N_37533,N_36042);
xnor U42508 (N_42508,N_35859,N_36431);
xnor U42509 (N_42509,N_35370,N_39347);
nor U42510 (N_42510,N_35344,N_37394);
nand U42511 (N_42511,N_36097,N_38363);
and U42512 (N_42512,N_35161,N_36651);
xnor U42513 (N_42513,N_38127,N_39905);
xor U42514 (N_42514,N_35364,N_37576);
or U42515 (N_42515,N_36672,N_37457);
nor U42516 (N_42516,N_39603,N_39670);
xnor U42517 (N_42517,N_39508,N_36288);
nor U42518 (N_42518,N_39153,N_39967);
and U42519 (N_42519,N_39398,N_37645);
nor U42520 (N_42520,N_39093,N_36743);
xnor U42521 (N_42521,N_37852,N_36984);
and U42522 (N_42522,N_39574,N_39034);
nor U42523 (N_42523,N_36320,N_39581);
nor U42524 (N_42524,N_35132,N_37108);
or U42525 (N_42525,N_35349,N_36172);
xnor U42526 (N_42526,N_36129,N_36239);
nand U42527 (N_42527,N_35205,N_36160);
or U42528 (N_42528,N_38578,N_36746);
and U42529 (N_42529,N_38608,N_38410);
nand U42530 (N_42530,N_38669,N_35061);
xnor U42531 (N_42531,N_36931,N_36180);
and U42532 (N_42532,N_37424,N_37957);
and U42533 (N_42533,N_36562,N_37647);
and U42534 (N_42534,N_37556,N_35490);
and U42535 (N_42535,N_39044,N_36229);
xnor U42536 (N_42536,N_35309,N_35850);
nand U42537 (N_42537,N_36251,N_35244);
xnor U42538 (N_42538,N_36646,N_38414);
or U42539 (N_42539,N_36644,N_39969);
and U42540 (N_42540,N_37329,N_35121);
xnor U42541 (N_42541,N_36822,N_36789);
xor U42542 (N_42542,N_39914,N_36975);
or U42543 (N_42543,N_36539,N_37778);
nor U42544 (N_42544,N_39991,N_38454);
nand U42545 (N_42545,N_36191,N_35873);
xnor U42546 (N_42546,N_38086,N_39021);
and U42547 (N_42547,N_38754,N_38766);
or U42548 (N_42548,N_37545,N_35079);
nor U42549 (N_42549,N_35942,N_39151);
nand U42550 (N_42550,N_36778,N_39189);
nor U42551 (N_42551,N_37826,N_35004);
or U42552 (N_42552,N_38685,N_35155);
xor U42553 (N_42553,N_38763,N_39617);
and U42554 (N_42554,N_37978,N_35203);
and U42555 (N_42555,N_36721,N_36802);
xor U42556 (N_42556,N_36124,N_39242);
and U42557 (N_42557,N_35214,N_37500);
or U42558 (N_42558,N_35658,N_36306);
nand U42559 (N_42559,N_36914,N_36131);
nand U42560 (N_42560,N_38309,N_35241);
or U42561 (N_42561,N_35967,N_35641);
or U42562 (N_42562,N_38983,N_37881);
or U42563 (N_42563,N_37901,N_39458);
xor U42564 (N_42564,N_35220,N_35924);
or U42565 (N_42565,N_37051,N_39568);
nand U42566 (N_42566,N_38522,N_38436);
nand U42567 (N_42567,N_35113,N_37077);
xnor U42568 (N_42568,N_38970,N_38167);
or U42569 (N_42569,N_36018,N_37687);
nor U42570 (N_42570,N_35944,N_35127);
and U42571 (N_42571,N_39420,N_36185);
nand U42572 (N_42572,N_37136,N_37929);
xor U42573 (N_42573,N_39499,N_39994);
xor U42574 (N_42574,N_37528,N_35972);
nand U42575 (N_42575,N_36512,N_37539);
xor U42576 (N_42576,N_35565,N_37321);
nand U42577 (N_42577,N_36157,N_37213);
nand U42578 (N_42578,N_35910,N_38221);
or U42579 (N_42579,N_35141,N_37676);
or U42580 (N_42580,N_36072,N_39500);
nand U42581 (N_42581,N_37785,N_38551);
nor U42582 (N_42582,N_39728,N_37087);
or U42583 (N_42583,N_37926,N_35609);
or U42584 (N_42584,N_35447,N_36068);
and U42585 (N_42585,N_36967,N_38983);
nand U42586 (N_42586,N_39627,N_39476);
and U42587 (N_42587,N_37118,N_36604);
nand U42588 (N_42588,N_37960,N_38417);
or U42589 (N_42589,N_38042,N_35407);
xnor U42590 (N_42590,N_37810,N_38019);
and U42591 (N_42591,N_38506,N_37205);
xor U42592 (N_42592,N_38730,N_39422);
xor U42593 (N_42593,N_35091,N_37827);
xor U42594 (N_42594,N_37741,N_39020);
and U42595 (N_42595,N_39953,N_36265);
nand U42596 (N_42596,N_35215,N_35660);
or U42597 (N_42597,N_36225,N_38226);
xor U42598 (N_42598,N_38717,N_37740);
nor U42599 (N_42599,N_36432,N_39446);
and U42600 (N_42600,N_37810,N_37993);
nor U42601 (N_42601,N_36153,N_36986);
xnor U42602 (N_42602,N_36480,N_36530);
nor U42603 (N_42603,N_37784,N_36947);
and U42604 (N_42604,N_35506,N_36344);
and U42605 (N_42605,N_36887,N_35493);
nor U42606 (N_42606,N_39725,N_35746);
nand U42607 (N_42607,N_36949,N_36263);
nor U42608 (N_42608,N_38852,N_37016);
nand U42609 (N_42609,N_38810,N_37974);
xor U42610 (N_42610,N_36421,N_35704);
or U42611 (N_42611,N_37194,N_37640);
nand U42612 (N_42612,N_37842,N_37280);
and U42613 (N_42613,N_38019,N_36943);
or U42614 (N_42614,N_38661,N_36515);
nand U42615 (N_42615,N_35756,N_35343);
nor U42616 (N_42616,N_36742,N_39115);
nand U42617 (N_42617,N_37126,N_37201);
nand U42618 (N_42618,N_38087,N_36412);
xnor U42619 (N_42619,N_36254,N_36985);
or U42620 (N_42620,N_37551,N_37507);
nor U42621 (N_42621,N_39364,N_36050);
or U42622 (N_42622,N_35596,N_39387);
and U42623 (N_42623,N_38201,N_37782);
and U42624 (N_42624,N_39413,N_38103);
or U42625 (N_42625,N_39428,N_36372);
nor U42626 (N_42626,N_37952,N_35066);
or U42627 (N_42627,N_39795,N_39357);
or U42628 (N_42628,N_39967,N_39646);
nand U42629 (N_42629,N_37281,N_35960);
xnor U42630 (N_42630,N_37587,N_35802);
nand U42631 (N_42631,N_37118,N_38921);
and U42632 (N_42632,N_37512,N_38856);
nand U42633 (N_42633,N_35251,N_36709);
nand U42634 (N_42634,N_38821,N_39412);
and U42635 (N_42635,N_35539,N_35688);
or U42636 (N_42636,N_35989,N_38434);
nor U42637 (N_42637,N_36371,N_39262);
or U42638 (N_42638,N_36708,N_36004);
xnor U42639 (N_42639,N_37527,N_38209);
or U42640 (N_42640,N_35816,N_37511);
and U42641 (N_42641,N_37580,N_36509);
xnor U42642 (N_42642,N_37502,N_36548);
nor U42643 (N_42643,N_38402,N_37765);
and U42644 (N_42644,N_35631,N_36946);
nor U42645 (N_42645,N_35622,N_38388);
nor U42646 (N_42646,N_36471,N_38233);
and U42647 (N_42647,N_37656,N_39589);
or U42648 (N_42648,N_37053,N_39839);
nor U42649 (N_42649,N_36876,N_38407);
nor U42650 (N_42650,N_37398,N_35816);
nor U42651 (N_42651,N_39246,N_36364);
nand U42652 (N_42652,N_39571,N_39971);
nand U42653 (N_42653,N_35202,N_36346);
xnor U42654 (N_42654,N_35527,N_36816);
nand U42655 (N_42655,N_39820,N_35385);
or U42656 (N_42656,N_39539,N_38611);
and U42657 (N_42657,N_35345,N_39874);
xor U42658 (N_42658,N_39260,N_39870);
xnor U42659 (N_42659,N_35262,N_39047);
nor U42660 (N_42660,N_35753,N_35042);
nand U42661 (N_42661,N_37247,N_35641);
nand U42662 (N_42662,N_35762,N_37914);
xnor U42663 (N_42663,N_37158,N_39183);
nor U42664 (N_42664,N_39362,N_36773);
nand U42665 (N_42665,N_35379,N_36148);
and U42666 (N_42666,N_38264,N_36496);
nor U42667 (N_42667,N_38409,N_36424);
nor U42668 (N_42668,N_35792,N_39411);
nor U42669 (N_42669,N_36113,N_39450);
or U42670 (N_42670,N_36497,N_37564);
nor U42671 (N_42671,N_37225,N_36340);
and U42672 (N_42672,N_39080,N_38122);
or U42673 (N_42673,N_36965,N_39510);
nand U42674 (N_42674,N_35644,N_38712);
nor U42675 (N_42675,N_37009,N_36143);
and U42676 (N_42676,N_36658,N_38193);
and U42677 (N_42677,N_38816,N_37821);
and U42678 (N_42678,N_39211,N_36566);
nand U42679 (N_42679,N_35644,N_37349);
nand U42680 (N_42680,N_39713,N_36164);
nor U42681 (N_42681,N_38868,N_35975);
or U42682 (N_42682,N_35838,N_37475);
xnor U42683 (N_42683,N_36202,N_35275);
nand U42684 (N_42684,N_35842,N_36207);
nand U42685 (N_42685,N_36850,N_35051);
xor U42686 (N_42686,N_35463,N_39660);
nand U42687 (N_42687,N_38349,N_37958);
xor U42688 (N_42688,N_35261,N_39839);
nor U42689 (N_42689,N_38821,N_38945);
xnor U42690 (N_42690,N_38868,N_38133);
or U42691 (N_42691,N_35828,N_35131);
nor U42692 (N_42692,N_37792,N_39329);
or U42693 (N_42693,N_39129,N_35522);
xnor U42694 (N_42694,N_38967,N_35918);
nand U42695 (N_42695,N_39200,N_35529);
and U42696 (N_42696,N_37752,N_35870);
or U42697 (N_42697,N_36026,N_37613);
nand U42698 (N_42698,N_39999,N_35204);
nand U42699 (N_42699,N_39073,N_36048);
nand U42700 (N_42700,N_39613,N_36734);
nor U42701 (N_42701,N_39557,N_39211);
or U42702 (N_42702,N_39014,N_36556);
or U42703 (N_42703,N_39754,N_37120);
and U42704 (N_42704,N_36861,N_37244);
or U42705 (N_42705,N_36169,N_36987);
or U42706 (N_42706,N_38273,N_35464);
xnor U42707 (N_42707,N_37240,N_38628);
nor U42708 (N_42708,N_38219,N_35797);
nor U42709 (N_42709,N_39144,N_38982);
and U42710 (N_42710,N_35089,N_39607);
and U42711 (N_42711,N_38218,N_36878);
and U42712 (N_42712,N_35411,N_36952);
nand U42713 (N_42713,N_35743,N_37985);
nor U42714 (N_42714,N_38541,N_38156);
nor U42715 (N_42715,N_35560,N_39351);
and U42716 (N_42716,N_38796,N_37495);
nor U42717 (N_42717,N_35745,N_36053);
and U42718 (N_42718,N_35186,N_35005);
nor U42719 (N_42719,N_39981,N_39294);
xnor U42720 (N_42720,N_38642,N_37217);
nand U42721 (N_42721,N_35124,N_38279);
xnor U42722 (N_42722,N_36295,N_38604);
or U42723 (N_42723,N_39963,N_36986);
xor U42724 (N_42724,N_39181,N_36604);
nand U42725 (N_42725,N_38771,N_38397);
xor U42726 (N_42726,N_37635,N_38284);
xnor U42727 (N_42727,N_38777,N_35943);
xnor U42728 (N_42728,N_38540,N_36691);
xnor U42729 (N_42729,N_39245,N_39391);
xor U42730 (N_42730,N_36446,N_37429);
and U42731 (N_42731,N_38885,N_36486);
and U42732 (N_42732,N_36950,N_39557);
nor U42733 (N_42733,N_37320,N_37975);
or U42734 (N_42734,N_37832,N_35142);
xor U42735 (N_42735,N_36380,N_39639);
nor U42736 (N_42736,N_37627,N_38911);
nor U42737 (N_42737,N_35160,N_35706);
or U42738 (N_42738,N_36298,N_36389);
and U42739 (N_42739,N_35867,N_36146);
xnor U42740 (N_42740,N_37144,N_37807);
xnor U42741 (N_42741,N_36471,N_38074);
nor U42742 (N_42742,N_36138,N_39832);
nor U42743 (N_42743,N_37618,N_37200);
or U42744 (N_42744,N_38695,N_38936);
nand U42745 (N_42745,N_39362,N_38072);
nand U42746 (N_42746,N_36857,N_35149);
and U42747 (N_42747,N_39806,N_38356);
xor U42748 (N_42748,N_39412,N_35032);
and U42749 (N_42749,N_36118,N_37697);
nand U42750 (N_42750,N_37940,N_36414);
or U42751 (N_42751,N_38125,N_36406);
and U42752 (N_42752,N_37563,N_38846);
nand U42753 (N_42753,N_37966,N_35070);
xnor U42754 (N_42754,N_36583,N_39387);
or U42755 (N_42755,N_39777,N_37377);
and U42756 (N_42756,N_37819,N_37380);
nor U42757 (N_42757,N_35456,N_36032);
and U42758 (N_42758,N_36869,N_36382);
and U42759 (N_42759,N_38878,N_35001);
or U42760 (N_42760,N_35498,N_35097);
or U42761 (N_42761,N_35760,N_35998);
nor U42762 (N_42762,N_38691,N_37782);
and U42763 (N_42763,N_35784,N_39921);
nand U42764 (N_42764,N_38033,N_36495);
and U42765 (N_42765,N_35874,N_37565);
or U42766 (N_42766,N_35175,N_36116);
or U42767 (N_42767,N_35075,N_35169);
or U42768 (N_42768,N_35773,N_35880);
and U42769 (N_42769,N_37464,N_36452);
nor U42770 (N_42770,N_38764,N_39798);
xor U42771 (N_42771,N_35153,N_37957);
nand U42772 (N_42772,N_38250,N_35153);
nand U42773 (N_42773,N_39748,N_36690);
xnor U42774 (N_42774,N_35377,N_39118);
and U42775 (N_42775,N_37987,N_35383);
and U42776 (N_42776,N_35747,N_35450);
and U42777 (N_42777,N_38715,N_36338);
nand U42778 (N_42778,N_36332,N_38828);
and U42779 (N_42779,N_37038,N_38253);
and U42780 (N_42780,N_38269,N_35031);
or U42781 (N_42781,N_35424,N_35978);
nor U42782 (N_42782,N_35829,N_36577);
or U42783 (N_42783,N_38011,N_38465);
nand U42784 (N_42784,N_38068,N_39573);
nor U42785 (N_42785,N_38460,N_38412);
or U42786 (N_42786,N_37382,N_39670);
nor U42787 (N_42787,N_37302,N_38002);
xor U42788 (N_42788,N_35217,N_36916);
nand U42789 (N_42789,N_35511,N_35671);
xnor U42790 (N_42790,N_38338,N_37086);
or U42791 (N_42791,N_37816,N_38731);
and U42792 (N_42792,N_39873,N_39556);
or U42793 (N_42793,N_38721,N_37941);
xor U42794 (N_42794,N_36549,N_38903);
and U42795 (N_42795,N_37765,N_38339);
and U42796 (N_42796,N_35916,N_39480);
xnor U42797 (N_42797,N_39308,N_36449);
nor U42798 (N_42798,N_39144,N_35512);
xor U42799 (N_42799,N_36573,N_35671);
nand U42800 (N_42800,N_39190,N_36633);
nand U42801 (N_42801,N_38909,N_35033);
xnor U42802 (N_42802,N_36554,N_38833);
xor U42803 (N_42803,N_36138,N_35439);
nand U42804 (N_42804,N_35892,N_38407);
or U42805 (N_42805,N_36747,N_35678);
xor U42806 (N_42806,N_39337,N_39991);
nor U42807 (N_42807,N_39727,N_39123);
nand U42808 (N_42808,N_39403,N_37190);
nand U42809 (N_42809,N_35055,N_35396);
and U42810 (N_42810,N_39284,N_36773);
nand U42811 (N_42811,N_36630,N_36691);
and U42812 (N_42812,N_38827,N_38339);
nand U42813 (N_42813,N_36050,N_35314);
nor U42814 (N_42814,N_37864,N_36825);
nand U42815 (N_42815,N_37382,N_36657);
xnor U42816 (N_42816,N_39553,N_35360);
xnor U42817 (N_42817,N_35792,N_35021);
nor U42818 (N_42818,N_36260,N_39764);
and U42819 (N_42819,N_38347,N_37987);
or U42820 (N_42820,N_35566,N_39721);
nand U42821 (N_42821,N_37808,N_39459);
nand U42822 (N_42822,N_36809,N_39352);
nor U42823 (N_42823,N_38289,N_37078);
or U42824 (N_42824,N_35058,N_39009);
xnor U42825 (N_42825,N_39688,N_39635);
or U42826 (N_42826,N_37560,N_36711);
and U42827 (N_42827,N_39261,N_35848);
nor U42828 (N_42828,N_39734,N_37365);
xor U42829 (N_42829,N_39460,N_37665);
xnor U42830 (N_42830,N_35696,N_35847);
xnor U42831 (N_42831,N_39037,N_39205);
xor U42832 (N_42832,N_39054,N_35583);
nor U42833 (N_42833,N_36000,N_38191);
nand U42834 (N_42834,N_37307,N_37106);
and U42835 (N_42835,N_37363,N_36177);
nand U42836 (N_42836,N_39421,N_36675);
xnor U42837 (N_42837,N_39542,N_37687);
and U42838 (N_42838,N_36209,N_39774);
and U42839 (N_42839,N_39443,N_36511);
xor U42840 (N_42840,N_36698,N_36922);
or U42841 (N_42841,N_36201,N_39360);
nor U42842 (N_42842,N_39732,N_39268);
or U42843 (N_42843,N_36573,N_38816);
xor U42844 (N_42844,N_39725,N_36532);
xnor U42845 (N_42845,N_36340,N_36313);
and U42846 (N_42846,N_39719,N_35659);
xnor U42847 (N_42847,N_36802,N_35912);
nand U42848 (N_42848,N_36068,N_39101);
or U42849 (N_42849,N_35324,N_35645);
nand U42850 (N_42850,N_36769,N_36170);
nand U42851 (N_42851,N_35326,N_38931);
and U42852 (N_42852,N_37432,N_38265);
nor U42853 (N_42853,N_38401,N_38604);
xnor U42854 (N_42854,N_38970,N_37900);
nand U42855 (N_42855,N_38493,N_37355);
xor U42856 (N_42856,N_37732,N_35791);
nand U42857 (N_42857,N_37298,N_39763);
nor U42858 (N_42858,N_36107,N_35073);
or U42859 (N_42859,N_39374,N_38349);
and U42860 (N_42860,N_38813,N_36147);
or U42861 (N_42861,N_35267,N_38732);
nand U42862 (N_42862,N_37256,N_39836);
and U42863 (N_42863,N_37733,N_38571);
nand U42864 (N_42864,N_37835,N_35524);
and U42865 (N_42865,N_39205,N_36764);
or U42866 (N_42866,N_37664,N_35641);
and U42867 (N_42867,N_38793,N_38130);
or U42868 (N_42868,N_38816,N_39685);
or U42869 (N_42869,N_36360,N_37135);
or U42870 (N_42870,N_37470,N_36323);
xnor U42871 (N_42871,N_38539,N_39760);
nor U42872 (N_42872,N_36016,N_35336);
nand U42873 (N_42873,N_36925,N_36184);
and U42874 (N_42874,N_35974,N_35521);
nor U42875 (N_42875,N_36691,N_37179);
xor U42876 (N_42876,N_38156,N_39300);
or U42877 (N_42877,N_36673,N_36450);
xor U42878 (N_42878,N_39157,N_35434);
or U42879 (N_42879,N_35332,N_37257);
nand U42880 (N_42880,N_38130,N_37298);
nor U42881 (N_42881,N_36360,N_39233);
nand U42882 (N_42882,N_35519,N_36130);
nor U42883 (N_42883,N_35488,N_35143);
nand U42884 (N_42884,N_36967,N_36472);
nand U42885 (N_42885,N_39564,N_37402);
nand U42886 (N_42886,N_37588,N_38178);
and U42887 (N_42887,N_38646,N_35592);
nand U42888 (N_42888,N_39042,N_36802);
nor U42889 (N_42889,N_35235,N_36868);
nand U42890 (N_42890,N_36367,N_37632);
or U42891 (N_42891,N_37789,N_38958);
or U42892 (N_42892,N_39093,N_36769);
or U42893 (N_42893,N_37255,N_38704);
nand U42894 (N_42894,N_39327,N_36512);
xnor U42895 (N_42895,N_37542,N_37098);
nand U42896 (N_42896,N_39174,N_36481);
or U42897 (N_42897,N_37313,N_37178);
nand U42898 (N_42898,N_37433,N_36159);
and U42899 (N_42899,N_37932,N_36850);
and U42900 (N_42900,N_37962,N_36609);
and U42901 (N_42901,N_35375,N_38444);
nand U42902 (N_42902,N_35205,N_37806);
nand U42903 (N_42903,N_37544,N_38299);
or U42904 (N_42904,N_39310,N_38059);
nor U42905 (N_42905,N_39038,N_35756);
and U42906 (N_42906,N_39399,N_36520);
nand U42907 (N_42907,N_37595,N_35762);
and U42908 (N_42908,N_37123,N_37507);
and U42909 (N_42909,N_35293,N_39963);
and U42910 (N_42910,N_35733,N_36695);
nand U42911 (N_42911,N_35588,N_39758);
nand U42912 (N_42912,N_36702,N_37674);
and U42913 (N_42913,N_36839,N_37113);
or U42914 (N_42914,N_35755,N_36261);
or U42915 (N_42915,N_39294,N_36246);
nor U42916 (N_42916,N_36031,N_37614);
nand U42917 (N_42917,N_37872,N_37707);
nand U42918 (N_42918,N_37712,N_35770);
nand U42919 (N_42919,N_37683,N_37915);
or U42920 (N_42920,N_37695,N_39638);
nand U42921 (N_42921,N_35490,N_36026);
nand U42922 (N_42922,N_35030,N_38295);
or U42923 (N_42923,N_39853,N_39938);
and U42924 (N_42924,N_37254,N_39255);
or U42925 (N_42925,N_36166,N_38901);
or U42926 (N_42926,N_35886,N_35821);
nor U42927 (N_42927,N_39520,N_36747);
nor U42928 (N_42928,N_37586,N_37516);
xor U42929 (N_42929,N_36234,N_39617);
and U42930 (N_42930,N_37899,N_36405);
nor U42931 (N_42931,N_35100,N_37397);
xor U42932 (N_42932,N_35280,N_37623);
and U42933 (N_42933,N_37348,N_35400);
nand U42934 (N_42934,N_36641,N_39383);
nand U42935 (N_42935,N_36313,N_36318);
xor U42936 (N_42936,N_35311,N_37228);
and U42937 (N_42937,N_38706,N_35387);
or U42938 (N_42938,N_35476,N_39708);
and U42939 (N_42939,N_35883,N_36621);
nor U42940 (N_42940,N_39767,N_38974);
nor U42941 (N_42941,N_36415,N_37711);
xor U42942 (N_42942,N_35045,N_37540);
or U42943 (N_42943,N_38264,N_36839);
xnor U42944 (N_42944,N_35130,N_37503);
xor U42945 (N_42945,N_37349,N_39707);
or U42946 (N_42946,N_35964,N_37715);
xnor U42947 (N_42947,N_36116,N_38935);
xnor U42948 (N_42948,N_35886,N_38406);
nor U42949 (N_42949,N_39226,N_36037);
nand U42950 (N_42950,N_36713,N_37672);
nor U42951 (N_42951,N_35043,N_37017);
nand U42952 (N_42952,N_39088,N_39659);
and U42953 (N_42953,N_38346,N_38298);
and U42954 (N_42954,N_36954,N_38755);
nand U42955 (N_42955,N_39708,N_37634);
or U42956 (N_42956,N_37280,N_36925);
xor U42957 (N_42957,N_39452,N_35255);
nor U42958 (N_42958,N_38316,N_35073);
xnor U42959 (N_42959,N_35282,N_39985);
nor U42960 (N_42960,N_36109,N_38922);
or U42961 (N_42961,N_37889,N_37989);
xnor U42962 (N_42962,N_35790,N_38303);
nand U42963 (N_42963,N_38712,N_38654);
and U42964 (N_42964,N_37606,N_37431);
xnor U42965 (N_42965,N_35971,N_35240);
xor U42966 (N_42966,N_36522,N_37772);
nand U42967 (N_42967,N_35793,N_37428);
nor U42968 (N_42968,N_38498,N_38243);
and U42969 (N_42969,N_37131,N_39243);
or U42970 (N_42970,N_35119,N_37870);
nand U42971 (N_42971,N_37140,N_35481);
and U42972 (N_42972,N_36559,N_35208);
xor U42973 (N_42973,N_38301,N_36923);
or U42974 (N_42974,N_37541,N_36223);
xnor U42975 (N_42975,N_37813,N_38732);
or U42976 (N_42976,N_39701,N_39529);
xnor U42977 (N_42977,N_37751,N_35792);
nor U42978 (N_42978,N_37506,N_39290);
nor U42979 (N_42979,N_39519,N_35519);
or U42980 (N_42980,N_39987,N_39495);
nor U42981 (N_42981,N_38246,N_37670);
or U42982 (N_42982,N_39417,N_37885);
and U42983 (N_42983,N_35825,N_35998);
or U42984 (N_42984,N_36926,N_35682);
nor U42985 (N_42985,N_35551,N_38200);
and U42986 (N_42986,N_39720,N_35509);
and U42987 (N_42987,N_38796,N_35230);
or U42988 (N_42988,N_38369,N_39662);
nand U42989 (N_42989,N_36040,N_36184);
nor U42990 (N_42990,N_36124,N_35942);
nor U42991 (N_42991,N_36015,N_35967);
nor U42992 (N_42992,N_39220,N_38530);
xor U42993 (N_42993,N_39222,N_36782);
and U42994 (N_42994,N_38298,N_35665);
xnor U42995 (N_42995,N_35478,N_38133);
and U42996 (N_42996,N_38364,N_36985);
nor U42997 (N_42997,N_36630,N_38873);
and U42998 (N_42998,N_35079,N_39239);
xnor U42999 (N_42999,N_39552,N_37079);
nor U43000 (N_43000,N_36498,N_36691);
or U43001 (N_43001,N_35902,N_37499);
or U43002 (N_43002,N_38833,N_38038);
and U43003 (N_43003,N_35035,N_39230);
and U43004 (N_43004,N_38358,N_39538);
and U43005 (N_43005,N_38548,N_37624);
and U43006 (N_43006,N_35214,N_39412);
and U43007 (N_43007,N_39658,N_39467);
or U43008 (N_43008,N_36890,N_38533);
and U43009 (N_43009,N_36389,N_36044);
and U43010 (N_43010,N_35740,N_37330);
or U43011 (N_43011,N_37281,N_37926);
and U43012 (N_43012,N_39448,N_37316);
xor U43013 (N_43013,N_35250,N_38087);
xor U43014 (N_43014,N_35432,N_37529);
nor U43015 (N_43015,N_38970,N_36856);
and U43016 (N_43016,N_38341,N_37175);
nand U43017 (N_43017,N_37700,N_38530);
nand U43018 (N_43018,N_35626,N_37552);
xor U43019 (N_43019,N_38424,N_35699);
xnor U43020 (N_43020,N_37692,N_37576);
xor U43021 (N_43021,N_35294,N_37103);
and U43022 (N_43022,N_39592,N_37881);
and U43023 (N_43023,N_37640,N_38523);
or U43024 (N_43024,N_36711,N_39342);
or U43025 (N_43025,N_39636,N_38187);
xnor U43026 (N_43026,N_35476,N_39623);
nor U43027 (N_43027,N_35931,N_38994);
nor U43028 (N_43028,N_39566,N_39710);
nor U43029 (N_43029,N_37398,N_36223);
nor U43030 (N_43030,N_37448,N_37325);
or U43031 (N_43031,N_37664,N_36417);
xor U43032 (N_43032,N_39347,N_37351);
or U43033 (N_43033,N_35732,N_37693);
nand U43034 (N_43034,N_36917,N_35348);
xnor U43035 (N_43035,N_36968,N_38928);
and U43036 (N_43036,N_38282,N_38534);
nor U43037 (N_43037,N_35911,N_35817);
or U43038 (N_43038,N_35054,N_38105);
or U43039 (N_43039,N_36148,N_38111);
or U43040 (N_43040,N_36983,N_37698);
nor U43041 (N_43041,N_35628,N_39945);
and U43042 (N_43042,N_35561,N_35753);
and U43043 (N_43043,N_38537,N_39122);
nand U43044 (N_43044,N_35759,N_35052);
and U43045 (N_43045,N_38936,N_36089);
nor U43046 (N_43046,N_37860,N_39740);
or U43047 (N_43047,N_35001,N_37133);
and U43048 (N_43048,N_35115,N_35004);
or U43049 (N_43049,N_38439,N_36464);
nand U43050 (N_43050,N_35068,N_37347);
nand U43051 (N_43051,N_38814,N_36457);
nand U43052 (N_43052,N_37771,N_38553);
and U43053 (N_43053,N_38137,N_39980);
nor U43054 (N_43054,N_35961,N_35924);
nor U43055 (N_43055,N_39745,N_39562);
and U43056 (N_43056,N_39336,N_36280);
nand U43057 (N_43057,N_36749,N_38444);
xnor U43058 (N_43058,N_39237,N_37250);
and U43059 (N_43059,N_36460,N_39792);
xnor U43060 (N_43060,N_36807,N_36197);
and U43061 (N_43061,N_37979,N_36441);
and U43062 (N_43062,N_38226,N_37004);
nor U43063 (N_43063,N_35582,N_36386);
nand U43064 (N_43064,N_36045,N_38325);
nand U43065 (N_43065,N_38666,N_35763);
xnor U43066 (N_43066,N_38784,N_35477);
nor U43067 (N_43067,N_38951,N_37948);
xor U43068 (N_43068,N_39229,N_36644);
and U43069 (N_43069,N_36240,N_35449);
or U43070 (N_43070,N_36505,N_37831);
nor U43071 (N_43071,N_37046,N_38481);
nand U43072 (N_43072,N_39074,N_39927);
and U43073 (N_43073,N_39061,N_35691);
nand U43074 (N_43074,N_35655,N_39669);
nor U43075 (N_43075,N_38566,N_36193);
nand U43076 (N_43076,N_37478,N_35903);
or U43077 (N_43077,N_37037,N_39747);
xor U43078 (N_43078,N_36158,N_39365);
and U43079 (N_43079,N_38704,N_38482);
xnor U43080 (N_43080,N_35581,N_39113);
or U43081 (N_43081,N_38553,N_39708);
or U43082 (N_43082,N_39175,N_37456);
nand U43083 (N_43083,N_35847,N_38032);
and U43084 (N_43084,N_38836,N_38478);
or U43085 (N_43085,N_39532,N_38542);
or U43086 (N_43086,N_37369,N_36391);
xnor U43087 (N_43087,N_36322,N_37129);
nand U43088 (N_43088,N_38847,N_39023);
or U43089 (N_43089,N_38814,N_36913);
and U43090 (N_43090,N_36525,N_36397);
or U43091 (N_43091,N_35783,N_37955);
nor U43092 (N_43092,N_39329,N_38370);
nor U43093 (N_43093,N_37643,N_36551);
or U43094 (N_43094,N_38102,N_36844);
xor U43095 (N_43095,N_35125,N_36506);
nor U43096 (N_43096,N_36939,N_37974);
nor U43097 (N_43097,N_39777,N_38113);
nor U43098 (N_43098,N_39871,N_39546);
or U43099 (N_43099,N_39113,N_38108);
or U43100 (N_43100,N_39363,N_38550);
xnor U43101 (N_43101,N_38614,N_35749);
nor U43102 (N_43102,N_36295,N_39151);
or U43103 (N_43103,N_35905,N_37872);
nand U43104 (N_43104,N_38756,N_37371);
nor U43105 (N_43105,N_36507,N_39768);
and U43106 (N_43106,N_37664,N_36695);
xnor U43107 (N_43107,N_35860,N_37701);
nand U43108 (N_43108,N_38868,N_38089);
nand U43109 (N_43109,N_38106,N_36738);
nand U43110 (N_43110,N_35747,N_39983);
or U43111 (N_43111,N_35851,N_37866);
xor U43112 (N_43112,N_36899,N_37894);
nand U43113 (N_43113,N_38591,N_37329);
and U43114 (N_43114,N_38819,N_36180);
and U43115 (N_43115,N_38060,N_39958);
nor U43116 (N_43116,N_35847,N_38583);
nand U43117 (N_43117,N_35799,N_38968);
nor U43118 (N_43118,N_38306,N_39194);
nand U43119 (N_43119,N_38520,N_39792);
nand U43120 (N_43120,N_39446,N_36589);
nor U43121 (N_43121,N_36161,N_35366);
nand U43122 (N_43122,N_38285,N_37454);
and U43123 (N_43123,N_35190,N_38288);
xnor U43124 (N_43124,N_35384,N_38377);
or U43125 (N_43125,N_35670,N_35526);
nor U43126 (N_43126,N_38176,N_36891);
xnor U43127 (N_43127,N_37571,N_35185);
xor U43128 (N_43128,N_39372,N_39864);
nor U43129 (N_43129,N_39215,N_39912);
nor U43130 (N_43130,N_35650,N_36982);
xnor U43131 (N_43131,N_37790,N_35456);
xor U43132 (N_43132,N_37701,N_35179);
xnor U43133 (N_43133,N_36368,N_37220);
or U43134 (N_43134,N_38866,N_38076);
xnor U43135 (N_43135,N_35784,N_39367);
nand U43136 (N_43136,N_37406,N_39523);
and U43137 (N_43137,N_39438,N_38672);
xor U43138 (N_43138,N_35302,N_35758);
nand U43139 (N_43139,N_35229,N_36421);
nand U43140 (N_43140,N_35124,N_35547);
xnor U43141 (N_43141,N_35691,N_36133);
nand U43142 (N_43142,N_35103,N_39728);
xnor U43143 (N_43143,N_35516,N_35096);
or U43144 (N_43144,N_35492,N_36669);
nand U43145 (N_43145,N_39481,N_35358);
or U43146 (N_43146,N_35960,N_36899);
or U43147 (N_43147,N_37322,N_38105);
or U43148 (N_43148,N_37530,N_36126);
nor U43149 (N_43149,N_35778,N_38530);
nor U43150 (N_43150,N_35083,N_39075);
nand U43151 (N_43151,N_39695,N_35854);
nor U43152 (N_43152,N_35705,N_39996);
and U43153 (N_43153,N_38972,N_37499);
nor U43154 (N_43154,N_38408,N_37974);
nor U43155 (N_43155,N_37122,N_35566);
and U43156 (N_43156,N_39360,N_38714);
nor U43157 (N_43157,N_37631,N_37955);
nand U43158 (N_43158,N_38799,N_37467);
nor U43159 (N_43159,N_37650,N_36239);
nand U43160 (N_43160,N_38827,N_38251);
nor U43161 (N_43161,N_39420,N_38644);
nand U43162 (N_43162,N_39227,N_39319);
and U43163 (N_43163,N_39875,N_36629);
nand U43164 (N_43164,N_38371,N_39235);
and U43165 (N_43165,N_37144,N_39607);
nor U43166 (N_43166,N_35932,N_35328);
nor U43167 (N_43167,N_37314,N_37451);
nand U43168 (N_43168,N_37656,N_38713);
nand U43169 (N_43169,N_36578,N_38264);
or U43170 (N_43170,N_38951,N_38538);
nor U43171 (N_43171,N_39069,N_38610);
and U43172 (N_43172,N_35748,N_36666);
xnor U43173 (N_43173,N_37248,N_38434);
nor U43174 (N_43174,N_38456,N_37976);
or U43175 (N_43175,N_38535,N_38084);
and U43176 (N_43176,N_36486,N_36503);
xnor U43177 (N_43177,N_36014,N_38690);
nand U43178 (N_43178,N_38361,N_35556);
nand U43179 (N_43179,N_38218,N_36657);
nor U43180 (N_43180,N_35937,N_39279);
nor U43181 (N_43181,N_37074,N_39781);
or U43182 (N_43182,N_38212,N_36341);
xor U43183 (N_43183,N_35786,N_36500);
and U43184 (N_43184,N_35808,N_37733);
xor U43185 (N_43185,N_35975,N_36772);
and U43186 (N_43186,N_37867,N_39630);
or U43187 (N_43187,N_38588,N_39234);
nand U43188 (N_43188,N_39897,N_38245);
xor U43189 (N_43189,N_36953,N_37664);
and U43190 (N_43190,N_37036,N_38616);
xor U43191 (N_43191,N_37879,N_39389);
nor U43192 (N_43192,N_39845,N_36204);
and U43193 (N_43193,N_35585,N_37601);
nand U43194 (N_43194,N_37179,N_36830);
or U43195 (N_43195,N_37993,N_37678);
or U43196 (N_43196,N_38805,N_37962);
xnor U43197 (N_43197,N_39639,N_39787);
nor U43198 (N_43198,N_36847,N_38104);
nand U43199 (N_43199,N_36835,N_39317);
or U43200 (N_43200,N_39521,N_39056);
or U43201 (N_43201,N_36518,N_37801);
xnor U43202 (N_43202,N_39423,N_36845);
xnor U43203 (N_43203,N_37463,N_39608);
or U43204 (N_43204,N_36581,N_37192);
nor U43205 (N_43205,N_38218,N_35948);
or U43206 (N_43206,N_37462,N_39326);
and U43207 (N_43207,N_37689,N_35795);
nor U43208 (N_43208,N_39844,N_36372);
nor U43209 (N_43209,N_35761,N_39295);
or U43210 (N_43210,N_37288,N_35128);
or U43211 (N_43211,N_35493,N_39900);
and U43212 (N_43212,N_35072,N_38062);
nand U43213 (N_43213,N_38364,N_36322);
xnor U43214 (N_43214,N_39238,N_35845);
xnor U43215 (N_43215,N_38814,N_36350);
nand U43216 (N_43216,N_37704,N_35766);
nor U43217 (N_43217,N_36072,N_39127);
nor U43218 (N_43218,N_35219,N_37922);
xor U43219 (N_43219,N_39044,N_37666);
nor U43220 (N_43220,N_36057,N_37795);
nor U43221 (N_43221,N_35818,N_35518);
xnor U43222 (N_43222,N_39946,N_38106);
nor U43223 (N_43223,N_38145,N_39814);
and U43224 (N_43224,N_39951,N_37513);
nand U43225 (N_43225,N_39136,N_39540);
xnor U43226 (N_43226,N_36744,N_35317);
and U43227 (N_43227,N_35389,N_35073);
or U43228 (N_43228,N_36339,N_35721);
xor U43229 (N_43229,N_35003,N_36723);
xor U43230 (N_43230,N_36246,N_38420);
and U43231 (N_43231,N_35589,N_36278);
xor U43232 (N_43232,N_36766,N_37823);
and U43233 (N_43233,N_39201,N_38608);
nand U43234 (N_43234,N_35182,N_37025);
nand U43235 (N_43235,N_38536,N_37010);
or U43236 (N_43236,N_36967,N_39160);
nand U43237 (N_43237,N_37539,N_37592);
nor U43238 (N_43238,N_36419,N_35960);
nand U43239 (N_43239,N_37207,N_36150);
and U43240 (N_43240,N_35404,N_36103);
xnor U43241 (N_43241,N_37336,N_37459);
and U43242 (N_43242,N_39609,N_39057);
or U43243 (N_43243,N_35710,N_39807);
or U43244 (N_43244,N_35002,N_37911);
nand U43245 (N_43245,N_35443,N_39236);
or U43246 (N_43246,N_35697,N_35291);
nand U43247 (N_43247,N_39841,N_35773);
and U43248 (N_43248,N_39703,N_39168);
and U43249 (N_43249,N_35843,N_39601);
nand U43250 (N_43250,N_36484,N_37200);
and U43251 (N_43251,N_35298,N_39880);
xnor U43252 (N_43252,N_38763,N_35420);
xor U43253 (N_43253,N_36839,N_38148);
nor U43254 (N_43254,N_39438,N_35053);
or U43255 (N_43255,N_37400,N_37254);
and U43256 (N_43256,N_37371,N_35751);
or U43257 (N_43257,N_37546,N_37688);
nand U43258 (N_43258,N_36912,N_37933);
xor U43259 (N_43259,N_36492,N_35877);
and U43260 (N_43260,N_39090,N_37370);
and U43261 (N_43261,N_39981,N_38180);
xor U43262 (N_43262,N_39575,N_39425);
or U43263 (N_43263,N_37261,N_38122);
nor U43264 (N_43264,N_36276,N_35256);
nand U43265 (N_43265,N_35444,N_38356);
nand U43266 (N_43266,N_37015,N_36936);
or U43267 (N_43267,N_38855,N_35958);
nand U43268 (N_43268,N_39087,N_37803);
or U43269 (N_43269,N_36989,N_38534);
xnor U43270 (N_43270,N_36521,N_39325);
nor U43271 (N_43271,N_38499,N_35775);
or U43272 (N_43272,N_35140,N_38318);
xnor U43273 (N_43273,N_38276,N_38876);
xor U43274 (N_43274,N_37024,N_38046);
or U43275 (N_43275,N_36526,N_37774);
nor U43276 (N_43276,N_37248,N_35281);
xnor U43277 (N_43277,N_38349,N_35422);
nor U43278 (N_43278,N_36093,N_35509);
and U43279 (N_43279,N_35693,N_35618);
xnor U43280 (N_43280,N_37949,N_39136);
xnor U43281 (N_43281,N_35904,N_38069);
or U43282 (N_43282,N_38981,N_38191);
nor U43283 (N_43283,N_35695,N_36689);
nand U43284 (N_43284,N_39855,N_37469);
nand U43285 (N_43285,N_36959,N_35075);
nor U43286 (N_43286,N_36825,N_36527);
nor U43287 (N_43287,N_37361,N_35841);
nand U43288 (N_43288,N_38339,N_39557);
xnor U43289 (N_43289,N_39887,N_35907);
and U43290 (N_43290,N_35260,N_36134);
xor U43291 (N_43291,N_35551,N_35724);
nor U43292 (N_43292,N_39376,N_37341);
and U43293 (N_43293,N_37750,N_39990);
and U43294 (N_43294,N_39010,N_35958);
or U43295 (N_43295,N_35660,N_39156);
xor U43296 (N_43296,N_37018,N_37095);
and U43297 (N_43297,N_37385,N_38600);
or U43298 (N_43298,N_36759,N_36959);
or U43299 (N_43299,N_37708,N_37084);
xor U43300 (N_43300,N_37521,N_37324);
nor U43301 (N_43301,N_35250,N_39583);
xor U43302 (N_43302,N_38183,N_37449);
and U43303 (N_43303,N_39422,N_36197);
nor U43304 (N_43304,N_36068,N_39190);
nor U43305 (N_43305,N_35831,N_37795);
nor U43306 (N_43306,N_37563,N_38169);
or U43307 (N_43307,N_35640,N_39832);
xnor U43308 (N_43308,N_39132,N_37741);
nand U43309 (N_43309,N_37103,N_37616);
xnor U43310 (N_43310,N_35762,N_39789);
or U43311 (N_43311,N_39424,N_39357);
and U43312 (N_43312,N_35287,N_39668);
nor U43313 (N_43313,N_35617,N_35923);
and U43314 (N_43314,N_35349,N_35653);
nor U43315 (N_43315,N_35741,N_36663);
and U43316 (N_43316,N_38500,N_38560);
or U43317 (N_43317,N_36518,N_35283);
nand U43318 (N_43318,N_37293,N_39847);
nor U43319 (N_43319,N_36875,N_36962);
and U43320 (N_43320,N_36544,N_38426);
nor U43321 (N_43321,N_38376,N_36992);
nand U43322 (N_43322,N_37344,N_38311);
and U43323 (N_43323,N_37776,N_38597);
and U43324 (N_43324,N_35385,N_39142);
nor U43325 (N_43325,N_35881,N_36361);
or U43326 (N_43326,N_38480,N_39943);
nor U43327 (N_43327,N_35331,N_38881);
nor U43328 (N_43328,N_38597,N_39644);
xor U43329 (N_43329,N_39990,N_39312);
or U43330 (N_43330,N_38125,N_36681);
and U43331 (N_43331,N_39728,N_36509);
xor U43332 (N_43332,N_35034,N_35525);
nor U43333 (N_43333,N_38569,N_36605);
nand U43334 (N_43334,N_39296,N_38542);
or U43335 (N_43335,N_35017,N_38768);
or U43336 (N_43336,N_39023,N_38206);
and U43337 (N_43337,N_38972,N_38188);
or U43338 (N_43338,N_35522,N_37929);
nand U43339 (N_43339,N_37123,N_35118);
or U43340 (N_43340,N_35714,N_38697);
xor U43341 (N_43341,N_38865,N_39879);
xnor U43342 (N_43342,N_39305,N_35240);
xnor U43343 (N_43343,N_37746,N_37244);
and U43344 (N_43344,N_38966,N_37183);
nor U43345 (N_43345,N_36359,N_38578);
nor U43346 (N_43346,N_37348,N_36121);
nand U43347 (N_43347,N_38896,N_36933);
and U43348 (N_43348,N_37807,N_35197);
xor U43349 (N_43349,N_39802,N_39535);
nand U43350 (N_43350,N_37909,N_36777);
or U43351 (N_43351,N_36494,N_37912);
or U43352 (N_43352,N_35284,N_35477);
nor U43353 (N_43353,N_35792,N_39802);
nand U43354 (N_43354,N_36024,N_39636);
nor U43355 (N_43355,N_39190,N_37956);
nor U43356 (N_43356,N_36925,N_38705);
and U43357 (N_43357,N_35060,N_36158);
xor U43358 (N_43358,N_38708,N_37870);
or U43359 (N_43359,N_36808,N_36113);
or U43360 (N_43360,N_35707,N_35325);
xor U43361 (N_43361,N_39366,N_36825);
or U43362 (N_43362,N_35443,N_37753);
nand U43363 (N_43363,N_39074,N_39178);
nand U43364 (N_43364,N_39843,N_36690);
xnor U43365 (N_43365,N_35757,N_36614);
nor U43366 (N_43366,N_35429,N_38643);
or U43367 (N_43367,N_39371,N_39415);
nor U43368 (N_43368,N_35302,N_37090);
or U43369 (N_43369,N_35180,N_36695);
xnor U43370 (N_43370,N_39591,N_35194);
or U43371 (N_43371,N_39264,N_37326);
xnor U43372 (N_43372,N_39494,N_35891);
or U43373 (N_43373,N_37645,N_36444);
or U43374 (N_43374,N_39932,N_37408);
or U43375 (N_43375,N_38487,N_37893);
nor U43376 (N_43376,N_37690,N_38076);
nor U43377 (N_43377,N_36469,N_36741);
nor U43378 (N_43378,N_37991,N_39680);
xor U43379 (N_43379,N_35888,N_38524);
nor U43380 (N_43380,N_37861,N_35743);
xor U43381 (N_43381,N_38955,N_36830);
or U43382 (N_43382,N_36523,N_38598);
and U43383 (N_43383,N_37489,N_39673);
nor U43384 (N_43384,N_37700,N_37149);
or U43385 (N_43385,N_39072,N_38815);
nand U43386 (N_43386,N_37512,N_39957);
xnor U43387 (N_43387,N_37478,N_38592);
nor U43388 (N_43388,N_35941,N_35788);
xnor U43389 (N_43389,N_35765,N_36768);
and U43390 (N_43390,N_38598,N_39946);
and U43391 (N_43391,N_35834,N_36715);
nor U43392 (N_43392,N_35963,N_37016);
and U43393 (N_43393,N_37238,N_36871);
or U43394 (N_43394,N_36220,N_39839);
or U43395 (N_43395,N_37659,N_39052);
or U43396 (N_43396,N_37968,N_38173);
nor U43397 (N_43397,N_35085,N_36468);
nor U43398 (N_43398,N_37403,N_37008);
nand U43399 (N_43399,N_38157,N_38319);
xnor U43400 (N_43400,N_36990,N_39159);
xor U43401 (N_43401,N_38280,N_35955);
xnor U43402 (N_43402,N_38555,N_37385);
or U43403 (N_43403,N_39121,N_35151);
or U43404 (N_43404,N_38905,N_37341);
or U43405 (N_43405,N_39699,N_37056);
nand U43406 (N_43406,N_37511,N_39841);
and U43407 (N_43407,N_38863,N_38367);
nand U43408 (N_43408,N_35038,N_37357);
nand U43409 (N_43409,N_37719,N_35128);
xnor U43410 (N_43410,N_36174,N_35073);
xnor U43411 (N_43411,N_39781,N_37380);
nand U43412 (N_43412,N_36363,N_36007);
xnor U43413 (N_43413,N_35748,N_37054);
xnor U43414 (N_43414,N_39592,N_35771);
xnor U43415 (N_43415,N_37803,N_36936);
or U43416 (N_43416,N_36257,N_35807);
and U43417 (N_43417,N_39505,N_35088);
nor U43418 (N_43418,N_36968,N_35163);
or U43419 (N_43419,N_35099,N_39662);
or U43420 (N_43420,N_36990,N_36486);
nor U43421 (N_43421,N_39038,N_35960);
nand U43422 (N_43422,N_36854,N_39070);
nand U43423 (N_43423,N_36259,N_37039);
xor U43424 (N_43424,N_36189,N_37878);
and U43425 (N_43425,N_37783,N_36776);
nand U43426 (N_43426,N_37254,N_35555);
nand U43427 (N_43427,N_39118,N_39370);
xnor U43428 (N_43428,N_37524,N_39774);
and U43429 (N_43429,N_36939,N_39957);
and U43430 (N_43430,N_38842,N_36125);
and U43431 (N_43431,N_39852,N_36003);
nor U43432 (N_43432,N_39084,N_39762);
or U43433 (N_43433,N_38129,N_37124);
and U43434 (N_43434,N_38118,N_39496);
nand U43435 (N_43435,N_37111,N_36482);
nor U43436 (N_43436,N_38155,N_35459);
nor U43437 (N_43437,N_35089,N_39422);
nor U43438 (N_43438,N_36335,N_36913);
nor U43439 (N_43439,N_37264,N_38296);
or U43440 (N_43440,N_37042,N_38033);
or U43441 (N_43441,N_35144,N_39558);
nor U43442 (N_43442,N_36806,N_37065);
or U43443 (N_43443,N_39243,N_39836);
xor U43444 (N_43444,N_37504,N_38352);
nor U43445 (N_43445,N_37761,N_38574);
and U43446 (N_43446,N_36274,N_36654);
and U43447 (N_43447,N_38005,N_37383);
nand U43448 (N_43448,N_35322,N_35097);
and U43449 (N_43449,N_37917,N_35651);
or U43450 (N_43450,N_39781,N_37139);
xor U43451 (N_43451,N_35753,N_37751);
and U43452 (N_43452,N_35840,N_38836);
nand U43453 (N_43453,N_37462,N_36261);
and U43454 (N_43454,N_35589,N_35161);
and U43455 (N_43455,N_36270,N_35449);
xor U43456 (N_43456,N_36674,N_37050);
and U43457 (N_43457,N_35483,N_35896);
and U43458 (N_43458,N_38036,N_39838);
nand U43459 (N_43459,N_37473,N_37398);
xnor U43460 (N_43460,N_35500,N_36647);
and U43461 (N_43461,N_39896,N_38996);
xor U43462 (N_43462,N_39471,N_35980);
xnor U43463 (N_43463,N_37154,N_35858);
nand U43464 (N_43464,N_37012,N_35429);
xor U43465 (N_43465,N_37297,N_37887);
xnor U43466 (N_43466,N_35518,N_38687);
nor U43467 (N_43467,N_37681,N_39504);
nor U43468 (N_43468,N_36183,N_37315);
or U43469 (N_43469,N_35040,N_39394);
and U43470 (N_43470,N_35478,N_39523);
nor U43471 (N_43471,N_35297,N_37442);
xor U43472 (N_43472,N_37320,N_39064);
and U43473 (N_43473,N_36728,N_37560);
nor U43474 (N_43474,N_36985,N_35541);
xnor U43475 (N_43475,N_38734,N_37336);
nand U43476 (N_43476,N_36968,N_38466);
nand U43477 (N_43477,N_37025,N_38071);
xnor U43478 (N_43478,N_39163,N_36128);
xor U43479 (N_43479,N_38047,N_38175);
and U43480 (N_43480,N_38740,N_37985);
nor U43481 (N_43481,N_39549,N_38051);
or U43482 (N_43482,N_35767,N_38064);
and U43483 (N_43483,N_35485,N_38442);
nor U43484 (N_43484,N_37998,N_37124);
nor U43485 (N_43485,N_37475,N_39035);
nor U43486 (N_43486,N_39531,N_36607);
nor U43487 (N_43487,N_39436,N_35806);
nor U43488 (N_43488,N_35075,N_39463);
nand U43489 (N_43489,N_38720,N_39215);
or U43490 (N_43490,N_37735,N_36745);
and U43491 (N_43491,N_36868,N_39896);
or U43492 (N_43492,N_36824,N_36186);
nor U43493 (N_43493,N_39147,N_39022);
nor U43494 (N_43494,N_35142,N_35324);
and U43495 (N_43495,N_36067,N_38486);
or U43496 (N_43496,N_36210,N_38204);
xor U43497 (N_43497,N_35928,N_38645);
nor U43498 (N_43498,N_36395,N_36305);
xnor U43499 (N_43499,N_37523,N_39521);
xnor U43500 (N_43500,N_37784,N_37150);
nand U43501 (N_43501,N_35528,N_38659);
nand U43502 (N_43502,N_39452,N_38632);
xnor U43503 (N_43503,N_38567,N_38557);
or U43504 (N_43504,N_37765,N_39965);
xnor U43505 (N_43505,N_35675,N_38716);
xnor U43506 (N_43506,N_39694,N_39234);
nand U43507 (N_43507,N_38971,N_39866);
nand U43508 (N_43508,N_39359,N_36246);
or U43509 (N_43509,N_36581,N_38522);
xor U43510 (N_43510,N_35279,N_37032);
xor U43511 (N_43511,N_38624,N_35452);
nor U43512 (N_43512,N_39051,N_36648);
or U43513 (N_43513,N_36902,N_38443);
and U43514 (N_43514,N_39152,N_38154);
nor U43515 (N_43515,N_35734,N_36532);
or U43516 (N_43516,N_37982,N_39678);
nand U43517 (N_43517,N_36939,N_35560);
nor U43518 (N_43518,N_36559,N_37286);
nand U43519 (N_43519,N_36898,N_35657);
and U43520 (N_43520,N_37150,N_36634);
and U43521 (N_43521,N_35016,N_39918);
xor U43522 (N_43522,N_38600,N_36740);
nor U43523 (N_43523,N_36337,N_39378);
xnor U43524 (N_43524,N_36992,N_39361);
nor U43525 (N_43525,N_37179,N_38108);
xor U43526 (N_43526,N_38585,N_36526);
xor U43527 (N_43527,N_36693,N_36222);
and U43528 (N_43528,N_38956,N_35669);
and U43529 (N_43529,N_35706,N_35637);
or U43530 (N_43530,N_37263,N_37091);
nor U43531 (N_43531,N_38370,N_38025);
and U43532 (N_43532,N_36057,N_39957);
and U43533 (N_43533,N_39775,N_36177);
nor U43534 (N_43534,N_39710,N_38447);
and U43535 (N_43535,N_38168,N_35736);
nand U43536 (N_43536,N_35897,N_39018);
xnor U43537 (N_43537,N_39044,N_39115);
nand U43538 (N_43538,N_37962,N_35983);
nor U43539 (N_43539,N_37686,N_35941);
or U43540 (N_43540,N_36278,N_39183);
or U43541 (N_43541,N_36740,N_39821);
nand U43542 (N_43542,N_36204,N_36131);
nand U43543 (N_43543,N_35010,N_38644);
or U43544 (N_43544,N_39418,N_37241);
nor U43545 (N_43545,N_35529,N_37493);
or U43546 (N_43546,N_36702,N_35137);
nand U43547 (N_43547,N_38755,N_36575);
nand U43548 (N_43548,N_38645,N_37528);
or U43549 (N_43549,N_38352,N_37755);
nor U43550 (N_43550,N_38689,N_38215);
nand U43551 (N_43551,N_39279,N_38516);
nand U43552 (N_43552,N_36340,N_38377);
nor U43553 (N_43553,N_38272,N_36626);
xnor U43554 (N_43554,N_39198,N_37807);
nor U43555 (N_43555,N_35400,N_37115);
or U43556 (N_43556,N_39524,N_39137);
nand U43557 (N_43557,N_39874,N_37935);
nand U43558 (N_43558,N_35990,N_37098);
xnor U43559 (N_43559,N_39174,N_35975);
xor U43560 (N_43560,N_37563,N_38882);
nor U43561 (N_43561,N_36254,N_39389);
and U43562 (N_43562,N_37190,N_39216);
nand U43563 (N_43563,N_35824,N_36813);
nand U43564 (N_43564,N_35389,N_39366);
or U43565 (N_43565,N_37457,N_35395);
or U43566 (N_43566,N_37853,N_36741);
nand U43567 (N_43567,N_38434,N_39722);
nand U43568 (N_43568,N_35595,N_39094);
xnor U43569 (N_43569,N_36223,N_39914);
xnor U43570 (N_43570,N_36997,N_37380);
xnor U43571 (N_43571,N_37116,N_36585);
xor U43572 (N_43572,N_35411,N_38770);
and U43573 (N_43573,N_39749,N_36196);
nor U43574 (N_43574,N_37680,N_35338);
and U43575 (N_43575,N_39461,N_39220);
or U43576 (N_43576,N_38371,N_39639);
and U43577 (N_43577,N_38281,N_36305);
nor U43578 (N_43578,N_36168,N_37376);
and U43579 (N_43579,N_37186,N_37414);
and U43580 (N_43580,N_35011,N_39134);
and U43581 (N_43581,N_38897,N_36672);
nand U43582 (N_43582,N_35740,N_36624);
or U43583 (N_43583,N_38398,N_38439);
nand U43584 (N_43584,N_36413,N_38991);
and U43585 (N_43585,N_39536,N_35581);
nand U43586 (N_43586,N_37684,N_36098);
or U43587 (N_43587,N_35089,N_37051);
nor U43588 (N_43588,N_36161,N_35331);
nand U43589 (N_43589,N_36077,N_36661);
xnor U43590 (N_43590,N_38820,N_37309);
and U43591 (N_43591,N_38525,N_36070);
or U43592 (N_43592,N_39499,N_39687);
or U43593 (N_43593,N_39435,N_37030);
nand U43594 (N_43594,N_39602,N_38309);
nand U43595 (N_43595,N_37865,N_38619);
xnor U43596 (N_43596,N_36902,N_37022);
and U43597 (N_43597,N_37768,N_35001);
nor U43598 (N_43598,N_36094,N_37130);
or U43599 (N_43599,N_36455,N_35624);
nor U43600 (N_43600,N_39992,N_36329);
nand U43601 (N_43601,N_36786,N_36950);
and U43602 (N_43602,N_36625,N_36615);
nand U43603 (N_43603,N_37583,N_39347);
and U43604 (N_43604,N_39501,N_35048);
xor U43605 (N_43605,N_39125,N_36588);
nand U43606 (N_43606,N_37815,N_37632);
nand U43607 (N_43607,N_36652,N_35981);
and U43608 (N_43608,N_35979,N_39055);
and U43609 (N_43609,N_39346,N_35098);
and U43610 (N_43610,N_37539,N_36438);
and U43611 (N_43611,N_39695,N_36051);
xnor U43612 (N_43612,N_35528,N_35357);
xor U43613 (N_43613,N_38259,N_39443);
nand U43614 (N_43614,N_37170,N_37827);
and U43615 (N_43615,N_37788,N_35519);
and U43616 (N_43616,N_37542,N_36155);
nor U43617 (N_43617,N_38312,N_35368);
xor U43618 (N_43618,N_39353,N_37374);
xnor U43619 (N_43619,N_36695,N_36162);
xor U43620 (N_43620,N_37413,N_39343);
nand U43621 (N_43621,N_38743,N_35761);
nor U43622 (N_43622,N_38883,N_37192);
nor U43623 (N_43623,N_35685,N_35488);
nand U43624 (N_43624,N_36257,N_37829);
or U43625 (N_43625,N_37732,N_37836);
nand U43626 (N_43626,N_36477,N_39990);
nor U43627 (N_43627,N_39203,N_39477);
and U43628 (N_43628,N_38405,N_38471);
and U43629 (N_43629,N_38106,N_38355);
nor U43630 (N_43630,N_35322,N_35005);
nand U43631 (N_43631,N_35030,N_39599);
and U43632 (N_43632,N_39660,N_37614);
nor U43633 (N_43633,N_35705,N_35382);
and U43634 (N_43634,N_36152,N_36523);
xnor U43635 (N_43635,N_38418,N_36185);
or U43636 (N_43636,N_36517,N_36975);
xnor U43637 (N_43637,N_36323,N_38451);
xor U43638 (N_43638,N_39904,N_37549);
xnor U43639 (N_43639,N_37912,N_37794);
and U43640 (N_43640,N_35782,N_38255);
xor U43641 (N_43641,N_39938,N_39948);
nand U43642 (N_43642,N_39940,N_38726);
and U43643 (N_43643,N_37436,N_39552);
or U43644 (N_43644,N_38132,N_35326);
nand U43645 (N_43645,N_35923,N_36326);
or U43646 (N_43646,N_38293,N_39332);
nand U43647 (N_43647,N_39649,N_38363);
and U43648 (N_43648,N_38123,N_38721);
xor U43649 (N_43649,N_38068,N_37091);
or U43650 (N_43650,N_38621,N_35896);
or U43651 (N_43651,N_36998,N_35817);
nand U43652 (N_43652,N_36244,N_38947);
nand U43653 (N_43653,N_38628,N_35474);
nand U43654 (N_43654,N_39375,N_35042);
or U43655 (N_43655,N_36359,N_36251);
or U43656 (N_43656,N_39004,N_39702);
nand U43657 (N_43657,N_37651,N_36126);
or U43658 (N_43658,N_35326,N_36501);
nor U43659 (N_43659,N_39465,N_36742);
xnor U43660 (N_43660,N_38857,N_37427);
nand U43661 (N_43661,N_37512,N_36617);
nand U43662 (N_43662,N_38938,N_36721);
and U43663 (N_43663,N_39957,N_35623);
and U43664 (N_43664,N_38890,N_39246);
nand U43665 (N_43665,N_37845,N_36281);
xnor U43666 (N_43666,N_35161,N_36561);
or U43667 (N_43667,N_38598,N_35926);
nand U43668 (N_43668,N_39758,N_37699);
and U43669 (N_43669,N_36824,N_37458);
and U43670 (N_43670,N_38396,N_36596);
or U43671 (N_43671,N_35923,N_38984);
or U43672 (N_43672,N_39435,N_39260);
xor U43673 (N_43673,N_39566,N_35256);
or U43674 (N_43674,N_38870,N_37401);
and U43675 (N_43675,N_35659,N_37281);
nand U43676 (N_43676,N_35769,N_35483);
and U43677 (N_43677,N_39385,N_36850);
or U43678 (N_43678,N_39202,N_37702);
nor U43679 (N_43679,N_35383,N_38764);
nand U43680 (N_43680,N_36856,N_39178);
nor U43681 (N_43681,N_37290,N_37585);
and U43682 (N_43682,N_37482,N_35188);
nor U43683 (N_43683,N_37081,N_39253);
nor U43684 (N_43684,N_38210,N_36141);
xor U43685 (N_43685,N_38298,N_35105);
and U43686 (N_43686,N_38602,N_39418);
and U43687 (N_43687,N_36512,N_39502);
nand U43688 (N_43688,N_39079,N_35548);
and U43689 (N_43689,N_37290,N_38192);
nand U43690 (N_43690,N_38605,N_35054);
nor U43691 (N_43691,N_35677,N_35495);
and U43692 (N_43692,N_38936,N_35693);
and U43693 (N_43693,N_39413,N_36986);
and U43694 (N_43694,N_36274,N_35086);
and U43695 (N_43695,N_39340,N_35118);
and U43696 (N_43696,N_35385,N_38046);
xnor U43697 (N_43697,N_39317,N_37045);
and U43698 (N_43698,N_35031,N_35844);
nor U43699 (N_43699,N_36471,N_35066);
nor U43700 (N_43700,N_38466,N_37324);
xor U43701 (N_43701,N_38403,N_39530);
nand U43702 (N_43702,N_35009,N_36691);
xor U43703 (N_43703,N_38938,N_37171);
xor U43704 (N_43704,N_39902,N_35675);
and U43705 (N_43705,N_37137,N_37672);
xnor U43706 (N_43706,N_37655,N_36807);
nor U43707 (N_43707,N_38526,N_37735);
or U43708 (N_43708,N_35200,N_35286);
and U43709 (N_43709,N_37979,N_39084);
nor U43710 (N_43710,N_38201,N_39542);
nand U43711 (N_43711,N_38230,N_39957);
and U43712 (N_43712,N_39238,N_37903);
xor U43713 (N_43713,N_37383,N_39281);
xor U43714 (N_43714,N_35948,N_38078);
and U43715 (N_43715,N_38453,N_39152);
or U43716 (N_43716,N_37834,N_36693);
nor U43717 (N_43717,N_37340,N_35220);
and U43718 (N_43718,N_37588,N_36598);
nand U43719 (N_43719,N_37767,N_39313);
or U43720 (N_43720,N_38776,N_37761);
and U43721 (N_43721,N_39886,N_35972);
nand U43722 (N_43722,N_39324,N_35597);
or U43723 (N_43723,N_37900,N_37376);
or U43724 (N_43724,N_36490,N_38057);
nand U43725 (N_43725,N_39242,N_35676);
or U43726 (N_43726,N_35856,N_38269);
nor U43727 (N_43727,N_37375,N_35211);
or U43728 (N_43728,N_35232,N_37854);
and U43729 (N_43729,N_36923,N_35464);
nand U43730 (N_43730,N_39848,N_39133);
nand U43731 (N_43731,N_38871,N_38669);
nor U43732 (N_43732,N_39313,N_36381);
xnor U43733 (N_43733,N_38877,N_36294);
or U43734 (N_43734,N_36070,N_38020);
nor U43735 (N_43735,N_38756,N_37726);
nand U43736 (N_43736,N_35955,N_35923);
or U43737 (N_43737,N_35608,N_36305);
and U43738 (N_43738,N_35033,N_37897);
or U43739 (N_43739,N_36745,N_38177);
xnor U43740 (N_43740,N_37092,N_39392);
xor U43741 (N_43741,N_35205,N_36913);
xor U43742 (N_43742,N_39237,N_38619);
or U43743 (N_43743,N_35836,N_38434);
nand U43744 (N_43744,N_39457,N_39355);
nor U43745 (N_43745,N_36236,N_36475);
or U43746 (N_43746,N_37037,N_35272);
and U43747 (N_43747,N_35257,N_36791);
nand U43748 (N_43748,N_36204,N_38643);
and U43749 (N_43749,N_35884,N_37947);
or U43750 (N_43750,N_37599,N_37235);
nand U43751 (N_43751,N_38632,N_35353);
and U43752 (N_43752,N_36869,N_38958);
nor U43753 (N_43753,N_38544,N_39465);
nor U43754 (N_43754,N_35365,N_38099);
or U43755 (N_43755,N_35241,N_38354);
xnor U43756 (N_43756,N_35451,N_35805);
or U43757 (N_43757,N_35494,N_35037);
or U43758 (N_43758,N_39541,N_38868);
nand U43759 (N_43759,N_39515,N_39127);
and U43760 (N_43760,N_36139,N_38839);
nand U43761 (N_43761,N_37056,N_38225);
nand U43762 (N_43762,N_36769,N_38141);
nor U43763 (N_43763,N_35209,N_37337);
and U43764 (N_43764,N_35495,N_36072);
xor U43765 (N_43765,N_36804,N_37556);
or U43766 (N_43766,N_37878,N_35753);
nor U43767 (N_43767,N_35796,N_36134);
or U43768 (N_43768,N_36901,N_37455);
or U43769 (N_43769,N_39848,N_37151);
nor U43770 (N_43770,N_38377,N_36834);
nand U43771 (N_43771,N_37693,N_39115);
xor U43772 (N_43772,N_35078,N_38576);
xnor U43773 (N_43773,N_38393,N_35307);
or U43774 (N_43774,N_38757,N_39923);
nor U43775 (N_43775,N_39414,N_37187);
or U43776 (N_43776,N_35212,N_36004);
nand U43777 (N_43777,N_37981,N_39826);
nand U43778 (N_43778,N_38135,N_38020);
or U43779 (N_43779,N_36463,N_36011);
nor U43780 (N_43780,N_39134,N_35398);
and U43781 (N_43781,N_39622,N_37662);
xor U43782 (N_43782,N_37759,N_39913);
nand U43783 (N_43783,N_35295,N_36140);
and U43784 (N_43784,N_39310,N_39954);
nand U43785 (N_43785,N_39364,N_38779);
nand U43786 (N_43786,N_39599,N_38913);
nand U43787 (N_43787,N_35755,N_35171);
nor U43788 (N_43788,N_36123,N_39119);
xor U43789 (N_43789,N_36841,N_37792);
nand U43790 (N_43790,N_38627,N_37038);
nor U43791 (N_43791,N_36291,N_37648);
xnor U43792 (N_43792,N_36033,N_39657);
or U43793 (N_43793,N_35207,N_39244);
nor U43794 (N_43794,N_35737,N_37542);
and U43795 (N_43795,N_35565,N_39483);
and U43796 (N_43796,N_39564,N_38885);
nor U43797 (N_43797,N_39932,N_36306);
nand U43798 (N_43798,N_35497,N_39336);
or U43799 (N_43799,N_39735,N_37296);
nor U43800 (N_43800,N_39442,N_39489);
nor U43801 (N_43801,N_39475,N_39219);
and U43802 (N_43802,N_39788,N_37319);
and U43803 (N_43803,N_37187,N_36444);
or U43804 (N_43804,N_35581,N_38356);
xor U43805 (N_43805,N_38145,N_35474);
or U43806 (N_43806,N_38452,N_36231);
nor U43807 (N_43807,N_36321,N_39254);
or U43808 (N_43808,N_36737,N_38673);
nand U43809 (N_43809,N_38514,N_37157);
xnor U43810 (N_43810,N_37612,N_38428);
nor U43811 (N_43811,N_39553,N_35439);
nor U43812 (N_43812,N_37446,N_39235);
xor U43813 (N_43813,N_39159,N_39127);
nand U43814 (N_43814,N_39229,N_35512);
xor U43815 (N_43815,N_36752,N_37064);
xnor U43816 (N_43816,N_37898,N_37118);
and U43817 (N_43817,N_35283,N_39134);
and U43818 (N_43818,N_36024,N_38267);
xnor U43819 (N_43819,N_37941,N_37432);
nand U43820 (N_43820,N_39196,N_37142);
and U43821 (N_43821,N_35940,N_36215);
and U43822 (N_43822,N_35083,N_38300);
or U43823 (N_43823,N_35208,N_36849);
xor U43824 (N_43824,N_37418,N_38997);
and U43825 (N_43825,N_38110,N_37489);
and U43826 (N_43826,N_36482,N_35093);
nor U43827 (N_43827,N_37263,N_37497);
and U43828 (N_43828,N_35336,N_36565);
nor U43829 (N_43829,N_39963,N_36417);
nand U43830 (N_43830,N_36897,N_35386);
nor U43831 (N_43831,N_36734,N_37703);
xor U43832 (N_43832,N_37729,N_37903);
nand U43833 (N_43833,N_38005,N_37500);
nand U43834 (N_43834,N_35985,N_37610);
nand U43835 (N_43835,N_38218,N_35265);
xor U43836 (N_43836,N_38183,N_35870);
nor U43837 (N_43837,N_39710,N_35476);
or U43838 (N_43838,N_39406,N_39850);
nor U43839 (N_43839,N_37202,N_35681);
and U43840 (N_43840,N_35486,N_36882);
or U43841 (N_43841,N_36907,N_35025);
xor U43842 (N_43842,N_37896,N_38611);
or U43843 (N_43843,N_37915,N_38274);
nand U43844 (N_43844,N_35993,N_39375);
or U43845 (N_43845,N_39351,N_39748);
xor U43846 (N_43846,N_36039,N_38879);
nor U43847 (N_43847,N_38396,N_35510);
and U43848 (N_43848,N_37732,N_35764);
xnor U43849 (N_43849,N_35425,N_39187);
or U43850 (N_43850,N_37726,N_38214);
xnor U43851 (N_43851,N_37007,N_37574);
or U43852 (N_43852,N_38451,N_38588);
xnor U43853 (N_43853,N_39293,N_36497);
and U43854 (N_43854,N_37068,N_36911);
xor U43855 (N_43855,N_39669,N_36149);
or U43856 (N_43856,N_37607,N_38274);
and U43857 (N_43857,N_38740,N_36240);
nor U43858 (N_43858,N_39562,N_36918);
or U43859 (N_43859,N_39695,N_35748);
nor U43860 (N_43860,N_35536,N_37135);
nor U43861 (N_43861,N_36451,N_37610);
or U43862 (N_43862,N_37440,N_38803);
nand U43863 (N_43863,N_37691,N_37031);
and U43864 (N_43864,N_38220,N_39011);
or U43865 (N_43865,N_39136,N_36667);
and U43866 (N_43866,N_35623,N_38953);
nand U43867 (N_43867,N_38969,N_39500);
xnor U43868 (N_43868,N_37600,N_36850);
nor U43869 (N_43869,N_37847,N_39215);
nand U43870 (N_43870,N_36739,N_39852);
and U43871 (N_43871,N_39878,N_36558);
or U43872 (N_43872,N_38229,N_38561);
and U43873 (N_43873,N_35052,N_36335);
or U43874 (N_43874,N_37618,N_37087);
nor U43875 (N_43875,N_39996,N_37088);
xnor U43876 (N_43876,N_39629,N_38692);
nor U43877 (N_43877,N_39950,N_39752);
or U43878 (N_43878,N_36945,N_35697);
and U43879 (N_43879,N_37136,N_39062);
and U43880 (N_43880,N_35298,N_35507);
xnor U43881 (N_43881,N_36421,N_37505);
and U43882 (N_43882,N_39602,N_35598);
nor U43883 (N_43883,N_38372,N_36428);
or U43884 (N_43884,N_39082,N_38741);
nand U43885 (N_43885,N_35432,N_38019);
xnor U43886 (N_43886,N_37652,N_37533);
and U43887 (N_43887,N_37270,N_35576);
and U43888 (N_43888,N_37672,N_36346);
nand U43889 (N_43889,N_36060,N_35442);
nand U43890 (N_43890,N_36237,N_36247);
nor U43891 (N_43891,N_39474,N_39025);
and U43892 (N_43892,N_37463,N_35091);
nor U43893 (N_43893,N_36030,N_36670);
nor U43894 (N_43894,N_37704,N_36614);
or U43895 (N_43895,N_35821,N_38330);
nand U43896 (N_43896,N_36620,N_37732);
xnor U43897 (N_43897,N_39414,N_38587);
xor U43898 (N_43898,N_38865,N_39904);
nor U43899 (N_43899,N_35479,N_38607);
and U43900 (N_43900,N_37831,N_35953);
nand U43901 (N_43901,N_37180,N_39888);
nand U43902 (N_43902,N_36564,N_35384);
nand U43903 (N_43903,N_36627,N_38909);
or U43904 (N_43904,N_38436,N_35316);
and U43905 (N_43905,N_39002,N_36057);
nor U43906 (N_43906,N_35921,N_39886);
nor U43907 (N_43907,N_35619,N_38123);
and U43908 (N_43908,N_38413,N_36909);
and U43909 (N_43909,N_37901,N_36266);
and U43910 (N_43910,N_39516,N_39629);
nor U43911 (N_43911,N_39361,N_36101);
and U43912 (N_43912,N_38111,N_38858);
and U43913 (N_43913,N_37910,N_38622);
nor U43914 (N_43914,N_39649,N_39412);
nor U43915 (N_43915,N_37170,N_37146);
xnor U43916 (N_43916,N_36159,N_35346);
xor U43917 (N_43917,N_38046,N_35831);
and U43918 (N_43918,N_35066,N_37615);
nand U43919 (N_43919,N_37369,N_36339);
nor U43920 (N_43920,N_39896,N_39318);
nor U43921 (N_43921,N_37274,N_39006);
xor U43922 (N_43922,N_37743,N_39841);
and U43923 (N_43923,N_37933,N_39205);
and U43924 (N_43924,N_35316,N_36895);
or U43925 (N_43925,N_38521,N_39465);
xor U43926 (N_43926,N_38772,N_37587);
xor U43927 (N_43927,N_37735,N_35591);
nor U43928 (N_43928,N_35857,N_35567);
xnor U43929 (N_43929,N_36306,N_35444);
or U43930 (N_43930,N_35832,N_36098);
nand U43931 (N_43931,N_36884,N_35519);
nand U43932 (N_43932,N_39908,N_35767);
nand U43933 (N_43933,N_39848,N_37035);
or U43934 (N_43934,N_39385,N_38536);
xnor U43935 (N_43935,N_35989,N_35523);
xor U43936 (N_43936,N_35479,N_36007);
and U43937 (N_43937,N_37658,N_36739);
or U43938 (N_43938,N_36387,N_38505);
nand U43939 (N_43939,N_38081,N_38007);
or U43940 (N_43940,N_36065,N_36464);
nor U43941 (N_43941,N_39164,N_36238);
nor U43942 (N_43942,N_36779,N_36584);
or U43943 (N_43943,N_35867,N_37402);
nor U43944 (N_43944,N_39537,N_37918);
nand U43945 (N_43945,N_35164,N_36793);
nand U43946 (N_43946,N_39157,N_35413);
nor U43947 (N_43947,N_36881,N_37203);
nand U43948 (N_43948,N_35500,N_37883);
nor U43949 (N_43949,N_37764,N_39844);
xnor U43950 (N_43950,N_35039,N_37029);
xor U43951 (N_43951,N_36922,N_38075);
nand U43952 (N_43952,N_39398,N_37594);
xor U43953 (N_43953,N_39120,N_37184);
nand U43954 (N_43954,N_39884,N_38593);
xnor U43955 (N_43955,N_39213,N_39921);
or U43956 (N_43956,N_38542,N_35365);
nor U43957 (N_43957,N_36070,N_35821);
nand U43958 (N_43958,N_36709,N_37002);
and U43959 (N_43959,N_39780,N_35191);
or U43960 (N_43960,N_35979,N_38672);
and U43961 (N_43961,N_36821,N_36966);
nor U43962 (N_43962,N_37080,N_39379);
nand U43963 (N_43963,N_39595,N_36114);
nand U43964 (N_43964,N_36143,N_36015);
xnor U43965 (N_43965,N_37795,N_39798);
or U43966 (N_43966,N_36123,N_39187);
or U43967 (N_43967,N_38684,N_35038);
nor U43968 (N_43968,N_39727,N_39904);
or U43969 (N_43969,N_36818,N_39720);
or U43970 (N_43970,N_37741,N_38589);
nand U43971 (N_43971,N_39416,N_36437);
and U43972 (N_43972,N_39318,N_38085);
or U43973 (N_43973,N_37943,N_36255);
or U43974 (N_43974,N_39005,N_37553);
or U43975 (N_43975,N_35179,N_38358);
nand U43976 (N_43976,N_38032,N_35646);
xnor U43977 (N_43977,N_36170,N_38012);
nor U43978 (N_43978,N_37928,N_35767);
xnor U43979 (N_43979,N_36525,N_37338);
or U43980 (N_43980,N_36962,N_38827);
xnor U43981 (N_43981,N_39785,N_36155);
nor U43982 (N_43982,N_37675,N_39866);
nand U43983 (N_43983,N_36528,N_35396);
and U43984 (N_43984,N_35361,N_39128);
nand U43985 (N_43985,N_36433,N_35496);
xor U43986 (N_43986,N_38967,N_35772);
nand U43987 (N_43987,N_39232,N_38290);
nor U43988 (N_43988,N_39128,N_35676);
xnor U43989 (N_43989,N_39869,N_38752);
nand U43990 (N_43990,N_36576,N_36680);
nor U43991 (N_43991,N_35416,N_36203);
and U43992 (N_43992,N_38248,N_39177);
nand U43993 (N_43993,N_36373,N_38026);
or U43994 (N_43994,N_36290,N_35666);
or U43995 (N_43995,N_36330,N_35814);
xnor U43996 (N_43996,N_39984,N_39529);
xnor U43997 (N_43997,N_37436,N_38483);
xnor U43998 (N_43998,N_35993,N_35493);
or U43999 (N_43999,N_38945,N_37727);
nor U44000 (N_44000,N_37429,N_37670);
or U44001 (N_44001,N_38036,N_37844);
nor U44002 (N_44002,N_36310,N_38148);
and U44003 (N_44003,N_35869,N_35231);
xor U44004 (N_44004,N_36974,N_37898);
xor U44005 (N_44005,N_38711,N_36642);
and U44006 (N_44006,N_39170,N_39166);
nand U44007 (N_44007,N_36372,N_36568);
nor U44008 (N_44008,N_37804,N_37228);
or U44009 (N_44009,N_38235,N_35639);
or U44010 (N_44010,N_36786,N_38104);
nand U44011 (N_44011,N_39127,N_36012);
xnor U44012 (N_44012,N_35232,N_36973);
and U44013 (N_44013,N_36556,N_36317);
xnor U44014 (N_44014,N_39022,N_39483);
nor U44015 (N_44015,N_38553,N_38970);
nor U44016 (N_44016,N_39449,N_39262);
nor U44017 (N_44017,N_38704,N_39159);
or U44018 (N_44018,N_37301,N_35021);
or U44019 (N_44019,N_36116,N_36361);
nor U44020 (N_44020,N_39423,N_37999);
or U44021 (N_44021,N_35068,N_38285);
or U44022 (N_44022,N_37498,N_35295);
and U44023 (N_44023,N_38840,N_37284);
or U44024 (N_44024,N_38551,N_35869);
xor U44025 (N_44025,N_36341,N_35971);
xnor U44026 (N_44026,N_39045,N_38773);
nand U44027 (N_44027,N_37392,N_38234);
nor U44028 (N_44028,N_37524,N_38127);
xnor U44029 (N_44029,N_39108,N_36076);
and U44030 (N_44030,N_37139,N_38603);
and U44031 (N_44031,N_38548,N_37762);
or U44032 (N_44032,N_39049,N_38118);
nand U44033 (N_44033,N_38107,N_39938);
and U44034 (N_44034,N_37256,N_38802);
xor U44035 (N_44035,N_35319,N_38833);
nand U44036 (N_44036,N_38053,N_39510);
xor U44037 (N_44037,N_37659,N_38988);
and U44038 (N_44038,N_35724,N_36273);
or U44039 (N_44039,N_35100,N_38889);
nor U44040 (N_44040,N_36015,N_39607);
nor U44041 (N_44041,N_38563,N_37866);
nand U44042 (N_44042,N_35946,N_37580);
nand U44043 (N_44043,N_39701,N_37359);
nand U44044 (N_44044,N_35016,N_36421);
nor U44045 (N_44045,N_37970,N_37696);
or U44046 (N_44046,N_37433,N_35056);
nand U44047 (N_44047,N_35739,N_35153);
nand U44048 (N_44048,N_37345,N_37539);
xnor U44049 (N_44049,N_37150,N_39942);
nor U44050 (N_44050,N_38062,N_37562);
nor U44051 (N_44051,N_37730,N_37497);
nor U44052 (N_44052,N_36776,N_36829);
or U44053 (N_44053,N_36894,N_37237);
nand U44054 (N_44054,N_39736,N_36021);
xnor U44055 (N_44055,N_37867,N_38730);
nand U44056 (N_44056,N_39726,N_35805);
nand U44057 (N_44057,N_36843,N_39835);
nor U44058 (N_44058,N_39382,N_37373);
and U44059 (N_44059,N_35464,N_38564);
and U44060 (N_44060,N_37968,N_36742);
or U44061 (N_44061,N_38268,N_38667);
and U44062 (N_44062,N_38795,N_35877);
nor U44063 (N_44063,N_39435,N_36457);
or U44064 (N_44064,N_36329,N_39018);
and U44065 (N_44065,N_35699,N_37257);
xor U44066 (N_44066,N_35069,N_36504);
and U44067 (N_44067,N_39541,N_36044);
nand U44068 (N_44068,N_38017,N_38709);
or U44069 (N_44069,N_37014,N_35214);
or U44070 (N_44070,N_37306,N_38733);
and U44071 (N_44071,N_37702,N_37974);
nand U44072 (N_44072,N_36754,N_38599);
and U44073 (N_44073,N_38150,N_36031);
or U44074 (N_44074,N_37330,N_35429);
and U44075 (N_44075,N_39218,N_39666);
or U44076 (N_44076,N_39515,N_35013);
or U44077 (N_44077,N_37435,N_39341);
nor U44078 (N_44078,N_36966,N_36707);
or U44079 (N_44079,N_37816,N_38685);
or U44080 (N_44080,N_38721,N_37896);
or U44081 (N_44081,N_36081,N_37363);
or U44082 (N_44082,N_35622,N_37949);
and U44083 (N_44083,N_36154,N_38092);
nor U44084 (N_44084,N_35549,N_38397);
or U44085 (N_44085,N_38007,N_38464);
xnor U44086 (N_44086,N_38573,N_38496);
or U44087 (N_44087,N_35884,N_38009);
nand U44088 (N_44088,N_37608,N_36983);
or U44089 (N_44089,N_37115,N_39792);
xnor U44090 (N_44090,N_35818,N_36829);
or U44091 (N_44091,N_36942,N_39602);
and U44092 (N_44092,N_35831,N_38073);
and U44093 (N_44093,N_36054,N_35631);
xnor U44094 (N_44094,N_36604,N_38514);
xnor U44095 (N_44095,N_37399,N_39113);
nand U44096 (N_44096,N_39725,N_39261);
or U44097 (N_44097,N_35304,N_35750);
xnor U44098 (N_44098,N_39538,N_35757);
or U44099 (N_44099,N_35831,N_37013);
and U44100 (N_44100,N_37224,N_37842);
nand U44101 (N_44101,N_39439,N_35636);
or U44102 (N_44102,N_35279,N_35020);
or U44103 (N_44103,N_38476,N_39665);
or U44104 (N_44104,N_39833,N_36180);
xnor U44105 (N_44105,N_39017,N_39344);
nor U44106 (N_44106,N_36163,N_36319);
nor U44107 (N_44107,N_36976,N_38598);
and U44108 (N_44108,N_36486,N_37089);
nand U44109 (N_44109,N_36060,N_38872);
or U44110 (N_44110,N_35700,N_36756);
nor U44111 (N_44111,N_38277,N_36934);
nand U44112 (N_44112,N_35002,N_36095);
nor U44113 (N_44113,N_38796,N_35932);
nand U44114 (N_44114,N_38379,N_37921);
nand U44115 (N_44115,N_35792,N_35995);
nand U44116 (N_44116,N_38331,N_38879);
nand U44117 (N_44117,N_36338,N_35073);
and U44118 (N_44118,N_37111,N_36505);
or U44119 (N_44119,N_36726,N_36107);
and U44120 (N_44120,N_35402,N_35734);
xnor U44121 (N_44121,N_37343,N_36325);
and U44122 (N_44122,N_35403,N_38448);
nor U44123 (N_44123,N_36821,N_36647);
xnor U44124 (N_44124,N_35526,N_39972);
and U44125 (N_44125,N_36513,N_36778);
and U44126 (N_44126,N_39412,N_37332);
and U44127 (N_44127,N_36609,N_35048);
nand U44128 (N_44128,N_39077,N_36874);
and U44129 (N_44129,N_39479,N_37064);
nor U44130 (N_44130,N_38945,N_39405);
xnor U44131 (N_44131,N_37177,N_37053);
nor U44132 (N_44132,N_36924,N_37059);
nand U44133 (N_44133,N_38324,N_35782);
and U44134 (N_44134,N_39828,N_38541);
and U44135 (N_44135,N_35299,N_35277);
nor U44136 (N_44136,N_38037,N_39998);
nor U44137 (N_44137,N_38039,N_39536);
and U44138 (N_44138,N_38570,N_37513);
xor U44139 (N_44139,N_37691,N_39786);
nand U44140 (N_44140,N_36159,N_37098);
nand U44141 (N_44141,N_39462,N_36490);
or U44142 (N_44142,N_37639,N_35212);
nor U44143 (N_44143,N_38925,N_35105);
nand U44144 (N_44144,N_35044,N_39194);
xor U44145 (N_44145,N_37465,N_35428);
nor U44146 (N_44146,N_37041,N_36851);
or U44147 (N_44147,N_37310,N_39479);
or U44148 (N_44148,N_39290,N_39416);
xor U44149 (N_44149,N_39788,N_39686);
xnor U44150 (N_44150,N_38779,N_38063);
nand U44151 (N_44151,N_38185,N_35506);
xnor U44152 (N_44152,N_35492,N_38246);
nand U44153 (N_44153,N_37674,N_39051);
nor U44154 (N_44154,N_38167,N_38158);
nor U44155 (N_44155,N_36800,N_37559);
and U44156 (N_44156,N_39892,N_35057);
nand U44157 (N_44157,N_36372,N_35017);
and U44158 (N_44158,N_35739,N_37393);
nor U44159 (N_44159,N_37969,N_36025);
nor U44160 (N_44160,N_35098,N_38077);
and U44161 (N_44161,N_39670,N_39499);
nor U44162 (N_44162,N_37244,N_37424);
and U44163 (N_44163,N_36871,N_35782);
or U44164 (N_44164,N_35987,N_37117);
xor U44165 (N_44165,N_37862,N_36528);
nor U44166 (N_44166,N_39034,N_37654);
nand U44167 (N_44167,N_37118,N_37899);
nand U44168 (N_44168,N_35623,N_38795);
xor U44169 (N_44169,N_38653,N_35898);
xnor U44170 (N_44170,N_38236,N_39220);
nand U44171 (N_44171,N_35329,N_38684);
and U44172 (N_44172,N_38755,N_39061);
and U44173 (N_44173,N_38581,N_35861);
nand U44174 (N_44174,N_36188,N_36373);
nor U44175 (N_44175,N_35047,N_38610);
nand U44176 (N_44176,N_38547,N_36886);
nor U44177 (N_44177,N_36294,N_37585);
and U44178 (N_44178,N_37220,N_37219);
nor U44179 (N_44179,N_39201,N_39483);
and U44180 (N_44180,N_35317,N_39464);
or U44181 (N_44181,N_36226,N_38405);
xor U44182 (N_44182,N_35865,N_37857);
or U44183 (N_44183,N_39045,N_35069);
nand U44184 (N_44184,N_35902,N_36801);
nor U44185 (N_44185,N_38856,N_37379);
nand U44186 (N_44186,N_36675,N_36581);
and U44187 (N_44187,N_38616,N_37725);
and U44188 (N_44188,N_35157,N_37659);
nand U44189 (N_44189,N_39385,N_38756);
nor U44190 (N_44190,N_37050,N_38901);
and U44191 (N_44191,N_36833,N_39331);
and U44192 (N_44192,N_36468,N_38261);
nand U44193 (N_44193,N_39157,N_38506);
nand U44194 (N_44194,N_37748,N_35116);
nand U44195 (N_44195,N_38800,N_37505);
nor U44196 (N_44196,N_35593,N_38349);
nor U44197 (N_44197,N_39067,N_36371);
nand U44198 (N_44198,N_39812,N_39295);
nor U44199 (N_44199,N_39266,N_36087);
and U44200 (N_44200,N_38752,N_36407);
or U44201 (N_44201,N_35900,N_38868);
xor U44202 (N_44202,N_36245,N_39170);
or U44203 (N_44203,N_35352,N_39249);
xnor U44204 (N_44204,N_35258,N_35423);
xnor U44205 (N_44205,N_38396,N_37286);
xor U44206 (N_44206,N_36770,N_38456);
nor U44207 (N_44207,N_36462,N_35937);
nand U44208 (N_44208,N_38171,N_37988);
or U44209 (N_44209,N_37005,N_35427);
and U44210 (N_44210,N_36759,N_38587);
or U44211 (N_44211,N_36224,N_37345);
and U44212 (N_44212,N_39985,N_35911);
or U44213 (N_44213,N_38392,N_38289);
and U44214 (N_44214,N_36363,N_37244);
xnor U44215 (N_44215,N_38886,N_36870);
nand U44216 (N_44216,N_35802,N_39368);
or U44217 (N_44217,N_39462,N_39605);
nor U44218 (N_44218,N_37367,N_36086);
or U44219 (N_44219,N_36021,N_38964);
or U44220 (N_44220,N_35506,N_35414);
and U44221 (N_44221,N_36739,N_37266);
and U44222 (N_44222,N_35260,N_39684);
nor U44223 (N_44223,N_36009,N_38562);
nand U44224 (N_44224,N_39042,N_39872);
nor U44225 (N_44225,N_37023,N_39621);
nand U44226 (N_44226,N_38170,N_35575);
nand U44227 (N_44227,N_35650,N_39807);
xor U44228 (N_44228,N_38071,N_35900);
nor U44229 (N_44229,N_37954,N_39153);
nor U44230 (N_44230,N_38272,N_36590);
or U44231 (N_44231,N_37591,N_36879);
nor U44232 (N_44232,N_35864,N_39480);
and U44233 (N_44233,N_36086,N_35796);
and U44234 (N_44234,N_36488,N_37635);
or U44235 (N_44235,N_36818,N_35619);
nand U44236 (N_44236,N_37092,N_36302);
nand U44237 (N_44237,N_36087,N_37286);
xor U44238 (N_44238,N_39623,N_39351);
or U44239 (N_44239,N_37148,N_36332);
or U44240 (N_44240,N_37868,N_39815);
or U44241 (N_44241,N_38055,N_38321);
xnor U44242 (N_44242,N_39363,N_38837);
nor U44243 (N_44243,N_36174,N_39094);
xnor U44244 (N_44244,N_36845,N_39925);
nor U44245 (N_44245,N_36076,N_38958);
or U44246 (N_44246,N_38534,N_38342);
nand U44247 (N_44247,N_37821,N_36240);
xnor U44248 (N_44248,N_39492,N_38586);
nand U44249 (N_44249,N_35039,N_35073);
xor U44250 (N_44250,N_39078,N_38792);
nor U44251 (N_44251,N_36722,N_36704);
or U44252 (N_44252,N_38513,N_36513);
nor U44253 (N_44253,N_38829,N_35828);
and U44254 (N_44254,N_39008,N_39739);
and U44255 (N_44255,N_37384,N_37783);
nor U44256 (N_44256,N_38780,N_39938);
or U44257 (N_44257,N_36321,N_39034);
nor U44258 (N_44258,N_37779,N_39545);
or U44259 (N_44259,N_39451,N_35375);
nor U44260 (N_44260,N_35748,N_39432);
xor U44261 (N_44261,N_35936,N_36550);
nand U44262 (N_44262,N_37702,N_35754);
nand U44263 (N_44263,N_37287,N_39937);
xnor U44264 (N_44264,N_35654,N_36826);
nand U44265 (N_44265,N_38299,N_39058);
or U44266 (N_44266,N_36454,N_37729);
or U44267 (N_44267,N_38073,N_38793);
nand U44268 (N_44268,N_37483,N_35124);
nand U44269 (N_44269,N_38659,N_39334);
or U44270 (N_44270,N_38918,N_38832);
nor U44271 (N_44271,N_38169,N_36875);
nor U44272 (N_44272,N_39079,N_37778);
xor U44273 (N_44273,N_38655,N_37942);
xor U44274 (N_44274,N_35183,N_37726);
xnor U44275 (N_44275,N_36314,N_38984);
nor U44276 (N_44276,N_39426,N_37915);
xor U44277 (N_44277,N_37228,N_37945);
or U44278 (N_44278,N_37916,N_37305);
and U44279 (N_44279,N_39090,N_36080);
or U44280 (N_44280,N_37178,N_37993);
or U44281 (N_44281,N_37341,N_35995);
nand U44282 (N_44282,N_38550,N_36545);
nand U44283 (N_44283,N_39453,N_39346);
xnor U44284 (N_44284,N_37024,N_38775);
and U44285 (N_44285,N_38173,N_35253);
nor U44286 (N_44286,N_36679,N_36240);
or U44287 (N_44287,N_38469,N_38341);
nor U44288 (N_44288,N_39427,N_37034);
nor U44289 (N_44289,N_39072,N_35504);
and U44290 (N_44290,N_37966,N_38028);
xor U44291 (N_44291,N_35973,N_35043);
nand U44292 (N_44292,N_35949,N_36637);
xnor U44293 (N_44293,N_39772,N_39055);
and U44294 (N_44294,N_38421,N_39276);
or U44295 (N_44295,N_35654,N_39308);
nor U44296 (N_44296,N_39241,N_36124);
nor U44297 (N_44297,N_39434,N_39591);
or U44298 (N_44298,N_36101,N_37536);
and U44299 (N_44299,N_38544,N_35604);
xnor U44300 (N_44300,N_39139,N_39717);
nor U44301 (N_44301,N_37550,N_36495);
nor U44302 (N_44302,N_39167,N_37719);
and U44303 (N_44303,N_38024,N_35050);
nor U44304 (N_44304,N_35325,N_38500);
nand U44305 (N_44305,N_39072,N_35408);
xnor U44306 (N_44306,N_39596,N_38759);
xor U44307 (N_44307,N_35953,N_39118);
or U44308 (N_44308,N_38344,N_35684);
nor U44309 (N_44309,N_38979,N_35927);
nor U44310 (N_44310,N_36650,N_39380);
nor U44311 (N_44311,N_39014,N_36831);
xnor U44312 (N_44312,N_35731,N_35079);
nor U44313 (N_44313,N_39983,N_36425);
and U44314 (N_44314,N_39043,N_39283);
xnor U44315 (N_44315,N_36037,N_36565);
and U44316 (N_44316,N_38774,N_35291);
nand U44317 (N_44317,N_38956,N_35011);
or U44318 (N_44318,N_36273,N_36588);
nand U44319 (N_44319,N_35922,N_38682);
or U44320 (N_44320,N_38267,N_38012);
and U44321 (N_44321,N_39597,N_37940);
xnor U44322 (N_44322,N_36220,N_35888);
or U44323 (N_44323,N_35195,N_39214);
and U44324 (N_44324,N_36566,N_39804);
and U44325 (N_44325,N_35214,N_38842);
and U44326 (N_44326,N_35026,N_39636);
and U44327 (N_44327,N_36426,N_37902);
and U44328 (N_44328,N_38176,N_37730);
and U44329 (N_44329,N_39689,N_36315);
xnor U44330 (N_44330,N_37117,N_38937);
xnor U44331 (N_44331,N_37685,N_36083);
nand U44332 (N_44332,N_37020,N_38488);
nand U44333 (N_44333,N_37212,N_38666);
or U44334 (N_44334,N_36674,N_35382);
nor U44335 (N_44335,N_35649,N_39532);
nand U44336 (N_44336,N_35571,N_37468);
and U44337 (N_44337,N_38352,N_36346);
nand U44338 (N_44338,N_35342,N_39655);
xor U44339 (N_44339,N_38931,N_35641);
nor U44340 (N_44340,N_39108,N_35414);
xnor U44341 (N_44341,N_37803,N_36397);
xor U44342 (N_44342,N_36850,N_38733);
nor U44343 (N_44343,N_38853,N_36078);
nor U44344 (N_44344,N_37301,N_36011);
nand U44345 (N_44345,N_36278,N_36534);
nand U44346 (N_44346,N_37270,N_39798);
and U44347 (N_44347,N_36952,N_37714);
or U44348 (N_44348,N_36994,N_37448);
and U44349 (N_44349,N_36568,N_38330);
and U44350 (N_44350,N_37459,N_37615);
xnor U44351 (N_44351,N_36936,N_36881);
nor U44352 (N_44352,N_39281,N_37413);
nor U44353 (N_44353,N_36652,N_37762);
nand U44354 (N_44354,N_38944,N_36132);
or U44355 (N_44355,N_35695,N_37941);
xor U44356 (N_44356,N_37760,N_38337);
or U44357 (N_44357,N_35868,N_36090);
and U44358 (N_44358,N_39047,N_36613);
nand U44359 (N_44359,N_36080,N_37130);
and U44360 (N_44360,N_35771,N_39737);
and U44361 (N_44361,N_38295,N_35955);
xor U44362 (N_44362,N_37145,N_37266);
and U44363 (N_44363,N_35807,N_35164);
nand U44364 (N_44364,N_36851,N_38928);
and U44365 (N_44365,N_36361,N_39068);
and U44366 (N_44366,N_36077,N_35952);
nor U44367 (N_44367,N_38792,N_35945);
nor U44368 (N_44368,N_37363,N_35066);
or U44369 (N_44369,N_38612,N_36871);
or U44370 (N_44370,N_37403,N_38632);
xnor U44371 (N_44371,N_38323,N_39815);
nand U44372 (N_44372,N_35648,N_37648);
nand U44373 (N_44373,N_39665,N_38943);
nor U44374 (N_44374,N_35910,N_35576);
nand U44375 (N_44375,N_39698,N_39114);
nand U44376 (N_44376,N_38084,N_35981);
or U44377 (N_44377,N_39334,N_39589);
or U44378 (N_44378,N_37003,N_38399);
xor U44379 (N_44379,N_36250,N_35817);
xnor U44380 (N_44380,N_37388,N_36083);
nand U44381 (N_44381,N_35673,N_35851);
and U44382 (N_44382,N_36932,N_36529);
and U44383 (N_44383,N_36858,N_38460);
nor U44384 (N_44384,N_35320,N_37999);
and U44385 (N_44385,N_35738,N_39191);
nand U44386 (N_44386,N_36701,N_39575);
xnor U44387 (N_44387,N_37011,N_37282);
and U44388 (N_44388,N_37362,N_35290);
xnor U44389 (N_44389,N_38602,N_39224);
xnor U44390 (N_44390,N_38575,N_35407);
or U44391 (N_44391,N_38864,N_35701);
xnor U44392 (N_44392,N_39493,N_37453);
nor U44393 (N_44393,N_37966,N_39078);
nor U44394 (N_44394,N_36250,N_37536);
and U44395 (N_44395,N_39188,N_36595);
nand U44396 (N_44396,N_37660,N_36873);
and U44397 (N_44397,N_35282,N_36519);
nand U44398 (N_44398,N_36182,N_38717);
xnor U44399 (N_44399,N_36594,N_37790);
or U44400 (N_44400,N_39855,N_38947);
and U44401 (N_44401,N_36962,N_38517);
nand U44402 (N_44402,N_37456,N_38818);
xnor U44403 (N_44403,N_37237,N_35181);
or U44404 (N_44404,N_36994,N_36723);
xnor U44405 (N_44405,N_37273,N_39585);
nor U44406 (N_44406,N_36467,N_38561);
xnor U44407 (N_44407,N_35363,N_35004);
nor U44408 (N_44408,N_39512,N_38579);
xor U44409 (N_44409,N_37417,N_36301);
nor U44410 (N_44410,N_35429,N_36783);
nand U44411 (N_44411,N_36221,N_38043);
and U44412 (N_44412,N_37555,N_38277);
and U44413 (N_44413,N_35598,N_37103);
nor U44414 (N_44414,N_36840,N_39225);
and U44415 (N_44415,N_39363,N_36345);
or U44416 (N_44416,N_39709,N_37106);
and U44417 (N_44417,N_37690,N_38138);
and U44418 (N_44418,N_38013,N_37810);
and U44419 (N_44419,N_39423,N_35315);
or U44420 (N_44420,N_39988,N_36146);
xor U44421 (N_44421,N_35586,N_37981);
or U44422 (N_44422,N_37842,N_39345);
xnor U44423 (N_44423,N_37393,N_35475);
and U44424 (N_44424,N_36557,N_39381);
xor U44425 (N_44425,N_38904,N_35897);
nor U44426 (N_44426,N_39515,N_36517);
or U44427 (N_44427,N_37946,N_36097);
nor U44428 (N_44428,N_36446,N_37043);
and U44429 (N_44429,N_38671,N_36487);
nand U44430 (N_44430,N_39856,N_36173);
and U44431 (N_44431,N_35262,N_36993);
xor U44432 (N_44432,N_38220,N_38763);
xor U44433 (N_44433,N_39881,N_36651);
xor U44434 (N_44434,N_36176,N_39452);
or U44435 (N_44435,N_35138,N_35716);
nand U44436 (N_44436,N_36743,N_37147);
and U44437 (N_44437,N_38252,N_37612);
xnor U44438 (N_44438,N_36845,N_36193);
nor U44439 (N_44439,N_37926,N_35104);
and U44440 (N_44440,N_37742,N_35962);
and U44441 (N_44441,N_39989,N_37812);
xnor U44442 (N_44442,N_35724,N_38471);
nor U44443 (N_44443,N_35920,N_37627);
xor U44444 (N_44444,N_36893,N_38921);
nor U44445 (N_44445,N_37374,N_38711);
or U44446 (N_44446,N_35412,N_39436);
or U44447 (N_44447,N_37828,N_36177);
nor U44448 (N_44448,N_39008,N_39432);
nand U44449 (N_44449,N_39118,N_38259);
nor U44450 (N_44450,N_38980,N_36480);
xnor U44451 (N_44451,N_35727,N_35644);
nand U44452 (N_44452,N_36629,N_39625);
and U44453 (N_44453,N_35445,N_36426);
nor U44454 (N_44454,N_39413,N_37846);
or U44455 (N_44455,N_35170,N_38547);
nor U44456 (N_44456,N_37833,N_35094);
and U44457 (N_44457,N_36405,N_39066);
xor U44458 (N_44458,N_39380,N_39445);
and U44459 (N_44459,N_38379,N_38882);
xnor U44460 (N_44460,N_39382,N_38678);
nand U44461 (N_44461,N_36620,N_36791);
xnor U44462 (N_44462,N_35142,N_38158);
nor U44463 (N_44463,N_39518,N_37135);
and U44464 (N_44464,N_37666,N_36684);
and U44465 (N_44465,N_39440,N_38468);
nor U44466 (N_44466,N_37434,N_38155);
or U44467 (N_44467,N_35679,N_37390);
xor U44468 (N_44468,N_35834,N_36067);
or U44469 (N_44469,N_37742,N_36971);
nand U44470 (N_44470,N_39430,N_36407);
nand U44471 (N_44471,N_37033,N_36085);
and U44472 (N_44472,N_36325,N_35624);
and U44473 (N_44473,N_36135,N_39308);
or U44474 (N_44474,N_39504,N_37133);
or U44475 (N_44475,N_38592,N_37916);
xnor U44476 (N_44476,N_35642,N_38646);
nor U44477 (N_44477,N_35891,N_37938);
or U44478 (N_44478,N_37628,N_36451);
and U44479 (N_44479,N_38328,N_35625);
nor U44480 (N_44480,N_37863,N_38834);
nand U44481 (N_44481,N_39117,N_35350);
or U44482 (N_44482,N_37810,N_38165);
and U44483 (N_44483,N_38079,N_36465);
xor U44484 (N_44484,N_39928,N_39858);
and U44485 (N_44485,N_36786,N_36248);
nand U44486 (N_44486,N_35273,N_36810);
nand U44487 (N_44487,N_38812,N_35190);
nor U44488 (N_44488,N_37072,N_37550);
and U44489 (N_44489,N_38390,N_38737);
xnor U44490 (N_44490,N_37490,N_37204);
or U44491 (N_44491,N_35555,N_39983);
nand U44492 (N_44492,N_35657,N_39088);
or U44493 (N_44493,N_37991,N_38518);
nand U44494 (N_44494,N_38587,N_39936);
nor U44495 (N_44495,N_37529,N_35160);
nor U44496 (N_44496,N_37481,N_39619);
and U44497 (N_44497,N_36073,N_38897);
or U44498 (N_44498,N_37808,N_36803);
nand U44499 (N_44499,N_38282,N_36228);
and U44500 (N_44500,N_36101,N_38584);
nand U44501 (N_44501,N_37266,N_37206);
nand U44502 (N_44502,N_39318,N_39359);
nor U44503 (N_44503,N_36528,N_37348);
nor U44504 (N_44504,N_38174,N_36071);
nand U44505 (N_44505,N_37034,N_36589);
or U44506 (N_44506,N_38950,N_36445);
or U44507 (N_44507,N_35508,N_35263);
nor U44508 (N_44508,N_37905,N_35542);
nand U44509 (N_44509,N_39879,N_36748);
xnor U44510 (N_44510,N_39724,N_38755);
nor U44511 (N_44511,N_35255,N_37969);
and U44512 (N_44512,N_37496,N_36952);
or U44513 (N_44513,N_39409,N_37148);
nor U44514 (N_44514,N_37551,N_39423);
nand U44515 (N_44515,N_36075,N_37267);
and U44516 (N_44516,N_38929,N_36108);
nand U44517 (N_44517,N_36636,N_39278);
xnor U44518 (N_44518,N_35373,N_36030);
xor U44519 (N_44519,N_38627,N_38665);
xnor U44520 (N_44520,N_39016,N_37863);
nor U44521 (N_44521,N_35990,N_38422);
nand U44522 (N_44522,N_36721,N_38467);
xnor U44523 (N_44523,N_38926,N_38540);
nand U44524 (N_44524,N_39635,N_35008);
nor U44525 (N_44525,N_37063,N_36063);
or U44526 (N_44526,N_37734,N_36511);
or U44527 (N_44527,N_36198,N_36243);
xnor U44528 (N_44528,N_35626,N_36857);
and U44529 (N_44529,N_36803,N_37394);
or U44530 (N_44530,N_36019,N_39921);
nor U44531 (N_44531,N_36416,N_36090);
nor U44532 (N_44532,N_36748,N_36566);
nand U44533 (N_44533,N_38493,N_39425);
and U44534 (N_44534,N_36218,N_39118);
nor U44535 (N_44535,N_38397,N_35735);
xnor U44536 (N_44536,N_36160,N_37202);
nor U44537 (N_44537,N_36833,N_36024);
and U44538 (N_44538,N_36136,N_35651);
nand U44539 (N_44539,N_37085,N_37475);
and U44540 (N_44540,N_36145,N_39162);
and U44541 (N_44541,N_35952,N_39729);
or U44542 (N_44542,N_35202,N_35299);
or U44543 (N_44543,N_38675,N_36801);
or U44544 (N_44544,N_36054,N_38810);
xor U44545 (N_44545,N_36896,N_36257);
nor U44546 (N_44546,N_37196,N_38349);
or U44547 (N_44547,N_35456,N_35791);
or U44548 (N_44548,N_38328,N_35959);
xor U44549 (N_44549,N_38823,N_35994);
or U44550 (N_44550,N_38921,N_38893);
nor U44551 (N_44551,N_35960,N_35228);
nor U44552 (N_44552,N_36015,N_37776);
and U44553 (N_44553,N_36671,N_37989);
nor U44554 (N_44554,N_38974,N_39668);
or U44555 (N_44555,N_35594,N_36138);
nor U44556 (N_44556,N_35620,N_39236);
or U44557 (N_44557,N_37190,N_37630);
and U44558 (N_44558,N_37256,N_38850);
nor U44559 (N_44559,N_35423,N_39370);
xnor U44560 (N_44560,N_39959,N_39339);
nor U44561 (N_44561,N_39496,N_36412);
nand U44562 (N_44562,N_38105,N_35602);
xor U44563 (N_44563,N_35706,N_37844);
and U44564 (N_44564,N_35380,N_37768);
nand U44565 (N_44565,N_36408,N_39974);
nor U44566 (N_44566,N_35121,N_35015);
nor U44567 (N_44567,N_38251,N_38399);
nand U44568 (N_44568,N_39291,N_35334);
and U44569 (N_44569,N_38943,N_37646);
or U44570 (N_44570,N_36704,N_35255);
nor U44571 (N_44571,N_39800,N_37611);
nand U44572 (N_44572,N_39682,N_37089);
nand U44573 (N_44573,N_38820,N_35906);
or U44574 (N_44574,N_36393,N_36308);
nand U44575 (N_44575,N_38599,N_36506);
xor U44576 (N_44576,N_38958,N_39025);
nand U44577 (N_44577,N_39569,N_39296);
or U44578 (N_44578,N_36290,N_38628);
xnor U44579 (N_44579,N_35031,N_39044);
and U44580 (N_44580,N_37115,N_35102);
nand U44581 (N_44581,N_35061,N_39179);
or U44582 (N_44582,N_37389,N_36865);
nor U44583 (N_44583,N_38824,N_35271);
xor U44584 (N_44584,N_39433,N_37931);
nand U44585 (N_44585,N_36612,N_35939);
nand U44586 (N_44586,N_37741,N_36826);
xor U44587 (N_44587,N_35908,N_35289);
or U44588 (N_44588,N_37950,N_35861);
xor U44589 (N_44589,N_37114,N_36078);
nor U44590 (N_44590,N_37575,N_38672);
nand U44591 (N_44591,N_36630,N_38001);
or U44592 (N_44592,N_36161,N_37424);
xnor U44593 (N_44593,N_38611,N_36811);
xnor U44594 (N_44594,N_38108,N_36944);
nand U44595 (N_44595,N_35388,N_37191);
nor U44596 (N_44596,N_39417,N_39056);
nand U44597 (N_44597,N_36300,N_39797);
nor U44598 (N_44598,N_36891,N_36884);
xor U44599 (N_44599,N_38433,N_37552);
or U44600 (N_44600,N_35862,N_36131);
nor U44601 (N_44601,N_38127,N_38337);
or U44602 (N_44602,N_36613,N_39484);
and U44603 (N_44603,N_37413,N_39156);
nor U44604 (N_44604,N_36232,N_38161);
xor U44605 (N_44605,N_39893,N_36866);
xor U44606 (N_44606,N_39762,N_37964);
and U44607 (N_44607,N_37305,N_39393);
nor U44608 (N_44608,N_37680,N_36081);
nand U44609 (N_44609,N_37204,N_36786);
nand U44610 (N_44610,N_39573,N_37980);
nand U44611 (N_44611,N_37964,N_35550);
nand U44612 (N_44612,N_35128,N_39159);
nor U44613 (N_44613,N_38121,N_37924);
and U44614 (N_44614,N_37530,N_39713);
xor U44615 (N_44615,N_36755,N_39424);
and U44616 (N_44616,N_38389,N_35308);
xnor U44617 (N_44617,N_38610,N_38471);
xnor U44618 (N_44618,N_36168,N_37079);
and U44619 (N_44619,N_39522,N_38626);
xnor U44620 (N_44620,N_35653,N_37013);
xnor U44621 (N_44621,N_37390,N_37588);
and U44622 (N_44622,N_38407,N_37748);
or U44623 (N_44623,N_39844,N_39472);
and U44624 (N_44624,N_37140,N_38590);
xnor U44625 (N_44625,N_36290,N_38075);
nor U44626 (N_44626,N_38379,N_37601);
nand U44627 (N_44627,N_39133,N_38235);
or U44628 (N_44628,N_39892,N_37650);
and U44629 (N_44629,N_35572,N_37274);
or U44630 (N_44630,N_39648,N_36544);
nor U44631 (N_44631,N_37164,N_36545);
or U44632 (N_44632,N_36958,N_35469);
and U44633 (N_44633,N_39653,N_38576);
nand U44634 (N_44634,N_35033,N_35491);
nand U44635 (N_44635,N_35170,N_37454);
nor U44636 (N_44636,N_36511,N_39607);
and U44637 (N_44637,N_36862,N_36938);
or U44638 (N_44638,N_39561,N_35511);
or U44639 (N_44639,N_36211,N_35877);
nand U44640 (N_44640,N_35763,N_37567);
nor U44641 (N_44641,N_36712,N_36124);
or U44642 (N_44642,N_37990,N_35732);
and U44643 (N_44643,N_38035,N_37908);
nor U44644 (N_44644,N_38206,N_39453);
and U44645 (N_44645,N_37365,N_36906);
nor U44646 (N_44646,N_36165,N_36481);
nand U44647 (N_44647,N_36722,N_35855);
and U44648 (N_44648,N_37461,N_38202);
xor U44649 (N_44649,N_36176,N_35314);
or U44650 (N_44650,N_37444,N_37894);
and U44651 (N_44651,N_36130,N_35416);
nor U44652 (N_44652,N_36926,N_38444);
and U44653 (N_44653,N_35165,N_38325);
nand U44654 (N_44654,N_38690,N_37893);
nand U44655 (N_44655,N_37042,N_38242);
xnor U44656 (N_44656,N_35778,N_35398);
nor U44657 (N_44657,N_39799,N_35450);
and U44658 (N_44658,N_38385,N_39512);
nor U44659 (N_44659,N_38192,N_35086);
nor U44660 (N_44660,N_39358,N_37535);
nor U44661 (N_44661,N_35538,N_37303);
xnor U44662 (N_44662,N_37457,N_35872);
xnor U44663 (N_44663,N_37545,N_38478);
xor U44664 (N_44664,N_38267,N_36794);
nor U44665 (N_44665,N_38819,N_38972);
nand U44666 (N_44666,N_35805,N_37354);
xnor U44667 (N_44667,N_35490,N_39482);
and U44668 (N_44668,N_36505,N_39681);
nand U44669 (N_44669,N_39526,N_39161);
xor U44670 (N_44670,N_36576,N_37767);
and U44671 (N_44671,N_37279,N_36099);
or U44672 (N_44672,N_37715,N_35756);
xor U44673 (N_44673,N_36118,N_38833);
and U44674 (N_44674,N_35589,N_38297);
nor U44675 (N_44675,N_39069,N_36712);
and U44676 (N_44676,N_39318,N_36372);
or U44677 (N_44677,N_37947,N_35336);
or U44678 (N_44678,N_39357,N_37209);
or U44679 (N_44679,N_39227,N_36549);
nand U44680 (N_44680,N_38213,N_38937);
and U44681 (N_44681,N_38588,N_36728);
nand U44682 (N_44682,N_37178,N_38705);
nor U44683 (N_44683,N_39540,N_39654);
or U44684 (N_44684,N_38734,N_37330);
or U44685 (N_44685,N_38490,N_39867);
and U44686 (N_44686,N_35061,N_36280);
xor U44687 (N_44687,N_35155,N_35047);
nor U44688 (N_44688,N_35827,N_37458);
or U44689 (N_44689,N_37689,N_36348);
and U44690 (N_44690,N_37856,N_35936);
nand U44691 (N_44691,N_37709,N_39777);
nand U44692 (N_44692,N_37079,N_38600);
xor U44693 (N_44693,N_37811,N_39562);
xor U44694 (N_44694,N_36644,N_36489);
xnor U44695 (N_44695,N_39605,N_38167);
nor U44696 (N_44696,N_35945,N_39206);
xor U44697 (N_44697,N_35555,N_35681);
xnor U44698 (N_44698,N_37077,N_36825);
or U44699 (N_44699,N_37375,N_38074);
nand U44700 (N_44700,N_38768,N_35116);
and U44701 (N_44701,N_37954,N_35559);
xor U44702 (N_44702,N_38070,N_39293);
nand U44703 (N_44703,N_36855,N_35532);
xor U44704 (N_44704,N_38133,N_35046);
or U44705 (N_44705,N_36553,N_38135);
or U44706 (N_44706,N_36222,N_36745);
and U44707 (N_44707,N_39017,N_38195);
and U44708 (N_44708,N_38508,N_38119);
nor U44709 (N_44709,N_39147,N_38900);
xnor U44710 (N_44710,N_36184,N_39105);
nor U44711 (N_44711,N_38954,N_37930);
nor U44712 (N_44712,N_37253,N_38663);
xor U44713 (N_44713,N_39261,N_35467);
or U44714 (N_44714,N_38797,N_37521);
nand U44715 (N_44715,N_38017,N_38994);
or U44716 (N_44716,N_36245,N_36487);
or U44717 (N_44717,N_39469,N_36594);
nand U44718 (N_44718,N_37252,N_39713);
nand U44719 (N_44719,N_38194,N_36549);
nand U44720 (N_44720,N_36835,N_37858);
nand U44721 (N_44721,N_36206,N_39869);
nand U44722 (N_44722,N_38449,N_38587);
or U44723 (N_44723,N_35913,N_39683);
nand U44724 (N_44724,N_39383,N_38033);
nand U44725 (N_44725,N_35937,N_36975);
xnor U44726 (N_44726,N_35991,N_35455);
and U44727 (N_44727,N_36366,N_36375);
nand U44728 (N_44728,N_35455,N_38313);
and U44729 (N_44729,N_35729,N_35968);
nand U44730 (N_44730,N_39948,N_35128);
or U44731 (N_44731,N_36010,N_35910);
nor U44732 (N_44732,N_36406,N_36788);
and U44733 (N_44733,N_37966,N_37104);
or U44734 (N_44734,N_36540,N_39480);
xnor U44735 (N_44735,N_35270,N_37972);
nor U44736 (N_44736,N_35939,N_38077);
nand U44737 (N_44737,N_35496,N_38975);
nor U44738 (N_44738,N_37715,N_37138);
and U44739 (N_44739,N_36378,N_37735);
xor U44740 (N_44740,N_38269,N_37750);
or U44741 (N_44741,N_39143,N_36276);
nand U44742 (N_44742,N_37285,N_39990);
and U44743 (N_44743,N_39145,N_38106);
nand U44744 (N_44744,N_35893,N_35078);
nor U44745 (N_44745,N_36921,N_36085);
and U44746 (N_44746,N_39234,N_39081);
and U44747 (N_44747,N_35361,N_35601);
or U44748 (N_44748,N_38303,N_39346);
nor U44749 (N_44749,N_36758,N_39302);
and U44750 (N_44750,N_36641,N_38806);
nand U44751 (N_44751,N_36704,N_37318);
xnor U44752 (N_44752,N_38813,N_38520);
nand U44753 (N_44753,N_39330,N_37837);
nand U44754 (N_44754,N_38579,N_37718);
nand U44755 (N_44755,N_39708,N_35626);
xor U44756 (N_44756,N_37387,N_37186);
xor U44757 (N_44757,N_39518,N_36131);
and U44758 (N_44758,N_39863,N_37878);
nor U44759 (N_44759,N_36153,N_37058);
nor U44760 (N_44760,N_39985,N_35798);
xnor U44761 (N_44761,N_35415,N_35305);
nand U44762 (N_44762,N_36218,N_35135);
nor U44763 (N_44763,N_36127,N_37683);
or U44764 (N_44764,N_37944,N_35094);
and U44765 (N_44765,N_35683,N_39647);
nor U44766 (N_44766,N_35283,N_37973);
nor U44767 (N_44767,N_36859,N_36457);
nand U44768 (N_44768,N_37610,N_37821);
xor U44769 (N_44769,N_39899,N_38032);
and U44770 (N_44770,N_36496,N_35685);
nor U44771 (N_44771,N_36761,N_36819);
nor U44772 (N_44772,N_38291,N_37355);
and U44773 (N_44773,N_36103,N_35579);
nor U44774 (N_44774,N_38977,N_36310);
or U44775 (N_44775,N_38697,N_37652);
nor U44776 (N_44776,N_36206,N_37657);
or U44777 (N_44777,N_36636,N_36691);
or U44778 (N_44778,N_37685,N_35268);
or U44779 (N_44779,N_35461,N_39206);
or U44780 (N_44780,N_35449,N_37400);
or U44781 (N_44781,N_37836,N_37247);
or U44782 (N_44782,N_39760,N_37471);
and U44783 (N_44783,N_37910,N_38096);
nor U44784 (N_44784,N_39154,N_35216);
xor U44785 (N_44785,N_35397,N_36685);
or U44786 (N_44786,N_39788,N_35197);
xor U44787 (N_44787,N_36319,N_35405);
xnor U44788 (N_44788,N_35707,N_39941);
xor U44789 (N_44789,N_35924,N_37329);
and U44790 (N_44790,N_36492,N_36094);
nand U44791 (N_44791,N_39987,N_38039);
nor U44792 (N_44792,N_38494,N_35632);
xor U44793 (N_44793,N_39156,N_39330);
and U44794 (N_44794,N_39351,N_37555);
and U44795 (N_44795,N_35157,N_35029);
or U44796 (N_44796,N_36848,N_38249);
and U44797 (N_44797,N_35069,N_38644);
xnor U44798 (N_44798,N_38536,N_37083);
xnor U44799 (N_44799,N_38969,N_35404);
nand U44800 (N_44800,N_37813,N_36249);
or U44801 (N_44801,N_37930,N_39640);
nand U44802 (N_44802,N_37476,N_39589);
xnor U44803 (N_44803,N_38376,N_39865);
nand U44804 (N_44804,N_35115,N_38220);
xnor U44805 (N_44805,N_38226,N_39164);
and U44806 (N_44806,N_39740,N_37041);
or U44807 (N_44807,N_35662,N_36107);
or U44808 (N_44808,N_39577,N_36699);
xnor U44809 (N_44809,N_36951,N_39660);
and U44810 (N_44810,N_36763,N_39162);
xor U44811 (N_44811,N_38266,N_39273);
nor U44812 (N_44812,N_39306,N_38582);
xor U44813 (N_44813,N_36862,N_37793);
xnor U44814 (N_44814,N_36470,N_35309);
xor U44815 (N_44815,N_37497,N_39525);
and U44816 (N_44816,N_38440,N_38401);
and U44817 (N_44817,N_36847,N_38959);
nand U44818 (N_44818,N_36058,N_38006);
xor U44819 (N_44819,N_38137,N_35936);
nand U44820 (N_44820,N_37848,N_35805);
nand U44821 (N_44821,N_37543,N_36750);
or U44822 (N_44822,N_35137,N_36094);
nor U44823 (N_44823,N_36522,N_36684);
nand U44824 (N_44824,N_36755,N_39351);
nand U44825 (N_44825,N_35102,N_36926);
or U44826 (N_44826,N_37516,N_39850);
nor U44827 (N_44827,N_38418,N_38210);
and U44828 (N_44828,N_36314,N_37622);
nor U44829 (N_44829,N_38414,N_36858);
nand U44830 (N_44830,N_38572,N_35442);
nand U44831 (N_44831,N_37410,N_37577);
nor U44832 (N_44832,N_35281,N_39303);
and U44833 (N_44833,N_38531,N_38566);
or U44834 (N_44834,N_36060,N_35830);
or U44835 (N_44835,N_36424,N_39254);
nor U44836 (N_44836,N_35206,N_37373);
and U44837 (N_44837,N_35216,N_35291);
nand U44838 (N_44838,N_37315,N_38066);
xnor U44839 (N_44839,N_35551,N_39535);
nor U44840 (N_44840,N_37587,N_38248);
xnor U44841 (N_44841,N_35209,N_35825);
nand U44842 (N_44842,N_39269,N_38354);
xor U44843 (N_44843,N_38509,N_36309);
and U44844 (N_44844,N_38883,N_35313);
xnor U44845 (N_44845,N_36071,N_37806);
nor U44846 (N_44846,N_37118,N_38089);
xnor U44847 (N_44847,N_38405,N_35446);
and U44848 (N_44848,N_35738,N_37397);
or U44849 (N_44849,N_36283,N_38707);
nor U44850 (N_44850,N_37297,N_39892);
nor U44851 (N_44851,N_38754,N_37037);
or U44852 (N_44852,N_39513,N_37188);
nor U44853 (N_44853,N_39721,N_38420);
xor U44854 (N_44854,N_38276,N_35249);
nand U44855 (N_44855,N_38787,N_38662);
xor U44856 (N_44856,N_37929,N_38997);
nand U44857 (N_44857,N_39302,N_36511);
and U44858 (N_44858,N_38468,N_37682);
and U44859 (N_44859,N_35633,N_35444);
nand U44860 (N_44860,N_35083,N_36780);
nor U44861 (N_44861,N_39046,N_36880);
nand U44862 (N_44862,N_36017,N_36397);
and U44863 (N_44863,N_38519,N_38614);
nor U44864 (N_44864,N_38656,N_38125);
or U44865 (N_44865,N_39612,N_36501);
nand U44866 (N_44866,N_35318,N_39246);
nor U44867 (N_44867,N_36581,N_36317);
xnor U44868 (N_44868,N_39412,N_39097);
xor U44869 (N_44869,N_38182,N_37206);
or U44870 (N_44870,N_39758,N_37887);
nor U44871 (N_44871,N_37545,N_35147);
nor U44872 (N_44872,N_35041,N_37386);
nor U44873 (N_44873,N_35811,N_38725);
and U44874 (N_44874,N_35531,N_37206);
nor U44875 (N_44875,N_39053,N_35147);
xor U44876 (N_44876,N_35931,N_37455);
and U44877 (N_44877,N_36980,N_35207);
nor U44878 (N_44878,N_37163,N_36294);
nor U44879 (N_44879,N_37240,N_35355);
and U44880 (N_44880,N_38361,N_38479);
xnor U44881 (N_44881,N_37992,N_39185);
xor U44882 (N_44882,N_39293,N_37953);
and U44883 (N_44883,N_35206,N_39378);
and U44884 (N_44884,N_39072,N_37869);
or U44885 (N_44885,N_36260,N_37340);
xnor U44886 (N_44886,N_38996,N_35963);
xnor U44887 (N_44887,N_36214,N_39135);
and U44888 (N_44888,N_35852,N_36958);
nor U44889 (N_44889,N_37446,N_35031);
or U44890 (N_44890,N_35758,N_35288);
xor U44891 (N_44891,N_36957,N_36203);
and U44892 (N_44892,N_39236,N_38872);
and U44893 (N_44893,N_36971,N_39358);
nor U44894 (N_44894,N_35751,N_35237);
nand U44895 (N_44895,N_38005,N_35151);
or U44896 (N_44896,N_36795,N_38525);
xor U44897 (N_44897,N_39911,N_35355);
or U44898 (N_44898,N_36793,N_39411);
nor U44899 (N_44899,N_39770,N_38872);
or U44900 (N_44900,N_39826,N_36962);
or U44901 (N_44901,N_38293,N_36037);
and U44902 (N_44902,N_36166,N_37070);
xor U44903 (N_44903,N_39751,N_35436);
nor U44904 (N_44904,N_39008,N_37783);
nand U44905 (N_44905,N_38417,N_38680);
and U44906 (N_44906,N_38059,N_36666);
xnor U44907 (N_44907,N_38270,N_38072);
xnor U44908 (N_44908,N_37233,N_36758);
nor U44909 (N_44909,N_36543,N_35754);
xor U44910 (N_44910,N_37696,N_38113);
and U44911 (N_44911,N_36360,N_38818);
nor U44912 (N_44912,N_38656,N_36235);
and U44913 (N_44913,N_39834,N_39631);
nand U44914 (N_44914,N_38234,N_38601);
and U44915 (N_44915,N_39449,N_36243);
nor U44916 (N_44916,N_37454,N_38668);
or U44917 (N_44917,N_36328,N_38529);
xnor U44918 (N_44918,N_36990,N_36746);
xnor U44919 (N_44919,N_35595,N_39236);
nand U44920 (N_44920,N_39643,N_35838);
nor U44921 (N_44921,N_36105,N_39257);
and U44922 (N_44922,N_36572,N_35570);
and U44923 (N_44923,N_39832,N_38854);
nand U44924 (N_44924,N_35517,N_38840);
nand U44925 (N_44925,N_39809,N_38168);
and U44926 (N_44926,N_38572,N_36520);
xnor U44927 (N_44927,N_38746,N_38194);
nor U44928 (N_44928,N_37679,N_37038);
and U44929 (N_44929,N_39062,N_39772);
xor U44930 (N_44930,N_37190,N_36458);
or U44931 (N_44931,N_36275,N_36377);
and U44932 (N_44932,N_39322,N_39683);
nand U44933 (N_44933,N_39065,N_36672);
xor U44934 (N_44934,N_39357,N_39925);
and U44935 (N_44935,N_37507,N_35360);
and U44936 (N_44936,N_37334,N_36753);
and U44937 (N_44937,N_38847,N_38304);
nand U44938 (N_44938,N_37698,N_35092);
nand U44939 (N_44939,N_35703,N_38437);
nand U44940 (N_44940,N_35462,N_35218);
nand U44941 (N_44941,N_38645,N_39992);
xor U44942 (N_44942,N_36141,N_35529);
or U44943 (N_44943,N_39455,N_36465);
nor U44944 (N_44944,N_35706,N_35662);
xnor U44945 (N_44945,N_39390,N_38825);
nor U44946 (N_44946,N_36373,N_39969);
nand U44947 (N_44947,N_39344,N_35313);
nor U44948 (N_44948,N_38791,N_35841);
nor U44949 (N_44949,N_35402,N_38549);
nand U44950 (N_44950,N_38249,N_39226);
or U44951 (N_44951,N_39672,N_35726);
and U44952 (N_44952,N_36253,N_35650);
nor U44953 (N_44953,N_36844,N_37185);
and U44954 (N_44954,N_38425,N_36909);
or U44955 (N_44955,N_38437,N_36162);
nand U44956 (N_44956,N_35519,N_37899);
or U44957 (N_44957,N_38145,N_39087);
nand U44958 (N_44958,N_38804,N_35095);
and U44959 (N_44959,N_38858,N_39922);
nand U44960 (N_44960,N_36612,N_39534);
and U44961 (N_44961,N_35664,N_36563);
or U44962 (N_44962,N_37777,N_38436);
and U44963 (N_44963,N_39547,N_39459);
nor U44964 (N_44964,N_38082,N_39003);
and U44965 (N_44965,N_35060,N_38154);
nand U44966 (N_44966,N_35649,N_36790);
nor U44967 (N_44967,N_39715,N_38965);
xor U44968 (N_44968,N_36881,N_36748);
xnor U44969 (N_44969,N_37138,N_36319);
xnor U44970 (N_44970,N_37234,N_36912);
nor U44971 (N_44971,N_35128,N_39226);
nor U44972 (N_44972,N_35797,N_38155);
nor U44973 (N_44973,N_35936,N_35461);
nand U44974 (N_44974,N_38670,N_37608);
nand U44975 (N_44975,N_35891,N_35081);
xnor U44976 (N_44976,N_39018,N_37475);
xor U44977 (N_44977,N_39737,N_37124);
nand U44978 (N_44978,N_37161,N_35162);
or U44979 (N_44979,N_36827,N_39730);
or U44980 (N_44980,N_35050,N_39814);
or U44981 (N_44981,N_39970,N_38359);
nand U44982 (N_44982,N_39907,N_39345);
nor U44983 (N_44983,N_36228,N_38144);
nand U44984 (N_44984,N_39146,N_38553);
nor U44985 (N_44985,N_37842,N_39727);
nand U44986 (N_44986,N_35284,N_37550);
and U44987 (N_44987,N_39910,N_39255);
or U44988 (N_44988,N_39703,N_39241);
nor U44989 (N_44989,N_38881,N_36839);
nor U44990 (N_44990,N_37650,N_36905);
nor U44991 (N_44991,N_38505,N_39593);
nor U44992 (N_44992,N_36685,N_37055);
xor U44993 (N_44993,N_37589,N_35419);
and U44994 (N_44994,N_38921,N_39547);
nand U44995 (N_44995,N_39653,N_39502);
nand U44996 (N_44996,N_38125,N_38885);
xor U44997 (N_44997,N_39730,N_38942);
or U44998 (N_44998,N_35219,N_35921);
nand U44999 (N_44999,N_39830,N_37887);
nand U45000 (N_45000,N_44284,N_44186);
nor U45001 (N_45001,N_41514,N_41957);
nor U45002 (N_45002,N_43431,N_44541);
and U45003 (N_45003,N_44322,N_42845);
or U45004 (N_45004,N_44778,N_41008);
nand U45005 (N_45005,N_44825,N_40659);
and U45006 (N_45006,N_43894,N_43146);
xor U45007 (N_45007,N_44496,N_42492);
or U45008 (N_45008,N_42884,N_42383);
nand U45009 (N_45009,N_40050,N_44391);
xor U45010 (N_45010,N_42323,N_43628);
xnor U45011 (N_45011,N_40208,N_43184);
nor U45012 (N_45012,N_41811,N_42665);
or U45013 (N_45013,N_43683,N_40997);
xnor U45014 (N_45014,N_41027,N_41639);
and U45015 (N_45015,N_42469,N_40733);
or U45016 (N_45016,N_42747,N_41462);
and U45017 (N_45017,N_41756,N_43285);
and U45018 (N_45018,N_42745,N_42029);
xnor U45019 (N_45019,N_43964,N_42703);
nor U45020 (N_45020,N_44439,N_42381);
and U45021 (N_45021,N_43823,N_40273);
and U45022 (N_45022,N_43825,N_42082);
or U45023 (N_45023,N_40213,N_42881);
xnor U45024 (N_45024,N_40024,N_42503);
or U45025 (N_45025,N_42481,N_41839);
or U45026 (N_45026,N_43452,N_41308);
and U45027 (N_45027,N_41647,N_40500);
nor U45028 (N_45028,N_42688,N_40847);
nor U45029 (N_45029,N_42890,N_43904);
and U45030 (N_45030,N_44207,N_42791);
and U45031 (N_45031,N_42192,N_42651);
and U45032 (N_45032,N_43138,N_44008);
xnor U45033 (N_45033,N_43317,N_41411);
nor U45034 (N_45034,N_44631,N_40547);
nor U45035 (N_45035,N_42604,N_41294);
xor U45036 (N_45036,N_43723,N_41498);
and U45037 (N_45037,N_42416,N_43831);
and U45038 (N_45038,N_40751,N_43172);
nor U45039 (N_45039,N_43185,N_44427);
xnor U45040 (N_45040,N_42773,N_41237);
and U45041 (N_45041,N_42310,N_44504);
or U45042 (N_45042,N_43795,N_43237);
and U45043 (N_45043,N_42853,N_43523);
nor U45044 (N_45044,N_40275,N_42558);
nand U45045 (N_45045,N_43705,N_43821);
nand U45046 (N_45046,N_44055,N_41450);
nand U45047 (N_45047,N_40940,N_40076);
or U45048 (N_45048,N_42030,N_43142);
nand U45049 (N_45049,N_41365,N_44232);
or U45050 (N_45050,N_43501,N_42893);
or U45051 (N_45051,N_40781,N_41396);
nand U45052 (N_45052,N_44144,N_41831);
or U45053 (N_45053,N_40414,N_40945);
nor U45054 (N_45054,N_40061,N_41429);
and U45055 (N_45055,N_43113,N_44355);
nand U45056 (N_45056,N_42339,N_42186);
and U45057 (N_45057,N_43847,N_40017);
nor U45058 (N_45058,N_43630,N_40140);
and U45059 (N_45059,N_40251,N_40191);
xnor U45060 (N_45060,N_44110,N_43245);
xnor U45061 (N_45061,N_41423,N_44585);
xnor U45062 (N_45062,N_42292,N_43033);
nor U45063 (N_45063,N_42107,N_41400);
nand U45064 (N_45064,N_42119,N_44195);
nor U45065 (N_45065,N_43416,N_40784);
nand U45066 (N_45066,N_40141,N_43855);
xor U45067 (N_45067,N_40156,N_41962);
or U45068 (N_45068,N_41246,N_40403);
xnor U45069 (N_45069,N_43277,N_42515);
xnor U45070 (N_45070,N_43366,N_41381);
nand U45071 (N_45071,N_40212,N_42054);
nor U45072 (N_45072,N_40676,N_40885);
or U45073 (N_45073,N_41527,N_41555);
or U45074 (N_45074,N_40052,N_43955);
or U45075 (N_45075,N_43058,N_40005);
or U45076 (N_45076,N_42157,N_43588);
xnor U45077 (N_45077,N_43256,N_43393);
xor U45078 (N_45078,N_44663,N_42818);
nor U45079 (N_45079,N_42647,N_44592);
or U45080 (N_45080,N_40016,N_41779);
or U45081 (N_45081,N_42353,N_41581);
nor U45082 (N_45082,N_42460,N_42790);
and U45083 (N_45083,N_42785,N_42440);
xor U45084 (N_45084,N_40905,N_40708);
nor U45085 (N_45085,N_42173,N_40485);
or U45086 (N_45086,N_40675,N_40133);
nor U45087 (N_45087,N_42780,N_41676);
xnor U45088 (N_45088,N_41889,N_40787);
nor U45089 (N_45089,N_40450,N_40132);
and U45090 (N_45090,N_44237,N_42073);
or U45091 (N_45091,N_43536,N_44224);
or U45092 (N_45092,N_44738,N_43260);
nand U45093 (N_45093,N_44529,N_41179);
nand U45094 (N_45094,N_44680,N_44539);
and U45095 (N_45095,N_42034,N_40755);
xor U45096 (N_45096,N_40672,N_41241);
xor U45097 (N_45097,N_44382,N_41263);
xor U45098 (N_45098,N_42587,N_44637);
xnor U45099 (N_45099,N_41573,N_42961);
and U45100 (N_45100,N_44040,N_41163);
or U45101 (N_45101,N_41594,N_41947);
or U45102 (N_45102,N_41229,N_40419);
nor U45103 (N_45103,N_42386,N_40601);
or U45104 (N_45104,N_44313,N_40070);
and U45105 (N_45105,N_41216,N_41976);
and U45106 (N_45106,N_44405,N_43215);
or U45107 (N_45107,N_40244,N_40286);
nand U45108 (N_45108,N_42354,N_43912);
xnor U45109 (N_45109,N_41517,N_43797);
or U45110 (N_45110,N_42530,N_40261);
nand U45111 (N_45111,N_43947,N_41002);
nor U45112 (N_45112,N_42538,N_43733);
and U45113 (N_45113,N_41844,N_42692);
and U45114 (N_45114,N_41678,N_40874);
or U45115 (N_45115,N_42768,N_42204);
and U45116 (N_45116,N_42283,N_44134);
nand U45117 (N_45117,N_40652,N_40510);
nor U45118 (N_45118,N_44448,N_44170);
and U45119 (N_45119,N_41507,N_42936);
xor U45120 (N_45120,N_41283,N_41218);
nand U45121 (N_45121,N_44797,N_41091);
nand U45122 (N_45122,N_42614,N_40346);
nor U45123 (N_45123,N_43875,N_42450);
nand U45124 (N_45124,N_40287,N_41410);
or U45125 (N_45125,N_44665,N_42738);
nor U45126 (N_45126,N_43364,N_43568);
nor U45127 (N_45127,N_41311,N_44905);
and U45128 (N_45128,N_41474,N_43540);
nor U45129 (N_45129,N_43150,N_43573);
nor U45130 (N_45130,N_41605,N_42001);
nand U45131 (N_45131,N_44594,N_41826);
or U45132 (N_45132,N_43608,N_42970);
and U45133 (N_45133,N_41539,N_41031);
xnor U45134 (N_45134,N_40706,N_43326);
nand U45135 (N_45135,N_44203,N_41035);
nand U45136 (N_45136,N_43755,N_44239);
nor U45137 (N_45137,N_44161,N_43669);
nor U45138 (N_45138,N_43133,N_42271);
xnor U45139 (N_45139,N_41136,N_42009);
or U45140 (N_45140,N_41439,N_42588);
nand U45141 (N_45141,N_41733,N_40267);
xor U45142 (N_45142,N_41285,N_41104);
nand U45143 (N_45143,N_41706,N_42687);
nor U45144 (N_45144,N_41821,N_42153);
xor U45145 (N_45145,N_41759,N_44095);
and U45146 (N_45146,N_43688,N_42570);
nor U45147 (N_45147,N_40084,N_40685);
nand U45148 (N_45148,N_44273,N_41387);
or U45149 (N_45149,N_44075,N_41330);
and U45150 (N_45150,N_44786,N_41312);
and U45151 (N_45151,N_43175,N_42227);
nor U45152 (N_45152,N_44987,N_44071);
or U45153 (N_45153,N_42096,N_43589);
and U45154 (N_45154,N_40085,N_40777);
nor U45155 (N_45155,N_44373,N_44544);
nand U45156 (N_45156,N_44029,N_41030);
nor U45157 (N_45157,N_42183,N_40556);
nand U45158 (N_45158,N_40219,N_41476);
or U45159 (N_45159,N_40724,N_40066);
or U45160 (N_45160,N_44137,N_44542);
nor U45161 (N_45161,N_43899,N_42546);
nor U45162 (N_45162,N_42049,N_41010);
nand U45163 (N_45163,N_41998,N_41258);
xor U45164 (N_45164,N_43808,N_42443);
nand U45165 (N_45165,N_44844,N_41481);
nor U45166 (N_45166,N_44012,N_44490);
and U45167 (N_45167,N_40987,N_43454);
and U45168 (N_45168,N_44475,N_44904);
xnor U45169 (N_45169,N_43958,N_44979);
and U45170 (N_45170,N_42796,N_43999);
nand U45171 (N_45171,N_41667,N_43293);
nor U45172 (N_45172,N_40971,N_42319);
or U45173 (N_45173,N_43753,N_42465);
xor U45174 (N_45174,N_43807,N_40009);
nor U45175 (N_45175,N_44160,N_42159);
and U45176 (N_45176,N_44622,N_40850);
nor U45177 (N_45177,N_40578,N_41337);
and U45178 (N_45178,N_43410,N_42721);
or U45179 (N_45179,N_41233,N_41026);
nor U45180 (N_45180,N_42100,N_44573);
and U45181 (N_45181,N_42594,N_42878);
nand U45182 (N_45182,N_42824,N_43168);
and U45183 (N_45183,N_41970,N_43141);
xnor U45184 (N_45184,N_40859,N_44822);
or U45185 (N_45185,N_43219,N_40211);
xor U45186 (N_45186,N_42591,N_40655);
and U45187 (N_45187,N_40505,N_40234);
nand U45188 (N_45188,N_44532,N_40362);
or U45189 (N_45189,N_40795,N_40875);
nand U45190 (N_45190,N_40923,N_41509);
nor U45191 (N_45191,N_42631,N_44106);
xnor U45192 (N_45192,N_42982,N_43974);
or U45193 (N_45193,N_44017,N_42912);
xnor U45194 (N_45194,N_42285,N_40598);
nand U45195 (N_45195,N_43457,N_41975);
xor U45196 (N_45196,N_41862,N_40792);
nor U45197 (N_45197,N_43673,N_41700);
nor U45198 (N_45198,N_40101,N_43076);
and U45199 (N_45199,N_41972,N_40677);
nor U45200 (N_45200,N_41428,N_44520);
or U45201 (N_45201,N_40355,N_44766);
xor U45202 (N_45202,N_43583,N_41252);
and U45203 (N_45203,N_41152,N_43828);
or U45204 (N_45204,N_43089,N_42811);
or U45205 (N_45205,N_43319,N_44768);
nand U45206 (N_45206,N_43681,N_40840);
nor U45207 (N_45207,N_44880,N_44846);
and U45208 (N_45208,N_40773,N_44831);
or U45209 (N_45209,N_44067,N_41460);
and U45210 (N_45210,N_43191,N_42307);
and U45211 (N_45211,N_40749,N_42777);
xor U45212 (N_45212,N_44376,N_40621);
xnor U45213 (N_45213,N_40680,N_43786);
nor U45214 (N_45214,N_42236,N_42012);
and U45215 (N_45215,N_43852,N_42041);
xnor U45216 (N_45216,N_40006,N_44903);
nor U45217 (N_45217,N_40092,N_40550);
or U45218 (N_45218,N_43982,N_40284);
and U45219 (N_45219,N_41720,N_43164);
xor U45220 (N_45220,N_41427,N_41684);
or U45221 (N_45221,N_44695,N_44320);
xnor U45222 (N_45222,N_41042,N_43477);
xnor U45223 (N_45223,N_41340,N_40469);
or U45224 (N_45224,N_40925,N_43476);
xnor U45225 (N_45225,N_40168,N_40742);
nor U45226 (N_45226,N_43144,N_44523);
nand U45227 (N_45227,N_42017,N_44257);
nand U45228 (N_45228,N_43617,N_43502);
or U45229 (N_45229,N_43928,N_40282);
or U45230 (N_45230,N_40171,N_40065);
or U45231 (N_45231,N_42543,N_44407);
and U45232 (N_45232,N_42166,N_40048);
nor U45233 (N_45233,N_43061,N_43937);
nand U45234 (N_45234,N_42962,N_43742);
nand U45235 (N_45235,N_43846,N_41589);
xnor U45236 (N_45236,N_43992,N_40838);
or U45237 (N_45237,N_42161,N_43814);
or U45238 (N_45238,N_42918,N_44128);
or U45239 (N_45239,N_43938,N_42331);
or U45240 (N_45240,N_41397,N_43396);
or U45241 (N_45241,N_41028,N_42060);
nor U45242 (N_45242,N_40280,N_40456);
nand U45243 (N_45243,N_42038,N_44025);
nor U45244 (N_45244,N_42028,N_40319);
nand U45245 (N_45245,N_44612,N_44117);
nor U45246 (N_45246,N_41897,N_42395);
nand U45247 (N_45247,N_41820,N_40074);
and U45248 (N_45248,N_41382,N_42684);
nand U45249 (N_45249,N_40643,N_43620);
nor U45250 (N_45250,N_40077,N_41398);
nor U45251 (N_45251,N_43322,N_43612);
nand U45252 (N_45252,N_40245,N_40563);
and U45253 (N_45253,N_44586,N_43386);
or U45254 (N_45254,N_43811,N_41632);
xor U45255 (N_45255,N_44083,N_41544);
and U45256 (N_45256,N_42170,N_43897);
and U45257 (N_45257,N_40153,N_41162);
xnor U45258 (N_45258,N_41658,N_41804);
nand U45259 (N_45259,N_41234,N_40623);
xor U45260 (N_45260,N_42830,N_42135);
nor U45261 (N_45261,N_40125,N_42812);
xor U45262 (N_45262,N_44020,N_40719);
nor U45263 (N_45263,N_44717,N_44621);
nand U45264 (N_45264,N_41540,N_44700);
and U45265 (N_45265,N_42939,N_43145);
or U45266 (N_45266,N_42122,N_42995);
xor U45267 (N_45267,N_44625,N_41682);
xnor U45268 (N_45268,N_44640,N_44891);
or U45269 (N_45269,N_41687,N_43662);
and U45270 (N_45270,N_42399,N_40809);
nor U45271 (N_45271,N_44261,N_41089);
and U45272 (N_45272,N_40767,N_42290);
or U45273 (N_45273,N_41023,N_40744);
or U45274 (N_45274,N_41139,N_43743);
or U45275 (N_45275,N_43445,N_44103);
nand U45276 (N_45276,N_41845,N_43806);
xor U45277 (N_45277,N_44009,N_43280);
and U45278 (N_45278,N_41742,N_40854);
or U45279 (N_45279,N_40455,N_44143);
xor U45280 (N_45280,N_40970,N_44919);
or U45281 (N_45281,N_41566,N_42441);
nor U45282 (N_45282,N_44792,N_44870);
xnor U45283 (N_45283,N_40797,N_42784);
or U45284 (N_45284,N_43702,N_41364);
and U45285 (N_45285,N_40917,N_40931);
nor U45286 (N_45286,N_41471,N_41932);
nor U45287 (N_45287,N_40754,N_44502);
nor U45288 (N_45288,N_40095,N_43016);
xnor U45289 (N_45289,N_43602,N_40493);
or U45290 (N_45290,N_44780,N_44352);
and U45291 (N_45291,N_43264,N_41933);
and U45292 (N_45292,N_41668,N_44740);
xor U45293 (N_45293,N_41121,N_41006);
nand U45294 (N_45294,N_43011,N_42882);
nor U45295 (N_45295,N_40040,N_44135);
and U45296 (N_45296,N_41444,N_42691);
nand U45297 (N_45297,N_40723,N_40207);
or U45298 (N_45298,N_40844,N_44166);
nor U45299 (N_45299,N_41865,N_41230);
and U45300 (N_45300,N_43923,N_40972);
nor U45301 (N_45301,N_40994,N_44847);
xnor U45302 (N_45302,N_43554,N_43817);
xor U45303 (N_45303,N_40349,N_44521);
and U45304 (N_45304,N_41570,N_40597);
nor U45305 (N_45305,N_42453,N_42915);
nor U45306 (N_45306,N_42193,N_43495);
nor U45307 (N_45307,N_40188,N_42902);
and U45308 (N_45308,N_40779,N_41590);
nor U45309 (N_45309,N_40879,N_41112);
nor U45310 (N_45310,N_44922,N_43105);
nand U45311 (N_45311,N_44397,N_41693);
and U45312 (N_45312,N_42904,N_44684);
nand U45313 (N_45313,N_43283,N_43380);
nand U45314 (N_45314,N_41871,N_42209);
nor U45315 (N_45315,N_44611,N_41881);
nand U45316 (N_45316,N_41604,N_41314);
and U45317 (N_45317,N_42827,N_41380);
nand U45318 (N_45318,N_44064,N_43359);
or U45319 (N_45319,N_43533,N_41105);
xor U45320 (N_45320,N_42212,N_41361);
xor U45321 (N_45321,N_40043,N_44887);
nor U45322 (N_45322,N_43367,N_43041);
and U45323 (N_45323,N_43547,N_41917);
and U45324 (N_45324,N_40574,N_44812);
or U45325 (N_45325,N_42118,N_42302);
xor U45326 (N_45326,N_42101,N_43179);
or U45327 (N_45327,N_42497,N_42771);
nand U45328 (N_45328,N_41817,N_42014);
nor U45329 (N_45329,N_43463,N_41090);
nand U45330 (N_45330,N_42948,N_40726);
and U45331 (N_45331,N_41313,N_44901);
nand U45332 (N_45332,N_43096,N_40262);
xor U45333 (N_45333,N_44330,N_41609);
and U45334 (N_45334,N_40696,N_44892);
nor U45335 (N_45335,N_41847,N_42396);
xor U45336 (N_45336,N_40806,N_41614);
xnor U45337 (N_45337,N_43009,N_44519);
or U45338 (N_45338,N_41188,N_44381);
xor U45339 (N_45339,N_40393,N_40487);
nor U45340 (N_45340,N_44824,N_44858);
or U45341 (N_45341,N_43751,N_40012);
and U45342 (N_45342,N_44947,N_43752);
nor U45343 (N_45343,N_43188,N_41446);
nand U45344 (N_45344,N_42756,N_40474);
and U45345 (N_45345,N_43344,N_42875);
nor U45346 (N_45346,N_44560,N_42356);
nor U45347 (N_45347,N_41046,N_43639);
or U45348 (N_45348,N_41711,N_42221);
xnor U45349 (N_45349,N_42284,N_40035);
nor U45350 (N_45350,N_41531,N_43767);
or U45351 (N_45351,N_43914,N_43353);
xor U45352 (N_45352,N_42211,N_42788);
nand U45353 (N_45353,N_41982,N_44327);
xor U45354 (N_45354,N_40134,N_40364);
and U45355 (N_45355,N_42770,N_40502);
xor U45356 (N_45356,N_43126,N_40446);
or U45357 (N_45357,N_40105,N_42522);
nand U45358 (N_45358,N_41209,N_41571);
nor U45359 (N_45359,N_41150,N_44527);
xnor U45360 (N_45360,N_40130,N_42261);
nand U45361 (N_45361,N_42398,N_44453);
xnor U45362 (N_45362,N_40409,N_40851);
xor U45363 (N_45363,N_43843,N_40072);
xnor U45364 (N_45364,N_43004,N_42114);
xnor U45365 (N_45365,N_41458,N_43400);
or U45366 (N_45366,N_40688,N_42218);
nor U45367 (N_45367,N_42749,N_41629);
nand U45368 (N_45368,N_42005,N_43235);
or U45369 (N_45369,N_44167,N_41920);
nor U45370 (N_45370,N_43804,N_43027);
or U45371 (N_45371,N_41611,N_43980);
and U45372 (N_45372,N_41015,N_44602);
or U45373 (N_45373,N_44256,N_44359);
and U45374 (N_45374,N_40051,N_41092);
or U45375 (N_45375,N_41926,N_43908);
or U45376 (N_45376,N_41558,N_40379);
and U45377 (N_45377,N_40570,N_44531);
or U45378 (N_45378,N_41383,N_43960);
or U45379 (N_45379,N_43844,N_44341);
xnor U45380 (N_45380,N_40762,N_42897);
and U45381 (N_45381,N_43835,N_41595);
xnor U45382 (N_45382,N_43613,N_40820);
xnor U45383 (N_45383,N_42722,N_44830);
or U45384 (N_45384,N_43882,N_40158);
and U45385 (N_45385,N_44654,N_41317);
or U45386 (N_45386,N_41094,N_40962);
nor U45387 (N_45387,N_43800,N_43167);
xnor U45388 (N_45388,N_43961,N_42701);
or U45389 (N_45389,N_43975,N_42240);
nand U45390 (N_45390,N_44368,N_44626);
or U45391 (N_45391,N_41224,N_44365);
nor U45392 (N_45392,N_44796,N_43092);
nand U45393 (N_45393,N_43887,N_44077);
or U45394 (N_45394,N_40067,N_42873);
and U45395 (N_45395,N_44535,N_42362);
or U45396 (N_45396,N_41637,N_41384);
nor U45397 (N_45397,N_42025,N_43050);
and U45398 (N_45398,N_41966,N_40712);
nor U45399 (N_45399,N_40057,N_40938);
or U45400 (N_45400,N_44482,N_41608);
and U45401 (N_45401,N_43713,N_43838);
or U45402 (N_45402,N_40124,N_40537);
xor U45403 (N_45403,N_44956,N_42855);
xnor U45404 (N_45404,N_41334,N_43719);
xor U45405 (N_45405,N_41022,N_42269);
or U45406 (N_45406,N_41786,N_41447);
nor U45407 (N_45407,N_40614,N_41520);
xor U45408 (N_45408,N_40624,N_42981);
and U45409 (N_45409,N_44484,N_42430);
or U45410 (N_45410,N_41085,N_44566);
nand U45411 (N_45411,N_41255,N_41004);
and U45412 (N_45412,N_44952,N_42489);
nor U45413 (N_45413,N_42867,N_40109);
xnor U45414 (N_45414,N_43068,N_40709);
and U45415 (N_45415,N_42693,N_44001);
xor U45416 (N_45416,N_40626,N_40571);
nor U45417 (N_45417,N_40169,N_40628);
and U45418 (N_45418,N_42582,N_41618);
and U45419 (N_45419,N_44210,N_41730);
nor U45420 (N_45420,N_40150,N_41561);
nor U45421 (N_45421,N_43212,N_43906);
and U45422 (N_45422,N_41991,N_42486);
nand U45423 (N_45423,N_43551,N_42808);
or U45424 (N_45424,N_44080,N_40663);
or U45425 (N_45425,N_41291,N_44028);
xor U45426 (N_45426,N_44929,N_40123);
nor U45427 (N_45427,N_44066,N_40195);
nor U45428 (N_45428,N_44877,N_41469);
or U45429 (N_45429,N_42454,N_44292);
or U45430 (N_45430,N_44297,N_44153);
or U45431 (N_45431,N_44006,N_43182);
nand U45432 (N_45432,N_41869,N_43842);
and U45433 (N_45433,N_41078,N_41784);
or U45434 (N_45434,N_42532,N_43075);
or U45435 (N_45435,N_41191,N_43840);
and U45436 (N_45436,N_42925,N_40525);
xnor U45437 (N_45437,N_40309,N_43097);
nor U45438 (N_45438,N_41117,N_43526);
nor U45439 (N_45439,N_40573,N_43066);
or U45440 (N_45440,N_43349,N_44866);
and U45441 (N_45441,N_41265,N_42868);
or U45442 (N_45442,N_41556,N_43519);
and U45443 (N_45443,N_41415,N_44146);
xnor U45444 (N_45444,N_41393,N_43429);
nor U45445 (N_45445,N_42955,N_43645);
nand U45446 (N_45446,N_43171,N_40428);
or U45447 (N_45447,N_44130,N_40426);
and U45448 (N_45448,N_43448,N_43790);
or U45449 (N_45449,N_44869,N_44282);
nor U45450 (N_45450,N_43864,N_42633);
nand U45451 (N_45451,N_43658,N_42407);
xnor U45452 (N_45452,N_41298,N_40293);
or U45453 (N_45453,N_41059,N_44666);
xnor U45454 (N_45454,N_40738,N_43606);
nand U45455 (N_45455,N_43370,N_43045);
xnor U45456 (N_45456,N_41955,N_40593);
xor U45457 (N_45457,N_40834,N_40839);
nor U45458 (N_45458,N_40461,N_43419);
nand U45459 (N_45459,N_42748,N_44940);
and U45460 (N_45460,N_42423,N_41177);
nand U45461 (N_45461,N_41119,N_40071);
or U45462 (N_45462,N_41009,N_43279);
xnor U45463 (N_45463,N_41494,N_40445);
nand U45464 (N_45464,N_42993,N_41882);
or U45465 (N_45465,N_44636,N_43181);
xor U45466 (N_45466,N_44641,N_41158);
nand U45467 (N_45467,N_42184,N_44015);
nor U45468 (N_45468,N_41038,N_42402);
nor U45469 (N_45469,N_43927,N_41407);
xnor U45470 (N_45470,N_41825,N_40265);
or U45471 (N_45471,N_43263,N_44081);
nand U45472 (N_45472,N_42552,N_40778);
xor U45473 (N_45473,N_43604,N_44315);
nand U45474 (N_45474,N_41208,N_42487);
nand U45475 (N_45475,N_40387,N_40898);
and U45476 (N_45476,N_41133,N_42632);
and U45477 (N_45477,N_42580,N_43365);
nor U45478 (N_45478,N_41727,N_44466);
nor U45479 (N_45479,N_42056,N_41025);
xor U45480 (N_45480,N_41783,N_44098);
nand U45481 (N_45481,N_41395,N_40538);
xor U45482 (N_45482,N_40668,N_42542);
xor U45483 (N_45483,N_42358,N_44305);
or U45484 (N_45484,N_43039,N_43701);
nand U45485 (N_45485,N_43581,N_41129);
and U45486 (N_45486,N_43640,N_41601);
or U45487 (N_45487,N_42348,N_40315);
or U45488 (N_45488,N_43692,N_42677);
xnor U45489 (N_45489,N_40681,N_41773);
nor U45490 (N_45490,N_44004,N_41401);
nand U45491 (N_45491,N_41369,N_44158);
nand U45492 (N_45492,N_44311,N_42368);
and U45493 (N_45493,N_42006,N_42710);
and U45494 (N_45494,N_44048,N_44245);
nand U45495 (N_45495,N_41463,N_43163);
nor U45496 (N_45496,N_40222,N_44708);
nand U45497 (N_45497,N_42507,N_42091);
and U45498 (N_45498,N_42513,N_42917);
nand U45499 (N_45499,N_44449,N_44115);
nand U45500 (N_45500,N_42380,N_43868);
and U45501 (N_45501,N_41378,N_40323);
or U45502 (N_45502,N_43836,N_42942);
and U45503 (N_45503,N_41748,N_41456);
and U45504 (N_45504,N_40477,N_40711);
and U45505 (N_45505,N_43030,N_44107);
and U45506 (N_45506,N_44968,N_42560);
nor U45507 (N_45507,N_44304,N_42820);
nor U45508 (N_45508,N_42197,N_42579);
nor U45509 (N_45509,N_43475,N_40475);
nand U45510 (N_45510,N_40555,N_41870);
and U45511 (N_45511,N_41522,N_41029);
and U45512 (N_45512,N_42104,N_41187);
xor U45513 (N_45513,N_41994,N_44455);
and U45514 (N_45514,N_41368,N_40317);
nand U45515 (N_45515,N_42244,N_41610);
nor U45516 (N_45516,N_44323,N_42879);
or U45517 (N_45517,N_44145,N_40625);
xor U45518 (N_45518,N_40482,N_40372);
nand U45519 (N_45519,N_44725,N_41050);
nor U45520 (N_45520,N_40196,N_42959);
nor U45521 (N_45521,N_41596,N_44745);
xnor U45522 (N_45522,N_44508,N_40772);
and U45523 (N_45523,N_42741,N_40263);
nand U45524 (N_45524,N_40545,N_44886);
xnor U45525 (N_45525,N_41436,N_42156);
nand U45526 (N_45526,N_44241,N_42922);
nor U45527 (N_45527,N_40551,N_44422);
and U45528 (N_45528,N_43447,N_44838);
nand U45529 (N_45529,N_42052,N_42121);
or U45530 (N_45530,N_42892,N_43470);
or U45531 (N_45531,N_43924,N_43538);
or U45532 (N_45532,N_41256,N_40025);
nor U45533 (N_45533,N_44412,N_41525);
nand U45534 (N_45534,N_43449,N_42535);
and U45535 (N_45535,N_41360,N_43085);
nor U45536 (N_45536,N_41355,N_40835);
and U45537 (N_45537,N_44347,N_42190);
and U45538 (N_45538,N_41140,N_43651);
and U45539 (N_45539,N_43761,N_41838);
nor U45540 (N_45540,N_40750,N_43521);
or U45541 (N_45541,N_41457,N_44335);
and U45542 (N_45542,N_41167,N_40370);
xor U45543 (N_45543,N_42128,N_44507);
or U45544 (N_45544,N_40277,N_43444);
and U45545 (N_45545,N_41816,N_44572);
and U45546 (N_45546,N_42679,N_40103);
nand U45547 (N_45547,N_42675,N_42180);
nor U45548 (N_45548,N_44599,N_42840);
xor U45549 (N_45549,N_42907,N_42470);
xnor U45550 (N_45550,N_40295,N_44606);
or U45551 (N_45551,N_40982,N_42013);
nor U45552 (N_45552,N_41836,N_40225);
nand U45553 (N_45553,N_40473,N_41983);
nor U45554 (N_45554,N_44154,N_43973);
or U45555 (N_45555,N_42123,N_44435);
nor U45556 (N_45556,N_42088,N_44171);
nor U45557 (N_45557,N_44360,N_41704);
or U45558 (N_45558,N_40517,N_40701);
and U45559 (N_45559,N_44235,N_44057);
and U45560 (N_45560,N_42814,N_41985);
and U45561 (N_45561,N_43491,N_41775);
or U45562 (N_45562,N_43472,N_43099);
or U45563 (N_45563,N_41842,N_44579);
nor U45564 (N_45564,N_41734,N_41519);
or U45565 (N_45565,N_42821,N_44113);
or U45566 (N_45566,N_42697,N_41532);
or U45567 (N_45567,N_40867,N_40585);
or U45568 (N_45568,N_43684,N_41095);
nand U45569 (N_45569,N_44809,N_44584);
or U45570 (N_45570,N_44789,N_40629);
nor U45571 (N_45571,N_44426,N_42142);
or U45572 (N_45572,N_41127,N_42646);
nand U45573 (N_45573,N_43848,N_40258);
xnor U45574 (N_45574,N_43439,N_40102);
xor U45575 (N_45575,N_44129,N_44236);
or U45576 (N_45576,N_42834,N_43471);
nor U45577 (N_45577,N_43910,N_42977);
and U45578 (N_45578,N_42850,N_44897);
nor U45579 (N_45579,N_44771,N_40320);
nor U45580 (N_45580,N_43822,N_40613);
xor U45581 (N_45581,N_41528,N_42531);
xnor U45582 (N_45582,N_40247,N_41675);
xor U45583 (N_45583,N_44215,N_41075);
or U45584 (N_45584,N_44724,N_40023);
and U45585 (N_45585,N_42394,N_43479);
or U45586 (N_45586,N_40091,N_40531);
nor U45587 (N_45587,N_42059,N_43919);
and U45588 (N_45588,N_40137,N_43120);
xnor U45589 (N_45589,N_41088,N_44138);
xnor U45590 (N_45590,N_41910,N_40694);
xor U45591 (N_45591,N_40638,N_43802);
nand U45592 (N_45592,N_41841,N_40968);
nor U45593 (N_45593,N_40999,N_42966);
nand U45594 (N_45594,N_40359,N_43321);
xor U45595 (N_45595,N_42643,N_44741);
or U45596 (N_45596,N_42355,N_44963);
and U45597 (N_45597,N_42509,N_44189);
nor U45598 (N_45598,N_44772,N_40451);
or U45599 (N_45599,N_43879,N_44743);
nor U45600 (N_45600,N_42410,N_41909);
or U45601 (N_45601,N_44421,N_41616);
and U45602 (N_45602,N_43854,N_43745);
nor U45603 (N_45603,N_43316,N_40314);
or U45604 (N_45604,N_43867,N_44336);
and U45605 (N_45605,N_40536,N_42268);
or U45606 (N_45606,N_44093,N_42895);
and U45607 (N_45607,N_43953,N_41343);
xnor U45608 (N_45608,N_42432,N_43655);
and U45609 (N_45609,N_41221,N_42564);
nor U45610 (N_45610,N_41214,N_41485);
nand U45611 (N_45611,N_43132,N_40044);
xnor U45612 (N_45612,N_41912,N_41689);
or U45613 (N_45613,N_42657,N_40543);
or U45614 (N_45614,N_40335,N_44733);
nor U45615 (N_45615,N_41818,N_43302);
nor U45616 (N_45616,N_44353,N_42984);
and U45617 (N_45617,N_42216,N_44744);
nand U45618 (N_45618,N_40794,N_40172);
nor U45619 (N_45619,N_41013,N_41770);
or U45620 (N_45620,N_41236,N_44881);
and U45621 (N_45621,N_40511,N_43275);
nand U45622 (N_45622,N_43273,N_43666);
nor U45623 (N_45623,N_41248,N_43818);
nand U45624 (N_45624,N_43567,N_44148);
and U45625 (N_45625,N_42593,N_40637);
and U45626 (N_45626,N_42719,N_41834);
and U45627 (N_45627,N_40649,N_40786);
nand U45628 (N_45628,N_42615,N_41416);
or U45629 (N_45629,N_42843,N_44111);
or U45630 (N_45630,N_43015,N_42999);
or U45631 (N_45631,N_40961,N_41275);
nand U45632 (N_45632,N_42662,N_44139);
nor U45633 (N_45633,N_44472,N_42143);
nor U45634 (N_45634,N_40181,N_43203);
nor U45635 (N_45635,N_41131,N_42466);
and U45636 (N_45636,N_44995,N_44460);
or U45637 (N_45637,N_44671,N_41625);
and U45638 (N_45638,N_43348,N_44127);
nor U45639 (N_45639,N_40978,N_44580);
nand U45640 (N_45640,N_43327,N_44902);
nor U45641 (N_45641,N_44934,N_41270);
and U45642 (N_45642,N_42200,N_40901);
or U45643 (N_45643,N_40807,N_42529);
nor U45644 (N_45644,N_43347,N_42630);
nand U45645 (N_45645,N_43710,N_44091);
nor U45646 (N_45646,N_42877,N_40471);
or U45647 (N_45647,N_41789,N_41587);
or U45648 (N_45648,N_44525,N_40506);
or U45649 (N_45649,N_42066,N_40241);
nor U45650 (N_45650,N_44773,N_44616);
and U45651 (N_45651,N_41358,N_42015);
xnor U45652 (N_45652,N_44343,N_44763);
nand U45653 (N_45653,N_42437,N_41741);
nor U45654 (N_45654,N_41079,N_43346);
nand U45655 (N_45655,N_41293,N_44370);
and U45656 (N_45656,N_44461,N_40392);
xor U45657 (N_45657,N_42753,N_44540);
or U45658 (N_45658,N_42795,N_40458);
or U45659 (N_45659,N_44072,N_40798);
and U45660 (N_45660,N_44634,N_41670);
and U45661 (N_45661,N_42734,N_40090);
nor U45662 (N_45662,N_41183,N_44874);
nand U45663 (N_45663,N_42590,N_42573);
or U45664 (N_45664,N_41545,N_44906);
xor U45665 (N_45665,N_44191,N_40768);
and U45666 (N_45666,N_44433,N_43632);
and U45667 (N_45667,N_42067,N_42829);
and U45668 (N_45668,N_41533,N_43861);
or U45669 (N_45669,N_41289,N_42496);
or U45670 (N_45670,N_41243,N_43909);
or U45671 (N_45671,N_41344,N_41327);
or U45672 (N_45672,N_40058,N_43622);
xnor U45673 (N_45673,N_42141,N_40460);
nor U45674 (N_45674,N_42731,N_43007);
nor U45675 (N_45675,N_40865,N_42562);
nor U45676 (N_45676,N_43805,N_43102);
xor U45677 (N_45677,N_41419,N_41707);
or U45678 (N_45678,N_42366,N_42783);
or U45679 (N_45679,N_42343,N_43839);
nand U45680 (N_45680,N_40200,N_41978);
xnor U45681 (N_45681,N_44562,N_44483);
or U45682 (N_45682,N_40868,N_44454);
nor U45683 (N_45683,N_42243,N_42299);
nand U45684 (N_45684,N_43920,N_44565);
nor U45685 (N_45685,N_42498,N_44999);
nor U45686 (N_45686,N_44664,N_44173);
nand U45687 (N_45687,N_41504,N_43417);
or U45688 (N_45688,N_41437,N_43351);
nor U45689 (N_45689,N_44737,N_43549);
and U45690 (N_45690,N_44800,N_43160);
nand U45691 (N_45691,N_40702,N_43791);
or U45692 (N_45692,N_40342,N_40882);
xor U45693 (N_45693,N_41796,N_42043);
xnor U45694 (N_45694,N_44985,N_43082);
nand U45695 (N_45695,N_43917,N_44469);
or U45696 (N_45696,N_43561,N_44047);
or U45697 (N_45697,N_41490,N_42168);
and U45698 (N_45698,N_42387,N_40412);
nor U45699 (N_45699,N_40311,N_40289);
and U45700 (N_45700,N_40499,N_43197);
xnor U45701 (N_45701,N_41200,N_42778);
nor U45702 (N_45702,N_44675,N_42518);
and U45703 (N_45703,N_42858,N_40045);
nor U45704 (N_45704,N_40609,N_40783);
nor U45705 (N_45705,N_42207,N_44765);
or U45706 (N_45706,N_42160,N_41426);
or U45707 (N_45707,N_41181,N_42282);
xnor U45708 (N_45708,N_43060,N_42844);
xnor U45709 (N_45709,N_43268,N_43399);
and U45710 (N_45710,N_40345,N_40488);
and U45711 (N_45711,N_44497,N_40237);
xor U45712 (N_45712,N_43156,N_44180);
xor U45713 (N_45713,N_41239,N_41630);
nand U45714 (N_45714,N_40399,N_44890);
xor U45715 (N_45715,N_40700,N_44705);
xor U45716 (N_45716,N_40306,N_43869);
nor U45717 (N_45717,N_42676,N_40895);
or U45718 (N_45718,N_44908,N_40226);
and U45719 (N_45719,N_41697,N_42613);
nand U45720 (N_45720,N_40728,N_42191);
xnor U45721 (N_45721,N_40018,N_44932);
xnor U45722 (N_45722,N_44198,N_41854);
xor U45723 (N_45723,N_40327,N_40953);
or U45724 (N_45724,N_44657,N_41352);
nand U45725 (N_45725,N_43716,N_43670);
and U45726 (N_45726,N_44392,N_42742);
nand U45727 (N_45727,N_43234,N_43930);
or U45728 (N_45728,N_41943,N_40337);
or U45729 (N_45729,N_42277,N_40100);
and U45730 (N_45730,N_41694,N_44679);
or U45731 (N_45731,N_42802,N_43070);
nand U45732 (N_45732,N_44011,N_43201);
or U45733 (N_45733,N_44769,N_41622);
and U45734 (N_45734,N_40167,N_42714);
nor U45735 (N_45735,N_43464,N_41705);
nand U45736 (N_45736,N_40804,N_40832);
nand U45737 (N_45737,N_43170,N_42374);
xnor U45738 (N_45738,N_40734,N_43345);
nand U45739 (N_45739,N_42103,N_43886);
xor U45740 (N_45740,N_41302,N_40926);
nand U45741 (N_45741,N_43726,N_40899);
or U45742 (N_45742,N_43569,N_44907);
xor U45743 (N_45743,N_41712,N_43434);
or U45744 (N_45744,N_42640,N_43504);
or U45745 (N_45745,N_41731,N_40695);
xor U45746 (N_45746,N_43783,N_43687);
or U45747 (N_45747,N_41692,N_42991);
nor U45748 (N_45748,N_42120,N_41351);
or U45749 (N_45749,N_42458,N_44718);
and U45750 (N_45750,N_43990,N_40697);
nor U45751 (N_45751,N_41999,N_44994);
and U45752 (N_45752,N_41192,N_41492);
nand U45753 (N_45753,N_40888,N_42149);
or U45754 (N_45754,N_41794,N_44648);
or U45755 (N_45755,N_41726,N_43269);
xnor U45756 (N_45756,N_42894,N_42233);
and U45757 (N_45757,N_44875,N_41472);
or U45758 (N_45758,N_40748,N_44536);
nand U45759 (N_45759,N_41728,N_41231);
and U45760 (N_45760,N_40030,N_40131);
xor U45761 (N_45761,N_43343,N_43428);
xor U45762 (N_45762,N_42899,N_42336);
nand U45763 (N_45763,N_43198,N_42935);
nor U45764 (N_45764,N_44321,N_41633);
nor U45765 (N_45765,N_44946,N_40769);
xor U45766 (N_45766,N_44471,N_40841);
nand U45767 (N_45767,N_42278,N_44563);
or U45768 (N_45768,N_43137,N_41944);
nor U45769 (N_45769,N_44410,N_44790);
nand U45770 (N_45770,N_44133,N_43063);
and U45771 (N_45771,N_43310,N_43545);
or U45772 (N_45772,N_40421,N_44545);
nor U45773 (N_45773,N_44799,N_43989);
xnor U45774 (N_45774,N_44231,N_43813);
xor U45775 (N_45775,N_44306,N_44140);
nand U45776 (N_45776,N_42406,N_41489);
xor U45777 (N_45777,N_44272,N_40752);
nor U45778 (N_45778,N_42313,N_41477);
nand U45779 (N_45779,N_44156,N_43468);
or U45780 (N_45780,N_40328,N_43338);
nand U45781 (N_45781,N_43278,N_41338);
or U45782 (N_45782,N_41500,N_40553);
nand U45783 (N_45783,N_42585,N_43407);
or U45784 (N_45784,N_42370,N_44016);
or U45785 (N_45785,N_41357,N_41128);
or U45786 (N_45786,N_42076,N_44604);
nor U45787 (N_45787,N_41433,N_44429);
and U45788 (N_45788,N_44953,N_41432);
or U45789 (N_45789,N_44693,N_40959);
or U45790 (N_45790,N_41767,N_43754);
and U45791 (N_45791,N_43271,N_42612);
xor U45792 (N_45792,N_40152,N_42473);
and U45793 (N_45793,N_42686,N_41452);
nand U45794 (N_45794,N_43331,N_43432);
nand U45795 (N_45795,N_40302,N_41116);
nand U45796 (N_45796,N_44958,N_42446);
or U45797 (N_45797,N_42956,N_41196);
nor U45798 (N_45798,N_43626,N_43426);
and U45799 (N_45799,N_43577,N_43384);
nand U45800 (N_45800,N_44157,N_40427);
nor U45801 (N_45801,N_42976,N_41564);
and U45802 (N_45802,N_43481,N_42077);
xor U45803 (N_45803,N_40823,N_44293);
nand U45804 (N_45804,N_43001,N_43314);
and U45805 (N_45805,N_41326,N_40089);
xnor U45806 (N_45806,N_41174,N_40270);
or U45807 (N_45807,N_42841,N_43225);
xnor U45808 (N_45808,N_40627,N_41677);
or U45809 (N_45809,N_43288,N_41223);
nor U45810 (N_45810,N_44325,N_43466);
nand U45811 (N_45811,N_41696,N_41389);
xor U45812 (N_45812,N_41860,N_44109);
nand U45813 (N_45813,N_42185,N_43941);
xor U45814 (N_45814,N_43305,N_44667);
and U45815 (N_45815,N_40897,N_42425);
and U45816 (N_45816,N_42295,N_40228);
and U45817 (N_45817,N_42545,N_40157);
xor U45818 (N_45818,N_43853,N_42384);
nor U45819 (N_45819,N_43676,N_42463);
nor U45820 (N_45820,N_40580,N_44759);
nand U45821 (N_45821,N_43884,N_44432);
xnor U45822 (N_45822,N_42092,N_44424);
or U45823 (N_45823,N_42228,N_44818);
nor U45824 (N_45824,N_44811,N_43773);
nand U45825 (N_45825,N_41956,N_44876);
nand U45826 (N_45826,N_43750,N_43730);
xor U45827 (N_45827,N_41572,N_41738);
xor U45828 (N_45828,N_43903,N_43173);
or U45829 (N_45829,N_41965,N_40941);
nand U45830 (N_45830,N_40159,N_42978);
nor U45831 (N_45831,N_40093,N_40980);
nor U45832 (N_45832,N_43252,N_44530);
nand U45833 (N_45833,N_41512,N_43155);
or U45834 (N_45834,N_43952,N_42696);
xor U45835 (N_45835,N_44265,N_41064);
and U45836 (N_45836,N_42373,N_42206);
or U45837 (N_45837,N_44685,N_42079);
or U45838 (N_45838,N_44959,N_42685);
and U45839 (N_45839,N_43451,N_42210);
nor U45840 (N_45840,N_43993,N_44914);
and U45841 (N_45841,N_43779,N_44013);
or U45842 (N_45842,N_44833,N_41894);
and U45843 (N_45843,N_43422,N_42774);
xor U45844 (N_45844,N_40249,N_43500);
nand U45845 (N_45845,N_43031,N_44163);
nand U45846 (N_45846,N_40604,N_42421);
nor U45847 (N_45847,N_43499,N_40986);
xnor U45848 (N_45848,N_40128,N_40444);
and U45849 (N_45849,N_43490,N_41109);
xnor U45850 (N_45850,N_44872,N_40206);
nand U45851 (N_45851,N_44997,N_42671);
nor U45852 (N_45852,N_42472,N_41690);
nand U45853 (N_45853,N_40022,N_43631);
nand U45854 (N_45854,N_41855,N_43210);
and U45855 (N_45855,N_43077,N_40060);
or U45856 (N_45856,N_44396,N_43888);
xnor U45857 (N_45857,N_43266,N_41065);
nor U45858 (N_45858,N_44068,N_43340);
nand U45859 (N_45859,N_43161,N_41863);
nand U45860 (N_45860,N_42305,N_42226);
xnor U45861 (N_45861,N_42549,N_42276);
and U45862 (N_45862,N_44713,N_41321);
and U45863 (N_45863,N_44205,N_44152);
nand U45864 (N_45864,N_41648,N_40960);
and U45865 (N_45865,N_44263,N_43441);
xor U45866 (N_45866,N_44318,N_40239);
nand U45867 (N_45867,N_40433,N_44894);
nand U45868 (N_45868,N_41425,N_43633);
and U45869 (N_45869,N_42968,N_44208);
and U45870 (N_45870,N_42254,N_43357);
nor U45871 (N_45871,N_44746,N_43409);
xnor U45872 (N_45872,N_40989,N_44136);
and U45873 (N_45873,N_40466,N_42106);
nor U45874 (N_45874,N_42085,N_41161);
or U45875 (N_45875,N_43979,N_40285);
xor U45876 (N_45876,N_41554,N_40992);
nor U45877 (N_45877,N_43560,N_41623);
nand U45878 (N_45878,N_44301,N_43574);
and U45879 (N_45879,N_40561,N_42567);
nand U45880 (N_45880,N_43580,N_40889);
xnor U45881 (N_45881,N_40610,N_42690);
nand U45882 (N_45882,N_40257,N_42642);
nor U45883 (N_45883,N_41762,N_42986);
nor U45884 (N_45884,N_42761,N_42095);
and U45885 (N_45885,N_40927,N_41631);
or U45886 (N_45886,N_42019,N_41971);
nor U45887 (N_45887,N_44577,N_43740);
or U45888 (N_45888,N_43611,N_43404);
nor U45889 (N_45889,N_44597,N_42847);
and U45890 (N_45890,N_41086,N_42933);
nor U45891 (N_45891,N_42435,N_44118);
nand U45892 (N_45892,N_44227,N_43377);
xnor U45893 (N_45893,N_41848,N_43100);
xnor U45894 (N_45894,N_41585,N_40544);
and U45895 (N_45895,N_42583,N_42635);
nor U45896 (N_45896,N_42883,N_44251);
and U45897 (N_45897,N_41274,N_40853);
xnor U45898 (N_45898,N_42832,N_40190);
or U45899 (N_45899,N_41930,N_40666);
or U45900 (N_45900,N_43487,N_40481);
nor U45901 (N_45901,N_40902,N_40526);
nor U45902 (N_45902,N_41548,N_42181);
and U45903 (N_45903,N_42152,N_43196);
or U45904 (N_45904,N_44669,N_40679);
nand U45905 (N_45905,N_41830,N_40596);
or U45906 (N_45906,N_42151,N_44250);
nor U45907 (N_45907,N_40231,N_44291);
or U45908 (N_45908,N_40117,N_44390);
nand U45909 (N_45909,N_42385,N_40338);
and U45910 (N_45910,N_42068,N_43000);
nand U45911 (N_45911,N_41284,N_42315);
xor U45912 (N_45912,N_42298,N_44961);
or U45913 (N_45913,N_40205,N_44441);
and U45914 (N_45914,N_41057,N_44558);
nor U45915 (N_45915,N_42113,N_41534);
xor U45916 (N_45916,N_43306,N_44638);
or U45917 (N_45917,N_43981,N_44854);
or U45918 (N_45918,N_42102,N_40232);
or U45919 (N_45919,N_43330,N_40532);
nand U45920 (N_45920,N_44417,N_43871);
nand U45921 (N_45921,N_44614,N_41315);
or U45922 (N_45922,N_40415,N_40647);
or U45923 (N_45923,N_41333,N_40432);
nand U45924 (N_45924,N_41781,N_41077);
nand U45925 (N_45925,N_41977,N_44885);
or U45926 (N_45926,N_41156,N_40942);
xnor U45927 (N_45927,N_40836,N_41699);
or U45928 (N_45928,N_43619,N_44379);
nand U45929 (N_45929,N_44921,N_44501);
or U45930 (N_45930,N_43292,N_43324);
nor U45931 (N_45931,N_44443,N_41264);
nand U45932 (N_45932,N_40653,N_41903);
nor U45933 (N_45933,N_44819,N_40846);
or U45934 (N_45934,N_40170,N_41964);
or U45935 (N_45935,N_40958,N_44300);
nand U45936 (N_45936,N_42263,N_42711);
and U45937 (N_45937,N_44190,N_42097);
nand U45938 (N_45938,N_44334,N_43239);
nand U45939 (N_45939,N_41959,N_44609);
nor U45940 (N_45940,N_42798,N_44755);
nor U45941 (N_45941,N_41137,N_41851);
xor U45942 (N_45942,N_40862,N_44258);
xnor U45943 (N_45943,N_44505,N_42889);
nand U45944 (N_45944,N_43388,N_43615);
nand U45945 (N_45945,N_41857,N_40453);
or U45946 (N_45946,N_44899,N_41996);
or U45947 (N_45947,N_43177,N_43553);
or U45948 (N_45948,N_44652,N_41405);
nand U45949 (N_45949,N_42508,N_44660);
and U45950 (N_45950,N_40431,N_41052);
xor U45951 (N_45951,N_42484,N_42972);
nand U45952 (N_45952,N_42169,N_42766);
nand U45953 (N_45953,N_40705,N_42055);
or U45954 (N_45954,N_44393,N_41755);
nor U45955 (N_45955,N_43770,N_44271);
nand U45956 (N_45956,N_42397,N_44088);
or U45957 (N_45957,N_42866,N_44656);
xor U45958 (N_45958,N_41888,N_41721);
and U45959 (N_45959,N_44931,N_44598);
nor U45960 (N_45960,N_44014,N_40478);
nand U45961 (N_45961,N_40549,N_44688);
nand U45962 (N_45962,N_42445,N_40704);
xnor U45963 (N_45963,N_42412,N_43704);
or U45964 (N_45964,N_41126,N_42351);
or U45965 (N_45965,N_41636,N_41082);
nor U45966 (N_45966,N_44528,N_40503);
nor U45967 (N_45967,N_43984,N_41599);
nand U45968 (N_45968,N_42188,N_42940);
and U45969 (N_45969,N_43788,N_43572);
or U45970 (N_45970,N_40080,N_43759);
nand U45971 (N_45971,N_41812,N_44785);
nor U45972 (N_45972,N_43548,N_43665);
or U45973 (N_45973,N_44554,N_42602);
and U45974 (N_45974,N_42932,N_43498);
nand U45975 (N_45975,N_43543,N_42350);
nand U45976 (N_45976,N_44911,N_40470);
nand U45977 (N_45977,N_40401,N_44229);
xnor U45978 (N_45978,N_41938,N_41827);
and U45979 (N_45979,N_43152,N_44864);
nor U45980 (N_45980,N_43402,N_44791);
and U45981 (N_45981,N_44462,N_43738);
or U45982 (N_45982,N_44925,N_42782);
or U45983 (N_45983,N_44843,N_43566);
nand U45984 (N_45984,N_42133,N_40594);
xor U45985 (N_45985,N_44731,N_40541);
xor U45986 (N_45986,N_43550,N_41579);
xor U45987 (N_45987,N_42375,N_43136);
and U45988 (N_45988,N_43274,N_40149);
or U45989 (N_45989,N_42806,N_42636);
and U45990 (N_45990,N_40693,N_40848);
xnor U45991 (N_45991,N_43647,N_43775);
or U45992 (N_45992,N_41778,N_44035);
or U45993 (N_45993,N_44620,N_42534);
nand U45994 (N_45994,N_44559,N_41798);
or U45995 (N_45995,N_42913,N_41143);
nor U45996 (N_45996,N_41717,N_40418);
xor U45997 (N_45997,N_41747,N_42495);
and U45998 (N_45998,N_41217,N_41530);
nand U45999 (N_45999,N_40161,N_40021);
xor U46000 (N_46000,N_44817,N_40671);
and U46001 (N_46001,N_43121,N_40407);
or U46002 (N_46002,N_40235,N_44867);
nand U46003 (N_46003,N_42249,N_44492);
and U46004 (N_46004,N_42259,N_41885);
and U46005 (N_46005,N_40640,N_43352);
nor U46006 (N_46006,N_40377,N_40985);
xor U46007 (N_46007,N_43148,N_41113);
nand U46008 (N_46008,N_40689,N_44970);
or U46009 (N_46009,N_41803,N_42131);
nor U46010 (N_46010,N_42051,N_40331);
xor U46011 (N_46011,N_43334,N_41560);
nor U46012 (N_46012,N_44416,N_44121);
or U46013 (N_46013,N_42712,N_40957);
nand U46014 (N_46014,N_44165,N_44342);
xnor U46015 (N_46015,N_42027,N_42480);
nand U46016 (N_46016,N_41454,N_40894);
and U46017 (N_46017,N_40173,N_44712);
xnor U46018 (N_46018,N_40199,N_41961);
nand U46019 (N_46019,N_40274,N_43959);
xnor U46020 (N_46020,N_43709,N_43677);
nor U46021 (N_46021,N_42303,N_42379);
and U46022 (N_46022,N_44246,N_43623);
and U46023 (N_46023,N_43391,N_41001);
nand U46024 (N_46024,N_44097,N_42946);
nor U46025 (N_46025,N_43360,N_43557);
nand U46026 (N_46026,N_40872,N_41250);
or U46027 (N_46027,N_41069,N_41479);
xnor U46028 (N_46028,N_40584,N_44211);
and U46029 (N_46029,N_41583,N_40615);
nand U46030 (N_46030,N_44557,N_43244);
or U46031 (N_46031,N_43270,N_43246);
or U46032 (N_46032,N_44590,N_40272);
nand U46033 (N_46033,N_40935,N_41048);
xnor U46034 (N_46034,N_42329,N_41628);
or U46035 (N_46035,N_42164,N_41176);
nor U46036 (N_46036,N_40771,N_40255);
xor U46037 (N_46037,N_44051,N_42500);
or U46038 (N_46038,N_44845,N_44623);
and U46039 (N_46039,N_43859,N_41204);
or U46040 (N_46040,N_43599,N_40464);
nor U46041 (N_46041,N_44303,N_44723);
and U46042 (N_46042,N_44248,N_44711);
nand U46043 (N_46043,N_40028,N_43644);
nand U46044 (N_46044,N_42111,N_44046);
nand U46045 (N_46045,N_43415,N_43827);
nand U46046 (N_46046,N_43870,N_43291);
xnor U46047 (N_46047,N_43725,N_43913);
and U46048 (N_46048,N_40062,N_40741);
nand U46049 (N_46049,N_40497,N_42167);
or U46050 (N_46050,N_42304,N_42150);
xnor U46051 (N_46051,N_43570,N_40998);
or U46052 (N_46052,N_42349,N_43935);
nor U46053 (N_46053,N_40243,N_42297);
or U46054 (N_46054,N_41543,N_43907);
or U46055 (N_46055,N_44916,N_41814);
nand U46056 (N_46056,N_44204,N_41182);
nand U46057 (N_46057,N_42176,N_41922);
nor U46058 (N_46058,N_43516,N_42835);
and U46059 (N_46059,N_41709,N_41806);
or U46060 (N_46060,N_43998,N_40657);
and U46061 (N_46061,N_40126,N_40566);
nor U46062 (N_46062,N_43496,N_43350);
xor U46063 (N_46063,N_41620,N_43022);
nor U46064 (N_46064,N_41319,N_44551);
and U46065 (N_46065,N_43739,N_40930);
nor U46066 (N_46066,N_42557,N_40260);
or U46067 (N_46067,N_41448,N_40996);
nor U46068 (N_46068,N_44225,N_40576);
xor U46069 (N_46069,N_43690,N_44810);
nor U46070 (N_46070,N_40670,N_40828);
or U46071 (N_46071,N_42376,N_43830);
xor U46072 (N_46072,N_42125,N_43591);
nand U46073 (N_46073,N_43064,N_40351);
nor U46074 (N_46074,N_43017,N_41624);
or U46075 (N_46075,N_42112,N_43460);
or U46076 (N_46076,N_44813,N_41899);
xor U46077 (N_46077,N_42527,N_43686);
nor U46078 (N_46078,N_42222,N_40281);
or U46079 (N_46079,N_43957,N_43486);
xnor U46080 (N_46080,N_42334,N_42219);
nor U46081 (N_46081,N_41654,N_40813);
and U46082 (N_46082,N_40644,N_44803);
and U46083 (N_46083,N_41296,N_42171);
or U46084 (N_46084,N_43315,N_40916);
and U46085 (N_46085,N_40861,N_42070);
nor U46086 (N_46086,N_40881,N_43354);
nor U46087 (N_46087,N_42891,N_41115);
nor U46088 (N_46088,N_44437,N_43986);
and U46089 (N_46089,N_43649,N_40368);
and U46090 (N_46090,N_44172,N_43228);
xnor U46091 (N_46091,N_44219,N_43931);
or U46092 (N_46092,N_42346,N_44059);
or U46093 (N_46093,N_43221,N_44689);
nand U46094 (N_46094,N_43242,N_40154);
or U46095 (N_46095,N_41280,N_43071);
xnor U46096 (N_46096,N_42822,N_44930);
and U46097 (N_46097,N_41244,N_40408);
nand U46098 (N_46098,N_41070,N_42652);
and U46099 (N_46099,N_42314,N_42816);
and U46100 (N_46100,N_44967,N_40533);
nand U46101 (N_46101,N_42856,N_43034);
and U46102 (N_46102,N_40454,N_43284);
and U46103 (N_46103,N_42571,N_40214);
nand U46104 (N_46104,N_42906,N_44398);
xor U46105 (N_46105,N_43130,N_40816);
nand U46106 (N_46106,N_44548,N_40799);
nand U46107 (N_46107,N_43988,N_40805);
nor U46108 (N_46108,N_40027,N_41936);
or U46109 (N_46109,N_44860,N_44169);
xnor U46110 (N_46110,N_44567,N_44734);
and U46111 (N_46111,N_44307,N_41649);
xor U46112 (N_46112,N_44513,N_44696);
nor U46113 (N_46113,N_42886,N_42525);
and U46114 (N_46114,N_43885,N_42953);
nor U46115 (N_46115,N_43057,N_43116);
xor U46116 (N_46116,N_44865,N_40939);
or U46117 (N_46117,N_43657,N_42540);
and U46118 (N_46118,N_40567,N_43387);
nor U46119 (N_46119,N_44131,N_40522);
xnor U46120 (N_46120,N_41995,N_43128);
nor U46121 (N_46121,N_41776,N_42032);
xnor U46122 (N_46122,N_40063,N_42062);
nor U46123 (N_46123,N_44105,N_44879);
xor U46124 (N_46124,N_44533,N_41765);
and U46125 (N_46125,N_41508,N_43300);
or U46126 (N_46126,N_40291,N_40082);
or U46127 (N_46127,N_44494,N_44056);
nor U46128 (N_46128,N_40946,N_43240);
xor U46129 (N_46129,N_44506,N_43021);
and U46130 (N_46130,N_44704,N_41904);
nand U46131 (N_46131,N_44383,N_41329);
and U46132 (N_46132,N_44310,N_43044);
xnor U46133 (N_46133,N_42997,N_42945);
nor U46134 (N_46134,N_41408,N_43503);
and U46135 (N_46135,N_40687,N_41565);
xnor U46136 (N_46136,N_44782,N_42324);
or U46137 (N_46137,N_44073,N_40296);
nor U46138 (N_46138,N_42493,N_42667);
or U46139 (N_46139,N_42229,N_44032);
nor U46140 (N_46140,N_40631,N_43098);
nand U46141 (N_46141,N_41076,N_44754);
and U46142 (N_46142,N_40928,N_42996);
nor U46143 (N_46143,N_44378,N_41210);
xnor U46144 (N_46144,N_43307,N_43826);
nor U46145 (N_46145,N_43950,N_41795);
nor U46146 (N_46146,N_43969,N_41799);
nand U46147 (N_46147,N_41304,N_40965);
and U46148 (N_46148,N_41574,N_42702);
nor U46149 (N_46149,N_43081,N_43267);
and U46150 (N_46150,N_41580,N_41646);
nand U46151 (N_46151,N_43760,N_43119);
xor U46152 (N_46152,N_40202,N_43978);
or U46153 (N_46153,N_40721,N_40120);
or U46154 (N_46154,N_43159,N_42848);
and U46155 (N_46155,N_42511,N_42266);
or U46156 (N_46156,N_40276,N_41377);
nor U46157 (N_46157,N_44069,N_42372);
or U46158 (N_46158,N_41184,N_44233);
or U46159 (N_46159,N_43012,N_42442);
or U46160 (N_46160,N_42554,N_43459);
and U46161 (N_46161,N_40046,N_42417);
nand U46162 (N_46162,N_44561,N_40189);
and U46163 (N_46163,N_40948,N_42488);
and U46164 (N_46164,N_41598,N_40053);
xnor U46165 (N_46165,N_43053,N_43834);
nand U46166 (N_46166,N_44851,N_43374);
nand U46167 (N_46167,N_40564,N_44200);
nand U46168 (N_46168,N_43008,N_41058);
nand U46169 (N_46169,N_42553,N_40645);
nand U46170 (N_46170,N_43794,N_41526);
or U46171 (N_46171,N_41849,N_44280);
nand U46172 (N_46172,N_40581,N_40508);
nor U46173 (N_46173,N_42779,N_44965);
and U46174 (N_46174,N_44801,N_44950);
nand U46175 (N_46175,N_43944,N_41931);
or U46176 (N_46176,N_44366,N_40402);
nand U46177 (N_46177,N_41215,N_43205);
nand U46178 (N_46178,N_43712,N_41641);
nor U46179 (N_46179,N_41220,N_40114);
nand U46180 (N_46180,N_44174,N_41371);
and U46181 (N_46181,N_41643,N_44619);
nor U46182 (N_46182,N_42618,N_42124);
nor U46183 (N_46183,N_40746,N_42528);
or U46184 (N_46184,N_41040,N_40187);
xor U46185 (N_46185,N_41242,N_41443);
nand U46186 (N_46186,N_40642,N_44406);
or U46187 (N_46187,N_41226,N_43512);
or U46188 (N_46188,N_40332,N_44464);
nand U46189 (N_46189,N_40984,N_40007);
or U46190 (N_46190,N_42165,N_42280);
nand U46191 (N_46191,N_44727,N_40011);
nor U46192 (N_46192,N_43883,N_42264);
nand U46193 (N_46193,N_43186,N_44823);
xor U46194 (N_46194,N_41635,N_40582);
xnor U46195 (N_46195,N_42831,N_44770);
or U46196 (N_46196,N_42232,N_43763);
nor U46197 (N_46197,N_42247,N_42215);
xnor U46198 (N_46198,N_41499,N_40929);
xor U46199 (N_46199,N_44589,N_41946);
nand U46200 (N_46200,N_40572,N_40634);
nand U46201 (N_46201,N_40185,N_43488);
and U46202 (N_46202,N_40483,N_42660);
nand U46203 (N_46203,N_44058,N_41468);
or U46204 (N_46204,N_41356,N_42872);
nor U46205 (N_46205,N_44984,N_42775);
xor U46206 (N_46206,N_41627,N_40020);
xnor U46207 (N_46207,N_43552,N_40796);
and U46208 (N_46208,N_42345,N_43213);
nor U46209 (N_46209,N_40824,N_44187);
xnor U46210 (N_46210,N_43525,N_41122);
and U46211 (N_46211,N_42109,N_42344);
nand U46212 (N_46212,N_41725,N_41044);
xor U46213 (N_46213,N_42920,N_44787);
nand U46214 (N_46214,N_40288,N_43295);
nand U46215 (N_46215,N_44568,N_44992);
nand U46216 (N_46216,N_44002,N_42499);
nor U46217 (N_46217,N_41099,N_44534);
or U46218 (N_46218,N_42610,N_44149);
nand U46219 (N_46219,N_40871,N_43900);
or U46220 (N_46220,N_42729,N_43943);
and U46221 (N_46221,N_41434,N_41645);
nor U46222 (N_46222,N_42036,N_40887);
nand U46223 (N_46223,N_44793,N_42584);
xnor U46224 (N_46224,N_41537,N_44070);
or U46225 (N_46225,N_43513,N_41211);
and U46226 (N_46226,N_44516,N_41370);
xnor U46227 (N_46227,N_41597,N_42126);
nor U46228 (N_46228,N_40325,N_43026);
nand U46229 (N_46229,N_44756,N_43427);
nor U46230 (N_46230,N_41203,N_40142);
xor U46231 (N_46231,N_42599,N_40107);
nor U46232 (N_46232,N_43397,N_40381);
nand U46233 (N_46233,N_42147,N_42720);
nand U46234 (N_46234,N_44762,N_44141);
and U46235 (N_46235,N_41385,N_41019);
xnor U46236 (N_46236,N_40417,N_42286);
nand U46237 (N_46237,N_44729,N_42144);
nor U46238 (N_46238,N_40641,N_43837);
nand U46239 (N_46239,N_44267,N_42318);
xor U46240 (N_46240,N_44295,N_43390);
xor U46241 (N_46241,N_40764,N_43140);
and U46242 (N_46242,N_43394,N_43771);
nor U46243 (N_46243,N_43659,N_43255);
xnor U46244 (N_46244,N_44617,N_44913);
and U46245 (N_46245,N_40562,N_40240);
xnor U46246 (N_46246,N_42736,N_44491);
and U46247 (N_46247,N_40479,N_44871);
xnor U46248 (N_46248,N_40227,N_40068);
nand U46249 (N_46249,N_41149,N_41679);
nand U46250 (N_46250,N_44912,N_43579);
nor U46251 (N_46251,N_43131,N_42267);
xor U46252 (N_46252,N_42026,N_40761);
or U46253 (N_46253,N_41607,N_40682);
xor U46254 (N_46254,N_41901,N_40801);
nor U46255 (N_46255,N_41399,N_41661);
and U46256 (N_46256,N_41130,N_42162);
nand U46257 (N_46257,N_40108,N_40618);
and U46258 (N_46258,N_44112,N_44100);
xnor U46259 (N_46259,N_40936,N_42581);
xnor U46260 (N_46260,N_40720,N_41166);
and U46261 (N_46261,N_44061,N_41170);
xnor U46262 (N_46262,N_42231,N_42512);
nand U46263 (N_46263,N_41718,N_40303);
xnor U46264 (N_46264,N_41417,N_43373);
nand U46265 (N_46265,N_40250,N_41638);
nor U46266 (N_46266,N_41132,N_40064);
nor U46267 (N_46267,N_43474,N_40520);
nand U46268 (N_46268,N_40560,N_42608);
nor U46269 (N_46269,N_40523,N_42401);
nand U46270 (N_46270,N_42042,N_44350);
or U46271 (N_46271,N_43724,N_41951);
or U46272 (N_46272,N_41012,N_41659);
nor U46273 (N_46273,N_41511,N_41164);
nand U46274 (N_46274,N_42246,N_42717);
xor U46275 (N_46275,N_41402,N_40354);
nand U46276 (N_46276,N_43530,N_41852);
or U46277 (N_46277,N_42022,N_41205);
nand U46278 (N_46278,N_44094,N_40651);
and U46279 (N_46279,N_43289,N_42408);
nand U46280 (N_46280,N_41238,N_44900);
or U46281 (N_46281,N_40763,N_43010);
nand U46282 (N_46282,N_42960,N_44000);
nor U46283 (N_46283,N_42340,N_40774);
nand U46284 (N_46284,N_43037,N_43694);
or U46285 (N_46285,N_43029,N_40612);
nand U46286 (N_46286,N_44550,N_43874);
nor U46287 (N_46287,N_42420,N_41051);
or U46288 (N_46288,N_40356,N_44053);
nor U46289 (N_46289,N_41041,N_44582);
or U46290 (N_46290,N_43216,N_43329);
xor U46291 (N_46291,N_43123,N_40914);
xor U46292 (N_46292,N_41060,N_40490);
or U46293 (N_46293,N_43294,N_41768);
or U46294 (N_46294,N_40122,N_44517);
xor U46295 (N_46295,N_44687,N_42826);
or U46296 (N_46296,N_44690,N_44380);
nor U46297 (N_46297,N_44150,N_40484);
nor U46298 (N_46298,N_42409,N_42195);
and U46299 (N_46299,N_42075,N_40852);
and U46300 (N_46300,N_44493,N_40220);
or U46301 (N_46301,N_43363,N_43243);
nor U46302 (N_46302,N_44884,N_41409);
or U46303 (N_46303,N_42090,N_43162);
or U46304 (N_46304,N_42089,N_43598);
xor U46305 (N_46305,N_42196,N_40856);
or U46306 (N_46306,N_40758,N_40782);
or U46307 (N_46307,N_42172,N_40203);
or U46308 (N_46308,N_40014,N_40699);
xnor U46309 (N_46309,N_41290,N_42094);
or U46310 (N_46310,N_43785,N_40436);
xnor U46311 (N_46311,N_42389,N_44197);
nor U46312 (N_46312,N_41171,N_44776);
xor U46313 (N_46313,N_43971,N_44101);
nand U46314 (N_46314,N_43065,N_41003);
or U46315 (N_46315,N_42105,N_42154);
and U46316 (N_46316,N_43593,N_42517);
or U46317 (N_46317,N_40732,N_40041);
nor U46318 (N_46318,N_44937,N_41896);
xor U46319 (N_46319,N_44451,N_42004);
nand U46320 (N_46320,N_41247,N_42949);
nor U46321 (N_46321,N_43780,N_40441);
nor U46322 (N_46322,N_40073,N_41461);
or U46323 (N_46323,N_41937,N_40155);
or U46324 (N_46324,N_42732,N_41207);
nand U46325 (N_46325,N_44085,N_42910);
nand U46326 (N_46326,N_42328,N_41886);
nand U46327 (N_46327,N_43335,N_44658);
and U46328 (N_46328,N_44452,N_42801);
and U46329 (N_46329,N_40383,N_40656);
nand U46330 (N_46330,N_41054,N_43590);
nand U46331 (N_46331,N_43565,N_40759);
and U46332 (N_46332,N_41503,N_44242);
nand U46333 (N_46333,N_41802,N_40817);
nand U46334 (N_46334,N_40290,N_40144);
xor U46335 (N_46335,N_44943,N_44691);
or U46336 (N_46336,N_44698,N_43336);
or U46337 (N_46337,N_41650,N_44119);
xnor U46338 (N_46338,N_44630,N_41754);
and U46339 (N_46339,N_43636,N_40439);
and U46340 (N_46340,N_44402,N_40396);
and U46341 (N_46341,N_40921,N_42964);
or U46342 (N_46342,N_40745,N_40557);
or U46343 (N_46343,N_40509,N_43616);
nand U46344 (N_46344,N_44775,N_40900);
and U46345 (N_46345,N_43208,N_40224);
nand U46346 (N_46346,N_42539,N_44479);
xor U46347 (N_46347,N_41497,N_42436);
nand U46348 (N_46348,N_41666,N_42911);
xnor U46349 (N_46349,N_42039,N_41536);
and U46350 (N_46350,N_43209,N_43091);
xor U46351 (N_46351,N_42220,N_41412);
nor U46352 (N_46352,N_44974,N_44978);
nor U46353 (N_46353,N_43539,N_41613);
nand U46354 (N_46354,N_44395,N_40731);
nand U46355 (N_46355,N_42422,N_42317);
and U46356 (N_46356,N_42134,N_43229);
nand U46357 (N_46357,N_42586,N_40391);
xor U46358 (N_46358,N_41626,N_41887);
xnor U46359 (N_46359,N_42980,N_44720);
nor U46360 (N_46360,N_42616,N_41011);
and U46361 (N_46361,N_42658,N_44503);
and U46362 (N_46362,N_42332,N_43997);
nand U46363 (N_46363,N_40238,N_42709);
or U46364 (N_46364,N_40736,N_42288);
and U46365 (N_46365,N_43749,N_43601);
or U46366 (N_46366,N_40112,N_43856);
xor U46367 (N_46367,N_41307,N_42975);
nor U46368 (N_46368,N_44287,N_42656);
nor U46369 (N_46369,N_40322,N_42898);
and U46370 (N_46370,N_42929,N_42787);
and U46371 (N_46371,N_44742,N_42382);
or U46372 (N_46372,N_43682,N_43165);
xor U46373 (N_46373,N_41257,N_42434);
or U46374 (N_46374,N_41893,N_40230);
and U46375 (N_46375,N_43151,N_42427);
and U46376 (N_46376,N_44386,N_42129);
or U46377 (N_46377,N_43259,N_43002);
nand U46378 (N_46378,N_41866,N_43456);
nor U46379 (N_46379,N_41375,N_40406);
xor U46380 (N_46380,N_44122,N_43972);
and U46381 (N_46381,N_44339,N_43921);
xor U46382 (N_46382,N_43093,N_44895);
nand U46383 (N_46383,N_44986,N_42462);
or U46384 (N_46384,N_41760,N_40692);
nor U46385 (N_46385,N_42859,N_42664);
nand U46386 (N_46386,N_41861,N_43638);
and U46387 (N_46387,N_44645,N_44975);
nand U46388 (N_46388,N_40947,N_42746);
or U46389 (N_46389,N_41141,N_43833);
nor U46390 (N_46390,N_44633,N_41061);
nor U46391 (N_46391,N_41792,N_44926);
xor U46392 (N_46392,N_44159,N_42916);
xor U46393 (N_46393,N_42035,N_44276);
nand U46394 (N_46394,N_42947,N_43174);
nor U46395 (N_46395,N_42326,N_44673);
and U46396 (N_46396,N_43693,N_42272);
nor U46397 (N_46397,N_44289,N_41880);
and U46398 (N_46398,N_41576,N_42255);
and U46399 (N_46399,N_41942,N_43582);
xnor U46400 (N_46400,N_42536,N_41934);
nand U46401 (N_46401,N_40269,N_40633);
nor U46402 (N_46402,N_40955,N_44514);
xnor U46403 (N_46403,N_43265,N_40632);
or U46404 (N_46404,N_43401,N_42807);
nand U46405 (N_46405,N_43873,N_43643);
xor U46406 (N_46406,N_41219,N_40518);
and U46407 (N_46407,N_40494,N_40864);
and U46408 (N_46408,N_42623,N_44319);
or U46409 (N_46409,N_44574,N_44728);
xnor U46410 (N_46410,N_40883,N_44126);
nor U46411 (N_46411,N_43241,N_43656);
xnor U46412 (N_46412,N_43918,N_44354);
xor U46413 (N_46413,N_43019,N_40893);
and U46414 (N_46414,N_44459,N_42944);
or U46415 (N_46415,N_44240,N_43803);
nand U46416 (N_46416,N_44228,N_40008);
or U46417 (N_46417,N_40630,N_40365);
nor U46418 (N_46418,N_44060,N_41593);
nor U46419 (N_46419,N_44511,N_44155);
xnor U46420 (N_46420,N_42400,N_41941);
xor U46421 (N_46421,N_42776,N_40603);
nor U46422 (N_46422,N_40491,N_41577);
and U46423 (N_46423,N_44092,N_41295);
nor U46424 (N_46424,N_40129,N_41453);
and U46425 (N_46425,N_42659,N_43575);
xor U46426 (N_46426,N_44344,N_41736);
xnor U46427 (N_46427,N_43111,N_43281);
nand U46428 (N_46428,N_41808,N_41683);
and U46429 (N_46429,N_42429,N_42550);
or U46430 (N_46430,N_42187,N_43299);
xor U46431 (N_46431,N_43084,N_42327);
nor U46432 (N_46432,N_42789,N_42598);
and U46433 (N_46433,N_44308,N_40336);
xnor U46434 (N_46434,N_40300,N_44552);
or U46435 (N_46435,N_40321,N_43403);
nor U46436 (N_46436,N_42338,N_42363);
xor U46437 (N_46437,N_41359,N_42083);
and U46438 (N_46438,N_44701,N_42253);
and U46439 (N_46439,N_40151,N_43369);
or U46440 (N_46440,N_40034,N_41877);
nor U46441 (N_46441,N_42464,N_42045);
nor U46442 (N_46442,N_40420,N_40298);
and U46443 (N_46443,N_40819,N_43276);
nand U46444 (N_46444,N_42057,N_40146);
or U46445 (N_46445,N_42951,N_44385);
nor U46446 (N_46446,N_40218,N_42033);
and U46447 (N_46447,N_42888,N_42260);
xnor U46448 (N_46448,N_43042,N_44487);
nor U46449 (N_46449,N_44848,N_42767);
xor U46450 (N_46450,N_40611,N_41074);
nand U46451 (N_46451,N_42600,N_41107);
xnor U46452 (N_46452,N_42617,N_42575);
nor U46453 (N_46453,N_41021,N_42467);
nand U46454 (N_46454,N_40529,N_41701);
or U46455 (N_46455,N_40789,N_42235);
nor U46456 (N_46456,N_40814,N_42682);
xor U46457 (N_46457,N_43443,N_41906);
xnor U46458 (N_46458,N_41081,N_43916);
and U46459 (N_46459,N_42198,N_44802);
nor U46460 (N_46460,N_40031,N_40937);
xnor U46461 (N_46461,N_41924,N_44340);
and U46462 (N_46462,N_43905,N_43358);
and U46463 (N_46463,N_42957,N_41043);
xnor U46464 (N_46464,N_40737,N_40397);
xnor U46465 (N_46465,N_42457,N_44935);
xnor U46466 (N_46466,N_42258,N_43597);
and U46467 (N_46467,N_44445,N_42438);
nand U46468 (N_46468,N_44185,N_42969);
xnor U46469 (N_46469,N_42739,N_43995);
xnor U46470 (N_46470,N_42504,N_41981);
nand U46471 (N_46471,N_40416,N_41421);
or U46472 (N_46472,N_41376,N_44674);
xor U46473 (N_46473,N_44019,N_40714);
nand U46474 (N_46474,N_43627,N_44998);
xnor U46475 (N_46475,N_43945,N_42238);
nand U46476 (N_46476,N_42718,N_43378);
and U46477 (N_46477,N_43052,N_43287);
and U46478 (N_46478,N_43450,N_44647);
nand U46479 (N_46479,N_42158,N_43368);
or U46480 (N_46480,N_42622,N_41567);
xor U46481 (N_46481,N_44910,N_43678);
or U46482 (N_46482,N_41815,N_43253);
xor U46483 (N_46483,N_40788,N_43183);
xor U46484 (N_46484,N_42670,N_41516);
or U46485 (N_46485,N_42116,N_41785);
xnor U46486 (N_46486,N_43634,N_42490);
or U46487 (N_46487,N_42248,N_43258);
or U46488 (N_46488,N_44735,N_42952);
and U46489 (N_46489,N_41603,N_42864);
or U46490 (N_46490,N_41518,N_43956);
and U46491 (N_46491,N_44212,N_44941);
nor U46492 (N_46492,N_40357,N_41740);
xor U46493 (N_46493,N_41824,N_40330);
nor U46494 (N_46494,N_42638,N_43465);
or U46495 (N_46495,N_43224,N_40587);
and U46496 (N_46496,N_40369,N_42182);
nor U46497 (N_46497,N_41146,N_41379);
and U46498 (N_46498,N_43187,N_43257);
nor U46499 (N_46499,N_40078,N_40339);
xor U46500 (N_46500,N_43532,N_44794);
nor U46501 (N_46501,N_40350,N_42653);
nor U46502 (N_46502,N_41108,N_43125);
nor U46503 (N_46503,N_44923,N_41406);
nor U46504 (N_46504,N_41671,N_42705);
or U46505 (N_46505,N_40995,N_42047);
and U46506 (N_46506,N_40343,N_42849);
nor U46507 (N_46507,N_44960,N_43493);
xor U46508 (N_46508,N_43731,N_43217);
nand U46509 (N_46509,N_44805,N_44581);
nand U46510 (N_46510,N_42213,N_41197);
and U46511 (N_46511,N_41487,N_42728);
and U46512 (N_46512,N_44601,N_44192);
nand U46513 (N_46513,N_44509,N_43789);
xor U46514 (N_46514,N_40678,N_43433);
nor U46515 (N_46515,N_40081,N_42044);
nand U46516 (N_46516,N_44538,N_41286);
nor U46517 (N_46517,N_42706,N_42800);
or U46518 (N_46518,N_42306,N_43055);
or U46519 (N_46519,N_44042,N_40825);
and U46520 (N_46520,N_40664,N_40448);
and U46521 (N_46521,N_44732,N_44299);
xnor U46522 (N_46522,N_40111,N_44179);
xor U46523 (N_46523,N_40857,N_40636);
nor U46524 (N_46524,N_42279,N_43765);
xnor U46525 (N_46525,N_42444,N_44419);
or U46526 (N_46526,N_41310,N_44951);
or U46527 (N_46527,N_41535,N_41455);
xor U46528 (N_46528,N_42842,N_40174);
or U46529 (N_46529,N_41222,N_40443);
xor U46530 (N_46530,N_41301,N_43675);
and U46531 (N_46531,N_42189,N_43824);
or U46532 (N_46532,N_42178,N_40821);
or U46533 (N_46533,N_40753,N_43103);
nor U46534 (N_46534,N_42388,N_41106);
nor U46535 (N_46535,N_44049,N_42419);
nor U46536 (N_46536,N_40943,N_44774);
nor U46537 (N_46537,N_43544,N_41588);
or U46538 (N_46538,N_40648,N_42093);
nand U46539 (N_46539,N_40512,N_42857);
xor U46540 (N_46540,N_42016,N_42672);
and U46541 (N_46541,N_43576,N_43629);
and U46542 (N_46542,N_41488,N_41478);
and U46543 (N_46543,N_41513,N_41260);
nand U46544 (N_46544,N_43562,N_41615);
nand U46545 (N_46545,N_40934,N_43079);
and U46546 (N_46546,N_43555,N_43251);
and U46547 (N_46547,N_40266,N_41992);
nor U46548 (N_46548,N_40118,N_41884);
and U46549 (N_46549,N_44243,N_43379);
nor U46550 (N_46550,N_41819,N_42146);
and U46551 (N_46551,N_40299,N_41790);
nand U46552 (N_46552,N_40831,N_41743);
xnor U46553 (N_46553,N_41269,N_43911);
xor U46554 (N_46554,N_42002,N_43110);
nand U46555 (N_46555,N_43799,N_41486);
nor U46556 (N_46556,N_44114,N_41032);
or U46557 (N_46557,N_44722,N_40870);
nor U46558 (N_46558,N_42148,N_42699);
and U46559 (N_46559,N_42287,N_43005);
xor U46560 (N_46560,N_41097,N_43756);
or U46561 (N_46561,N_43112,N_40449);
or U46562 (N_46562,N_40099,N_40569);
and U46563 (N_46563,N_41619,N_44369);
or U46564 (N_46564,N_43522,N_40599);
nand U46565 (N_46565,N_41953,N_43028);
nor U46566 (N_46566,N_42139,N_42342);
nor U46567 (N_46567,N_41788,N_44798);
and U46568 (N_46568,N_41691,N_44132);
or U46569 (N_46569,N_42698,N_40577);
nor U46570 (N_46570,N_40667,N_44372);
nand U46571 (N_46571,N_43654,N_40347);
xor U46572 (N_46572,N_42793,N_40283);
and U46573 (N_46573,N_42452,N_44213);
xnor U46574 (N_46574,N_43517,N_41080);
nor U46575 (N_46575,N_44591,N_43696);
and U46576 (N_46576,N_42786,N_44326);
xor U46577 (N_46577,N_43509,N_43762);
and U46578 (N_46578,N_44863,N_43609);
xnor U46579 (N_46579,N_44418,N_40358);
or U46580 (N_46580,N_43564,N_43193);
nor U46581 (N_46581,N_44607,N_44230);
nand U46582 (N_46582,N_44337,N_40457);
nor U46583 (N_46583,N_44726,N_41921);
or U46584 (N_46584,N_41559,N_41729);
or U46585 (N_46585,N_42011,N_41431);
and U46586 (N_46586,N_44288,N_44333);
nor U46587 (N_46587,N_44668,N_41470);
nand U46588 (N_46588,N_42994,N_44835);
or U46589 (N_46589,N_42958,N_44332);
or U46590 (N_46590,N_44966,N_40308);
nor U46591 (N_46591,N_44945,N_41805);
nand U46592 (N_46592,N_43698,N_40259);
nor U46593 (N_46593,N_41979,N_44054);
xnor U46594 (N_46594,N_41963,N_42828);
and U46595 (N_46595,N_44027,N_42069);
and U46596 (N_46596,N_41173,N_43946);
and U46597 (N_46597,N_41342,N_43054);
nor U46598 (N_46598,N_41160,N_40373);
xnor U46599 (N_46599,N_41935,N_41653);
xnor U46600 (N_46600,N_41723,N_44486);
or U46601 (N_46601,N_40869,N_44578);
xnor U46602 (N_46602,N_44031,N_41056);
nand U46603 (N_46603,N_42794,N_43375);
xor U46604 (N_46604,N_43962,N_44760);
nand U46605 (N_46605,N_41053,N_41363);
or U46606 (N_46606,N_42322,N_44981);
xor U46607 (N_46607,N_44356,N_42669);
or U46608 (N_46608,N_43087,N_43664);
nor U46609 (N_46609,N_40467,N_44749);
or U46610 (N_46610,N_43003,N_42202);
and U46611 (N_46611,N_44222,N_42474);
xnor U46612 (N_46612,N_43238,N_41037);
or U46613 (N_46613,N_43841,N_43423);
nand U46614 (N_46614,N_42475,N_43192);
nor U46615 (N_46615,N_44764,N_41016);
nor U46616 (N_46616,N_41144,N_41473);
xnor U46617 (N_46617,N_41505,N_44747);
xor U46618 (N_46618,N_43866,N_43455);
nand U46619 (N_46619,N_43134,N_40911);
and U46620 (N_46620,N_41418,N_43714);
xnor U46621 (N_46621,N_42377,N_43206);
or U46622 (N_46622,N_42641,N_44627);
xnor U46623 (N_46623,N_44290,N_44537);
and U46624 (N_46624,N_41644,N_41868);
xor U46625 (N_46625,N_41617,N_43809);
nor U46626 (N_46626,N_44037,N_44361);
xor U46627 (N_46627,N_41282,N_44714);
nor U46628 (N_46628,N_42403,N_44022);
nand U46629 (N_46629,N_40115,N_41902);
nor U46630 (N_46630,N_42637,N_40143);
xnor U46631 (N_46631,N_43489,N_41348);
nand U46632 (N_46632,N_43505,N_40059);
or U46633 (N_46633,N_41206,N_44837);
or U46634 (N_46634,N_43497,N_40684);
nor U46635 (N_46635,N_44345,N_42574);
xnor U46636 (N_46636,N_44182,N_44882);
nor U46637 (N_46637,N_41634,N_41480);
nand U46638 (N_46638,N_41125,N_43865);
nor U46639 (N_46639,N_43596,N_40515);
nor U46640 (N_46640,N_42426,N_44678);
or U46641 (N_46641,N_44162,N_41325);
xnor U46642 (N_46642,N_41822,N_41774);
and U46643 (N_46643,N_42825,N_44102);
nand U46644 (N_46644,N_41120,N_42245);
xnor U46645 (N_46645,N_42880,N_41563);
and U46646 (N_46646,N_42797,N_42449);
or U46647 (N_46647,N_44522,N_42360);
xor U46648 (N_46648,N_44255,N_43746);
xor U46649 (N_46649,N_44524,N_43768);
and U46650 (N_46650,N_40447,N_43361);
xnor U46651 (N_46651,N_42364,N_44247);
and U46652 (N_46652,N_41550,N_42815);
or U46653 (N_46653,N_42296,N_41063);
xnor U46654 (N_46654,N_43858,N_41354);
nor U46655 (N_46655,N_41737,N_41201);
or U46656 (N_46656,N_40348,N_42471);
or U46657 (N_46657,N_42592,N_43072);
nor U46658 (N_46658,N_40710,N_44183);
nand U46659 (N_46659,N_40333,N_40884);
nand U46660 (N_46660,N_40292,N_42024);
or U46661 (N_46661,N_44605,N_40915);
xor U46662 (N_46662,N_40691,N_44852);
nor U46663 (N_46663,N_44260,N_44030);
or U46664 (N_46664,N_42681,N_42257);
nor U46665 (N_46665,N_44613,N_41318);
or U46666 (N_46666,N_40747,N_43313);
or U46667 (N_46667,N_40162,N_43067);
or U46668 (N_46668,N_44430,N_40908);
nor U46669 (N_46669,N_41404,N_44181);
and U46670 (N_46670,N_41175,N_40776);
nand U46671 (N_46671,N_40912,N_42485);
nor U46672 (N_46672,N_44672,N_43018);
or U46673 (N_46673,N_42700,N_41189);
xnor U46674 (N_46674,N_41165,N_43337);
nand U46675 (N_46675,N_44883,N_41039);
or U46676 (N_46676,N_40329,N_41749);
or U46677 (N_46677,N_44957,N_43325);
xnor U46678 (N_46678,N_44214,N_40530);
xnor U46679 (N_46679,N_43135,N_44977);
and U46680 (N_46680,N_41757,N_42589);
xor U46681 (N_46681,N_44226,N_43954);
and U46682 (N_46682,N_43437,N_41997);
nor U46683 (N_46683,N_40891,N_44815);
xnor U46684 (N_46684,N_41496,N_42896);
xor U46685 (N_46685,N_40554,N_42179);
and U46686 (N_46686,N_41276,N_40964);
xor U46687 (N_46687,N_42155,N_43878);
nor U46688 (N_46688,N_41394,N_42274);
or U46689 (N_46689,N_44346,N_43482);
nand U46690 (N_46690,N_43051,N_40371);
xor U46691 (N_46691,N_42804,N_44703);
xnor U46692 (N_46692,N_41110,N_40312);
nor U46693 (N_46693,N_41714,N_41722);
or U46694 (N_46694,N_41303,N_40944);
xor U46695 (N_46695,N_42927,N_41169);
nand U46696 (N_46696,N_44686,N_44104);
xnor U46697 (N_46697,N_40588,N_42411);
nor U46698 (N_46698,N_44962,N_40589);
nand U46699 (N_46699,N_44988,N_41515);
and U46700 (N_46700,N_41542,N_43211);
nand U46701 (N_46701,N_41606,N_44549);
nor U46702 (N_46702,N_40552,N_42448);
nor U46703 (N_46703,N_42838,N_40780);
xor U46704 (N_46704,N_44062,N_44357);
nand U46705 (N_46705,N_42250,N_43207);
nand U46706 (N_46706,N_41652,N_43782);
or U46707 (N_46707,N_43385,N_43074);
and U46708 (N_46708,N_42803,N_41898);
nand U46709 (N_46709,N_44827,N_40608);
xnor U46710 (N_46710,N_44555,N_44495);
nand U46711 (N_46711,N_41907,N_42256);
nor U46712 (N_46712,N_41271,N_42242);
nor U46713 (N_46713,N_40534,N_43948);
and U46714 (N_46714,N_44176,N_42763);
nor U46715 (N_46715,N_44428,N_40198);
nand U46716 (N_46716,N_40878,N_42468);
nor U46717 (N_46717,N_44856,N_44716);
or U46718 (N_46718,N_42439,N_41309);
nand U46719 (N_46719,N_42201,N_40812);
nand U46720 (N_46720,N_43862,N_43769);
nand U46721 (N_46721,N_42846,N_42074);
nand U46722 (N_46722,N_43901,N_41073);
and U46723 (N_46723,N_40686,N_43442);
xor U46724 (N_46724,N_44849,N_43934);
and U46725 (N_46725,N_44853,N_41185);
xnor U46726 (N_46726,N_41202,N_44832);
nor U46727 (N_46727,N_41299,N_43963);
nor U46728 (N_46728,N_40698,N_40810);
and U46729 (N_46729,N_41850,N_44298);
nand U46730 (N_46730,N_42502,N_41253);
nand U46731 (N_46731,N_41305,N_41232);
or U46732 (N_46732,N_43332,N_40318);
nor U46733 (N_46733,N_43896,N_42456);
nand U46734 (N_46734,N_42597,N_43966);
or U46735 (N_46735,N_44052,N_40760);
nand U46736 (N_46736,N_41430,N_43915);
or U46737 (N_46737,N_42482,N_42817);
or U46738 (N_46738,N_41083,N_41791);
nand U46739 (N_46739,N_44283,N_42533);
or U46740 (N_46740,N_44108,N_44063);
nor U46741 (N_46741,N_42424,N_42003);
nand U46742 (N_46742,N_40367,N_43653);
nand U46743 (N_46743,N_41297,N_40877);
and U46744 (N_46744,N_44442,N_43845);
nand U46745 (N_46745,N_41986,N_42526);
and U46746 (N_46746,N_41367,N_42098);
nand U46747 (N_46747,N_41087,N_41751);
nand U46748 (N_46748,N_44938,N_43936);
xor U46749 (N_46749,N_44547,N_44371);
xnor U46750 (N_46750,N_44216,N_40619);
and U46751 (N_46751,N_41249,N_42627);
and U46752 (N_46752,N_44036,N_41523);
and U46753 (N_46753,N_41451,N_40210);
nor U46754 (N_46754,N_40600,N_42359);
nand U46755 (N_46755,N_40462,N_43524);
or U46756 (N_46756,N_40138,N_42072);
nor U46757 (N_46757,N_40056,N_44954);
and U46758 (N_46758,N_40661,N_41148);
and U46759 (N_46759,N_40163,N_40192);
xor U46760 (N_46760,N_40438,N_41828);
and U46761 (N_46761,N_43176,N_40389);
xnor U46762 (N_46762,N_40818,N_43721);
and U46763 (N_46763,N_42743,N_42117);
xor U46764 (N_46764,N_41323,N_43515);
xor U46765 (N_46765,N_44120,N_44269);
nor U46766 (N_46766,N_41716,N_44043);
nor U46767 (N_46767,N_43013,N_41466);
and U46768 (N_46768,N_44481,N_44889);
nand U46769 (N_46769,N_44005,N_40830);
xor U46770 (N_46770,N_40622,N_44828);
nor U46771 (N_46771,N_44404,N_43801);
nand U46772 (N_46772,N_41883,N_43541);
xnor U46773 (N_46773,N_43587,N_40425);
nor U46774 (N_46774,N_42735,N_40434);
or U46775 (N_46775,N_44644,N_40519);
nor U46776 (N_46776,N_40390,N_40489);
or U46777 (N_46777,N_40662,N_41193);
xor U46778 (N_46778,N_41698,N_40180);
nand U46779 (N_46779,N_41034,N_44661);
nand U46780 (N_46780,N_43940,N_41673);
and U46781 (N_46781,N_41782,N_43494);
nor U46782 (N_46782,N_44444,N_44259);
nand U46783 (N_46783,N_41988,N_42730);
and U46784 (N_46784,N_41777,N_44972);
xnor U46785 (N_46785,N_42990,N_43727);
or U46786 (N_46786,N_40424,N_42137);
nand U46787 (N_46787,N_40843,N_42931);
and U46788 (N_46788,N_41681,N_43610);
and U46789 (N_46789,N_42683,N_41872);
nand U46790 (N_46790,N_44850,N_41801);
xor U46791 (N_46791,N_41967,N_41928);
or U46792 (N_46792,N_44710,N_43312);
or U46793 (N_46793,N_40440,N_43406);
xor U46794 (N_46794,N_41272,N_40858);
nand U46795 (N_46795,N_40340,N_43558);
nor U46796 (N_46796,N_41155,N_42751);
or U46797 (N_46797,N_44089,N_42854);
or U46798 (N_46798,N_42224,N_44349);
or U46799 (N_46799,N_44928,N_42080);
nand U46800 (N_46800,N_41702,N_41769);
xor U46801 (N_46801,N_42037,N_43382);
nor U46802 (N_46802,N_43458,N_41047);
nand U46803 (N_46803,N_41688,N_41339);
xor U46804 (N_46804,N_42241,N_42760);
nand U46805 (N_46805,N_43850,N_42365);
or U46806 (N_46806,N_41502,N_43876);
nand U46807 (N_46807,N_42301,N_41987);
or U46808 (N_46808,N_43792,N_42565);
or U46809 (N_46809,N_42548,N_41068);
or U46810 (N_46810,N_42887,N_43106);
xnor U46811 (N_46811,N_44650,N_44164);
and U46812 (N_46812,N_43741,N_41800);
nand U46813 (N_46813,N_42876,N_41602);
and U46814 (N_46814,N_41036,N_44600);
nand U46815 (N_46815,N_43663,N_43511);
xnor U46816 (N_46816,N_44659,N_42433);
and U46817 (N_46817,N_41118,N_43983);
xnor U46818 (N_46818,N_42937,N_40590);
nand U46819 (N_46819,N_40826,N_43025);
xor U46820 (N_46820,N_43642,N_44116);
nand U46821 (N_46821,N_41663,N_42516);
xor U46822 (N_46822,N_42163,N_43614);
and U46823 (N_46823,N_42654,N_41665);
or U46824 (N_46824,N_40054,N_41018);
and U46825 (N_46825,N_40376,N_40949);
or U46826 (N_46826,N_44915,N_43829);
or U46827 (N_46827,N_40665,N_43362);
or U46828 (N_46828,N_42666,N_42566);
or U46829 (N_46829,N_41464,N_43985);
xnor U46830 (N_46830,N_43650,N_42556);
xnor U46831 (N_46831,N_43090,N_40003);
or U46832 (N_46832,N_42405,N_43040);
and U46833 (N_46833,N_42727,N_44990);
nor U46834 (N_46834,N_41927,N_42905);
nand U46835 (N_46835,N_43679,N_40969);
or U46836 (N_46836,N_43605,N_43124);
or U46837 (N_46837,N_42048,N_41391);
nor U46838 (N_46838,N_41199,N_44050);
and U46839 (N_46839,N_44194,N_40106);
nor U46840 (N_46840,N_40366,N_42764);
or U46841 (N_46841,N_41413,N_41324);
xnor U46842 (N_46842,N_43699,N_44653);
nand U46843 (N_46843,N_41066,N_43080);
or U46844 (N_46844,N_41190,N_42217);
or U46845 (N_46845,N_42031,N_40913);
or U46846 (N_46846,N_41719,N_42606);
xnor U46847 (N_46847,N_42928,N_41578);
xnor U46848 (N_46848,N_42765,N_41680);
nand U46849 (N_46849,N_42281,N_42725);
xnor U46850 (N_46850,N_44515,N_44807);
nand U46851 (N_46851,N_43571,N_44896);
nand U46852 (N_46852,N_44821,N_41891);
and U46853 (N_46853,N_41422,N_40876);
xor U46854 (N_46854,N_42568,N_42239);
and U46855 (N_46855,N_42695,N_43478);
or U46856 (N_46856,N_41662,N_40217);
xor U46857 (N_46857,N_42595,N_44003);
and U46858 (N_46858,N_41328,N_40951);
nand U46859 (N_46859,N_44593,N_44655);
or U46860 (N_46860,N_43949,N_42010);
nor U46861 (N_46861,N_42645,N_44457);
nand U46862 (N_46862,N_40873,N_41660);
or U46863 (N_46863,N_40221,N_42862);
nor U46864 (N_46864,N_41445,N_44779);
nor U46865 (N_46865,N_44588,N_40558);
or U46866 (N_46866,N_41235,N_43059);
xor U46867 (N_46867,N_40001,N_43421);
nor U46868 (N_46868,N_42461,N_40242);
or U46869 (N_46869,N_41656,N_42715);
nand U46870 (N_46870,N_44363,N_44629);
and U46871 (N_46871,N_40148,N_40658);
and U46872 (N_46872,N_42930,N_43250);
or U46873 (N_46873,N_40435,N_40026);
nor U46874 (N_46874,N_40246,N_40166);
xnor U46875 (N_46875,N_44757,N_43195);
nand U46876 (N_46876,N_43236,N_43661);
and U46877 (N_46877,N_40495,N_44087);
nand U46878 (N_46878,N_43863,N_43339);
nor U46879 (N_46879,N_40236,N_43889);
nor U46880 (N_46880,N_44024,N_41228);
xor U46881 (N_46881,N_40620,N_42750);
xor U46882 (N_46882,N_44618,N_40886);
or U46883 (N_46883,N_41708,N_44624);
and U46884 (N_46884,N_41251,N_41168);
nand U46885 (N_46885,N_44748,N_44178);
or U46886 (N_46886,N_44576,N_44411);
nor U46887 (N_46887,N_41669,N_40098);
nor U46888 (N_46888,N_44434,N_42262);
nor U46889 (N_46889,N_40394,N_43297);
and U46890 (N_46890,N_43248,N_41350);
and U46891 (N_46891,N_42860,N_43718);
xor U46892 (N_46892,N_40880,N_40979);
xor U46893 (N_46893,N_41245,N_42625);
nand U46894 (N_46894,N_41501,N_43618);
xor U46895 (N_46895,N_43190,N_44991);
nor U46896 (N_46896,N_44670,N_42628);
xor U46897 (N_46897,N_42823,N_42987);
nand U46898 (N_46898,N_44209,N_42431);
or U46899 (N_46899,N_42943,N_41793);
or U46900 (N_46900,N_43038,N_44408);
nor U46901 (N_46901,N_40540,N_41142);
and U46902 (N_46902,N_42335,N_40516);
and U46903 (N_46903,N_42251,N_42293);
and U46904 (N_46904,N_41546,N_44399);
and U46905 (N_46905,N_44175,N_42762);
nand U46906 (N_46906,N_43223,N_40575);
nand U46907 (N_46907,N_43073,N_44898);
xnor U46908 (N_46908,N_40579,N_41923);
nor U46909 (N_46909,N_44078,N_42836);
and U46910 (N_46910,N_44694,N_44431);
and U46911 (N_46911,N_44044,N_44309);
nand U46912 (N_46912,N_40036,N_40083);
xnor U46913 (N_46913,N_43996,N_40808);
xor U46914 (N_46914,N_41911,N_44596);
nor U46915 (N_46915,N_40413,N_42661);
and U46916 (N_46916,N_40423,N_44784);
or U46917 (N_46917,N_40904,N_40104);
xor U46918 (N_46918,N_43624,N_40715);
or U46919 (N_46919,N_44403,N_41908);
and U46920 (N_46920,N_44570,N_43200);
or U46921 (N_46921,N_42799,N_44697);
and U46922 (N_46922,N_41948,N_43722);
nor U46923 (N_46923,N_41374,N_42923);
xnor U46924 (N_46924,N_41438,N_42230);
nor U46925 (N_46925,N_43301,N_44820);
xor U46926 (N_46926,N_44277,N_42752);
nor U46927 (N_46927,N_42914,N_44364);
nor U46928 (N_46928,N_44281,N_42781);
nor U46929 (N_46929,N_44808,N_41157);
or U46930 (N_46930,N_42626,N_43506);
nor U46931 (N_46931,N_41858,N_43109);
and U46932 (N_46932,N_40378,N_42341);
and U46933 (N_46933,N_43508,N_40088);
nand U46934 (N_46934,N_43232,N_44266);
xnor U46935 (N_46935,N_41875,N_41529);
nand U46936 (N_46936,N_44316,N_44168);
or U46937 (N_46937,N_41750,N_43233);
nor U46938 (N_46938,N_43514,N_43290);
nor U46939 (N_46939,N_43467,N_44855);
nor U46940 (N_46940,N_42634,N_41744);
or U46941 (N_46941,N_43411,N_40639);
nand U46942 (N_46942,N_43893,N_40975);
nor U46943 (N_46943,N_44317,N_40548);
and U46944 (N_46944,N_40429,N_40145);
and U46945 (N_46945,N_41005,N_40410);
or U46946 (N_46946,N_43318,N_41840);
nor U46947 (N_46947,N_44234,N_44996);
nand U46948 (N_46948,N_40361,N_44041);
nor U46949 (N_46949,N_40592,N_40452);
nand U46950 (N_46950,N_43671,N_40673);
and U46951 (N_46951,N_40725,N_40713);
nor U46952 (N_46952,N_40204,N_42451);
xnor U46953 (N_46953,N_44400,N_41483);
xor U46954 (N_46954,N_40271,N_42415);
nand U46955 (N_46955,N_42603,N_44646);
and U46956 (N_46956,N_43776,N_40363);
and U46957 (N_46957,N_42624,N_44351);
and U46958 (N_46958,N_41491,N_40183);
nand U46959 (N_46959,N_42214,N_44478);
nand U46960 (N_46960,N_42347,N_40004);
or U46961 (N_46961,N_42369,N_42521);
nand U46962 (N_46962,N_41809,N_41287);
nand U46963 (N_46963,N_41990,N_40903);
nor U46964 (N_46964,N_43872,N_40305);
nor U46965 (N_46965,N_40983,N_41262);
and U46966 (N_46966,N_41642,N_41925);
or U46967 (N_46967,N_43672,N_42885);
nand U46968 (N_46968,N_44993,N_44518);
and U46969 (N_46969,N_41913,N_43881);
xor U46970 (N_46970,N_41475,N_43395);
nand U46971 (N_46971,N_40616,N_43720);
and U46972 (N_46972,N_43942,N_44498);
and U46973 (N_46973,N_41093,N_42863);
and U46974 (N_46974,N_44446,N_44254);
or U46975 (N_46975,N_43356,N_42275);
and U46976 (N_46976,N_43078,N_44084);
xnor U46977 (N_46977,N_42639,N_43392);
nor U46978 (N_46978,N_43425,N_42537);
xor U46979 (N_46979,N_42805,N_42974);
and U46980 (N_46980,N_40165,N_40197);
or U46981 (N_46981,N_41346,N_43711);
nand U46982 (N_46982,N_44389,N_40015);
and U46983 (N_46983,N_44415,N_43689);
nand U46984 (N_46984,N_42404,N_44338);
nand U46985 (N_46985,N_40501,N_43118);
nor U46986 (N_46986,N_40254,N_44920);
nand U46987 (N_46987,N_44783,N_44034);
nand U46988 (N_46988,N_40400,N_42050);
and U46989 (N_46989,N_44409,N_43286);
or U46990 (N_46990,N_44949,N_42950);
nor U46991 (N_46991,N_41154,N_40480);
or U46992 (N_46992,N_41772,N_43898);
and U46993 (N_46993,N_42596,N_43734);
nand U46994 (N_46994,N_43646,N_40294);
nor U46995 (N_46995,N_40683,N_43926);
or U46996 (N_46996,N_40136,N_41254);
nand U46997 (N_46997,N_42413,N_42724);
nor U46998 (N_46998,N_42312,N_42601);
nand U46999 (N_46999,N_43860,N_41362);
xnor U47000 (N_47000,N_41552,N_40186);
and U47001 (N_47001,N_40119,N_43729);
xor U47002 (N_47002,N_42145,N_42607);
xor U47003 (N_47003,N_40504,N_41172);
nand U47004 (N_47004,N_43424,N_41071);
and U47005 (N_47005,N_44976,N_41919);
xor U47006 (N_47006,N_41195,N_41746);
xnor U47007 (N_47007,N_43674,N_43122);
or U47008 (N_47008,N_42459,N_41441);
nand U47009 (N_47009,N_43892,N_42576);
and U47010 (N_47010,N_41151,N_43272);
xor U47011 (N_47011,N_40386,N_44761);
and U47012 (N_47012,N_40793,N_41306);
or U47013 (N_47013,N_43891,N_43129);
xor U47014 (N_47014,N_43178,N_42673);
xnor U47015 (N_47015,N_40950,N_41390);
nor U47016 (N_47016,N_40967,N_42110);
nand U47017 (N_47017,N_43976,N_43520);
xor U47018 (N_47018,N_41178,N_44682);
xnor U47019 (N_47019,N_44840,N_41194);
nand U47020 (N_47020,N_41916,N_44147);
and U47021 (N_47021,N_40094,N_44470);
and U47022 (N_47022,N_42674,N_42544);
xor U47023 (N_47023,N_40583,N_41974);
xnor U47024 (N_47024,N_44023,N_43056);
or U47025 (N_47025,N_43095,N_43062);
or U47026 (N_47026,N_40209,N_41114);
nor U47027 (N_47027,N_40690,N_42852);
xor U47028 (N_47028,N_42479,N_42208);
nor U47029 (N_47029,N_40730,N_43226);
nand U47030 (N_47030,N_41780,N_40860);
and U47031 (N_47031,N_42393,N_44499);
and U47032 (N_47032,N_40039,N_43323);
or U47033 (N_47033,N_42273,N_43529);
nand U47034 (N_47034,N_41879,N_44942);
nand U47035 (N_47035,N_41102,N_44595);
nor U47036 (N_47036,N_43139,N_41878);
nand U47037 (N_47037,N_43204,N_40079);
or U47038 (N_47038,N_43700,N_42921);
and U47039 (N_47039,N_41685,N_42733);
nand U47040 (N_47040,N_42979,N_44859);
xor U47041 (N_47041,N_40437,N_43218);
nor U47042 (N_47042,N_40635,N_41890);
and U47043 (N_47043,N_40442,N_43832);
or U47044 (N_47044,N_44841,N_44564);
nor U47045 (N_47045,N_43169,N_44425);
xor U47046 (N_47046,N_44692,N_42265);
nor U47047 (N_47047,N_41950,N_41227);
and U47048 (N_47048,N_44074,N_42992);
or U47049 (N_47049,N_42561,N_42740);
nand U47050 (N_47050,N_43014,N_44377);
and U47051 (N_47051,N_42418,N_42523);
xor U47052 (N_47052,N_42021,N_40956);
and U47053 (N_47053,N_44936,N_44485);
nand U47054 (N_47054,N_41958,N_42175);
xnor U47055 (N_47055,N_44328,N_40385);
and U47056 (N_47056,N_42678,N_41984);
or U47057 (N_47057,N_43032,N_40264);
and U47058 (N_47058,N_41752,N_43024);
xor U47059 (N_47059,N_41180,N_44868);
or U47060 (N_47060,N_44489,N_43376);
or U47061 (N_47061,N_43214,N_43586);
nand U47062 (N_47062,N_41837,N_43559);
nand U47063 (N_47063,N_44202,N_42758);
nor U47064 (N_47064,N_43227,N_43006);
and U47065 (N_47065,N_44546,N_43043);
or U47066 (N_47066,N_43341,N_43735);
or U47067 (N_47067,N_43262,N_43691);
nor U47068 (N_47068,N_42174,N_43812);
and U47069 (N_47069,N_42371,N_43117);
xnor U47070 (N_47070,N_41366,N_41745);
nor U47071 (N_47071,N_44220,N_40388);
or U47072 (N_47072,N_44583,N_42061);
or U47073 (N_47073,N_42064,N_40038);
nand U47074 (N_47074,N_42559,N_41213);
xor U47075 (N_47075,N_43652,N_41198);
nand U47076 (N_47076,N_42520,N_42046);
and U47077 (N_47077,N_44862,N_42547);
or U47078 (N_47078,N_41703,N_41484);
nand U47079 (N_47079,N_41547,N_40845);
and U47080 (N_47080,N_40833,N_42352);
and U47081 (N_47081,N_43787,N_40791);
or U47082 (N_47082,N_42869,N_41686);
or U47083 (N_47083,N_40892,N_41292);
or U47084 (N_47084,N_41764,N_41763);
nor U47085 (N_47085,N_42291,N_41273);
nand U47086 (N_47086,N_40360,N_44603);
or U47087 (N_47087,N_40472,N_40486);
nor U47088 (N_47088,N_43309,N_41724);
or U47089 (N_47089,N_42203,N_43635);
xor U47090 (N_47090,N_41138,N_42578);
or U47091 (N_47091,N_42483,N_44367);
xnor U47092 (N_47092,N_41873,N_40785);
xnor U47093 (N_47093,N_43708,N_41278);
or U47094 (N_47094,N_41813,N_43127);
nand U47095 (N_47095,N_42476,N_44777);
nand U47096 (N_47096,N_43254,N_41084);
nand U47097 (N_47097,N_40716,N_41582);
or U47098 (N_47098,N_43697,N_43757);
xor U47099 (N_47099,N_42330,N_44752);
or U47100 (N_47100,N_40316,N_42234);
nand U47101 (N_47101,N_44816,N_42938);
or U47102 (N_47102,N_41674,N_40802);
nand U47103 (N_47103,N_42967,N_44018);
or U47104 (N_47104,N_44980,N_44569);
or U47105 (N_47105,N_42563,N_42744);
and U47106 (N_47106,N_43585,N_40029);
nor U47107 (N_47107,N_44253,N_44302);
and U47108 (N_47108,N_41960,N_42971);
nor U47109 (N_47109,N_43311,N_42108);
or U47110 (N_47110,N_42087,N_41186);
and U47111 (N_47111,N_44249,N_40977);
nor U47112 (N_47112,N_41266,N_42871);
or U47113 (N_47113,N_44296,N_41062);
xor U47114 (N_47114,N_40013,N_40055);
and U47115 (N_47115,N_42071,N_43461);
and U47116 (N_47116,N_41753,N_40800);
and U47117 (N_47117,N_44124,N_42136);
or U47118 (N_47118,N_40404,N_43108);
nor U47119 (N_47119,N_42983,N_40920);
nand U47120 (N_47120,N_44375,N_44188);
or U47121 (N_47121,N_40954,N_41715);
and U47122 (N_47122,N_43732,N_43902);
nand U47123 (N_47123,N_40248,N_41562);
and U47124 (N_47124,N_42270,N_43977);
and U47125 (N_47125,N_43880,N_44939);
or U47126 (N_47126,N_43158,N_43320);
nor U47127 (N_47127,N_44039,N_41657);
nand U47128 (N_47128,N_41969,N_40010);
nand U47129 (N_47129,N_40591,N_43199);
nand U47130 (N_47130,N_44238,N_44767);
xnor U47131 (N_47131,N_42138,N_41874);
nand U47132 (N_47132,N_42926,N_44473);
nand U47133 (N_47133,N_44683,N_42792);
and U47134 (N_47134,N_43261,N_40922);
and U47135 (N_47135,N_43563,N_42337);
or U47136 (N_47136,N_43381,N_44223);
or U47137 (N_47137,N_44480,N_41843);
and U47138 (N_47138,N_41300,N_40827);
and U47139 (N_47139,N_42316,N_44458);
and U47140 (N_47140,N_40743,N_40513);
xnor U47141 (N_47141,N_40803,N_41905);
nand U47142 (N_47142,N_44781,N_41281);
and U47143 (N_47143,N_43625,N_41017);
and U47144 (N_47144,N_40002,N_40411);
nor U47145 (N_47145,N_41915,N_44270);
and U47146 (N_47146,N_42308,N_41045);
nor U47147 (N_47147,N_43744,N_40086);
and U47148 (N_47148,N_40514,N_42605);
nor U47149 (N_47149,N_40463,N_40307);
xor U47150 (N_47150,N_43154,N_40974);
and U47151 (N_47151,N_42963,N_41900);
or U47152 (N_47152,N_40465,N_41414);
nor U47153 (N_47153,N_44969,N_42294);
and U47154 (N_47154,N_40047,N_43668);
nand U47155 (N_47155,N_43778,N_44861);
nor U47156 (N_47156,N_44447,N_40539);
or U47157 (N_47157,N_43816,N_42713);
or U47158 (N_47158,N_40918,N_40595);
nand U47159 (N_47159,N_44151,N_43772);
or U47160 (N_47160,N_40324,N_41758);
or U47161 (N_47161,N_43736,N_44252);
nor U47162 (N_47162,N_40607,N_44394);
or U47163 (N_47163,N_41420,N_42655);
and U47164 (N_47164,N_42909,N_42620);
xnor U47165 (N_47165,N_41072,N_40605);
nand U47166 (N_47166,N_43592,N_43398);
xnor U47167 (N_47167,N_40193,N_43987);
xnor U47168 (N_47168,N_40032,N_43877);
nand U47169 (N_47169,N_41279,N_43180);
nor U47170 (N_47170,N_42078,N_41940);
and U47171 (N_47171,N_43680,N_43114);
or U47172 (N_47172,N_42839,N_41823);
nand U47173 (N_47173,N_42081,N_43798);
or U47174 (N_47174,N_41929,N_40739);
xnor U47175 (N_47175,N_40310,N_42833);
and U47176 (N_47176,N_44751,N_44436);
nor U47177 (N_47177,N_41373,N_40991);
xor U47178 (N_47178,N_42428,N_41124);
or U47179 (N_47179,N_40546,N_43355);
xor U47180 (N_47180,N_40405,N_40952);
xnor U47181 (N_47181,N_42737,N_44278);
nand U47182 (N_47182,N_44476,N_41864);
nor U47183 (N_47183,N_43929,N_44099);
xnor U47184 (N_47184,N_40304,N_44465);
and U47185 (N_47185,N_41949,N_42754);
xor U47186 (N_47186,N_42491,N_43371);
xor U47187 (N_47187,N_40542,N_43994);
nor U47188 (N_47188,N_42477,N_41100);
nand U47189 (N_47189,N_40973,N_41797);
nor U47190 (N_47190,N_42577,N_43922);
nand U47191 (N_47191,N_42694,N_44463);
xor U47192 (N_47192,N_41521,N_44526);
nor U47193 (N_47193,N_44971,N_43104);
or U47194 (N_47194,N_42086,N_43546);
or U47195 (N_47195,N_40135,N_42140);
xor U47196 (N_47196,N_42668,N_43420);
nand U47197 (N_47197,N_40492,N_41568);
or U47198 (N_47198,N_44873,N_41524);
xnor U47199 (N_47199,N_43584,N_42494);
nand U47200 (N_47200,N_43637,N_41225);
nand U47201 (N_47201,N_43047,N_42759);
and U47202 (N_47202,N_44615,N_43107);
xor U47203 (N_47203,N_43695,N_42813);
nand U47204 (N_47204,N_43484,N_43535);
or U47205 (N_47205,N_43932,N_40422);
or U47206 (N_47206,N_40674,N_40344);
and U47207 (N_47207,N_44467,N_40087);
or U47208 (N_47208,N_44221,N_43412);
and U47209 (N_47209,N_43890,N_40019);
xor U47210 (N_47210,N_40194,N_44468);
or U47211 (N_47211,N_44217,N_40496);
nor U47212 (N_47212,N_44553,N_44587);
and U47213 (N_47213,N_44677,N_41553);
xnor U47214 (N_47214,N_44927,N_40735);
xnor U47215 (N_47215,N_40770,N_43793);
nand U47216 (N_47216,N_42225,N_41096);
or U47217 (N_47217,N_43147,N_44651);
xnor U47218 (N_47218,N_44983,N_40910);
xnor U47219 (N_47219,N_44010,N_41651);
nand U47220 (N_47220,N_42390,N_44184);
and U47221 (N_47221,N_41055,N_42648);
or U47222 (N_47222,N_43405,N_43796);
or U47223 (N_47223,N_43485,N_40815);
xnor U47224 (N_47224,N_40765,N_42555);
nand U47225 (N_47225,N_40988,N_44955);
xor U47226 (N_47226,N_43389,N_40527);
and U47227 (N_47227,N_41465,N_44142);
or U47228 (N_47228,N_43230,N_40790);
and U47229 (N_47229,N_44721,N_44888);
nor U47230 (N_47230,N_43820,N_41347);
and U47231 (N_47231,N_42008,N_43247);
nor U47232 (N_47232,N_41101,N_43849);
nor U47233 (N_47233,N_43815,N_41735);
nor U47234 (N_47234,N_44982,N_42378);
or U47235 (N_47235,N_44414,N_43595);
nor U47236 (N_47236,N_40507,N_42901);
nand U47237 (N_47237,N_41829,N_41123);
xor U47238 (N_47238,N_41134,N_40775);
nand U47239 (N_47239,N_42455,N_43462);
nor U47240 (N_47240,N_44065,N_41538);
or U47241 (N_47241,N_40096,N_42223);
or U47242 (N_47242,N_40113,N_41557);
nand U47243 (N_47243,N_43023,N_41449);
and U47244 (N_47244,N_42723,N_42861);
and U47245 (N_47245,N_40459,N_43968);
nand U47246 (N_47246,N_44639,N_40160);
or U47247 (N_47247,N_41007,N_43784);
or U47248 (N_47248,N_43453,N_43446);
or U47249 (N_47249,N_41695,N_41098);
and U47250 (N_47250,N_40498,N_40981);
and U47251 (N_47251,N_40382,N_40565);
nand U47252 (N_47252,N_40334,N_41993);
or U47253 (N_47253,N_41954,N_44199);
xor U47254 (N_47254,N_43083,N_42644);
nor U47255 (N_47255,N_40907,N_44201);
or U47256 (N_47256,N_41442,N_43621);
and U47257 (N_47257,N_43715,N_42053);
and U47258 (N_47258,N_44358,N_41067);
nor U47259 (N_47259,N_42519,N_44279);
nand U47260 (N_47260,N_43492,N_44836);
and U47261 (N_47261,N_40223,N_42127);
nand U47262 (N_47262,N_44438,N_42704);
nand U47263 (N_47263,N_42988,N_44699);
xor U47264 (N_47264,N_43748,N_40353);
nand U47265 (N_47265,N_44362,N_41586);
nand U47266 (N_47266,N_41261,N_41482);
xor U47267 (N_47267,N_43967,N_44268);
nand U47268 (N_47268,N_40890,N_44893);
nor U47269 (N_47269,N_43528,N_41259);
and U47270 (N_47270,N_43115,N_44795);
or U47271 (N_47271,N_43527,N_42810);
nand U47272 (N_47272,N_41495,N_43438);
nand U47273 (N_47273,N_42757,N_42924);
xnor U47274 (N_47274,N_44324,N_43094);
nor U47275 (N_47275,N_43308,N_40837);
or U47276 (N_47276,N_41968,N_42908);
nand U47277 (N_47277,N_40722,N_41541);
xnor U47278 (N_47278,N_41859,N_40669);
and U47279 (N_47279,N_43220,N_42063);
or U47280 (N_47280,N_40229,N_44702);
nand U47281 (N_47281,N_41153,N_44948);
nor U47282 (N_47282,N_44989,N_44096);
xor U47283 (N_47283,N_44079,N_44331);
and U47284 (N_47284,N_42361,N_42965);
xor U47285 (N_47285,N_43328,N_44715);
and U47286 (N_47286,N_41810,N_42541);
nor U47287 (N_47287,N_43020,N_42680);
nand U47288 (N_47288,N_40476,N_43933);
or U47289 (N_47289,N_44123,N_44206);
or U47290 (N_47290,N_43282,N_43048);
nor U47291 (N_47291,N_41591,N_40177);
nand U47292 (N_47292,N_42510,N_40740);
nand U47293 (N_47293,N_44788,N_41939);
or U47294 (N_47294,N_41832,N_44575);
nor U47295 (N_47295,N_42020,N_42447);
or U47296 (N_47296,N_44021,N_42973);
nand U47297 (N_47297,N_44401,N_43660);
nor U47298 (N_47298,N_41000,N_44177);
nor U47299 (N_47299,N_40375,N_41549);
nor U47300 (N_47300,N_42391,N_40069);
xnor U47301 (N_47301,N_42252,N_44082);
nand U47302 (N_47302,N_41575,N_41332);
nand U47303 (N_47303,N_42874,N_40384);
or U47304 (N_47304,N_41973,N_43143);
xnor U47305 (N_47305,N_42040,N_42367);
xnor U47306 (N_47306,N_44635,N_40855);
or U47307 (N_47307,N_44262,N_41592);
nand U47308 (N_47308,N_44973,N_44086);
xnor U47309 (N_47309,N_43641,N_42205);
and U47310 (N_47310,N_43537,N_42058);
xor U47311 (N_47311,N_41600,N_43166);
and U47312 (N_47312,N_42989,N_44730);
xor U47313 (N_47313,N_43578,N_40602);
and U47314 (N_47314,N_41392,N_41853);
nand U47315 (N_47315,N_40184,N_41020);
nand U47316 (N_47316,N_40849,N_44286);
nand U47317 (N_47317,N_40201,N_42478);
nand U47318 (N_47318,N_40042,N_42769);
nand U47319 (N_47319,N_42954,N_44709);
nand U47320 (N_47320,N_43296,N_42708);
or U47321 (N_47321,N_42084,N_44384);
nor U47322 (N_47322,N_44076,N_40559);
and U47323 (N_47323,N_42837,N_43194);
nor U47324 (N_47324,N_43430,N_40646);
or U47325 (N_47325,N_43542,N_44026);
nand U47326 (N_47326,N_42934,N_43440);
nor U47327 (N_47327,N_43857,N_44374);
or U47328 (N_47328,N_42065,N_41341);
nand U47329 (N_47329,N_43342,N_42689);
xnor U47330 (N_47330,N_44750,N_40729);
xnor U47331 (N_47331,N_41945,N_41145);
and U47332 (N_47332,N_42199,N_43991);
nor U47333 (N_47333,N_43483,N_43189);
nor U47334 (N_47334,N_41388,N_43069);
or U47335 (N_47335,N_41621,N_43436);
nand U47336 (N_47336,N_40650,N_44125);
nor U47337 (N_47337,N_41980,N_44312);
xnor U47338 (N_47338,N_41147,N_43101);
nor U47339 (N_47339,N_41551,N_43049);
xor U47340 (N_47340,N_44736,N_44842);
xor U47341 (N_47341,N_42414,N_44285);
nor U47342 (N_47342,N_44806,N_43473);
nand U47343 (N_47343,N_43758,N_40268);
and U47344 (N_47344,N_40175,N_41833);
nor U47345 (N_47345,N_40097,N_40842);
xnor U47346 (N_47346,N_42194,N_40164);
or U47347 (N_47347,N_41493,N_44878);
and U47348 (N_47348,N_44440,N_43925);
or U47349 (N_47349,N_41440,N_42321);
xor U47350 (N_47350,N_42919,N_40037);
nand U47351 (N_47351,N_41024,N_40178);
and U47352 (N_47352,N_43480,N_44420);
nor U47353 (N_47353,N_41664,N_41892);
nand U47354 (N_47354,N_41732,N_43157);
nor U47355 (N_47355,N_40147,N_43408);
and U47356 (N_47356,N_44839,N_40822);
nor U47357 (N_47357,N_41267,N_44264);
nor U47358 (N_47358,N_43685,N_43035);
and U47359 (N_47359,N_43036,N_44834);
or U47360 (N_47360,N_40252,N_41277);
xor U47361 (N_47361,N_44857,N_43435);
or U47362 (N_47362,N_43970,N_43249);
xor U47363 (N_47363,N_41506,N_44348);
xnor U47364 (N_47364,N_41739,N_44329);
xor U47365 (N_47365,N_42572,N_40654);
nand U47366 (N_47366,N_40906,N_44814);
nor U47367 (N_47367,N_40301,N_40756);
or U47368 (N_47368,N_42132,N_43728);
xnor U47369 (N_47369,N_43222,N_44387);
nand U47370 (N_47370,N_43600,N_41761);
nor U47371 (N_47371,N_42941,N_43819);
and U47372 (N_47372,N_40919,N_41459);
or U47373 (N_47373,N_43648,N_42505);
xnor U47374 (N_47374,N_41672,N_44909);
nand U47375 (N_47375,N_44510,N_42000);
nor U47376 (N_47376,N_42320,N_40176);
and U47377 (N_47377,N_43667,N_41316);
nand U47378 (N_47378,N_41349,N_43766);
nand U47379 (N_47379,N_44045,N_44758);
nor U47380 (N_47380,N_40121,N_40000);
xnor U47381 (N_47381,N_44933,N_40909);
nor U47382 (N_47382,N_40707,N_40617);
nor U47383 (N_47383,N_41510,N_43088);
nor U47384 (N_47384,N_40966,N_42998);
nand U47385 (N_47385,N_43304,N_42663);
and U47386 (N_47386,N_42524,N_43153);
or U47387 (N_47387,N_40233,N_43510);
nor U47388 (N_47388,N_42551,N_43594);
and U47389 (N_47389,N_44944,N_43939);
nand U47390 (N_47390,N_44804,N_44719);
and U47391 (N_47391,N_41710,N_40075);
and U47392 (N_47392,N_42569,N_42611);
nor U47393 (N_47393,N_42007,N_40116);
nor U47394 (N_47394,N_41372,N_40182);
or U47395 (N_47395,N_40718,N_43372);
nand U47396 (N_47396,N_41111,N_41655);
nand U47397 (N_47397,N_40586,N_41335);
nor U47398 (N_47398,N_44196,N_43046);
nor U47399 (N_47399,N_42621,N_44218);
nand U47400 (N_47400,N_44090,N_40179);
nand U47401 (N_47401,N_41353,N_43202);
or U47402 (N_47402,N_40727,N_44543);
xnor U47403 (N_47403,N_43231,N_41103);
or U47404 (N_47404,N_43413,N_43851);
or U47405 (N_47405,N_42309,N_44917);
and U47406 (N_47406,N_44314,N_44628);
and U47407 (N_47407,N_43717,N_40326);
and U47408 (N_47408,N_44477,N_43534);
and U47409 (N_47409,N_42311,N_42900);
nor U47410 (N_47410,N_41386,N_42851);
nand U47411 (N_47411,N_40757,N_41914);
and U47412 (N_47412,N_40521,N_44244);
or U47413 (N_47413,N_40380,N_40395);
xnor U47414 (N_47414,N_43298,N_40963);
xor U47415 (N_47415,N_40528,N_44676);
nor U47416 (N_47416,N_41288,N_42870);
nor U47417 (N_47417,N_42772,N_44707);
xnor U47418 (N_47418,N_41424,N_43149);
and U47419 (N_47419,N_43895,N_40976);
nor U47420 (N_47420,N_43333,N_41336);
xnor U47421 (N_47421,N_41240,N_40110);
and U47422 (N_47422,N_40215,N_42023);
xnor U47423 (N_47423,N_41345,N_42501);
nand U47424 (N_47424,N_42716,N_40568);
nor U47425 (N_47425,N_43737,N_43810);
nor U47426 (N_47426,N_44924,N_42514);
and U47427 (N_47427,N_40468,N_43764);
xor U47428 (N_47428,N_41846,N_44275);
xor U47429 (N_47429,N_44038,N_44632);
and U47430 (N_47430,N_40933,N_42177);
xnor U47431 (N_47431,N_44294,N_43965);
or U47432 (N_47432,N_40033,N_44706);
xor U47433 (N_47433,N_41835,N_40717);
nor U47434 (N_47434,N_43414,N_43531);
nand U47435 (N_47435,N_44274,N_41918);
and U47436 (N_47436,N_43607,N_42755);
nor U47437 (N_47437,N_44642,N_41435);
xor U47438 (N_47438,N_44033,N_41895);
and U47439 (N_47439,N_40430,N_42325);
or U47440 (N_47440,N_42333,N_44571);
and U47441 (N_47441,N_41867,N_43747);
nor U47442 (N_47442,N_41640,N_44964);
and U47443 (N_47443,N_42357,N_42650);
nand U47444 (N_47444,N_41952,N_42392);
xnor U47445 (N_47445,N_40993,N_41787);
and U47446 (N_47446,N_40524,N_44556);
or U47447 (N_47447,N_42985,N_42300);
or U47448 (N_47448,N_40297,N_42707);
and U47449 (N_47449,N_42130,N_41569);
and U47450 (N_47450,N_43086,N_40535);
and U47451 (N_47451,N_41807,N_44500);
or U47452 (N_47452,N_41989,N_44610);
and U47453 (N_47453,N_41135,N_40139);
or U47454 (N_47454,N_44662,N_42629);
or U47455 (N_47455,N_42289,N_40829);
xnor U47456 (N_47456,N_42018,N_41766);
nand U47457 (N_47457,N_44456,N_40279);
xor U47458 (N_47458,N_40896,N_44450);
nor U47459 (N_47459,N_41268,N_42099);
nand U47460 (N_47460,N_44488,N_41771);
nor U47461 (N_47461,N_44608,N_44826);
nor U47462 (N_47462,N_41876,N_41014);
and U47463 (N_47463,N_43777,N_40811);
or U47464 (N_47464,N_42649,N_40660);
or U47465 (N_47465,N_40216,N_40606);
nand U47466 (N_47466,N_40127,N_43518);
xnor U47467 (N_47467,N_42865,N_43383);
nor U47468 (N_47468,N_44193,N_42809);
or U47469 (N_47469,N_41033,N_40253);
xnor U47470 (N_47470,N_40990,N_42903);
nor U47471 (N_47471,N_41331,N_44643);
or U47472 (N_47472,N_44739,N_44829);
and U47473 (N_47473,N_41612,N_43418);
or U47474 (N_47474,N_44512,N_40766);
nor U47475 (N_47475,N_43774,N_43507);
and U47476 (N_47476,N_42237,N_44918);
xnor U47477 (N_47477,N_40863,N_42506);
nor U47478 (N_47478,N_44423,N_40374);
nand U47479 (N_47479,N_40352,N_42726);
nand U47480 (N_47480,N_44753,N_41856);
and U47481 (N_47481,N_44007,N_41467);
nand U47482 (N_47482,N_40924,N_44681);
and U47483 (N_47483,N_40341,N_43469);
nand U47484 (N_47484,N_42619,N_42819);
xnor U47485 (N_47485,N_40313,N_43303);
nor U47486 (N_47486,N_42115,N_41322);
xnor U47487 (N_47487,N_40256,N_40703);
and U47488 (N_47488,N_41584,N_44474);
or U47489 (N_47489,N_41320,N_43706);
nor U47490 (N_47490,N_42609,N_44649);
or U47491 (N_47491,N_43603,N_40866);
nand U47492 (N_47492,N_43707,N_40049);
nor U47493 (N_47493,N_43703,N_40398);
nand U47494 (N_47494,N_43556,N_41403);
nor U47495 (N_47495,N_44388,N_41159);
nand U47496 (N_47496,N_41049,N_41713);
and U47497 (N_47497,N_43951,N_40278);
nand U47498 (N_47498,N_43781,N_44413);
and U47499 (N_47499,N_40932,N_41212);
nand U47500 (N_47500,N_40792,N_42016);
nand U47501 (N_47501,N_44756,N_40776);
nand U47502 (N_47502,N_41485,N_43045);
and U47503 (N_47503,N_44586,N_43141);
nor U47504 (N_47504,N_41194,N_43134);
or U47505 (N_47505,N_40623,N_41266);
or U47506 (N_47506,N_43969,N_42255);
or U47507 (N_47507,N_41104,N_40715);
nand U47508 (N_47508,N_40010,N_41964);
nand U47509 (N_47509,N_43662,N_44014);
nand U47510 (N_47510,N_43261,N_44847);
or U47511 (N_47511,N_44841,N_44017);
nor U47512 (N_47512,N_42435,N_43097);
nand U47513 (N_47513,N_41521,N_43409);
xnor U47514 (N_47514,N_40409,N_40576);
xnor U47515 (N_47515,N_42184,N_40888);
nand U47516 (N_47516,N_43202,N_44611);
and U47517 (N_47517,N_44860,N_42039);
nand U47518 (N_47518,N_43953,N_42993);
xor U47519 (N_47519,N_43129,N_40903);
nor U47520 (N_47520,N_41338,N_43163);
nor U47521 (N_47521,N_40458,N_41313);
nor U47522 (N_47522,N_44283,N_44609);
and U47523 (N_47523,N_41159,N_44360);
nor U47524 (N_47524,N_43036,N_43864);
nand U47525 (N_47525,N_42808,N_41389);
nor U47526 (N_47526,N_44442,N_42025);
or U47527 (N_47527,N_41234,N_43390);
nor U47528 (N_47528,N_42062,N_42672);
nor U47529 (N_47529,N_40213,N_41440);
nand U47530 (N_47530,N_40345,N_42479);
nor U47531 (N_47531,N_41237,N_41366);
or U47532 (N_47532,N_44273,N_43900);
xor U47533 (N_47533,N_42002,N_44502);
xor U47534 (N_47534,N_40686,N_41546);
nor U47535 (N_47535,N_41793,N_42495);
nor U47536 (N_47536,N_44535,N_42501);
nor U47537 (N_47537,N_43434,N_43833);
or U47538 (N_47538,N_41247,N_40839);
and U47539 (N_47539,N_44471,N_43644);
nand U47540 (N_47540,N_42810,N_41238);
and U47541 (N_47541,N_43034,N_43811);
nand U47542 (N_47542,N_43831,N_44166);
and U47543 (N_47543,N_42801,N_40185);
or U47544 (N_47544,N_40857,N_41397);
and U47545 (N_47545,N_40753,N_44806);
xnor U47546 (N_47546,N_41158,N_44639);
xor U47547 (N_47547,N_42891,N_42712);
or U47548 (N_47548,N_44039,N_42100);
nand U47549 (N_47549,N_40574,N_43482);
or U47550 (N_47550,N_41597,N_42639);
nand U47551 (N_47551,N_40675,N_41697);
xor U47552 (N_47552,N_43883,N_42278);
and U47553 (N_47553,N_40194,N_44765);
nor U47554 (N_47554,N_41501,N_42600);
xnor U47555 (N_47555,N_41188,N_44209);
nand U47556 (N_47556,N_42776,N_41064);
xnor U47557 (N_47557,N_42893,N_42901);
or U47558 (N_47558,N_44463,N_44274);
xnor U47559 (N_47559,N_43655,N_43310);
xnor U47560 (N_47560,N_41254,N_42465);
and U47561 (N_47561,N_40870,N_44234);
xnor U47562 (N_47562,N_42897,N_40806);
nor U47563 (N_47563,N_43626,N_41255);
or U47564 (N_47564,N_42181,N_44075);
and U47565 (N_47565,N_41738,N_42870);
nand U47566 (N_47566,N_40467,N_42078);
nand U47567 (N_47567,N_40548,N_41535);
xor U47568 (N_47568,N_43882,N_40462);
xnor U47569 (N_47569,N_41235,N_43372);
nand U47570 (N_47570,N_42487,N_44318);
xor U47571 (N_47571,N_41344,N_40270);
xnor U47572 (N_47572,N_40094,N_42235);
xnor U47573 (N_47573,N_43564,N_44657);
nor U47574 (N_47574,N_41142,N_44494);
nand U47575 (N_47575,N_42228,N_41789);
nor U47576 (N_47576,N_44082,N_44642);
nand U47577 (N_47577,N_42222,N_44651);
nand U47578 (N_47578,N_42958,N_41257);
nand U47579 (N_47579,N_42345,N_43150);
or U47580 (N_47580,N_40832,N_42884);
nor U47581 (N_47581,N_40612,N_41680);
or U47582 (N_47582,N_43469,N_44579);
or U47583 (N_47583,N_44141,N_42949);
or U47584 (N_47584,N_42392,N_42379);
xnor U47585 (N_47585,N_41521,N_43757);
and U47586 (N_47586,N_40281,N_42280);
nand U47587 (N_47587,N_42706,N_43972);
or U47588 (N_47588,N_44810,N_41205);
xor U47589 (N_47589,N_41794,N_44908);
and U47590 (N_47590,N_41671,N_40868);
nor U47591 (N_47591,N_44570,N_41341);
nor U47592 (N_47592,N_42549,N_41712);
nor U47593 (N_47593,N_41166,N_42207);
nor U47594 (N_47594,N_41905,N_44600);
and U47595 (N_47595,N_41968,N_42558);
nand U47596 (N_47596,N_40426,N_40017);
nor U47597 (N_47597,N_41506,N_40116);
and U47598 (N_47598,N_42465,N_42316);
or U47599 (N_47599,N_42620,N_42630);
and U47600 (N_47600,N_42906,N_40446);
or U47601 (N_47601,N_40224,N_40698);
nor U47602 (N_47602,N_43667,N_40277);
nor U47603 (N_47603,N_41282,N_43793);
xnor U47604 (N_47604,N_41105,N_44000);
or U47605 (N_47605,N_41485,N_41864);
and U47606 (N_47606,N_40819,N_40131);
nor U47607 (N_47607,N_43442,N_43294);
nor U47608 (N_47608,N_43806,N_44865);
nor U47609 (N_47609,N_43061,N_44952);
or U47610 (N_47610,N_44316,N_43611);
and U47611 (N_47611,N_41230,N_42845);
or U47612 (N_47612,N_43461,N_41441);
nand U47613 (N_47613,N_43370,N_40715);
nand U47614 (N_47614,N_42630,N_40192);
nand U47615 (N_47615,N_43021,N_43940);
xor U47616 (N_47616,N_40727,N_42579);
or U47617 (N_47617,N_43706,N_40113);
nand U47618 (N_47618,N_40685,N_40459);
or U47619 (N_47619,N_44346,N_42285);
nor U47620 (N_47620,N_41261,N_40484);
nand U47621 (N_47621,N_43207,N_42929);
or U47622 (N_47622,N_44195,N_41727);
xor U47623 (N_47623,N_44148,N_43919);
xnor U47624 (N_47624,N_40190,N_44559);
nand U47625 (N_47625,N_40984,N_42508);
or U47626 (N_47626,N_41581,N_43032);
nand U47627 (N_47627,N_43549,N_40292);
nand U47628 (N_47628,N_41240,N_40743);
nor U47629 (N_47629,N_43035,N_41854);
or U47630 (N_47630,N_42562,N_44095);
xor U47631 (N_47631,N_40467,N_40234);
and U47632 (N_47632,N_41020,N_44709);
and U47633 (N_47633,N_43329,N_41980);
and U47634 (N_47634,N_43969,N_40005);
nor U47635 (N_47635,N_40930,N_44022);
and U47636 (N_47636,N_42882,N_43137);
xor U47637 (N_47637,N_40427,N_43922);
xnor U47638 (N_47638,N_40589,N_44723);
nor U47639 (N_47639,N_42803,N_43018);
nand U47640 (N_47640,N_41181,N_42361);
or U47641 (N_47641,N_42327,N_43893);
xnor U47642 (N_47642,N_43041,N_44362);
and U47643 (N_47643,N_44747,N_42656);
and U47644 (N_47644,N_42470,N_42484);
nand U47645 (N_47645,N_44883,N_40551);
nand U47646 (N_47646,N_44570,N_44648);
or U47647 (N_47647,N_44819,N_40383);
or U47648 (N_47648,N_41766,N_43576);
or U47649 (N_47649,N_43986,N_40032);
and U47650 (N_47650,N_41772,N_41344);
nand U47651 (N_47651,N_42859,N_43717);
and U47652 (N_47652,N_40198,N_40997);
xnor U47653 (N_47653,N_41622,N_40605);
or U47654 (N_47654,N_40284,N_40683);
and U47655 (N_47655,N_42254,N_41845);
nand U47656 (N_47656,N_43210,N_42912);
or U47657 (N_47657,N_44881,N_41927);
xnor U47658 (N_47658,N_41872,N_42451);
nand U47659 (N_47659,N_43990,N_41190);
and U47660 (N_47660,N_40156,N_43425);
xor U47661 (N_47661,N_43196,N_42003);
nor U47662 (N_47662,N_41559,N_41496);
nor U47663 (N_47663,N_43211,N_44450);
or U47664 (N_47664,N_40141,N_42738);
xor U47665 (N_47665,N_44288,N_43138);
or U47666 (N_47666,N_44321,N_44871);
and U47667 (N_47667,N_41660,N_44276);
xnor U47668 (N_47668,N_43328,N_43019);
and U47669 (N_47669,N_41353,N_42390);
xnor U47670 (N_47670,N_40910,N_41578);
nor U47671 (N_47671,N_44621,N_44121);
or U47672 (N_47672,N_43941,N_40836);
xnor U47673 (N_47673,N_44417,N_42675);
xor U47674 (N_47674,N_41128,N_40956);
xnor U47675 (N_47675,N_42328,N_40812);
or U47676 (N_47676,N_44089,N_40615);
and U47677 (N_47677,N_40487,N_44465);
and U47678 (N_47678,N_44852,N_43944);
or U47679 (N_47679,N_44783,N_44154);
nand U47680 (N_47680,N_44153,N_40493);
xor U47681 (N_47681,N_42918,N_43187);
nor U47682 (N_47682,N_40042,N_41798);
and U47683 (N_47683,N_40689,N_40063);
xor U47684 (N_47684,N_43126,N_41748);
nand U47685 (N_47685,N_41439,N_42825);
nand U47686 (N_47686,N_42442,N_42511);
nand U47687 (N_47687,N_40378,N_43395);
xnor U47688 (N_47688,N_44235,N_42999);
or U47689 (N_47689,N_42655,N_40987);
or U47690 (N_47690,N_42112,N_41052);
xor U47691 (N_47691,N_41495,N_43317);
and U47692 (N_47692,N_42829,N_40216);
and U47693 (N_47693,N_42545,N_41154);
xor U47694 (N_47694,N_43628,N_43255);
or U47695 (N_47695,N_43364,N_43565);
xnor U47696 (N_47696,N_43579,N_44743);
xnor U47697 (N_47697,N_40628,N_40173);
nor U47698 (N_47698,N_41782,N_41535);
or U47699 (N_47699,N_44392,N_41042);
and U47700 (N_47700,N_44688,N_41623);
nor U47701 (N_47701,N_43393,N_40026);
nand U47702 (N_47702,N_44180,N_41668);
and U47703 (N_47703,N_44933,N_44591);
xor U47704 (N_47704,N_40065,N_44513);
or U47705 (N_47705,N_40151,N_41186);
and U47706 (N_47706,N_42809,N_44256);
and U47707 (N_47707,N_41476,N_42784);
nand U47708 (N_47708,N_41584,N_42691);
nor U47709 (N_47709,N_44393,N_41416);
or U47710 (N_47710,N_44888,N_43062);
and U47711 (N_47711,N_40689,N_40122);
xnor U47712 (N_47712,N_41257,N_44733);
and U47713 (N_47713,N_43292,N_40196);
nand U47714 (N_47714,N_44353,N_44454);
or U47715 (N_47715,N_42207,N_44924);
or U47716 (N_47716,N_43164,N_41488);
and U47717 (N_47717,N_41747,N_44396);
nand U47718 (N_47718,N_42957,N_44658);
xor U47719 (N_47719,N_44054,N_40338);
or U47720 (N_47720,N_40794,N_42631);
nor U47721 (N_47721,N_40849,N_41461);
nand U47722 (N_47722,N_42374,N_44919);
nor U47723 (N_47723,N_43201,N_42025);
xnor U47724 (N_47724,N_44868,N_41505);
and U47725 (N_47725,N_40549,N_41022);
nand U47726 (N_47726,N_41366,N_42579);
xor U47727 (N_47727,N_41685,N_43333);
xnor U47728 (N_47728,N_40167,N_41850);
and U47729 (N_47729,N_40141,N_42861);
nand U47730 (N_47730,N_40404,N_43492);
nor U47731 (N_47731,N_42970,N_42838);
or U47732 (N_47732,N_40781,N_42800);
nor U47733 (N_47733,N_42639,N_40620);
and U47734 (N_47734,N_44253,N_44577);
xnor U47735 (N_47735,N_43885,N_40147);
nand U47736 (N_47736,N_44562,N_44918);
xor U47737 (N_47737,N_41123,N_41365);
nand U47738 (N_47738,N_44637,N_42659);
or U47739 (N_47739,N_41711,N_42129);
xnor U47740 (N_47740,N_40083,N_43573);
and U47741 (N_47741,N_40244,N_44673);
or U47742 (N_47742,N_40719,N_41337);
or U47743 (N_47743,N_42630,N_42643);
and U47744 (N_47744,N_41232,N_42782);
or U47745 (N_47745,N_42781,N_43636);
xor U47746 (N_47746,N_40795,N_41336);
or U47747 (N_47747,N_40058,N_41402);
or U47748 (N_47748,N_44801,N_43334);
and U47749 (N_47749,N_43360,N_44376);
nor U47750 (N_47750,N_42113,N_43828);
and U47751 (N_47751,N_42997,N_42996);
or U47752 (N_47752,N_41188,N_44548);
xnor U47753 (N_47753,N_41807,N_42718);
nand U47754 (N_47754,N_44454,N_41182);
xnor U47755 (N_47755,N_44090,N_40198);
and U47756 (N_47756,N_42996,N_40565);
nor U47757 (N_47757,N_44168,N_44851);
and U47758 (N_47758,N_43200,N_42570);
nand U47759 (N_47759,N_41310,N_44147);
and U47760 (N_47760,N_44463,N_44215);
or U47761 (N_47761,N_41576,N_43018);
or U47762 (N_47762,N_41766,N_42289);
xor U47763 (N_47763,N_41738,N_40702);
or U47764 (N_47764,N_40373,N_42726);
nor U47765 (N_47765,N_40964,N_42863);
nor U47766 (N_47766,N_40874,N_41698);
nand U47767 (N_47767,N_40434,N_44626);
and U47768 (N_47768,N_44422,N_44420);
or U47769 (N_47769,N_40926,N_41042);
nand U47770 (N_47770,N_44508,N_40967);
or U47771 (N_47771,N_41976,N_43377);
or U47772 (N_47772,N_40111,N_43345);
nand U47773 (N_47773,N_43268,N_40610);
xnor U47774 (N_47774,N_40287,N_42637);
nor U47775 (N_47775,N_42165,N_44924);
xor U47776 (N_47776,N_40345,N_41899);
nand U47777 (N_47777,N_41773,N_42950);
xor U47778 (N_47778,N_44710,N_41150);
or U47779 (N_47779,N_44587,N_42085);
and U47780 (N_47780,N_41116,N_43541);
and U47781 (N_47781,N_40523,N_44725);
nand U47782 (N_47782,N_40230,N_44051);
or U47783 (N_47783,N_43921,N_42158);
xor U47784 (N_47784,N_44086,N_41538);
and U47785 (N_47785,N_44516,N_43440);
nor U47786 (N_47786,N_41296,N_42341);
nor U47787 (N_47787,N_43212,N_43982);
nor U47788 (N_47788,N_40317,N_40635);
or U47789 (N_47789,N_44296,N_42890);
xor U47790 (N_47790,N_40437,N_43022);
and U47791 (N_47791,N_41478,N_41219);
nand U47792 (N_47792,N_43562,N_41393);
and U47793 (N_47793,N_44835,N_42506);
or U47794 (N_47794,N_42057,N_42500);
nor U47795 (N_47795,N_43566,N_41412);
nor U47796 (N_47796,N_41107,N_41562);
and U47797 (N_47797,N_41930,N_43310);
nor U47798 (N_47798,N_41750,N_44739);
or U47799 (N_47799,N_42065,N_41462);
xor U47800 (N_47800,N_44292,N_41203);
nor U47801 (N_47801,N_42073,N_44426);
xor U47802 (N_47802,N_42619,N_44697);
or U47803 (N_47803,N_44620,N_42542);
xor U47804 (N_47804,N_40032,N_40257);
nand U47805 (N_47805,N_41466,N_40853);
and U47806 (N_47806,N_44629,N_42334);
nand U47807 (N_47807,N_40229,N_41588);
nor U47808 (N_47808,N_44050,N_44891);
nor U47809 (N_47809,N_42793,N_42799);
xnor U47810 (N_47810,N_41688,N_44206);
nor U47811 (N_47811,N_43912,N_40689);
and U47812 (N_47812,N_42245,N_44004);
nand U47813 (N_47813,N_44944,N_41040);
nor U47814 (N_47814,N_42758,N_42173);
or U47815 (N_47815,N_44332,N_44726);
nor U47816 (N_47816,N_44535,N_44550);
nor U47817 (N_47817,N_43961,N_40169);
or U47818 (N_47818,N_42307,N_41002);
or U47819 (N_47819,N_44488,N_41810);
nor U47820 (N_47820,N_42106,N_41111);
and U47821 (N_47821,N_40256,N_40852);
and U47822 (N_47822,N_42803,N_43879);
and U47823 (N_47823,N_40065,N_42247);
nand U47824 (N_47824,N_43053,N_41732);
and U47825 (N_47825,N_41133,N_42728);
nor U47826 (N_47826,N_40288,N_44194);
nor U47827 (N_47827,N_41460,N_40351);
xnor U47828 (N_47828,N_42319,N_40557);
nor U47829 (N_47829,N_41284,N_41023);
nor U47830 (N_47830,N_42367,N_40077);
xnor U47831 (N_47831,N_40074,N_43145);
nand U47832 (N_47832,N_43415,N_40797);
or U47833 (N_47833,N_41022,N_41502);
nor U47834 (N_47834,N_44591,N_41311);
nor U47835 (N_47835,N_43277,N_42268);
xnor U47836 (N_47836,N_40664,N_40434);
nor U47837 (N_47837,N_43108,N_43488);
nand U47838 (N_47838,N_43425,N_44848);
or U47839 (N_47839,N_42084,N_43562);
nor U47840 (N_47840,N_41503,N_44729);
nand U47841 (N_47841,N_43490,N_42912);
or U47842 (N_47842,N_44643,N_42659);
nor U47843 (N_47843,N_40878,N_40213);
nor U47844 (N_47844,N_43654,N_40355);
and U47845 (N_47845,N_42006,N_43334);
nor U47846 (N_47846,N_44257,N_44550);
and U47847 (N_47847,N_40945,N_40764);
and U47848 (N_47848,N_40293,N_40568);
xnor U47849 (N_47849,N_44109,N_41693);
nand U47850 (N_47850,N_44386,N_42367);
or U47851 (N_47851,N_40162,N_42913);
xor U47852 (N_47852,N_44485,N_40540);
xnor U47853 (N_47853,N_43588,N_43002);
and U47854 (N_47854,N_40771,N_42486);
and U47855 (N_47855,N_40159,N_44089);
nand U47856 (N_47856,N_44486,N_40878);
nor U47857 (N_47857,N_42246,N_40586);
and U47858 (N_47858,N_44814,N_43362);
xnor U47859 (N_47859,N_44373,N_40504);
or U47860 (N_47860,N_41908,N_44014);
nor U47861 (N_47861,N_42048,N_43091);
or U47862 (N_47862,N_43955,N_43933);
and U47863 (N_47863,N_44719,N_43632);
and U47864 (N_47864,N_40702,N_40012);
xnor U47865 (N_47865,N_40348,N_42310);
nor U47866 (N_47866,N_40080,N_42425);
xor U47867 (N_47867,N_40656,N_42400);
or U47868 (N_47868,N_40487,N_40745);
or U47869 (N_47869,N_44587,N_40475);
nor U47870 (N_47870,N_44514,N_41143);
xnor U47871 (N_47871,N_43355,N_44083);
nand U47872 (N_47872,N_40269,N_40433);
and U47873 (N_47873,N_44565,N_44185);
nand U47874 (N_47874,N_43397,N_41392);
or U47875 (N_47875,N_44797,N_41481);
or U47876 (N_47876,N_43837,N_43140);
or U47877 (N_47877,N_43628,N_43873);
nand U47878 (N_47878,N_42088,N_41150);
and U47879 (N_47879,N_41327,N_43328);
nor U47880 (N_47880,N_42890,N_42850);
nand U47881 (N_47881,N_43110,N_44807);
nand U47882 (N_47882,N_44205,N_44342);
or U47883 (N_47883,N_40802,N_40436);
nand U47884 (N_47884,N_43943,N_44682);
xnor U47885 (N_47885,N_43043,N_40952);
nor U47886 (N_47886,N_43845,N_42249);
or U47887 (N_47887,N_41911,N_42801);
and U47888 (N_47888,N_40021,N_40309);
xor U47889 (N_47889,N_41397,N_42999);
nand U47890 (N_47890,N_41670,N_41936);
nand U47891 (N_47891,N_44500,N_42196);
or U47892 (N_47892,N_42531,N_41155);
nor U47893 (N_47893,N_44976,N_42585);
xor U47894 (N_47894,N_41756,N_40727);
nor U47895 (N_47895,N_41388,N_42298);
nand U47896 (N_47896,N_40884,N_43406);
nor U47897 (N_47897,N_41812,N_42791);
nand U47898 (N_47898,N_41198,N_44513);
or U47899 (N_47899,N_44596,N_40393);
xor U47900 (N_47900,N_43414,N_42109);
or U47901 (N_47901,N_41614,N_40759);
nor U47902 (N_47902,N_43807,N_41211);
and U47903 (N_47903,N_41233,N_43310);
or U47904 (N_47904,N_41354,N_41904);
xor U47905 (N_47905,N_44585,N_43212);
xor U47906 (N_47906,N_44352,N_43085);
nand U47907 (N_47907,N_42513,N_44433);
and U47908 (N_47908,N_40132,N_41676);
nand U47909 (N_47909,N_41762,N_40433);
and U47910 (N_47910,N_40978,N_41964);
nor U47911 (N_47911,N_40180,N_44308);
nor U47912 (N_47912,N_40342,N_41097);
and U47913 (N_47913,N_41750,N_44709);
or U47914 (N_47914,N_44369,N_42282);
or U47915 (N_47915,N_41595,N_43969);
xnor U47916 (N_47916,N_40875,N_44638);
or U47917 (N_47917,N_42021,N_42870);
nand U47918 (N_47918,N_42928,N_41706);
nand U47919 (N_47919,N_40699,N_40298);
xor U47920 (N_47920,N_40258,N_44182);
nor U47921 (N_47921,N_43252,N_42597);
xor U47922 (N_47922,N_41253,N_43438);
nand U47923 (N_47923,N_40904,N_40609);
nor U47924 (N_47924,N_40511,N_42717);
xor U47925 (N_47925,N_40670,N_43059);
or U47926 (N_47926,N_41873,N_42902);
nand U47927 (N_47927,N_44230,N_42080);
or U47928 (N_47928,N_40996,N_44071);
and U47929 (N_47929,N_44784,N_40126);
and U47930 (N_47930,N_41013,N_44197);
or U47931 (N_47931,N_41895,N_42007);
nand U47932 (N_47932,N_40508,N_42252);
and U47933 (N_47933,N_44621,N_42704);
xnor U47934 (N_47934,N_40552,N_44905);
xnor U47935 (N_47935,N_44432,N_44848);
nand U47936 (N_47936,N_41839,N_40541);
and U47937 (N_47937,N_42804,N_40327);
nor U47938 (N_47938,N_41679,N_41292);
or U47939 (N_47939,N_43724,N_44197);
nor U47940 (N_47940,N_40335,N_40375);
nor U47941 (N_47941,N_43912,N_43739);
xnor U47942 (N_47942,N_44337,N_42007);
or U47943 (N_47943,N_42982,N_40007);
nor U47944 (N_47944,N_40607,N_44105);
nand U47945 (N_47945,N_44546,N_42813);
and U47946 (N_47946,N_40937,N_42331);
nor U47947 (N_47947,N_41934,N_43712);
xnor U47948 (N_47948,N_43217,N_40843);
and U47949 (N_47949,N_43927,N_44136);
or U47950 (N_47950,N_42769,N_42906);
nor U47951 (N_47951,N_41183,N_42930);
and U47952 (N_47952,N_43822,N_44156);
xnor U47953 (N_47953,N_41033,N_40839);
xor U47954 (N_47954,N_44182,N_40025);
xnor U47955 (N_47955,N_44790,N_42285);
nand U47956 (N_47956,N_40110,N_43158);
or U47957 (N_47957,N_41678,N_42545);
or U47958 (N_47958,N_42883,N_42017);
and U47959 (N_47959,N_41291,N_43176);
or U47960 (N_47960,N_44411,N_43656);
nand U47961 (N_47961,N_44499,N_40501);
nand U47962 (N_47962,N_41119,N_40893);
xnor U47963 (N_47963,N_44316,N_40210);
or U47964 (N_47964,N_44951,N_42863);
xnor U47965 (N_47965,N_42343,N_42992);
nand U47966 (N_47966,N_44820,N_41227);
xor U47967 (N_47967,N_43700,N_44131);
xor U47968 (N_47968,N_43655,N_42755);
xnor U47969 (N_47969,N_41155,N_44849);
xor U47970 (N_47970,N_44241,N_42576);
or U47971 (N_47971,N_41227,N_44275);
nand U47972 (N_47972,N_40255,N_41003);
nand U47973 (N_47973,N_44534,N_40503);
or U47974 (N_47974,N_43321,N_44232);
nor U47975 (N_47975,N_43648,N_44298);
nor U47976 (N_47976,N_41947,N_40403);
nand U47977 (N_47977,N_44793,N_42868);
nor U47978 (N_47978,N_44229,N_41673);
or U47979 (N_47979,N_40385,N_43872);
xor U47980 (N_47980,N_40703,N_44536);
or U47981 (N_47981,N_43147,N_42289);
nor U47982 (N_47982,N_42015,N_40907);
xnor U47983 (N_47983,N_40234,N_41711);
or U47984 (N_47984,N_43054,N_40382);
or U47985 (N_47985,N_43122,N_41468);
nor U47986 (N_47986,N_43957,N_41951);
xnor U47987 (N_47987,N_43217,N_42854);
xor U47988 (N_47988,N_44378,N_41392);
or U47989 (N_47989,N_42099,N_44603);
nand U47990 (N_47990,N_42773,N_42558);
or U47991 (N_47991,N_44346,N_44273);
or U47992 (N_47992,N_44270,N_44147);
xnor U47993 (N_47993,N_41690,N_42297);
and U47994 (N_47994,N_40325,N_44140);
xor U47995 (N_47995,N_40183,N_43145);
nor U47996 (N_47996,N_41568,N_44439);
nor U47997 (N_47997,N_44083,N_40984);
nand U47998 (N_47998,N_44036,N_43631);
or U47999 (N_47999,N_40164,N_44913);
xnor U48000 (N_48000,N_44375,N_42354);
or U48001 (N_48001,N_40990,N_42527);
xnor U48002 (N_48002,N_43873,N_43650);
xor U48003 (N_48003,N_42565,N_44399);
or U48004 (N_48004,N_40197,N_42686);
and U48005 (N_48005,N_43444,N_40778);
xnor U48006 (N_48006,N_43932,N_41346);
nand U48007 (N_48007,N_42167,N_44405);
xnor U48008 (N_48008,N_40434,N_41527);
or U48009 (N_48009,N_42544,N_42666);
xor U48010 (N_48010,N_43633,N_44402);
and U48011 (N_48011,N_41456,N_41325);
nor U48012 (N_48012,N_42098,N_42853);
and U48013 (N_48013,N_42339,N_43681);
xor U48014 (N_48014,N_42621,N_44791);
xnor U48015 (N_48015,N_41731,N_43847);
and U48016 (N_48016,N_40514,N_41273);
xnor U48017 (N_48017,N_44306,N_42819);
nand U48018 (N_48018,N_44295,N_44515);
nand U48019 (N_48019,N_41540,N_40807);
nand U48020 (N_48020,N_41773,N_44664);
nand U48021 (N_48021,N_41417,N_44782);
and U48022 (N_48022,N_41792,N_42810);
nor U48023 (N_48023,N_43901,N_43099);
nand U48024 (N_48024,N_43984,N_43287);
xnor U48025 (N_48025,N_44327,N_44567);
nor U48026 (N_48026,N_43918,N_41601);
or U48027 (N_48027,N_44883,N_44389);
xor U48028 (N_48028,N_43933,N_44601);
nor U48029 (N_48029,N_41591,N_40204);
or U48030 (N_48030,N_42255,N_42397);
or U48031 (N_48031,N_44161,N_40936);
nand U48032 (N_48032,N_42938,N_40878);
and U48033 (N_48033,N_40641,N_41705);
nor U48034 (N_48034,N_41078,N_40227);
or U48035 (N_48035,N_42895,N_44381);
xor U48036 (N_48036,N_41249,N_41027);
nor U48037 (N_48037,N_41640,N_43328);
nand U48038 (N_48038,N_40569,N_41128);
and U48039 (N_48039,N_42048,N_42139);
xnor U48040 (N_48040,N_40215,N_40686);
nor U48041 (N_48041,N_42148,N_41758);
xnor U48042 (N_48042,N_40870,N_44840);
nor U48043 (N_48043,N_43999,N_42409);
xnor U48044 (N_48044,N_40490,N_42494);
xnor U48045 (N_48045,N_41009,N_41501);
nand U48046 (N_48046,N_42754,N_40059);
nand U48047 (N_48047,N_43048,N_41258);
nand U48048 (N_48048,N_44865,N_40942);
nand U48049 (N_48049,N_41654,N_44356);
nor U48050 (N_48050,N_42339,N_44428);
or U48051 (N_48051,N_43801,N_44698);
nand U48052 (N_48052,N_42346,N_44662);
xor U48053 (N_48053,N_41235,N_41299);
or U48054 (N_48054,N_44793,N_41771);
or U48055 (N_48055,N_43162,N_42503);
nor U48056 (N_48056,N_41483,N_42540);
nand U48057 (N_48057,N_42726,N_44142);
nand U48058 (N_48058,N_44962,N_42647);
and U48059 (N_48059,N_41852,N_43997);
nand U48060 (N_48060,N_44908,N_43074);
nor U48061 (N_48061,N_40085,N_41059);
nand U48062 (N_48062,N_42215,N_44998);
nand U48063 (N_48063,N_40230,N_43620);
nor U48064 (N_48064,N_43636,N_41838);
nor U48065 (N_48065,N_44362,N_44015);
nor U48066 (N_48066,N_41776,N_43915);
nor U48067 (N_48067,N_40086,N_41057);
nor U48068 (N_48068,N_40962,N_44480);
nor U48069 (N_48069,N_42181,N_40581);
nand U48070 (N_48070,N_42735,N_43751);
or U48071 (N_48071,N_43704,N_41585);
nor U48072 (N_48072,N_44746,N_40044);
and U48073 (N_48073,N_41937,N_44869);
xnor U48074 (N_48074,N_42361,N_42329);
and U48075 (N_48075,N_43239,N_40438);
or U48076 (N_48076,N_40069,N_43614);
or U48077 (N_48077,N_43864,N_41033);
and U48078 (N_48078,N_41322,N_40259);
and U48079 (N_48079,N_43308,N_40099);
nand U48080 (N_48080,N_43132,N_42380);
xnor U48081 (N_48081,N_44532,N_42374);
nor U48082 (N_48082,N_42348,N_40125);
or U48083 (N_48083,N_40860,N_43113);
xor U48084 (N_48084,N_40018,N_40976);
xor U48085 (N_48085,N_42497,N_41245);
or U48086 (N_48086,N_43319,N_41166);
or U48087 (N_48087,N_40740,N_43362);
xnor U48088 (N_48088,N_41470,N_40216);
nor U48089 (N_48089,N_42719,N_44889);
and U48090 (N_48090,N_42014,N_43212);
or U48091 (N_48091,N_40452,N_44279);
and U48092 (N_48092,N_41537,N_41062);
xnor U48093 (N_48093,N_43006,N_42404);
or U48094 (N_48094,N_41624,N_40947);
xor U48095 (N_48095,N_43833,N_41924);
nand U48096 (N_48096,N_41880,N_43004);
xor U48097 (N_48097,N_42882,N_44484);
nor U48098 (N_48098,N_42760,N_43795);
xor U48099 (N_48099,N_41054,N_44108);
nand U48100 (N_48100,N_43679,N_43891);
nand U48101 (N_48101,N_42336,N_40742);
nand U48102 (N_48102,N_41798,N_43478);
nor U48103 (N_48103,N_41465,N_43175);
or U48104 (N_48104,N_42680,N_41092);
or U48105 (N_48105,N_43876,N_44827);
nand U48106 (N_48106,N_42789,N_40545);
nand U48107 (N_48107,N_40791,N_42602);
or U48108 (N_48108,N_40293,N_42200);
or U48109 (N_48109,N_44921,N_40873);
or U48110 (N_48110,N_43129,N_41547);
nand U48111 (N_48111,N_44824,N_43269);
nor U48112 (N_48112,N_41940,N_43404);
xnor U48113 (N_48113,N_40443,N_42119);
and U48114 (N_48114,N_43826,N_44884);
nor U48115 (N_48115,N_41994,N_43022);
or U48116 (N_48116,N_44093,N_41019);
and U48117 (N_48117,N_44750,N_40318);
nor U48118 (N_48118,N_40959,N_44018);
xor U48119 (N_48119,N_41595,N_42406);
and U48120 (N_48120,N_43136,N_43042);
or U48121 (N_48121,N_40605,N_43988);
xnor U48122 (N_48122,N_43098,N_41843);
or U48123 (N_48123,N_40327,N_42186);
xnor U48124 (N_48124,N_42210,N_40146);
xor U48125 (N_48125,N_43538,N_44287);
or U48126 (N_48126,N_42413,N_40449);
and U48127 (N_48127,N_42646,N_40061);
or U48128 (N_48128,N_44716,N_42493);
nand U48129 (N_48129,N_41168,N_40259);
or U48130 (N_48130,N_40877,N_44459);
or U48131 (N_48131,N_42998,N_42817);
nor U48132 (N_48132,N_42392,N_42344);
nand U48133 (N_48133,N_41280,N_43106);
nand U48134 (N_48134,N_44734,N_41227);
nand U48135 (N_48135,N_44837,N_43867);
nand U48136 (N_48136,N_41196,N_40585);
nand U48137 (N_48137,N_44078,N_44693);
nor U48138 (N_48138,N_42343,N_41183);
or U48139 (N_48139,N_43034,N_42132);
nor U48140 (N_48140,N_41917,N_40494);
nand U48141 (N_48141,N_42949,N_43872);
nor U48142 (N_48142,N_44478,N_40261);
nor U48143 (N_48143,N_41470,N_43148);
xor U48144 (N_48144,N_42289,N_44746);
nor U48145 (N_48145,N_40419,N_43785);
nor U48146 (N_48146,N_42701,N_43198);
or U48147 (N_48147,N_42703,N_44008);
or U48148 (N_48148,N_41167,N_43737);
and U48149 (N_48149,N_42401,N_43517);
or U48150 (N_48150,N_42788,N_41663);
nand U48151 (N_48151,N_43029,N_42712);
nor U48152 (N_48152,N_43897,N_44782);
or U48153 (N_48153,N_43391,N_40772);
and U48154 (N_48154,N_44082,N_44482);
xor U48155 (N_48155,N_43463,N_42863);
xor U48156 (N_48156,N_42446,N_40883);
and U48157 (N_48157,N_44161,N_41250);
and U48158 (N_48158,N_43996,N_43200);
nor U48159 (N_48159,N_44623,N_41646);
nand U48160 (N_48160,N_42670,N_40194);
or U48161 (N_48161,N_40149,N_40295);
and U48162 (N_48162,N_41061,N_40360);
or U48163 (N_48163,N_41092,N_40288);
and U48164 (N_48164,N_40122,N_40804);
nor U48165 (N_48165,N_40307,N_44581);
xor U48166 (N_48166,N_43856,N_44435);
and U48167 (N_48167,N_44854,N_40320);
and U48168 (N_48168,N_41504,N_44615);
or U48169 (N_48169,N_41300,N_44966);
nor U48170 (N_48170,N_40458,N_44805);
or U48171 (N_48171,N_40133,N_43094);
xor U48172 (N_48172,N_40818,N_41443);
xnor U48173 (N_48173,N_40338,N_41305);
or U48174 (N_48174,N_43291,N_43657);
or U48175 (N_48175,N_40651,N_41986);
nand U48176 (N_48176,N_43757,N_41803);
or U48177 (N_48177,N_40242,N_43896);
or U48178 (N_48178,N_44757,N_43741);
or U48179 (N_48179,N_44120,N_41575);
xor U48180 (N_48180,N_43342,N_40692);
and U48181 (N_48181,N_42166,N_40305);
xnor U48182 (N_48182,N_40411,N_41255);
and U48183 (N_48183,N_40274,N_40314);
and U48184 (N_48184,N_43941,N_40366);
or U48185 (N_48185,N_44095,N_44417);
nand U48186 (N_48186,N_40322,N_43975);
and U48187 (N_48187,N_42756,N_43091);
and U48188 (N_48188,N_42833,N_40896);
nand U48189 (N_48189,N_44824,N_41944);
xnor U48190 (N_48190,N_40337,N_42003);
xor U48191 (N_48191,N_41053,N_43078);
xnor U48192 (N_48192,N_42662,N_43210);
nor U48193 (N_48193,N_43483,N_41693);
nand U48194 (N_48194,N_43170,N_42605);
or U48195 (N_48195,N_40398,N_42582);
or U48196 (N_48196,N_42011,N_44667);
nand U48197 (N_48197,N_43199,N_41758);
nand U48198 (N_48198,N_44510,N_41871);
nand U48199 (N_48199,N_41289,N_43884);
and U48200 (N_48200,N_41594,N_41744);
and U48201 (N_48201,N_43396,N_41058);
and U48202 (N_48202,N_42931,N_41036);
nor U48203 (N_48203,N_43365,N_40771);
nand U48204 (N_48204,N_44810,N_43108);
and U48205 (N_48205,N_42113,N_43126);
or U48206 (N_48206,N_40039,N_40835);
nand U48207 (N_48207,N_40428,N_42406);
and U48208 (N_48208,N_40151,N_42435);
and U48209 (N_48209,N_40093,N_43393);
nor U48210 (N_48210,N_42540,N_42902);
nor U48211 (N_48211,N_41644,N_40911);
nand U48212 (N_48212,N_44192,N_42986);
nor U48213 (N_48213,N_41258,N_41037);
and U48214 (N_48214,N_40059,N_42686);
or U48215 (N_48215,N_44231,N_44999);
and U48216 (N_48216,N_42523,N_40178);
xnor U48217 (N_48217,N_43219,N_43155);
or U48218 (N_48218,N_40754,N_40939);
and U48219 (N_48219,N_41143,N_41957);
nor U48220 (N_48220,N_44672,N_40983);
and U48221 (N_48221,N_40648,N_40578);
nand U48222 (N_48222,N_41625,N_41462);
or U48223 (N_48223,N_42014,N_41558);
nor U48224 (N_48224,N_41988,N_43148);
xnor U48225 (N_48225,N_42410,N_40400);
or U48226 (N_48226,N_43416,N_44479);
or U48227 (N_48227,N_42625,N_40155);
xor U48228 (N_48228,N_43628,N_43005);
nor U48229 (N_48229,N_40240,N_43251);
nand U48230 (N_48230,N_42490,N_43597);
or U48231 (N_48231,N_42093,N_44879);
and U48232 (N_48232,N_44031,N_40825);
nand U48233 (N_48233,N_42447,N_42796);
and U48234 (N_48234,N_40981,N_40245);
nor U48235 (N_48235,N_42052,N_43436);
nand U48236 (N_48236,N_44703,N_44920);
or U48237 (N_48237,N_40312,N_42554);
nor U48238 (N_48238,N_44043,N_42265);
or U48239 (N_48239,N_41906,N_42051);
nor U48240 (N_48240,N_42601,N_42646);
nor U48241 (N_48241,N_44163,N_40826);
nor U48242 (N_48242,N_44988,N_40226);
and U48243 (N_48243,N_44201,N_42462);
nor U48244 (N_48244,N_44159,N_44899);
nor U48245 (N_48245,N_40725,N_41125);
or U48246 (N_48246,N_44168,N_40730);
nor U48247 (N_48247,N_44648,N_40290);
nor U48248 (N_48248,N_42694,N_41820);
xnor U48249 (N_48249,N_41448,N_44038);
and U48250 (N_48250,N_44648,N_44229);
xnor U48251 (N_48251,N_43370,N_44968);
or U48252 (N_48252,N_41074,N_44325);
nor U48253 (N_48253,N_42640,N_44613);
and U48254 (N_48254,N_43562,N_41638);
nand U48255 (N_48255,N_41302,N_40577);
nand U48256 (N_48256,N_41289,N_44941);
nand U48257 (N_48257,N_42211,N_43697);
nand U48258 (N_48258,N_42134,N_44570);
xor U48259 (N_48259,N_40276,N_40038);
and U48260 (N_48260,N_43779,N_40562);
or U48261 (N_48261,N_41394,N_42995);
and U48262 (N_48262,N_43526,N_43373);
nand U48263 (N_48263,N_40921,N_43318);
xor U48264 (N_48264,N_42455,N_42512);
xnor U48265 (N_48265,N_43816,N_44069);
nand U48266 (N_48266,N_43699,N_43540);
nor U48267 (N_48267,N_42821,N_44574);
or U48268 (N_48268,N_42786,N_41378);
or U48269 (N_48269,N_43347,N_40358);
or U48270 (N_48270,N_43239,N_41551);
or U48271 (N_48271,N_40722,N_41795);
nor U48272 (N_48272,N_44303,N_41952);
xor U48273 (N_48273,N_43384,N_43197);
nor U48274 (N_48274,N_40627,N_40617);
xnor U48275 (N_48275,N_41386,N_41638);
nand U48276 (N_48276,N_43951,N_43929);
nand U48277 (N_48277,N_43056,N_44558);
xor U48278 (N_48278,N_43842,N_41521);
and U48279 (N_48279,N_44724,N_42197);
nand U48280 (N_48280,N_41140,N_42009);
nor U48281 (N_48281,N_42296,N_43532);
and U48282 (N_48282,N_44868,N_43265);
and U48283 (N_48283,N_42476,N_41458);
or U48284 (N_48284,N_43871,N_43708);
nand U48285 (N_48285,N_43843,N_41077);
xor U48286 (N_48286,N_40623,N_43634);
nand U48287 (N_48287,N_40687,N_43252);
nor U48288 (N_48288,N_43239,N_42207);
xnor U48289 (N_48289,N_40637,N_43240);
and U48290 (N_48290,N_41427,N_40269);
or U48291 (N_48291,N_43338,N_41808);
and U48292 (N_48292,N_44475,N_40199);
nor U48293 (N_48293,N_42802,N_44015);
and U48294 (N_48294,N_43277,N_43142);
or U48295 (N_48295,N_41160,N_42347);
or U48296 (N_48296,N_40654,N_43908);
xor U48297 (N_48297,N_42860,N_43005);
or U48298 (N_48298,N_40123,N_44657);
or U48299 (N_48299,N_44575,N_44749);
nor U48300 (N_48300,N_44421,N_42295);
nand U48301 (N_48301,N_41263,N_42430);
xor U48302 (N_48302,N_44486,N_44185);
nand U48303 (N_48303,N_40896,N_40403);
nand U48304 (N_48304,N_43742,N_43713);
nand U48305 (N_48305,N_43256,N_44597);
or U48306 (N_48306,N_41068,N_42331);
nand U48307 (N_48307,N_43262,N_44774);
xor U48308 (N_48308,N_42969,N_42399);
nor U48309 (N_48309,N_44168,N_42407);
nand U48310 (N_48310,N_43121,N_41737);
nor U48311 (N_48311,N_41397,N_40500);
xnor U48312 (N_48312,N_43482,N_40610);
xnor U48313 (N_48313,N_44315,N_42125);
xnor U48314 (N_48314,N_43991,N_43786);
nor U48315 (N_48315,N_43639,N_43832);
or U48316 (N_48316,N_42343,N_41084);
and U48317 (N_48317,N_40856,N_44193);
nand U48318 (N_48318,N_43311,N_43578);
nor U48319 (N_48319,N_44051,N_44459);
xnor U48320 (N_48320,N_44527,N_40276);
xnor U48321 (N_48321,N_40349,N_43099);
or U48322 (N_48322,N_40479,N_43589);
xor U48323 (N_48323,N_40267,N_42686);
and U48324 (N_48324,N_41817,N_43814);
and U48325 (N_48325,N_43211,N_44116);
nor U48326 (N_48326,N_43242,N_43762);
nor U48327 (N_48327,N_43270,N_41519);
nor U48328 (N_48328,N_41996,N_44654);
xnor U48329 (N_48329,N_42556,N_41324);
or U48330 (N_48330,N_41843,N_42604);
and U48331 (N_48331,N_42344,N_43605);
nor U48332 (N_48332,N_42469,N_42311);
nor U48333 (N_48333,N_41540,N_43115);
or U48334 (N_48334,N_43842,N_43344);
nand U48335 (N_48335,N_41646,N_40444);
and U48336 (N_48336,N_44860,N_43947);
nand U48337 (N_48337,N_42736,N_42538);
xnor U48338 (N_48338,N_44404,N_44385);
or U48339 (N_48339,N_43851,N_40556);
nand U48340 (N_48340,N_42482,N_40447);
xor U48341 (N_48341,N_41257,N_43598);
xor U48342 (N_48342,N_43892,N_41801);
nor U48343 (N_48343,N_42101,N_40983);
and U48344 (N_48344,N_41458,N_44352);
nand U48345 (N_48345,N_44841,N_44398);
and U48346 (N_48346,N_42686,N_42653);
nor U48347 (N_48347,N_41440,N_40981);
or U48348 (N_48348,N_44628,N_41210);
nand U48349 (N_48349,N_40789,N_43474);
and U48350 (N_48350,N_40984,N_40057);
and U48351 (N_48351,N_42989,N_40003);
nand U48352 (N_48352,N_44607,N_44525);
and U48353 (N_48353,N_41737,N_41433);
nand U48354 (N_48354,N_42695,N_40924);
or U48355 (N_48355,N_42421,N_44506);
and U48356 (N_48356,N_42422,N_42880);
nand U48357 (N_48357,N_40601,N_43277);
nand U48358 (N_48358,N_44940,N_40120);
nor U48359 (N_48359,N_44540,N_41090);
xor U48360 (N_48360,N_41557,N_42236);
or U48361 (N_48361,N_40964,N_44178);
and U48362 (N_48362,N_40538,N_41474);
or U48363 (N_48363,N_44802,N_43115);
and U48364 (N_48364,N_41696,N_44816);
nand U48365 (N_48365,N_41175,N_43291);
nor U48366 (N_48366,N_40229,N_43570);
and U48367 (N_48367,N_43498,N_43160);
nor U48368 (N_48368,N_43848,N_41695);
and U48369 (N_48369,N_40795,N_40223);
xnor U48370 (N_48370,N_43899,N_40488);
and U48371 (N_48371,N_40831,N_42959);
nor U48372 (N_48372,N_41966,N_42233);
and U48373 (N_48373,N_42017,N_41997);
or U48374 (N_48374,N_43917,N_43127);
and U48375 (N_48375,N_40619,N_40429);
and U48376 (N_48376,N_40337,N_40805);
or U48377 (N_48377,N_41579,N_43171);
and U48378 (N_48378,N_43468,N_42043);
xnor U48379 (N_48379,N_43370,N_42305);
and U48380 (N_48380,N_42991,N_41205);
or U48381 (N_48381,N_41252,N_44447);
xor U48382 (N_48382,N_42412,N_44753);
xnor U48383 (N_48383,N_41283,N_44058);
or U48384 (N_48384,N_43954,N_44095);
nand U48385 (N_48385,N_41513,N_42191);
or U48386 (N_48386,N_44385,N_43734);
xnor U48387 (N_48387,N_41450,N_40777);
xnor U48388 (N_48388,N_44747,N_41199);
nand U48389 (N_48389,N_43207,N_42707);
nand U48390 (N_48390,N_42104,N_41290);
nor U48391 (N_48391,N_42737,N_43140);
or U48392 (N_48392,N_43663,N_44696);
and U48393 (N_48393,N_43011,N_41377);
xnor U48394 (N_48394,N_41061,N_42795);
nor U48395 (N_48395,N_40034,N_41496);
nor U48396 (N_48396,N_44151,N_42900);
nor U48397 (N_48397,N_40885,N_41005);
or U48398 (N_48398,N_42164,N_44868);
nand U48399 (N_48399,N_42042,N_40648);
or U48400 (N_48400,N_40120,N_41603);
or U48401 (N_48401,N_41099,N_42361);
and U48402 (N_48402,N_41661,N_44506);
or U48403 (N_48403,N_41091,N_40289);
xor U48404 (N_48404,N_40774,N_44540);
and U48405 (N_48405,N_43029,N_41355);
xnor U48406 (N_48406,N_42073,N_42897);
or U48407 (N_48407,N_44359,N_41708);
nor U48408 (N_48408,N_41525,N_44602);
nand U48409 (N_48409,N_40738,N_43752);
xor U48410 (N_48410,N_40930,N_41846);
xor U48411 (N_48411,N_40806,N_41515);
and U48412 (N_48412,N_40926,N_44121);
or U48413 (N_48413,N_42699,N_42293);
and U48414 (N_48414,N_44691,N_41914);
and U48415 (N_48415,N_41380,N_41344);
nor U48416 (N_48416,N_44520,N_43488);
or U48417 (N_48417,N_42584,N_42092);
and U48418 (N_48418,N_40610,N_43588);
nand U48419 (N_48419,N_43852,N_43200);
and U48420 (N_48420,N_41910,N_42557);
xnor U48421 (N_48421,N_43149,N_41767);
xnor U48422 (N_48422,N_44089,N_40942);
xor U48423 (N_48423,N_43501,N_44749);
and U48424 (N_48424,N_42028,N_40669);
or U48425 (N_48425,N_40693,N_43394);
and U48426 (N_48426,N_44889,N_40850);
nand U48427 (N_48427,N_41368,N_44821);
nand U48428 (N_48428,N_41973,N_41000);
or U48429 (N_48429,N_44384,N_40880);
nand U48430 (N_48430,N_41847,N_40605);
nand U48431 (N_48431,N_41384,N_41830);
and U48432 (N_48432,N_42144,N_44318);
or U48433 (N_48433,N_41133,N_43539);
and U48434 (N_48434,N_42558,N_43853);
or U48435 (N_48435,N_43783,N_40216);
or U48436 (N_48436,N_41549,N_41938);
and U48437 (N_48437,N_41172,N_41558);
and U48438 (N_48438,N_44880,N_44695);
nand U48439 (N_48439,N_40307,N_42025);
nor U48440 (N_48440,N_44425,N_44063);
nand U48441 (N_48441,N_41417,N_41142);
nand U48442 (N_48442,N_40798,N_40523);
or U48443 (N_48443,N_43412,N_43034);
nor U48444 (N_48444,N_44557,N_41804);
nand U48445 (N_48445,N_41611,N_44292);
and U48446 (N_48446,N_42235,N_41662);
and U48447 (N_48447,N_43166,N_40576);
nand U48448 (N_48448,N_43911,N_40866);
nor U48449 (N_48449,N_43654,N_42781);
or U48450 (N_48450,N_40428,N_43801);
nor U48451 (N_48451,N_40384,N_42974);
nand U48452 (N_48452,N_40695,N_41102);
nor U48453 (N_48453,N_43738,N_43864);
and U48454 (N_48454,N_43193,N_40557);
and U48455 (N_48455,N_40451,N_43611);
nand U48456 (N_48456,N_44247,N_44394);
or U48457 (N_48457,N_43158,N_43061);
nor U48458 (N_48458,N_44348,N_40985);
or U48459 (N_48459,N_43050,N_44851);
xnor U48460 (N_48460,N_40707,N_40702);
or U48461 (N_48461,N_43361,N_42748);
xnor U48462 (N_48462,N_41554,N_40190);
and U48463 (N_48463,N_41225,N_41427);
nand U48464 (N_48464,N_42293,N_40071);
nor U48465 (N_48465,N_43654,N_41955);
nor U48466 (N_48466,N_41356,N_42523);
nor U48467 (N_48467,N_44995,N_43586);
nand U48468 (N_48468,N_43517,N_41422);
or U48469 (N_48469,N_40886,N_42351);
xor U48470 (N_48470,N_44281,N_43608);
nor U48471 (N_48471,N_41651,N_43407);
nor U48472 (N_48472,N_42384,N_43734);
or U48473 (N_48473,N_42537,N_40644);
xnor U48474 (N_48474,N_42993,N_40719);
nor U48475 (N_48475,N_41021,N_40925);
nor U48476 (N_48476,N_43632,N_43331);
and U48477 (N_48477,N_43707,N_43912);
nand U48478 (N_48478,N_42069,N_44245);
or U48479 (N_48479,N_43908,N_41498);
and U48480 (N_48480,N_41201,N_41978);
nor U48481 (N_48481,N_42602,N_42054);
nor U48482 (N_48482,N_42645,N_41399);
or U48483 (N_48483,N_43615,N_43394);
nor U48484 (N_48484,N_42991,N_44158);
and U48485 (N_48485,N_41844,N_40338);
xor U48486 (N_48486,N_43240,N_43110);
nand U48487 (N_48487,N_40626,N_41946);
xor U48488 (N_48488,N_41274,N_40454);
xor U48489 (N_48489,N_40804,N_42681);
or U48490 (N_48490,N_42106,N_41785);
xnor U48491 (N_48491,N_44497,N_43673);
and U48492 (N_48492,N_42332,N_44294);
xnor U48493 (N_48493,N_41067,N_43205);
nor U48494 (N_48494,N_40677,N_43026);
nand U48495 (N_48495,N_41252,N_40276);
and U48496 (N_48496,N_42118,N_44151);
and U48497 (N_48497,N_40926,N_43230);
nor U48498 (N_48498,N_41089,N_44922);
nand U48499 (N_48499,N_41386,N_41830);
nor U48500 (N_48500,N_44459,N_42035);
nand U48501 (N_48501,N_44717,N_44221);
or U48502 (N_48502,N_42859,N_44097);
or U48503 (N_48503,N_43526,N_44824);
or U48504 (N_48504,N_41770,N_44626);
xnor U48505 (N_48505,N_41747,N_40274);
nand U48506 (N_48506,N_42262,N_43340);
and U48507 (N_48507,N_42859,N_43973);
nor U48508 (N_48508,N_42107,N_43386);
nor U48509 (N_48509,N_42526,N_40006);
and U48510 (N_48510,N_43785,N_42687);
and U48511 (N_48511,N_40647,N_41113);
nand U48512 (N_48512,N_40210,N_44540);
or U48513 (N_48513,N_40506,N_43356);
xnor U48514 (N_48514,N_41156,N_44032);
nor U48515 (N_48515,N_43562,N_42192);
xor U48516 (N_48516,N_40654,N_44832);
xnor U48517 (N_48517,N_44145,N_43237);
nor U48518 (N_48518,N_44142,N_42025);
nand U48519 (N_48519,N_41388,N_41397);
and U48520 (N_48520,N_40694,N_40155);
or U48521 (N_48521,N_43740,N_41118);
xnor U48522 (N_48522,N_41637,N_42815);
xnor U48523 (N_48523,N_42194,N_42353);
nor U48524 (N_48524,N_41329,N_42751);
and U48525 (N_48525,N_41209,N_44112);
nand U48526 (N_48526,N_40194,N_43360);
and U48527 (N_48527,N_40434,N_42191);
nand U48528 (N_48528,N_42524,N_44373);
nand U48529 (N_48529,N_41020,N_43518);
xnor U48530 (N_48530,N_43245,N_42362);
nor U48531 (N_48531,N_43543,N_42540);
and U48532 (N_48532,N_43225,N_41798);
or U48533 (N_48533,N_44453,N_44784);
or U48534 (N_48534,N_41070,N_41681);
nor U48535 (N_48535,N_43968,N_41247);
xor U48536 (N_48536,N_41171,N_42095);
and U48537 (N_48537,N_43479,N_41169);
xor U48538 (N_48538,N_44543,N_44726);
xnor U48539 (N_48539,N_44856,N_41374);
xnor U48540 (N_48540,N_41329,N_43382);
nor U48541 (N_48541,N_41768,N_41499);
nor U48542 (N_48542,N_42743,N_43075);
or U48543 (N_48543,N_40450,N_41808);
nor U48544 (N_48544,N_44561,N_43591);
xnor U48545 (N_48545,N_40307,N_43799);
or U48546 (N_48546,N_44341,N_41926);
xnor U48547 (N_48547,N_42219,N_42095);
xnor U48548 (N_48548,N_41443,N_44561);
nor U48549 (N_48549,N_41857,N_41237);
nand U48550 (N_48550,N_40336,N_43046);
and U48551 (N_48551,N_42468,N_43903);
and U48552 (N_48552,N_44121,N_40349);
and U48553 (N_48553,N_43375,N_41559);
and U48554 (N_48554,N_41307,N_44424);
nor U48555 (N_48555,N_42526,N_44915);
nand U48556 (N_48556,N_40746,N_42656);
or U48557 (N_48557,N_41531,N_42357);
nor U48558 (N_48558,N_42381,N_40882);
nor U48559 (N_48559,N_43650,N_40044);
or U48560 (N_48560,N_44435,N_41281);
and U48561 (N_48561,N_42416,N_43675);
nand U48562 (N_48562,N_41711,N_43226);
nand U48563 (N_48563,N_40076,N_43678);
nand U48564 (N_48564,N_43736,N_41877);
nor U48565 (N_48565,N_40846,N_41689);
and U48566 (N_48566,N_44582,N_40046);
xnor U48567 (N_48567,N_41413,N_43729);
nor U48568 (N_48568,N_41619,N_43730);
nand U48569 (N_48569,N_42837,N_44959);
and U48570 (N_48570,N_41075,N_41259);
nor U48571 (N_48571,N_42993,N_42488);
xor U48572 (N_48572,N_40097,N_42298);
nand U48573 (N_48573,N_41253,N_43312);
xor U48574 (N_48574,N_43993,N_42655);
xor U48575 (N_48575,N_43154,N_41290);
nand U48576 (N_48576,N_40921,N_41456);
nor U48577 (N_48577,N_44507,N_44484);
xnor U48578 (N_48578,N_41114,N_43245);
nor U48579 (N_48579,N_40085,N_41702);
or U48580 (N_48580,N_41822,N_42879);
or U48581 (N_48581,N_40197,N_44165);
nand U48582 (N_48582,N_43586,N_44472);
nor U48583 (N_48583,N_42471,N_40999);
nand U48584 (N_48584,N_42047,N_42293);
nor U48585 (N_48585,N_40753,N_40751);
and U48586 (N_48586,N_44220,N_40213);
or U48587 (N_48587,N_44919,N_41446);
xor U48588 (N_48588,N_43982,N_43432);
nand U48589 (N_48589,N_43811,N_43355);
nor U48590 (N_48590,N_40307,N_41293);
nand U48591 (N_48591,N_41626,N_41054);
xnor U48592 (N_48592,N_40249,N_44485);
xnor U48593 (N_48593,N_40268,N_43228);
nor U48594 (N_48594,N_41686,N_40810);
nor U48595 (N_48595,N_42911,N_40155);
and U48596 (N_48596,N_42865,N_44586);
nand U48597 (N_48597,N_44946,N_43517);
and U48598 (N_48598,N_43194,N_43709);
and U48599 (N_48599,N_40754,N_42460);
nand U48600 (N_48600,N_42762,N_44759);
xor U48601 (N_48601,N_40338,N_43894);
and U48602 (N_48602,N_44625,N_42177);
and U48603 (N_48603,N_43844,N_41168);
or U48604 (N_48604,N_44208,N_44592);
xor U48605 (N_48605,N_43528,N_40497);
and U48606 (N_48606,N_42715,N_42353);
nand U48607 (N_48607,N_43642,N_40707);
xor U48608 (N_48608,N_42942,N_41807);
and U48609 (N_48609,N_41426,N_42437);
and U48610 (N_48610,N_40376,N_40103);
nor U48611 (N_48611,N_43013,N_43393);
or U48612 (N_48612,N_44257,N_44127);
or U48613 (N_48613,N_43454,N_41340);
or U48614 (N_48614,N_40137,N_43088);
nand U48615 (N_48615,N_41300,N_42476);
or U48616 (N_48616,N_42974,N_44933);
xnor U48617 (N_48617,N_40405,N_40510);
xor U48618 (N_48618,N_44198,N_42599);
nor U48619 (N_48619,N_40792,N_43366);
and U48620 (N_48620,N_40614,N_41242);
nand U48621 (N_48621,N_44091,N_42175);
nor U48622 (N_48622,N_44760,N_41644);
xnor U48623 (N_48623,N_42160,N_43532);
xnor U48624 (N_48624,N_42365,N_40252);
and U48625 (N_48625,N_41663,N_44561);
xnor U48626 (N_48626,N_44788,N_41494);
and U48627 (N_48627,N_41764,N_41070);
or U48628 (N_48628,N_44518,N_44931);
or U48629 (N_48629,N_43804,N_42729);
xor U48630 (N_48630,N_44116,N_40195);
nor U48631 (N_48631,N_42553,N_42418);
nor U48632 (N_48632,N_40367,N_43542);
and U48633 (N_48633,N_44108,N_40957);
xnor U48634 (N_48634,N_40612,N_43383);
xor U48635 (N_48635,N_40802,N_41126);
and U48636 (N_48636,N_42394,N_40497);
and U48637 (N_48637,N_41418,N_42476);
and U48638 (N_48638,N_41995,N_44001);
xnor U48639 (N_48639,N_40653,N_44275);
and U48640 (N_48640,N_42647,N_44773);
and U48641 (N_48641,N_40535,N_40389);
or U48642 (N_48642,N_43703,N_40460);
and U48643 (N_48643,N_44849,N_43487);
and U48644 (N_48644,N_42216,N_40814);
nor U48645 (N_48645,N_42641,N_41107);
nor U48646 (N_48646,N_40004,N_41664);
or U48647 (N_48647,N_40798,N_42195);
nand U48648 (N_48648,N_40355,N_40545);
or U48649 (N_48649,N_41916,N_43629);
nor U48650 (N_48650,N_40197,N_42275);
or U48651 (N_48651,N_41907,N_43620);
nor U48652 (N_48652,N_40967,N_41322);
xor U48653 (N_48653,N_42101,N_42719);
xor U48654 (N_48654,N_41220,N_43713);
nand U48655 (N_48655,N_41784,N_44579);
nor U48656 (N_48656,N_41806,N_41365);
nand U48657 (N_48657,N_42698,N_42563);
nand U48658 (N_48658,N_41288,N_40688);
nor U48659 (N_48659,N_41972,N_43183);
nor U48660 (N_48660,N_43425,N_41320);
nor U48661 (N_48661,N_43829,N_42839);
xor U48662 (N_48662,N_42705,N_41328);
xor U48663 (N_48663,N_41927,N_42453);
xnor U48664 (N_48664,N_41167,N_44000);
xor U48665 (N_48665,N_42208,N_40819);
or U48666 (N_48666,N_44307,N_41836);
nand U48667 (N_48667,N_40059,N_40530);
xor U48668 (N_48668,N_41915,N_41438);
nor U48669 (N_48669,N_42879,N_43437);
nand U48670 (N_48670,N_41005,N_42849);
nand U48671 (N_48671,N_40372,N_44062);
and U48672 (N_48672,N_40507,N_44748);
nand U48673 (N_48673,N_41611,N_43866);
nor U48674 (N_48674,N_43448,N_44142);
or U48675 (N_48675,N_41210,N_41653);
nor U48676 (N_48676,N_44761,N_41266);
nand U48677 (N_48677,N_41935,N_40519);
nor U48678 (N_48678,N_40826,N_43835);
and U48679 (N_48679,N_44230,N_41510);
nand U48680 (N_48680,N_44246,N_44967);
nand U48681 (N_48681,N_44836,N_40482);
and U48682 (N_48682,N_40725,N_44481);
and U48683 (N_48683,N_40636,N_41476);
nor U48684 (N_48684,N_40120,N_40284);
and U48685 (N_48685,N_41273,N_44382);
nor U48686 (N_48686,N_43139,N_41987);
or U48687 (N_48687,N_44923,N_43053);
or U48688 (N_48688,N_44328,N_44265);
or U48689 (N_48689,N_44279,N_40694);
nor U48690 (N_48690,N_40162,N_40033);
nand U48691 (N_48691,N_41992,N_44014);
or U48692 (N_48692,N_41913,N_40000);
xnor U48693 (N_48693,N_41201,N_40813);
and U48694 (N_48694,N_40491,N_40871);
and U48695 (N_48695,N_41729,N_40643);
xnor U48696 (N_48696,N_44263,N_40448);
nand U48697 (N_48697,N_41848,N_43144);
nor U48698 (N_48698,N_41666,N_42737);
nor U48699 (N_48699,N_40309,N_41276);
or U48700 (N_48700,N_40194,N_44888);
and U48701 (N_48701,N_41421,N_41966);
and U48702 (N_48702,N_41119,N_43329);
xor U48703 (N_48703,N_41942,N_43030);
and U48704 (N_48704,N_40423,N_40401);
and U48705 (N_48705,N_40389,N_40531);
xnor U48706 (N_48706,N_43491,N_42882);
and U48707 (N_48707,N_44254,N_42490);
nor U48708 (N_48708,N_43048,N_43921);
or U48709 (N_48709,N_42973,N_40299);
nor U48710 (N_48710,N_44898,N_42578);
or U48711 (N_48711,N_43570,N_43457);
nor U48712 (N_48712,N_42260,N_43000);
nor U48713 (N_48713,N_41623,N_40114);
and U48714 (N_48714,N_40838,N_44419);
and U48715 (N_48715,N_43176,N_42965);
xor U48716 (N_48716,N_40067,N_42689);
nand U48717 (N_48717,N_40697,N_43725);
or U48718 (N_48718,N_41168,N_40044);
xnor U48719 (N_48719,N_40344,N_42329);
or U48720 (N_48720,N_43899,N_44093);
xor U48721 (N_48721,N_44329,N_40715);
or U48722 (N_48722,N_44565,N_44277);
nor U48723 (N_48723,N_44049,N_41917);
and U48724 (N_48724,N_41791,N_44379);
and U48725 (N_48725,N_43472,N_44370);
and U48726 (N_48726,N_42794,N_43898);
or U48727 (N_48727,N_40539,N_44849);
nand U48728 (N_48728,N_40536,N_43008);
and U48729 (N_48729,N_43470,N_44411);
xnor U48730 (N_48730,N_44113,N_42868);
nand U48731 (N_48731,N_44115,N_44729);
nor U48732 (N_48732,N_40678,N_42235);
nor U48733 (N_48733,N_41308,N_42712);
nand U48734 (N_48734,N_40941,N_42797);
or U48735 (N_48735,N_40160,N_44924);
nand U48736 (N_48736,N_40490,N_40657);
or U48737 (N_48737,N_44318,N_43418);
or U48738 (N_48738,N_41313,N_41498);
and U48739 (N_48739,N_42956,N_41266);
nor U48740 (N_48740,N_40053,N_43444);
nand U48741 (N_48741,N_40549,N_44646);
xnor U48742 (N_48742,N_42160,N_40871);
nor U48743 (N_48743,N_41328,N_42459);
xnor U48744 (N_48744,N_41396,N_43598);
or U48745 (N_48745,N_44607,N_42934);
xnor U48746 (N_48746,N_44440,N_41959);
nand U48747 (N_48747,N_40098,N_40812);
and U48748 (N_48748,N_42346,N_42331);
and U48749 (N_48749,N_40550,N_43680);
and U48750 (N_48750,N_44953,N_42737);
or U48751 (N_48751,N_42105,N_43700);
nand U48752 (N_48752,N_41008,N_42561);
nor U48753 (N_48753,N_42290,N_41910);
and U48754 (N_48754,N_40853,N_42222);
and U48755 (N_48755,N_42307,N_41372);
and U48756 (N_48756,N_42011,N_42727);
nor U48757 (N_48757,N_40474,N_41154);
and U48758 (N_48758,N_44018,N_42956);
and U48759 (N_48759,N_41651,N_42006);
xnor U48760 (N_48760,N_44785,N_42896);
and U48761 (N_48761,N_43134,N_41140);
xnor U48762 (N_48762,N_40058,N_40062);
and U48763 (N_48763,N_40535,N_41499);
and U48764 (N_48764,N_42807,N_40598);
nand U48765 (N_48765,N_41522,N_40576);
xor U48766 (N_48766,N_41356,N_44759);
nand U48767 (N_48767,N_40688,N_40054);
nand U48768 (N_48768,N_42249,N_41524);
xnor U48769 (N_48769,N_42678,N_42385);
or U48770 (N_48770,N_40242,N_41504);
and U48771 (N_48771,N_41707,N_42163);
xor U48772 (N_48772,N_43151,N_43417);
or U48773 (N_48773,N_43695,N_40753);
xnor U48774 (N_48774,N_43342,N_40294);
or U48775 (N_48775,N_44133,N_42253);
xnor U48776 (N_48776,N_41636,N_40441);
or U48777 (N_48777,N_41088,N_41807);
nor U48778 (N_48778,N_43433,N_44316);
nand U48779 (N_48779,N_40283,N_41132);
and U48780 (N_48780,N_42434,N_43302);
nor U48781 (N_48781,N_43476,N_43112);
and U48782 (N_48782,N_43648,N_42972);
and U48783 (N_48783,N_43049,N_44260);
and U48784 (N_48784,N_42603,N_41618);
xor U48785 (N_48785,N_43597,N_41444);
nand U48786 (N_48786,N_44258,N_40859);
xor U48787 (N_48787,N_41844,N_41889);
nand U48788 (N_48788,N_41833,N_42506);
nor U48789 (N_48789,N_44756,N_44536);
nand U48790 (N_48790,N_42225,N_41058);
xor U48791 (N_48791,N_42160,N_40976);
nand U48792 (N_48792,N_41287,N_42386);
xnor U48793 (N_48793,N_40013,N_41955);
or U48794 (N_48794,N_41275,N_42789);
xnor U48795 (N_48795,N_41174,N_44284);
xor U48796 (N_48796,N_43581,N_42375);
nand U48797 (N_48797,N_44042,N_40546);
or U48798 (N_48798,N_43567,N_41324);
or U48799 (N_48799,N_44542,N_44515);
nand U48800 (N_48800,N_42558,N_43921);
nand U48801 (N_48801,N_43780,N_43746);
and U48802 (N_48802,N_40126,N_41710);
or U48803 (N_48803,N_44939,N_41464);
and U48804 (N_48804,N_44210,N_43389);
nor U48805 (N_48805,N_40595,N_42640);
or U48806 (N_48806,N_41735,N_40828);
xor U48807 (N_48807,N_43081,N_41077);
nand U48808 (N_48808,N_41973,N_43425);
or U48809 (N_48809,N_42341,N_40985);
or U48810 (N_48810,N_41346,N_43563);
xor U48811 (N_48811,N_41136,N_44625);
or U48812 (N_48812,N_40807,N_42845);
xnor U48813 (N_48813,N_40055,N_41127);
nor U48814 (N_48814,N_42030,N_43550);
and U48815 (N_48815,N_44430,N_43983);
nor U48816 (N_48816,N_41807,N_43258);
and U48817 (N_48817,N_43337,N_43416);
and U48818 (N_48818,N_43704,N_41734);
xor U48819 (N_48819,N_44901,N_44142);
and U48820 (N_48820,N_41735,N_42615);
or U48821 (N_48821,N_40743,N_42581);
and U48822 (N_48822,N_40583,N_40731);
or U48823 (N_48823,N_43900,N_41752);
xor U48824 (N_48824,N_42987,N_43061);
xnor U48825 (N_48825,N_42190,N_43894);
nor U48826 (N_48826,N_40387,N_42502);
nand U48827 (N_48827,N_40693,N_44982);
or U48828 (N_48828,N_40813,N_43125);
or U48829 (N_48829,N_42800,N_42177);
or U48830 (N_48830,N_42649,N_42356);
or U48831 (N_48831,N_43518,N_43740);
or U48832 (N_48832,N_40132,N_44990);
and U48833 (N_48833,N_40335,N_41537);
xor U48834 (N_48834,N_41148,N_42675);
xor U48835 (N_48835,N_41331,N_41133);
nand U48836 (N_48836,N_42630,N_44331);
and U48837 (N_48837,N_42587,N_42923);
and U48838 (N_48838,N_43717,N_41764);
and U48839 (N_48839,N_40944,N_44584);
nor U48840 (N_48840,N_44039,N_43566);
and U48841 (N_48841,N_41396,N_40128);
nand U48842 (N_48842,N_41768,N_42121);
nor U48843 (N_48843,N_40205,N_40754);
nor U48844 (N_48844,N_44728,N_43775);
and U48845 (N_48845,N_41361,N_43508);
nor U48846 (N_48846,N_40748,N_44425);
and U48847 (N_48847,N_40373,N_44434);
and U48848 (N_48848,N_43810,N_42277);
nor U48849 (N_48849,N_43944,N_43160);
or U48850 (N_48850,N_43898,N_41218);
xor U48851 (N_48851,N_40622,N_42538);
or U48852 (N_48852,N_41039,N_44369);
xor U48853 (N_48853,N_40224,N_44300);
nand U48854 (N_48854,N_40336,N_44955);
xor U48855 (N_48855,N_40789,N_40032);
xnor U48856 (N_48856,N_43530,N_43671);
nor U48857 (N_48857,N_42245,N_41020);
xnor U48858 (N_48858,N_41363,N_43036);
nor U48859 (N_48859,N_44662,N_40525);
xnor U48860 (N_48860,N_43974,N_41628);
and U48861 (N_48861,N_42919,N_42385);
or U48862 (N_48862,N_44770,N_43414);
and U48863 (N_48863,N_41046,N_42516);
and U48864 (N_48864,N_42948,N_43507);
nand U48865 (N_48865,N_42559,N_40243);
nand U48866 (N_48866,N_41048,N_43292);
xnor U48867 (N_48867,N_41708,N_41928);
nor U48868 (N_48868,N_41227,N_43797);
nand U48869 (N_48869,N_42243,N_40100);
and U48870 (N_48870,N_41963,N_44650);
xor U48871 (N_48871,N_40120,N_44301);
nand U48872 (N_48872,N_42754,N_44825);
nand U48873 (N_48873,N_41323,N_43560);
or U48874 (N_48874,N_42353,N_42970);
and U48875 (N_48875,N_42620,N_44948);
nand U48876 (N_48876,N_43012,N_43412);
and U48877 (N_48877,N_42581,N_40105);
xnor U48878 (N_48878,N_44118,N_42755);
nor U48879 (N_48879,N_42094,N_43542);
and U48880 (N_48880,N_43955,N_42388);
nor U48881 (N_48881,N_43403,N_42648);
nand U48882 (N_48882,N_43573,N_43331);
nand U48883 (N_48883,N_44636,N_43556);
nor U48884 (N_48884,N_42266,N_44298);
xnor U48885 (N_48885,N_44876,N_42771);
or U48886 (N_48886,N_43181,N_42810);
and U48887 (N_48887,N_41876,N_41939);
nand U48888 (N_48888,N_43382,N_40222);
nand U48889 (N_48889,N_41938,N_44256);
nor U48890 (N_48890,N_42347,N_44108);
nor U48891 (N_48891,N_40429,N_41129);
and U48892 (N_48892,N_44797,N_43224);
nor U48893 (N_48893,N_41102,N_44785);
or U48894 (N_48894,N_44905,N_43231);
and U48895 (N_48895,N_43449,N_42945);
xnor U48896 (N_48896,N_43676,N_43619);
and U48897 (N_48897,N_44789,N_40128);
nand U48898 (N_48898,N_44469,N_40711);
nor U48899 (N_48899,N_42622,N_42533);
nand U48900 (N_48900,N_44792,N_40379);
nand U48901 (N_48901,N_44748,N_41072);
nor U48902 (N_48902,N_43549,N_43081);
and U48903 (N_48903,N_43209,N_42223);
and U48904 (N_48904,N_40919,N_42891);
nor U48905 (N_48905,N_42961,N_44829);
xnor U48906 (N_48906,N_44052,N_41337);
or U48907 (N_48907,N_43551,N_44705);
xor U48908 (N_48908,N_41050,N_41885);
nand U48909 (N_48909,N_44646,N_42347);
xor U48910 (N_48910,N_42866,N_43922);
nor U48911 (N_48911,N_43407,N_44136);
or U48912 (N_48912,N_43750,N_40756);
or U48913 (N_48913,N_40178,N_44998);
nor U48914 (N_48914,N_44567,N_42467);
xor U48915 (N_48915,N_44552,N_44044);
or U48916 (N_48916,N_40252,N_40942);
or U48917 (N_48917,N_44008,N_41411);
nor U48918 (N_48918,N_42675,N_40319);
and U48919 (N_48919,N_40512,N_40277);
nand U48920 (N_48920,N_40011,N_42681);
nand U48921 (N_48921,N_41025,N_43142);
nor U48922 (N_48922,N_42447,N_40473);
xor U48923 (N_48923,N_40042,N_44522);
or U48924 (N_48924,N_44944,N_44212);
nor U48925 (N_48925,N_43612,N_43663);
xnor U48926 (N_48926,N_42857,N_42255);
nor U48927 (N_48927,N_41829,N_41155);
nor U48928 (N_48928,N_40656,N_44634);
and U48929 (N_48929,N_42626,N_42640);
xor U48930 (N_48930,N_41264,N_42100);
nand U48931 (N_48931,N_43779,N_40501);
or U48932 (N_48932,N_43598,N_42302);
xor U48933 (N_48933,N_42654,N_40653);
or U48934 (N_48934,N_40602,N_43976);
or U48935 (N_48935,N_43331,N_43700);
nor U48936 (N_48936,N_41094,N_41093);
and U48937 (N_48937,N_40834,N_40242);
nand U48938 (N_48938,N_44325,N_40960);
or U48939 (N_48939,N_44346,N_40487);
xor U48940 (N_48940,N_44476,N_43362);
and U48941 (N_48941,N_42972,N_40966);
nor U48942 (N_48942,N_44613,N_43663);
xor U48943 (N_48943,N_41820,N_44719);
nor U48944 (N_48944,N_40582,N_44122);
and U48945 (N_48945,N_42188,N_40231);
nand U48946 (N_48946,N_41212,N_41497);
xor U48947 (N_48947,N_41879,N_42632);
and U48948 (N_48948,N_42442,N_43930);
and U48949 (N_48949,N_43417,N_40954);
xnor U48950 (N_48950,N_43609,N_41837);
nor U48951 (N_48951,N_40655,N_42667);
and U48952 (N_48952,N_42231,N_42888);
xor U48953 (N_48953,N_42011,N_44664);
nand U48954 (N_48954,N_43435,N_42206);
and U48955 (N_48955,N_40507,N_44491);
and U48956 (N_48956,N_43963,N_40726);
or U48957 (N_48957,N_44219,N_40490);
xor U48958 (N_48958,N_42202,N_44805);
xor U48959 (N_48959,N_42696,N_43223);
or U48960 (N_48960,N_40579,N_43438);
or U48961 (N_48961,N_44260,N_40568);
or U48962 (N_48962,N_43597,N_40333);
xor U48963 (N_48963,N_42562,N_41720);
or U48964 (N_48964,N_41888,N_43803);
and U48965 (N_48965,N_41539,N_44880);
nor U48966 (N_48966,N_40097,N_42488);
or U48967 (N_48967,N_43796,N_44140);
nor U48968 (N_48968,N_42617,N_41275);
and U48969 (N_48969,N_44482,N_44263);
nand U48970 (N_48970,N_44482,N_43509);
and U48971 (N_48971,N_44089,N_41328);
xnor U48972 (N_48972,N_42605,N_40279);
nand U48973 (N_48973,N_43268,N_43961);
xnor U48974 (N_48974,N_40470,N_42790);
nand U48975 (N_48975,N_40902,N_43376);
nor U48976 (N_48976,N_42222,N_41522);
xor U48977 (N_48977,N_44892,N_44086);
xor U48978 (N_48978,N_40141,N_40015);
nand U48979 (N_48979,N_44273,N_41060);
and U48980 (N_48980,N_40536,N_44479);
and U48981 (N_48981,N_40480,N_43635);
nand U48982 (N_48982,N_44141,N_42904);
nand U48983 (N_48983,N_41471,N_44424);
xnor U48984 (N_48984,N_44716,N_43256);
xor U48985 (N_48985,N_41108,N_44581);
nand U48986 (N_48986,N_40251,N_41898);
nand U48987 (N_48987,N_43676,N_42795);
nand U48988 (N_48988,N_43697,N_43765);
xor U48989 (N_48989,N_42201,N_43658);
nand U48990 (N_48990,N_44690,N_40821);
or U48991 (N_48991,N_43730,N_42768);
xnor U48992 (N_48992,N_41472,N_43810);
xnor U48993 (N_48993,N_41256,N_43314);
nand U48994 (N_48994,N_41529,N_43048);
nand U48995 (N_48995,N_41684,N_40220);
xnor U48996 (N_48996,N_43823,N_41066);
or U48997 (N_48997,N_41872,N_44152);
or U48998 (N_48998,N_41007,N_41437);
nor U48999 (N_48999,N_42671,N_42849);
xnor U49000 (N_49000,N_42465,N_44655);
xnor U49001 (N_49001,N_42673,N_40944);
xor U49002 (N_49002,N_41506,N_40812);
nor U49003 (N_49003,N_43278,N_43774);
xor U49004 (N_49004,N_40070,N_42830);
nand U49005 (N_49005,N_44364,N_40888);
nand U49006 (N_49006,N_42028,N_41653);
and U49007 (N_49007,N_44595,N_43856);
or U49008 (N_49008,N_44805,N_43698);
or U49009 (N_49009,N_44567,N_42012);
nor U49010 (N_49010,N_41493,N_41731);
nand U49011 (N_49011,N_43246,N_41504);
xnor U49012 (N_49012,N_43990,N_44787);
or U49013 (N_49013,N_40704,N_43863);
nand U49014 (N_49014,N_41821,N_41607);
or U49015 (N_49015,N_42866,N_42383);
nand U49016 (N_49016,N_42544,N_44313);
xnor U49017 (N_49017,N_43239,N_43057);
or U49018 (N_49018,N_44808,N_42653);
nand U49019 (N_49019,N_41339,N_41225);
nand U49020 (N_49020,N_41390,N_44544);
or U49021 (N_49021,N_41832,N_43377);
or U49022 (N_49022,N_42680,N_40534);
xor U49023 (N_49023,N_40798,N_42422);
or U49024 (N_49024,N_44152,N_41842);
and U49025 (N_49025,N_43119,N_43008);
nand U49026 (N_49026,N_44397,N_44574);
nand U49027 (N_49027,N_42264,N_40238);
or U49028 (N_49028,N_44514,N_44620);
or U49029 (N_49029,N_41402,N_41576);
and U49030 (N_49030,N_40068,N_41894);
xnor U49031 (N_49031,N_44450,N_44362);
xnor U49032 (N_49032,N_40631,N_44802);
xnor U49033 (N_49033,N_42928,N_43828);
and U49034 (N_49034,N_41814,N_43835);
nor U49035 (N_49035,N_42930,N_43684);
nor U49036 (N_49036,N_41323,N_43137);
xnor U49037 (N_49037,N_42610,N_44671);
xnor U49038 (N_49038,N_40125,N_44049);
nand U49039 (N_49039,N_40915,N_43156);
and U49040 (N_49040,N_44760,N_43725);
and U49041 (N_49041,N_40817,N_44272);
or U49042 (N_49042,N_40887,N_43030);
nand U49043 (N_49043,N_44056,N_43798);
or U49044 (N_49044,N_40512,N_42431);
nor U49045 (N_49045,N_41075,N_41768);
nor U49046 (N_49046,N_41208,N_44323);
nor U49047 (N_49047,N_44224,N_43669);
nand U49048 (N_49048,N_40468,N_42365);
nand U49049 (N_49049,N_44556,N_41765);
or U49050 (N_49050,N_42720,N_42207);
nand U49051 (N_49051,N_42653,N_43390);
xnor U49052 (N_49052,N_43677,N_44536);
or U49053 (N_49053,N_41632,N_41290);
or U49054 (N_49054,N_43087,N_41832);
nor U49055 (N_49055,N_41915,N_41368);
or U49056 (N_49056,N_40094,N_44371);
nand U49057 (N_49057,N_44737,N_43935);
or U49058 (N_49058,N_41106,N_44269);
nor U49059 (N_49059,N_44815,N_40911);
nor U49060 (N_49060,N_40936,N_43338);
xnor U49061 (N_49061,N_42004,N_42875);
nor U49062 (N_49062,N_40088,N_41516);
xor U49063 (N_49063,N_42167,N_42217);
nor U49064 (N_49064,N_41105,N_43911);
nand U49065 (N_49065,N_44986,N_43625);
nand U49066 (N_49066,N_42250,N_42801);
xnor U49067 (N_49067,N_41437,N_44261);
nor U49068 (N_49068,N_43590,N_41049);
or U49069 (N_49069,N_43088,N_42539);
nand U49070 (N_49070,N_40387,N_43258);
or U49071 (N_49071,N_40359,N_43651);
xnor U49072 (N_49072,N_41605,N_41956);
or U49073 (N_49073,N_43382,N_40014);
and U49074 (N_49074,N_40330,N_44028);
and U49075 (N_49075,N_42631,N_41892);
and U49076 (N_49076,N_40109,N_43465);
nand U49077 (N_49077,N_44999,N_41218);
nand U49078 (N_49078,N_40004,N_43957);
nand U49079 (N_49079,N_42847,N_42049);
nand U49080 (N_49080,N_40021,N_43984);
or U49081 (N_49081,N_41709,N_42064);
nand U49082 (N_49082,N_41426,N_44400);
nand U49083 (N_49083,N_43714,N_42394);
or U49084 (N_49084,N_41020,N_43266);
nor U49085 (N_49085,N_42328,N_42124);
nand U49086 (N_49086,N_41461,N_41509);
or U49087 (N_49087,N_42129,N_42854);
and U49088 (N_49088,N_42630,N_41153);
xor U49089 (N_49089,N_42736,N_41440);
xor U49090 (N_49090,N_42983,N_41503);
nand U49091 (N_49091,N_40127,N_40501);
xor U49092 (N_49092,N_40028,N_41075);
xnor U49093 (N_49093,N_40538,N_41172);
nor U49094 (N_49094,N_43778,N_40246);
nor U49095 (N_49095,N_43029,N_42815);
nand U49096 (N_49096,N_40795,N_40399);
xnor U49097 (N_49097,N_42237,N_43454);
and U49098 (N_49098,N_40186,N_40391);
xor U49099 (N_49099,N_41207,N_41518);
and U49100 (N_49100,N_40104,N_41199);
xnor U49101 (N_49101,N_43801,N_43653);
xnor U49102 (N_49102,N_42286,N_41253);
nand U49103 (N_49103,N_44362,N_44481);
or U49104 (N_49104,N_43137,N_43260);
nand U49105 (N_49105,N_41018,N_44177);
xnor U49106 (N_49106,N_44762,N_41687);
nor U49107 (N_49107,N_44269,N_43388);
nand U49108 (N_49108,N_44142,N_44992);
xor U49109 (N_49109,N_43149,N_41989);
xor U49110 (N_49110,N_42917,N_40308);
or U49111 (N_49111,N_44598,N_41884);
nand U49112 (N_49112,N_42610,N_43275);
nor U49113 (N_49113,N_40874,N_40869);
nor U49114 (N_49114,N_40302,N_41614);
nor U49115 (N_49115,N_40462,N_42141);
xor U49116 (N_49116,N_44221,N_44321);
nand U49117 (N_49117,N_44176,N_43226);
or U49118 (N_49118,N_41886,N_41523);
xnor U49119 (N_49119,N_43281,N_43451);
or U49120 (N_49120,N_44963,N_44187);
nor U49121 (N_49121,N_40655,N_41698);
and U49122 (N_49122,N_43038,N_43897);
nand U49123 (N_49123,N_41085,N_42851);
nor U49124 (N_49124,N_41286,N_40598);
nor U49125 (N_49125,N_44790,N_43702);
and U49126 (N_49126,N_42539,N_43384);
xnor U49127 (N_49127,N_44328,N_41196);
nand U49128 (N_49128,N_40276,N_43747);
nor U49129 (N_49129,N_40439,N_42044);
or U49130 (N_49130,N_44695,N_40625);
and U49131 (N_49131,N_42981,N_44313);
nor U49132 (N_49132,N_40995,N_43585);
nor U49133 (N_49133,N_40324,N_40594);
xnor U49134 (N_49134,N_43784,N_43415);
xor U49135 (N_49135,N_43859,N_44117);
and U49136 (N_49136,N_44566,N_41932);
nor U49137 (N_49137,N_41310,N_43096);
or U49138 (N_49138,N_43276,N_44825);
xor U49139 (N_49139,N_44259,N_41765);
nand U49140 (N_49140,N_41245,N_43281);
or U49141 (N_49141,N_41138,N_42184);
xor U49142 (N_49142,N_40330,N_42131);
or U49143 (N_49143,N_44466,N_40292);
nor U49144 (N_49144,N_44315,N_44899);
or U49145 (N_49145,N_43686,N_42448);
or U49146 (N_49146,N_43517,N_44499);
nand U49147 (N_49147,N_42063,N_44737);
nand U49148 (N_49148,N_41494,N_43294);
and U49149 (N_49149,N_42304,N_43596);
or U49150 (N_49150,N_41972,N_43136);
nand U49151 (N_49151,N_44240,N_43742);
xnor U49152 (N_49152,N_44179,N_41972);
nand U49153 (N_49153,N_42577,N_44422);
or U49154 (N_49154,N_43512,N_41023);
or U49155 (N_49155,N_43287,N_44989);
nor U49156 (N_49156,N_41717,N_43058);
nand U49157 (N_49157,N_42132,N_41795);
nor U49158 (N_49158,N_41918,N_43023);
nand U49159 (N_49159,N_41168,N_43860);
xnor U49160 (N_49160,N_44255,N_40008);
xor U49161 (N_49161,N_42185,N_42962);
or U49162 (N_49162,N_41244,N_43320);
xnor U49163 (N_49163,N_41836,N_43014);
nor U49164 (N_49164,N_42750,N_44009);
and U49165 (N_49165,N_43608,N_44486);
nand U49166 (N_49166,N_41709,N_44579);
xor U49167 (N_49167,N_43633,N_41935);
and U49168 (N_49168,N_43419,N_43167);
and U49169 (N_49169,N_41556,N_42991);
xor U49170 (N_49170,N_43284,N_40085);
nand U49171 (N_49171,N_42602,N_43008);
nor U49172 (N_49172,N_43516,N_41685);
or U49173 (N_49173,N_42503,N_43418);
nor U49174 (N_49174,N_44097,N_42327);
and U49175 (N_49175,N_40601,N_42304);
nor U49176 (N_49176,N_44298,N_41558);
xor U49177 (N_49177,N_44569,N_42783);
xor U49178 (N_49178,N_44489,N_42485);
and U49179 (N_49179,N_43903,N_42935);
xor U49180 (N_49180,N_44983,N_40145);
nand U49181 (N_49181,N_41983,N_40505);
or U49182 (N_49182,N_42485,N_42423);
xor U49183 (N_49183,N_44661,N_41359);
nand U49184 (N_49184,N_41338,N_40277);
xor U49185 (N_49185,N_40604,N_44076);
xor U49186 (N_49186,N_43772,N_43985);
or U49187 (N_49187,N_40141,N_40304);
or U49188 (N_49188,N_40759,N_42768);
xor U49189 (N_49189,N_43058,N_44238);
xor U49190 (N_49190,N_40986,N_40823);
and U49191 (N_49191,N_41422,N_43458);
xor U49192 (N_49192,N_41598,N_43354);
and U49193 (N_49193,N_44834,N_43293);
xor U49194 (N_49194,N_43589,N_40744);
or U49195 (N_49195,N_42061,N_41246);
nand U49196 (N_49196,N_42629,N_43254);
and U49197 (N_49197,N_44945,N_42071);
xnor U49198 (N_49198,N_41347,N_41250);
or U49199 (N_49199,N_42859,N_43238);
and U49200 (N_49200,N_44416,N_44589);
and U49201 (N_49201,N_41903,N_40006);
xor U49202 (N_49202,N_44941,N_44504);
or U49203 (N_49203,N_41137,N_43696);
nor U49204 (N_49204,N_41253,N_44418);
nand U49205 (N_49205,N_40046,N_44378);
nor U49206 (N_49206,N_40631,N_40335);
or U49207 (N_49207,N_43890,N_42881);
nor U49208 (N_49208,N_42215,N_42966);
and U49209 (N_49209,N_40253,N_43634);
and U49210 (N_49210,N_40827,N_42837);
and U49211 (N_49211,N_41259,N_41774);
nor U49212 (N_49212,N_44038,N_41878);
or U49213 (N_49213,N_42135,N_44660);
or U49214 (N_49214,N_40808,N_44077);
and U49215 (N_49215,N_42804,N_43025);
nor U49216 (N_49216,N_44884,N_40317);
xnor U49217 (N_49217,N_42863,N_41086);
xnor U49218 (N_49218,N_41488,N_44329);
nand U49219 (N_49219,N_42672,N_40637);
nor U49220 (N_49220,N_40999,N_44703);
xnor U49221 (N_49221,N_44215,N_44551);
nor U49222 (N_49222,N_43094,N_42677);
or U49223 (N_49223,N_40547,N_42414);
and U49224 (N_49224,N_41343,N_44240);
nand U49225 (N_49225,N_42801,N_41521);
or U49226 (N_49226,N_42924,N_44380);
nor U49227 (N_49227,N_40811,N_43110);
or U49228 (N_49228,N_41210,N_44247);
or U49229 (N_49229,N_44103,N_41961);
xnor U49230 (N_49230,N_43757,N_42590);
nor U49231 (N_49231,N_42850,N_43803);
nor U49232 (N_49232,N_43846,N_42288);
xnor U49233 (N_49233,N_44068,N_40512);
nor U49234 (N_49234,N_43504,N_43702);
xor U49235 (N_49235,N_42630,N_40542);
xor U49236 (N_49236,N_43081,N_41641);
nor U49237 (N_49237,N_44835,N_41900);
nor U49238 (N_49238,N_40873,N_40369);
nor U49239 (N_49239,N_43093,N_41006);
and U49240 (N_49240,N_41490,N_43648);
or U49241 (N_49241,N_40796,N_43946);
and U49242 (N_49242,N_41810,N_40382);
or U49243 (N_49243,N_44405,N_40456);
or U49244 (N_49244,N_43576,N_43291);
xnor U49245 (N_49245,N_41965,N_44656);
nand U49246 (N_49246,N_40839,N_40812);
nor U49247 (N_49247,N_42923,N_41332);
nor U49248 (N_49248,N_40966,N_44254);
or U49249 (N_49249,N_43648,N_44943);
nand U49250 (N_49250,N_42762,N_43699);
or U49251 (N_49251,N_43023,N_42516);
or U49252 (N_49252,N_43447,N_41769);
nand U49253 (N_49253,N_43395,N_42111);
or U49254 (N_49254,N_43438,N_40786);
xor U49255 (N_49255,N_42664,N_43814);
nor U49256 (N_49256,N_44904,N_43277);
and U49257 (N_49257,N_43510,N_44928);
or U49258 (N_49258,N_41801,N_43770);
xnor U49259 (N_49259,N_40793,N_40558);
nand U49260 (N_49260,N_43929,N_44096);
or U49261 (N_49261,N_43097,N_40858);
nand U49262 (N_49262,N_44452,N_40396);
or U49263 (N_49263,N_41876,N_42227);
nand U49264 (N_49264,N_44026,N_41017);
and U49265 (N_49265,N_43735,N_41978);
nor U49266 (N_49266,N_40793,N_42511);
xor U49267 (N_49267,N_44754,N_44903);
or U49268 (N_49268,N_44861,N_40051);
nand U49269 (N_49269,N_40213,N_43223);
nand U49270 (N_49270,N_40726,N_43585);
nor U49271 (N_49271,N_43487,N_43282);
nor U49272 (N_49272,N_43727,N_41616);
nand U49273 (N_49273,N_44894,N_43942);
and U49274 (N_49274,N_42152,N_40111);
nor U49275 (N_49275,N_40845,N_42046);
xnor U49276 (N_49276,N_42594,N_43607);
nand U49277 (N_49277,N_44995,N_40113);
or U49278 (N_49278,N_41864,N_40914);
or U49279 (N_49279,N_40899,N_43581);
nand U49280 (N_49280,N_42915,N_42736);
nor U49281 (N_49281,N_41247,N_44259);
and U49282 (N_49282,N_42712,N_40436);
and U49283 (N_49283,N_42932,N_44009);
and U49284 (N_49284,N_41228,N_42038);
nor U49285 (N_49285,N_43379,N_41580);
nand U49286 (N_49286,N_40535,N_41804);
xor U49287 (N_49287,N_41687,N_44267);
and U49288 (N_49288,N_40272,N_41939);
and U49289 (N_49289,N_40850,N_42237);
xnor U49290 (N_49290,N_40632,N_41791);
and U49291 (N_49291,N_41476,N_43804);
nand U49292 (N_49292,N_42209,N_43761);
or U49293 (N_49293,N_41573,N_41160);
and U49294 (N_49294,N_44283,N_41252);
nand U49295 (N_49295,N_40865,N_44325);
and U49296 (N_49296,N_42468,N_44609);
nor U49297 (N_49297,N_40444,N_41857);
nand U49298 (N_49298,N_41994,N_43748);
or U49299 (N_49299,N_41761,N_40586);
and U49300 (N_49300,N_42021,N_43086);
or U49301 (N_49301,N_41085,N_44740);
nor U49302 (N_49302,N_42920,N_42349);
xor U49303 (N_49303,N_41201,N_40499);
xnor U49304 (N_49304,N_44445,N_44214);
xor U49305 (N_49305,N_43908,N_43347);
nor U49306 (N_49306,N_40726,N_41132);
nor U49307 (N_49307,N_41346,N_40287);
nand U49308 (N_49308,N_40255,N_42168);
nand U49309 (N_49309,N_43676,N_42310);
and U49310 (N_49310,N_40350,N_44630);
nor U49311 (N_49311,N_44889,N_40478);
nand U49312 (N_49312,N_44334,N_40507);
nand U49313 (N_49313,N_40866,N_41463);
nor U49314 (N_49314,N_41894,N_40331);
nand U49315 (N_49315,N_40099,N_43575);
xor U49316 (N_49316,N_43877,N_44785);
nor U49317 (N_49317,N_40048,N_40490);
nor U49318 (N_49318,N_41268,N_40934);
xor U49319 (N_49319,N_40915,N_44510);
and U49320 (N_49320,N_42504,N_41435);
nor U49321 (N_49321,N_40135,N_44668);
and U49322 (N_49322,N_43302,N_42085);
or U49323 (N_49323,N_40118,N_41449);
or U49324 (N_49324,N_43141,N_40568);
xnor U49325 (N_49325,N_44775,N_42865);
nor U49326 (N_49326,N_44362,N_41166);
or U49327 (N_49327,N_40903,N_43836);
and U49328 (N_49328,N_40152,N_42163);
nand U49329 (N_49329,N_44898,N_40126);
nand U49330 (N_49330,N_44984,N_42226);
or U49331 (N_49331,N_43377,N_40698);
nand U49332 (N_49332,N_44027,N_42536);
nand U49333 (N_49333,N_42848,N_40527);
xor U49334 (N_49334,N_43938,N_41134);
nand U49335 (N_49335,N_41921,N_43401);
and U49336 (N_49336,N_40157,N_40118);
and U49337 (N_49337,N_42276,N_40586);
and U49338 (N_49338,N_41220,N_40746);
and U49339 (N_49339,N_42465,N_40067);
xnor U49340 (N_49340,N_44682,N_42581);
and U49341 (N_49341,N_42601,N_41576);
xnor U49342 (N_49342,N_44611,N_42123);
or U49343 (N_49343,N_44244,N_43243);
nor U49344 (N_49344,N_44200,N_41000);
nand U49345 (N_49345,N_43524,N_43109);
and U49346 (N_49346,N_43785,N_41865);
nor U49347 (N_49347,N_44831,N_41697);
or U49348 (N_49348,N_40431,N_44460);
or U49349 (N_49349,N_43592,N_44602);
nor U49350 (N_49350,N_43739,N_44833);
nand U49351 (N_49351,N_42782,N_41153);
xnor U49352 (N_49352,N_44021,N_41052);
nor U49353 (N_49353,N_42227,N_41128);
nor U49354 (N_49354,N_44058,N_43049);
and U49355 (N_49355,N_44454,N_44433);
nand U49356 (N_49356,N_40507,N_43157);
or U49357 (N_49357,N_44580,N_41109);
or U49358 (N_49358,N_44573,N_40348);
nand U49359 (N_49359,N_40194,N_40776);
or U49360 (N_49360,N_40273,N_44673);
nand U49361 (N_49361,N_40494,N_44358);
xor U49362 (N_49362,N_42166,N_42765);
or U49363 (N_49363,N_42346,N_40430);
nor U49364 (N_49364,N_42259,N_41099);
nor U49365 (N_49365,N_40927,N_44500);
and U49366 (N_49366,N_41023,N_40404);
nand U49367 (N_49367,N_42874,N_42537);
or U49368 (N_49368,N_41507,N_43698);
and U49369 (N_49369,N_44072,N_42578);
xnor U49370 (N_49370,N_41271,N_41805);
nor U49371 (N_49371,N_42049,N_43859);
nor U49372 (N_49372,N_40432,N_44949);
nor U49373 (N_49373,N_41188,N_40296);
nor U49374 (N_49374,N_40952,N_44068);
nand U49375 (N_49375,N_44569,N_44918);
nor U49376 (N_49376,N_42564,N_44153);
nor U49377 (N_49377,N_42841,N_44010);
nand U49378 (N_49378,N_42869,N_41251);
and U49379 (N_49379,N_42959,N_41799);
xnor U49380 (N_49380,N_42932,N_40172);
xnor U49381 (N_49381,N_40330,N_41295);
xor U49382 (N_49382,N_44007,N_43618);
nor U49383 (N_49383,N_41762,N_42456);
or U49384 (N_49384,N_42099,N_40632);
or U49385 (N_49385,N_44528,N_40207);
nor U49386 (N_49386,N_44886,N_42028);
nor U49387 (N_49387,N_41829,N_44237);
or U49388 (N_49388,N_44037,N_40521);
xnor U49389 (N_49389,N_44184,N_41424);
and U49390 (N_49390,N_42534,N_44505);
or U49391 (N_49391,N_44171,N_43600);
nor U49392 (N_49392,N_42639,N_40159);
and U49393 (N_49393,N_44791,N_43420);
nor U49394 (N_49394,N_40672,N_44175);
and U49395 (N_49395,N_44856,N_44675);
and U49396 (N_49396,N_42367,N_42370);
and U49397 (N_49397,N_41859,N_41197);
or U49398 (N_49398,N_43929,N_44352);
nor U49399 (N_49399,N_41536,N_43006);
nand U49400 (N_49400,N_40743,N_40519);
nand U49401 (N_49401,N_41016,N_40647);
or U49402 (N_49402,N_41086,N_40868);
and U49403 (N_49403,N_42057,N_43426);
xnor U49404 (N_49404,N_40808,N_40917);
xnor U49405 (N_49405,N_44617,N_41185);
nand U49406 (N_49406,N_43706,N_44365);
xnor U49407 (N_49407,N_44774,N_43087);
or U49408 (N_49408,N_43214,N_44359);
or U49409 (N_49409,N_42552,N_41047);
and U49410 (N_49410,N_41863,N_44825);
or U49411 (N_49411,N_43986,N_41947);
xor U49412 (N_49412,N_43806,N_41993);
or U49413 (N_49413,N_43148,N_40939);
or U49414 (N_49414,N_43049,N_40283);
nor U49415 (N_49415,N_41517,N_41509);
or U49416 (N_49416,N_42314,N_41441);
nand U49417 (N_49417,N_44466,N_40235);
nand U49418 (N_49418,N_41229,N_42349);
and U49419 (N_49419,N_41364,N_43416);
or U49420 (N_49420,N_43246,N_41961);
nor U49421 (N_49421,N_44849,N_40625);
xor U49422 (N_49422,N_42387,N_42161);
or U49423 (N_49423,N_41415,N_43515);
or U49424 (N_49424,N_41955,N_43410);
xor U49425 (N_49425,N_43499,N_41669);
nand U49426 (N_49426,N_40046,N_44778);
xnor U49427 (N_49427,N_40885,N_44501);
or U49428 (N_49428,N_40926,N_44716);
or U49429 (N_49429,N_41297,N_40446);
xnor U49430 (N_49430,N_41284,N_42314);
nand U49431 (N_49431,N_42488,N_44286);
xnor U49432 (N_49432,N_42584,N_41773);
and U49433 (N_49433,N_40283,N_44982);
xnor U49434 (N_49434,N_43028,N_40250);
or U49435 (N_49435,N_40758,N_44485);
nand U49436 (N_49436,N_40009,N_43493);
xor U49437 (N_49437,N_44031,N_40461);
nand U49438 (N_49438,N_40237,N_44369);
nand U49439 (N_49439,N_43247,N_44446);
nand U49440 (N_49440,N_42661,N_43180);
and U49441 (N_49441,N_42443,N_44885);
or U49442 (N_49442,N_40374,N_44219);
nor U49443 (N_49443,N_40848,N_40826);
or U49444 (N_49444,N_43221,N_43534);
nor U49445 (N_49445,N_44478,N_41515);
nor U49446 (N_49446,N_40683,N_42264);
xnor U49447 (N_49447,N_40692,N_41161);
xnor U49448 (N_49448,N_44200,N_43959);
nor U49449 (N_49449,N_40801,N_43789);
xor U49450 (N_49450,N_43239,N_42156);
and U49451 (N_49451,N_43803,N_42857);
and U49452 (N_49452,N_41808,N_42207);
nor U49453 (N_49453,N_43445,N_42897);
xnor U49454 (N_49454,N_41205,N_41727);
or U49455 (N_49455,N_41269,N_41721);
nor U49456 (N_49456,N_41136,N_41750);
nand U49457 (N_49457,N_41530,N_40288);
xor U49458 (N_49458,N_40100,N_44145);
xor U49459 (N_49459,N_41545,N_40522);
nor U49460 (N_49460,N_44122,N_42052);
nand U49461 (N_49461,N_43316,N_40659);
and U49462 (N_49462,N_40719,N_43285);
and U49463 (N_49463,N_44871,N_42603);
or U49464 (N_49464,N_40447,N_44061);
nor U49465 (N_49465,N_43404,N_42465);
xnor U49466 (N_49466,N_42695,N_43433);
nor U49467 (N_49467,N_41425,N_40771);
xor U49468 (N_49468,N_42553,N_43457);
xnor U49469 (N_49469,N_42487,N_44183);
nand U49470 (N_49470,N_43029,N_40595);
or U49471 (N_49471,N_41779,N_40941);
or U49472 (N_49472,N_42611,N_41676);
and U49473 (N_49473,N_42687,N_40934);
nor U49474 (N_49474,N_40940,N_43748);
xnor U49475 (N_49475,N_42823,N_43258);
xnor U49476 (N_49476,N_44189,N_40197);
xor U49477 (N_49477,N_43828,N_43300);
xnor U49478 (N_49478,N_40273,N_43930);
nand U49479 (N_49479,N_41247,N_42710);
nand U49480 (N_49480,N_42644,N_40674);
and U49481 (N_49481,N_44935,N_43845);
nor U49482 (N_49482,N_43159,N_42177);
nor U49483 (N_49483,N_41660,N_42972);
xor U49484 (N_49484,N_43689,N_43544);
nand U49485 (N_49485,N_43653,N_40090);
nand U49486 (N_49486,N_40810,N_44887);
xnor U49487 (N_49487,N_41331,N_40970);
nand U49488 (N_49488,N_42051,N_42949);
or U49489 (N_49489,N_43506,N_44179);
and U49490 (N_49490,N_41511,N_42422);
and U49491 (N_49491,N_41570,N_40114);
nor U49492 (N_49492,N_41088,N_44990);
and U49493 (N_49493,N_44156,N_41873);
nor U49494 (N_49494,N_44156,N_41474);
and U49495 (N_49495,N_41957,N_41083);
or U49496 (N_49496,N_44050,N_44542);
nand U49497 (N_49497,N_42540,N_44845);
nor U49498 (N_49498,N_42961,N_42749);
nand U49499 (N_49499,N_40233,N_44248);
nor U49500 (N_49500,N_42975,N_41319);
nor U49501 (N_49501,N_40943,N_43103);
or U49502 (N_49502,N_42471,N_40977);
xnor U49503 (N_49503,N_42140,N_42868);
or U49504 (N_49504,N_41968,N_43767);
nor U49505 (N_49505,N_41706,N_44578);
xnor U49506 (N_49506,N_42535,N_44739);
or U49507 (N_49507,N_41695,N_42218);
and U49508 (N_49508,N_43694,N_40907);
and U49509 (N_49509,N_43260,N_41183);
or U49510 (N_49510,N_40858,N_44179);
or U49511 (N_49511,N_44136,N_41228);
nand U49512 (N_49512,N_43207,N_42676);
nor U49513 (N_49513,N_42006,N_43446);
and U49514 (N_49514,N_41081,N_40797);
nor U49515 (N_49515,N_44351,N_43462);
or U49516 (N_49516,N_44820,N_40548);
nor U49517 (N_49517,N_44394,N_43377);
nand U49518 (N_49518,N_42743,N_44854);
and U49519 (N_49519,N_42923,N_41139);
or U49520 (N_49520,N_41930,N_40077);
xnor U49521 (N_49521,N_41098,N_43483);
or U49522 (N_49522,N_43939,N_44617);
xor U49523 (N_49523,N_41266,N_43547);
and U49524 (N_49524,N_42975,N_42172);
nand U49525 (N_49525,N_41532,N_40770);
nor U49526 (N_49526,N_41893,N_42462);
and U49527 (N_49527,N_40489,N_44291);
nor U49528 (N_49528,N_43379,N_42682);
nand U49529 (N_49529,N_44342,N_43717);
nor U49530 (N_49530,N_41483,N_40437);
xnor U49531 (N_49531,N_41341,N_41414);
nor U49532 (N_49532,N_43660,N_41535);
nand U49533 (N_49533,N_44808,N_44883);
and U49534 (N_49534,N_44653,N_43587);
nor U49535 (N_49535,N_43574,N_42875);
nor U49536 (N_49536,N_44336,N_43971);
nand U49537 (N_49537,N_40562,N_42592);
nor U49538 (N_49538,N_41357,N_42920);
and U49539 (N_49539,N_44036,N_41081);
nor U49540 (N_49540,N_44202,N_42607);
nand U49541 (N_49541,N_42945,N_42681);
nor U49542 (N_49542,N_43517,N_40605);
and U49543 (N_49543,N_42483,N_42706);
or U49544 (N_49544,N_44274,N_44108);
and U49545 (N_49545,N_40526,N_44200);
or U49546 (N_49546,N_41302,N_44774);
and U49547 (N_49547,N_43143,N_43293);
or U49548 (N_49548,N_41786,N_44519);
xor U49549 (N_49549,N_44084,N_41297);
or U49550 (N_49550,N_41841,N_44962);
or U49551 (N_49551,N_43857,N_40712);
xnor U49552 (N_49552,N_44174,N_44426);
nor U49553 (N_49553,N_42815,N_44198);
or U49554 (N_49554,N_41906,N_44452);
and U49555 (N_49555,N_43239,N_42945);
or U49556 (N_49556,N_41355,N_40151);
nand U49557 (N_49557,N_42227,N_42986);
nor U49558 (N_49558,N_43380,N_40502);
xor U49559 (N_49559,N_42704,N_42438);
or U49560 (N_49560,N_41748,N_40905);
and U49561 (N_49561,N_43270,N_41681);
or U49562 (N_49562,N_43945,N_41451);
or U49563 (N_49563,N_42814,N_40963);
and U49564 (N_49564,N_41809,N_44766);
nand U49565 (N_49565,N_42226,N_43267);
or U49566 (N_49566,N_44353,N_40543);
nor U49567 (N_49567,N_40826,N_41741);
and U49568 (N_49568,N_42175,N_40512);
xor U49569 (N_49569,N_44369,N_44256);
nor U49570 (N_49570,N_43302,N_43961);
and U49571 (N_49571,N_42170,N_40979);
nand U49572 (N_49572,N_41060,N_41026);
and U49573 (N_49573,N_40486,N_44928);
nor U49574 (N_49574,N_44831,N_40030);
nand U49575 (N_49575,N_41204,N_42817);
xor U49576 (N_49576,N_42707,N_42710);
or U49577 (N_49577,N_44775,N_44809);
or U49578 (N_49578,N_40378,N_42621);
nor U49579 (N_49579,N_43715,N_40437);
xnor U49580 (N_49580,N_40525,N_42553);
nand U49581 (N_49581,N_42184,N_41650);
and U49582 (N_49582,N_42619,N_41192);
and U49583 (N_49583,N_42240,N_40739);
nand U49584 (N_49584,N_43750,N_41435);
nand U49585 (N_49585,N_44236,N_44583);
and U49586 (N_49586,N_44248,N_42039);
nor U49587 (N_49587,N_40431,N_44192);
nand U49588 (N_49588,N_42195,N_43968);
or U49589 (N_49589,N_41003,N_40017);
xor U49590 (N_49590,N_44400,N_44795);
nor U49591 (N_49591,N_42655,N_44378);
nor U49592 (N_49592,N_41575,N_44317);
and U49593 (N_49593,N_43802,N_43339);
or U49594 (N_49594,N_43443,N_44519);
nor U49595 (N_49595,N_40844,N_40224);
xor U49596 (N_49596,N_43625,N_43916);
or U49597 (N_49597,N_40881,N_42481);
and U49598 (N_49598,N_41407,N_41418);
nand U49599 (N_49599,N_44928,N_44732);
or U49600 (N_49600,N_40670,N_42006);
nand U49601 (N_49601,N_40658,N_42443);
nand U49602 (N_49602,N_44082,N_41471);
nor U49603 (N_49603,N_42656,N_41321);
nor U49604 (N_49604,N_42461,N_40275);
nor U49605 (N_49605,N_43435,N_41908);
or U49606 (N_49606,N_41257,N_44427);
and U49607 (N_49607,N_40244,N_42229);
or U49608 (N_49608,N_42791,N_43876);
and U49609 (N_49609,N_41003,N_41064);
and U49610 (N_49610,N_40871,N_41638);
and U49611 (N_49611,N_44269,N_41590);
xnor U49612 (N_49612,N_44217,N_43497);
and U49613 (N_49613,N_42072,N_41644);
and U49614 (N_49614,N_42895,N_42831);
xor U49615 (N_49615,N_42034,N_44344);
nand U49616 (N_49616,N_40219,N_41557);
xnor U49617 (N_49617,N_40696,N_41819);
and U49618 (N_49618,N_44895,N_41361);
or U49619 (N_49619,N_44430,N_43755);
nor U49620 (N_49620,N_44462,N_41585);
nand U49621 (N_49621,N_42952,N_42247);
and U49622 (N_49622,N_44825,N_44907);
nor U49623 (N_49623,N_41584,N_40340);
and U49624 (N_49624,N_40078,N_43963);
or U49625 (N_49625,N_44629,N_44967);
or U49626 (N_49626,N_44844,N_43035);
and U49627 (N_49627,N_41866,N_44543);
and U49628 (N_49628,N_41659,N_44333);
nor U49629 (N_49629,N_44439,N_42026);
xnor U49630 (N_49630,N_41982,N_42687);
nand U49631 (N_49631,N_42592,N_43099);
or U49632 (N_49632,N_44934,N_44166);
nand U49633 (N_49633,N_40051,N_41363);
nor U49634 (N_49634,N_43377,N_40436);
and U49635 (N_49635,N_42314,N_40547);
nand U49636 (N_49636,N_41863,N_42353);
nand U49637 (N_49637,N_40869,N_43209);
nand U49638 (N_49638,N_41725,N_43042);
and U49639 (N_49639,N_44383,N_41379);
xnor U49640 (N_49640,N_43156,N_43147);
or U49641 (N_49641,N_42120,N_43538);
nor U49642 (N_49642,N_42880,N_42759);
and U49643 (N_49643,N_41042,N_41585);
nor U49644 (N_49644,N_40647,N_44115);
nor U49645 (N_49645,N_42826,N_44051);
nand U49646 (N_49646,N_43037,N_41931);
xnor U49647 (N_49647,N_41360,N_44978);
and U49648 (N_49648,N_41708,N_44514);
nand U49649 (N_49649,N_40644,N_43530);
or U49650 (N_49650,N_42575,N_41752);
or U49651 (N_49651,N_41228,N_40146);
and U49652 (N_49652,N_41716,N_40960);
nand U49653 (N_49653,N_43912,N_40888);
and U49654 (N_49654,N_41748,N_44192);
nand U49655 (N_49655,N_41951,N_40641);
and U49656 (N_49656,N_44791,N_43181);
nand U49657 (N_49657,N_42562,N_41503);
and U49658 (N_49658,N_44675,N_44265);
and U49659 (N_49659,N_44026,N_43225);
nand U49660 (N_49660,N_41997,N_41950);
xor U49661 (N_49661,N_41344,N_42698);
or U49662 (N_49662,N_41243,N_42102);
and U49663 (N_49663,N_40833,N_40176);
nand U49664 (N_49664,N_44650,N_40380);
nor U49665 (N_49665,N_44923,N_42221);
nor U49666 (N_49666,N_42483,N_41318);
xor U49667 (N_49667,N_41926,N_43636);
xor U49668 (N_49668,N_42878,N_44540);
or U49669 (N_49669,N_41885,N_40011);
xor U49670 (N_49670,N_43712,N_40073);
nor U49671 (N_49671,N_41821,N_40445);
or U49672 (N_49672,N_44980,N_44357);
nor U49673 (N_49673,N_43364,N_43855);
and U49674 (N_49674,N_44637,N_43152);
xor U49675 (N_49675,N_42041,N_40858);
xor U49676 (N_49676,N_41252,N_42433);
xnor U49677 (N_49677,N_44288,N_40510);
and U49678 (N_49678,N_43637,N_43628);
and U49679 (N_49679,N_42652,N_42486);
xor U49680 (N_49680,N_41954,N_44198);
xnor U49681 (N_49681,N_40511,N_41705);
nor U49682 (N_49682,N_43417,N_40338);
xnor U49683 (N_49683,N_42161,N_43825);
xnor U49684 (N_49684,N_44745,N_43658);
nor U49685 (N_49685,N_44039,N_43139);
and U49686 (N_49686,N_43507,N_44715);
nor U49687 (N_49687,N_43965,N_41229);
xnor U49688 (N_49688,N_44710,N_42509);
xor U49689 (N_49689,N_43735,N_43953);
nand U49690 (N_49690,N_44476,N_43299);
xor U49691 (N_49691,N_40746,N_40587);
nor U49692 (N_49692,N_42607,N_42420);
nand U49693 (N_49693,N_42721,N_43486);
nor U49694 (N_49694,N_42034,N_40682);
nor U49695 (N_49695,N_41534,N_41396);
xor U49696 (N_49696,N_43925,N_41623);
nand U49697 (N_49697,N_41022,N_44917);
nand U49698 (N_49698,N_40487,N_42666);
and U49699 (N_49699,N_41897,N_42995);
nor U49700 (N_49700,N_41036,N_42860);
xor U49701 (N_49701,N_41030,N_43133);
and U49702 (N_49702,N_44097,N_40422);
or U49703 (N_49703,N_42498,N_42150);
and U49704 (N_49704,N_40256,N_40142);
or U49705 (N_49705,N_41453,N_41865);
and U49706 (N_49706,N_43801,N_41021);
nand U49707 (N_49707,N_44091,N_42747);
nand U49708 (N_49708,N_44339,N_44123);
and U49709 (N_49709,N_41963,N_44033);
xnor U49710 (N_49710,N_40963,N_43782);
nor U49711 (N_49711,N_42797,N_41468);
nand U49712 (N_49712,N_43329,N_42619);
xnor U49713 (N_49713,N_41652,N_40297);
nor U49714 (N_49714,N_42057,N_42775);
or U49715 (N_49715,N_44300,N_42061);
nor U49716 (N_49716,N_40333,N_40733);
nand U49717 (N_49717,N_43643,N_43027);
and U49718 (N_49718,N_41790,N_42382);
xnor U49719 (N_49719,N_43569,N_40895);
xnor U49720 (N_49720,N_43649,N_43091);
xnor U49721 (N_49721,N_42557,N_40958);
or U49722 (N_49722,N_41537,N_41484);
and U49723 (N_49723,N_41801,N_41788);
xnor U49724 (N_49724,N_43046,N_44516);
or U49725 (N_49725,N_40954,N_40176);
nand U49726 (N_49726,N_44536,N_42500);
or U49727 (N_49727,N_41112,N_41617);
or U49728 (N_49728,N_40848,N_43218);
nor U49729 (N_49729,N_44459,N_44826);
nand U49730 (N_49730,N_40018,N_44990);
xnor U49731 (N_49731,N_40417,N_42818);
and U49732 (N_49732,N_43811,N_40929);
nand U49733 (N_49733,N_44217,N_40208);
nand U49734 (N_49734,N_40349,N_42040);
nand U49735 (N_49735,N_40696,N_42389);
nand U49736 (N_49736,N_44084,N_43209);
and U49737 (N_49737,N_42691,N_44894);
nor U49738 (N_49738,N_40209,N_43663);
xnor U49739 (N_49739,N_42311,N_44143);
xnor U49740 (N_49740,N_43986,N_40110);
xnor U49741 (N_49741,N_41162,N_44339);
and U49742 (N_49742,N_44303,N_41140);
nor U49743 (N_49743,N_42194,N_40155);
nor U49744 (N_49744,N_42553,N_42395);
nand U49745 (N_49745,N_44253,N_44649);
xnor U49746 (N_49746,N_41252,N_40154);
xor U49747 (N_49747,N_41446,N_43712);
xor U49748 (N_49748,N_44069,N_43887);
nor U49749 (N_49749,N_41763,N_40688);
nand U49750 (N_49750,N_42588,N_44753);
and U49751 (N_49751,N_42112,N_42430);
or U49752 (N_49752,N_41784,N_43431);
xor U49753 (N_49753,N_44282,N_43027);
and U49754 (N_49754,N_42367,N_42056);
or U49755 (N_49755,N_40796,N_40488);
nor U49756 (N_49756,N_41906,N_41776);
or U49757 (N_49757,N_44839,N_43585);
xnor U49758 (N_49758,N_44010,N_43432);
or U49759 (N_49759,N_44742,N_44026);
nor U49760 (N_49760,N_43720,N_41428);
or U49761 (N_49761,N_40061,N_40822);
xor U49762 (N_49762,N_41167,N_40946);
or U49763 (N_49763,N_44818,N_42264);
nand U49764 (N_49764,N_41937,N_43285);
or U49765 (N_49765,N_40935,N_42528);
nor U49766 (N_49766,N_40508,N_43967);
nand U49767 (N_49767,N_44689,N_44986);
nand U49768 (N_49768,N_43336,N_40625);
xor U49769 (N_49769,N_41489,N_41731);
or U49770 (N_49770,N_44720,N_43853);
nor U49771 (N_49771,N_43848,N_44966);
nor U49772 (N_49772,N_42457,N_44262);
nor U49773 (N_49773,N_41484,N_41281);
nor U49774 (N_49774,N_42069,N_44545);
or U49775 (N_49775,N_42454,N_40102);
nand U49776 (N_49776,N_44150,N_44786);
nand U49777 (N_49777,N_43056,N_41493);
nand U49778 (N_49778,N_40013,N_41382);
nor U49779 (N_49779,N_40073,N_44752);
nand U49780 (N_49780,N_42281,N_42248);
or U49781 (N_49781,N_42226,N_42249);
and U49782 (N_49782,N_43755,N_41415);
nor U49783 (N_49783,N_41240,N_42670);
or U49784 (N_49784,N_41907,N_43712);
and U49785 (N_49785,N_42557,N_44550);
and U49786 (N_49786,N_41555,N_41629);
nor U49787 (N_49787,N_41546,N_42447);
nand U49788 (N_49788,N_43605,N_41710);
nor U49789 (N_49789,N_44356,N_43087);
nand U49790 (N_49790,N_42307,N_43729);
and U49791 (N_49791,N_44074,N_43690);
or U49792 (N_49792,N_43703,N_44719);
and U49793 (N_49793,N_43113,N_40653);
and U49794 (N_49794,N_40221,N_43364);
nand U49795 (N_49795,N_40778,N_43145);
nor U49796 (N_49796,N_42101,N_43735);
or U49797 (N_49797,N_40577,N_43238);
xor U49798 (N_49798,N_44833,N_44877);
xor U49799 (N_49799,N_40403,N_44952);
nand U49800 (N_49800,N_44865,N_41279);
xor U49801 (N_49801,N_42347,N_42032);
or U49802 (N_49802,N_40209,N_40978);
nand U49803 (N_49803,N_44271,N_40792);
xnor U49804 (N_49804,N_44960,N_43876);
and U49805 (N_49805,N_43009,N_40331);
or U49806 (N_49806,N_42318,N_44725);
or U49807 (N_49807,N_41985,N_40872);
nand U49808 (N_49808,N_42951,N_44178);
nor U49809 (N_49809,N_42088,N_43400);
xor U49810 (N_49810,N_40750,N_44548);
and U49811 (N_49811,N_43970,N_40605);
and U49812 (N_49812,N_43808,N_40340);
nand U49813 (N_49813,N_42968,N_42458);
xnor U49814 (N_49814,N_44577,N_40278);
xnor U49815 (N_49815,N_41825,N_41263);
xor U49816 (N_49816,N_41241,N_42994);
nor U49817 (N_49817,N_40374,N_42069);
nor U49818 (N_49818,N_41650,N_40136);
xnor U49819 (N_49819,N_44127,N_43207);
and U49820 (N_49820,N_44139,N_40263);
or U49821 (N_49821,N_44439,N_44232);
nor U49822 (N_49822,N_43887,N_41619);
nand U49823 (N_49823,N_40576,N_44194);
nor U49824 (N_49824,N_41095,N_41673);
and U49825 (N_49825,N_42504,N_41349);
nand U49826 (N_49826,N_41667,N_43045);
nand U49827 (N_49827,N_44627,N_43051);
nor U49828 (N_49828,N_40103,N_43691);
or U49829 (N_49829,N_44737,N_44215);
nand U49830 (N_49830,N_41676,N_40188);
nand U49831 (N_49831,N_44171,N_41503);
nand U49832 (N_49832,N_41028,N_41887);
or U49833 (N_49833,N_44145,N_42815);
or U49834 (N_49834,N_41009,N_41138);
nand U49835 (N_49835,N_40705,N_44650);
or U49836 (N_49836,N_44140,N_43802);
and U49837 (N_49837,N_40662,N_44631);
and U49838 (N_49838,N_42983,N_41820);
nor U49839 (N_49839,N_42930,N_43610);
xnor U49840 (N_49840,N_43725,N_40093);
xor U49841 (N_49841,N_41370,N_42882);
and U49842 (N_49842,N_41089,N_43572);
or U49843 (N_49843,N_44563,N_44042);
and U49844 (N_49844,N_44308,N_40736);
or U49845 (N_49845,N_41456,N_44765);
nand U49846 (N_49846,N_44543,N_40032);
and U49847 (N_49847,N_42858,N_40983);
nor U49848 (N_49848,N_42292,N_43081);
or U49849 (N_49849,N_42748,N_40795);
nand U49850 (N_49850,N_41130,N_40865);
or U49851 (N_49851,N_43553,N_40182);
and U49852 (N_49852,N_44726,N_40805);
and U49853 (N_49853,N_40793,N_41721);
xor U49854 (N_49854,N_43137,N_41048);
and U49855 (N_49855,N_40926,N_41522);
or U49856 (N_49856,N_43881,N_40176);
or U49857 (N_49857,N_43826,N_44387);
or U49858 (N_49858,N_40550,N_41992);
nor U49859 (N_49859,N_44281,N_42022);
nor U49860 (N_49860,N_41903,N_43921);
nor U49861 (N_49861,N_43390,N_41196);
or U49862 (N_49862,N_44709,N_42031);
nor U49863 (N_49863,N_41941,N_44987);
nor U49864 (N_49864,N_40394,N_40035);
nand U49865 (N_49865,N_40322,N_43331);
nand U49866 (N_49866,N_43728,N_43798);
nand U49867 (N_49867,N_41048,N_40585);
nand U49868 (N_49868,N_44912,N_43644);
and U49869 (N_49869,N_42615,N_40666);
nor U49870 (N_49870,N_44037,N_43656);
xnor U49871 (N_49871,N_43713,N_42987);
or U49872 (N_49872,N_41247,N_43842);
or U49873 (N_49873,N_43859,N_42378);
nor U49874 (N_49874,N_43296,N_44447);
nor U49875 (N_49875,N_41608,N_44968);
and U49876 (N_49876,N_40523,N_41915);
or U49877 (N_49877,N_40393,N_44607);
and U49878 (N_49878,N_42307,N_40919);
nor U49879 (N_49879,N_44459,N_43278);
or U49880 (N_49880,N_42728,N_41378);
and U49881 (N_49881,N_44129,N_42083);
xor U49882 (N_49882,N_40279,N_42978);
or U49883 (N_49883,N_40427,N_41039);
and U49884 (N_49884,N_44708,N_41124);
and U49885 (N_49885,N_43078,N_44199);
nor U49886 (N_49886,N_41595,N_42970);
and U49887 (N_49887,N_42658,N_42842);
or U49888 (N_49888,N_41444,N_42837);
xor U49889 (N_49889,N_43592,N_43008);
nor U49890 (N_49890,N_40878,N_42705);
and U49891 (N_49891,N_41125,N_42382);
xnor U49892 (N_49892,N_42757,N_40498);
xor U49893 (N_49893,N_42031,N_43763);
nand U49894 (N_49894,N_44112,N_40023);
xor U49895 (N_49895,N_42761,N_41825);
nor U49896 (N_49896,N_40686,N_43589);
xnor U49897 (N_49897,N_42700,N_41542);
xnor U49898 (N_49898,N_44547,N_44404);
xnor U49899 (N_49899,N_40186,N_44412);
nor U49900 (N_49900,N_40157,N_44222);
or U49901 (N_49901,N_43283,N_42085);
and U49902 (N_49902,N_40339,N_41835);
xnor U49903 (N_49903,N_43603,N_43267);
nor U49904 (N_49904,N_44639,N_42113);
or U49905 (N_49905,N_41283,N_40273);
xnor U49906 (N_49906,N_43123,N_41745);
or U49907 (N_49907,N_40374,N_40494);
xnor U49908 (N_49908,N_41368,N_44906);
and U49909 (N_49909,N_41318,N_43528);
xnor U49910 (N_49910,N_41292,N_41209);
nand U49911 (N_49911,N_44400,N_43245);
nor U49912 (N_49912,N_44122,N_40961);
and U49913 (N_49913,N_41404,N_44269);
and U49914 (N_49914,N_43986,N_42878);
and U49915 (N_49915,N_40290,N_44501);
nand U49916 (N_49916,N_44917,N_44923);
nand U49917 (N_49917,N_43253,N_42583);
nor U49918 (N_49918,N_42209,N_42760);
nand U49919 (N_49919,N_41110,N_41252);
or U49920 (N_49920,N_43044,N_44270);
nand U49921 (N_49921,N_41618,N_44502);
nor U49922 (N_49922,N_42183,N_43834);
or U49923 (N_49923,N_44872,N_41874);
and U49924 (N_49924,N_40270,N_40340);
nand U49925 (N_49925,N_40157,N_41578);
nor U49926 (N_49926,N_44646,N_43252);
nor U49927 (N_49927,N_44117,N_41166);
nor U49928 (N_49928,N_44183,N_42352);
xnor U49929 (N_49929,N_41323,N_43993);
xor U49930 (N_49930,N_42616,N_44600);
nor U49931 (N_49931,N_42330,N_41241);
nand U49932 (N_49932,N_43296,N_44025);
nor U49933 (N_49933,N_40014,N_40837);
nor U49934 (N_49934,N_43890,N_44848);
and U49935 (N_49935,N_43997,N_44095);
nor U49936 (N_49936,N_43041,N_40918);
or U49937 (N_49937,N_44386,N_40267);
xnor U49938 (N_49938,N_43261,N_42272);
xor U49939 (N_49939,N_41852,N_44744);
nand U49940 (N_49940,N_43025,N_40185);
nor U49941 (N_49941,N_44832,N_40128);
nand U49942 (N_49942,N_43460,N_44524);
nor U49943 (N_49943,N_44996,N_41033);
nand U49944 (N_49944,N_42493,N_42557);
nand U49945 (N_49945,N_43677,N_40419);
xor U49946 (N_49946,N_43410,N_40221);
nand U49947 (N_49947,N_43710,N_43981);
nand U49948 (N_49948,N_42266,N_42991);
or U49949 (N_49949,N_44166,N_44557);
and U49950 (N_49950,N_42861,N_42758);
or U49951 (N_49951,N_42626,N_40636);
or U49952 (N_49952,N_42789,N_41508);
xnor U49953 (N_49953,N_42577,N_42654);
nor U49954 (N_49954,N_40334,N_41992);
nor U49955 (N_49955,N_42974,N_43325);
xnor U49956 (N_49956,N_42167,N_44006);
nor U49957 (N_49957,N_44576,N_42964);
and U49958 (N_49958,N_40572,N_43416);
and U49959 (N_49959,N_44652,N_41564);
nand U49960 (N_49960,N_42461,N_43507);
and U49961 (N_49961,N_40494,N_42491);
or U49962 (N_49962,N_44572,N_40801);
and U49963 (N_49963,N_43720,N_43926);
nand U49964 (N_49964,N_41088,N_43525);
and U49965 (N_49965,N_42754,N_42445);
xor U49966 (N_49966,N_42579,N_42614);
xnor U49967 (N_49967,N_44832,N_42841);
nand U49968 (N_49968,N_40202,N_43986);
nor U49969 (N_49969,N_43285,N_42612);
nand U49970 (N_49970,N_43819,N_44951);
nor U49971 (N_49971,N_40011,N_44423);
nor U49972 (N_49972,N_40314,N_40430);
and U49973 (N_49973,N_41282,N_42954);
or U49974 (N_49974,N_42721,N_43226);
nand U49975 (N_49975,N_42861,N_40893);
xor U49976 (N_49976,N_40463,N_42836);
nor U49977 (N_49977,N_42624,N_40272);
xor U49978 (N_49978,N_40021,N_44157);
or U49979 (N_49979,N_40565,N_40421);
nor U49980 (N_49980,N_42972,N_42097);
nand U49981 (N_49981,N_42822,N_42002);
xnor U49982 (N_49982,N_41195,N_41948);
nand U49983 (N_49983,N_41893,N_42525);
nor U49984 (N_49984,N_43034,N_43632);
xor U49985 (N_49985,N_40260,N_41563);
and U49986 (N_49986,N_40367,N_42692);
xnor U49987 (N_49987,N_42000,N_44767);
or U49988 (N_49988,N_44214,N_44107);
and U49989 (N_49989,N_44297,N_44782);
nor U49990 (N_49990,N_40965,N_41163);
and U49991 (N_49991,N_43390,N_44041);
and U49992 (N_49992,N_41196,N_43603);
xnor U49993 (N_49993,N_41852,N_44061);
or U49994 (N_49994,N_41674,N_40913);
nor U49995 (N_49995,N_42525,N_40474);
xnor U49996 (N_49996,N_41369,N_43592);
and U49997 (N_49997,N_40664,N_40526);
and U49998 (N_49998,N_42265,N_42212);
xnor U49999 (N_49999,N_44160,N_43546);
xor UO_0 (O_0,N_47461,N_48918);
nor UO_1 (O_1,N_45590,N_45530);
nor UO_2 (O_2,N_47626,N_49124);
xor UO_3 (O_3,N_46700,N_45688);
and UO_4 (O_4,N_46963,N_48207);
nor UO_5 (O_5,N_47121,N_47023);
or UO_6 (O_6,N_46585,N_48663);
xnor UO_7 (O_7,N_48622,N_48959);
and UO_8 (O_8,N_46240,N_47340);
or UO_9 (O_9,N_48670,N_48773);
or UO_10 (O_10,N_45242,N_48742);
or UO_11 (O_11,N_49704,N_49994);
or UO_12 (O_12,N_48493,N_47689);
and UO_13 (O_13,N_46468,N_49983);
nand UO_14 (O_14,N_46413,N_49791);
xor UO_15 (O_15,N_45396,N_45108);
and UO_16 (O_16,N_48549,N_45989);
or UO_17 (O_17,N_46673,N_48821);
and UO_18 (O_18,N_46458,N_49629);
nand UO_19 (O_19,N_46844,N_49497);
nor UO_20 (O_20,N_45320,N_48151);
or UO_21 (O_21,N_46698,N_47156);
nor UO_22 (O_22,N_46613,N_48180);
nor UO_23 (O_23,N_46017,N_46467);
and UO_24 (O_24,N_47552,N_47111);
or UO_25 (O_25,N_45425,N_49584);
nor UO_26 (O_26,N_45114,N_47840);
xor UO_27 (O_27,N_45604,N_47754);
and UO_28 (O_28,N_48417,N_46560);
nor UO_29 (O_29,N_47845,N_47183);
or UO_30 (O_30,N_45823,N_46184);
or UO_31 (O_31,N_45469,N_48406);
and UO_32 (O_32,N_45915,N_49128);
xor UO_33 (O_33,N_49831,N_46833);
or UO_34 (O_34,N_46480,N_48097);
or UO_35 (O_35,N_45283,N_46367);
and UO_36 (O_36,N_46397,N_46211);
or UO_37 (O_37,N_46845,N_48708);
and UO_38 (O_38,N_45843,N_49502);
and UO_39 (O_39,N_49751,N_45079);
and UO_40 (O_40,N_49323,N_49859);
and UO_41 (O_41,N_46869,N_47791);
nand UO_42 (O_42,N_45642,N_45326);
and UO_43 (O_43,N_47787,N_46427);
and UO_44 (O_44,N_46137,N_47057);
nand UO_45 (O_45,N_49238,N_48788);
xnor UO_46 (O_46,N_45875,N_45908);
or UO_47 (O_47,N_45676,N_47602);
or UO_48 (O_48,N_49771,N_45446);
nor UO_49 (O_49,N_48226,N_49800);
and UO_50 (O_50,N_49869,N_48601);
nand UO_51 (O_51,N_49550,N_46263);
nand UO_52 (O_52,N_45312,N_48771);
xnor UO_53 (O_53,N_48929,N_47694);
or UO_54 (O_54,N_49820,N_46054);
or UO_55 (O_55,N_45775,N_47661);
nor UO_56 (O_56,N_49273,N_48634);
nand UO_57 (O_57,N_46549,N_45551);
nor UO_58 (O_58,N_49557,N_48319);
xor UO_59 (O_59,N_49946,N_49554);
and UO_60 (O_60,N_49640,N_45541);
and UO_61 (O_61,N_45089,N_49900);
xor UO_62 (O_62,N_45390,N_46862);
or UO_63 (O_63,N_49190,N_46841);
nand UO_64 (O_64,N_46766,N_48184);
xor UO_65 (O_65,N_47529,N_47677);
or UO_66 (O_66,N_46260,N_48351);
xor UO_67 (O_67,N_48341,N_45923);
xnor UO_68 (O_68,N_49913,N_46813);
nor UO_69 (O_69,N_48290,N_46547);
and UO_70 (O_70,N_49438,N_45419);
and UO_71 (O_71,N_48761,N_47394);
and UO_72 (O_72,N_46393,N_45757);
and UO_73 (O_73,N_49740,N_46164);
or UO_74 (O_74,N_49732,N_47317);
nor UO_75 (O_75,N_49226,N_45005);
nor UO_76 (O_76,N_49218,N_46364);
and UO_77 (O_77,N_47707,N_47886);
nand UO_78 (O_78,N_47733,N_45076);
xnor UO_79 (O_79,N_48695,N_45494);
and UO_80 (O_80,N_49999,N_49018);
nand UO_81 (O_81,N_46569,N_45232);
xor UO_82 (O_82,N_47204,N_49169);
xor UO_83 (O_83,N_48669,N_49693);
nor UO_84 (O_84,N_47187,N_46695);
xnor UO_85 (O_85,N_47166,N_46207);
nand UO_86 (O_86,N_46274,N_45934);
nand UO_87 (O_87,N_49102,N_49283);
and UO_88 (O_88,N_49329,N_49464);
or UO_89 (O_89,N_48727,N_46190);
and UO_90 (O_90,N_45095,N_46471);
and UO_91 (O_91,N_49403,N_45481);
nand UO_92 (O_92,N_48537,N_46681);
nand UO_93 (O_93,N_46913,N_49523);
or UO_94 (O_94,N_48216,N_48912);
or UO_95 (O_95,N_48814,N_45796);
xor UO_96 (O_96,N_48600,N_46511);
nand UO_97 (O_97,N_49490,N_47700);
xnor UO_98 (O_98,N_49370,N_46677);
nand UO_99 (O_99,N_48352,N_49394);
nand UO_100 (O_100,N_46734,N_49798);
and UO_101 (O_101,N_47087,N_45547);
nand UO_102 (O_102,N_45834,N_45088);
xnor UO_103 (O_103,N_45714,N_47920);
and UO_104 (O_104,N_48135,N_48752);
or UO_105 (O_105,N_47100,N_45392);
and UO_106 (O_106,N_49970,N_47654);
or UO_107 (O_107,N_49173,N_47369);
nand UO_108 (O_108,N_45622,N_49929);
xnor UO_109 (O_109,N_48443,N_47022);
or UO_110 (O_110,N_46665,N_48222);
nor UO_111 (O_111,N_49980,N_45281);
xnor UO_112 (O_112,N_45080,N_47887);
and UO_113 (O_113,N_45240,N_49996);
and UO_114 (O_114,N_48577,N_46988);
and UO_115 (O_115,N_49690,N_48423);
or UO_116 (O_116,N_46252,N_48598);
nand UO_117 (O_117,N_48468,N_49585);
and UO_118 (O_118,N_45030,N_47199);
or UO_119 (O_119,N_48705,N_45962);
and UO_120 (O_120,N_48532,N_49728);
nand UO_121 (O_121,N_46842,N_46289);
nor UO_122 (O_122,N_48125,N_47160);
nand UO_123 (O_123,N_46118,N_45053);
nand UO_124 (O_124,N_47193,N_48426);
nand UO_125 (O_125,N_48115,N_46646);
or UO_126 (O_126,N_48697,N_48270);
nor UO_127 (O_127,N_46788,N_46243);
nand UO_128 (O_128,N_46902,N_47486);
xnor UO_129 (O_129,N_49140,N_49504);
xor UO_130 (O_130,N_48173,N_46683);
and UO_131 (O_131,N_49434,N_46120);
nand UO_132 (O_132,N_45776,N_46564);
nand UO_133 (O_133,N_47447,N_46571);
nor UO_134 (O_134,N_45206,N_45637);
or UO_135 (O_135,N_45580,N_48466);
nand UO_136 (O_136,N_48242,N_47641);
and UO_137 (O_137,N_45851,N_47348);
and UO_138 (O_138,N_46708,N_47370);
xor UO_139 (O_139,N_45857,N_45701);
or UO_140 (O_140,N_45393,N_47083);
and UO_141 (O_141,N_47667,N_46326);
or UO_142 (O_142,N_49953,N_49799);
nand UO_143 (O_143,N_49042,N_47969);
and UO_144 (O_144,N_46702,N_49269);
or UO_145 (O_145,N_49471,N_49565);
xnor UO_146 (O_146,N_47429,N_46524);
xor UO_147 (O_147,N_45485,N_49427);
and UO_148 (O_148,N_49902,N_48172);
nand UO_149 (O_149,N_49657,N_49308);
xor UO_150 (O_150,N_48344,N_47567);
nand UO_151 (O_151,N_49944,N_47477);
and UO_152 (O_152,N_46596,N_49373);
nand UO_153 (O_153,N_46155,N_45391);
xnor UO_154 (O_154,N_45606,N_48256);
nand UO_155 (O_155,N_47028,N_45286);
nor UO_156 (O_156,N_47625,N_49883);
nor UO_157 (O_157,N_45598,N_48595);
nand UO_158 (O_158,N_48698,N_48220);
or UO_159 (O_159,N_46610,N_49296);
xnor UO_160 (O_160,N_47851,N_47263);
nand UO_161 (O_161,N_46238,N_47511);
xor UO_162 (O_162,N_48690,N_48464);
nor UO_163 (O_163,N_47206,N_47467);
nor UO_164 (O_164,N_49611,N_46691);
and UO_165 (O_165,N_45723,N_46738);
or UO_166 (O_166,N_48396,N_49223);
xnor UO_167 (O_167,N_47118,N_48283);
nor UO_168 (O_168,N_49833,N_48413);
or UO_169 (O_169,N_47462,N_49749);
nand UO_170 (O_170,N_47926,N_47381);
nor UO_171 (O_171,N_47101,N_49166);
and UO_172 (O_172,N_46023,N_45204);
nand UO_173 (O_173,N_45815,N_47765);
or UO_174 (O_174,N_45090,N_49162);
nor UO_175 (O_175,N_49267,N_46523);
nand UO_176 (O_176,N_46705,N_49988);
or UO_177 (O_177,N_45929,N_48904);
nor UO_178 (O_178,N_46457,N_46945);
and UO_179 (O_179,N_48185,N_47088);
and UO_180 (O_180,N_45795,N_49627);
nand UO_181 (O_181,N_45837,N_45895);
and UO_182 (O_182,N_47656,N_46455);
xor UO_183 (O_183,N_47725,N_45236);
and UO_184 (O_184,N_46772,N_48903);
nand UO_185 (O_185,N_47908,N_47227);
or UO_186 (O_186,N_46218,N_46215);
and UO_187 (O_187,N_46386,N_47323);
nand UO_188 (O_188,N_48093,N_48853);
and UO_189 (O_189,N_48559,N_45996);
xor UO_190 (O_190,N_47863,N_48524);
nor UO_191 (O_191,N_45632,N_47616);
or UO_192 (O_192,N_49286,N_49915);
nand UO_193 (O_193,N_48244,N_49463);
xnor UO_194 (O_194,N_48806,N_46831);
nor UO_195 (O_195,N_45174,N_45129);
and UO_196 (O_196,N_45615,N_47386);
xnor UO_197 (O_197,N_49414,N_45533);
nand UO_198 (O_198,N_47113,N_46855);
nand UO_199 (O_199,N_45462,N_45522);
nand UO_200 (O_200,N_47294,N_46961);
or UO_201 (O_201,N_45133,N_47251);
nand UO_202 (O_202,N_48069,N_45909);
or UO_203 (O_203,N_47195,N_48931);
xor UO_204 (O_204,N_48016,N_48816);
nor UO_205 (O_205,N_48593,N_45683);
or UO_206 (O_206,N_45461,N_48714);
nor UO_207 (O_207,N_46509,N_48123);
xnor UO_208 (O_208,N_49802,N_45715);
nor UO_209 (O_209,N_48612,N_46548);
or UO_210 (O_210,N_47321,N_49577);
nor UO_211 (O_211,N_48741,N_45704);
xor UO_212 (O_212,N_48512,N_47419);
nor UO_213 (O_213,N_48022,N_46892);
or UO_214 (O_214,N_48334,N_47893);
or UO_215 (O_215,N_46601,N_47871);
nor UO_216 (O_216,N_48001,N_45948);
or UO_217 (O_217,N_49251,N_45060);
nor UO_218 (O_218,N_45819,N_48840);
nor UO_219 (O_219,N_47485,N_46929);
or UO_220 (O_220,N_46608,N_46958);
or UO_221 (O_221,N_45488,N_49816);
or UO_222 (O_222,N_45428,N_45433);
and UO_223 (O_223,N_49422,N_46568);
nor UO_224 (O_224,N_48322,N_49324);
or UO_225 (O_225,N_48553,N_46586);
nor UO_226 (O_226,N_46345,N_46553);
or UO_227 (O_227,N_49404,N_48178);
and UO_228 (O_228,N_48809,N_48602);
nor UO_229 (O_229,N_46410,N_49663);
and UO_230 (O_230,N_45557,N_46246);
nand UO_231 (O_231,N_49266,N_49193);
nand UO_232 (O_232,N_45262,N_47001);
or UO_233 (O_233,N_48040,N_45781);
nor UO_234 (O_234,N_45453,N_48101);
or UO_235 (O_235,N_45752,N_49770);
nor UO_236 (O_236,N_49436,N_48990);
nor UO_237 (O_237,N_46755,N_45142);
and UO_238 (O_238,N_45051,N_45324);
xnor UO_239 (O_239,N_49142,N_45317);
or UO_240 (O_240,N_48041,N_49048);
or UO_241 (O_241,N_47766,N_45057);
xnor UO_242 (O_242,N_48848,N_45859);
xor UO_243 (O_243,N_47012,N_49756);
or UO_244 (O_244,N_49753,N_48203);
nand UO_245 (O_245,N_45542,N_49220);
nand UO_246 (O_246,N_46461,N_46031);
nand UO_247 (O_247,N_48960,N_48765);
nor UO_248 (O_248,N_46911,N_48150);
nand UO_249 (O_249,N_46329,N_46485);
nand UO_250 (O_250,N_49551,N_45917);
nand UO_251 (O_251,N_49790,N_49315);
nand UO_252 (O_252,N_49846,N_45639);
or UO_253 (O_253,N_45046,N_45126);
xor UO_254 (O_254,N_46948,N_48868);
xnor UO_255 (O_255,N_45071,N_45749);
xnor UO_256 (O_256,N_49407,N_45650);
or UO_257 (O_257,N_47723,N_49121);
nand UO_258 (O_258,N_47789,N_49104);
xnor UO_259 (O_259,N_49393,N_45944);
nor UO_260 (O_260,N_46998,N_49651);
and UO_261 (O_261,N_49194,N_49763);
xnor UO_262 (O_262,N_46394,N_47997);
xor UO_263 (O_263,N_47421,N_47412);
nor UO_264 (O_264,N_45573,N_49325);
and UO_265 (O_265,N_45018,N_47049);
nor UO_266 (O_266,N_49467,N_49845);
xor UO_267 (O_267,N_46332,N_45685);
xor UO_268 (O_268,N_46498,N_48358);
xor UO_269 (O_269,N_49090,N_47438);
or UO_270 (O_270,N_47543,N_47579);
and UO_271 (O_271,N_46968,N_45986);
and UO_272 (O_272,N_48120,N_45282);
nor UO_273 (O_273,N_48228,N_46551);
and UO_274 (O_274,N_45828,N_47705);
xor UO_275 (O_275,N_47962,N_49475);
nand UO_276 (O_276,N_48521,N_49503);
or UO_277 (O_277,N_48709,N_48455);
nor UO_278 (O_278,N_45487,N_48168);
and UO_279 (O_279,N_46850,N_47722);
nor UO_280 (O_280,N_49524,N_45531);
or UO_281 (O_281,N_46521,N_49012);
xor UO_282 (O_282,N_48935,N_48199);
nor UO_283 (O_283,N_46133,N_45904);
nand UO_284 (O_284,N_45212,N_49945);
xor UO_285 (O_285,N_46465,N_47141);
xor UO_286 (O_286,N_46436,N_47878);
or UO_287 (O_287,N_49884,N_49950);
nor UO_288 (O_288,N_45896,N_47210);
nor UO_289 (O_289,N_48003,N_45653);
and UO_290 (O_290,N_48643,N_47937);
nand UO_291 (O_291,N_47152,N_46769);
or UO_292 (O_292,N_48749,N_48425);
or UO_293 (O_293,N_48099,N_47054);
nand UO_294 (O_294,N_47663,N_47848);
and UO_295 (O_295,N_48673,N_49256);
and UO_296 (O_296,N_49293,N_45926);
xnor UO_297 (O_297,N_46007,N_46213);
xor UO_298 (O_298,N_49781,N_49589);
and UO_299 (O_299,N_46527,N_48649);
nor UO_300 (O_300,N_47856,N_46113);
nand UO_301 (O_301,N_46905,N_49113);
and UO_302 (O_302,N_49973,N_46577);
and UO_303 (O_303,N_47683,N_49862);
and UO_304 (O_304,N_47885,N_48143);
or UO_305 (O_305,N_45786,N_48900);
or UO_306 (O_306,N_49865,N_47933);
nand UO_307 (O_307,N_48799,N_49499);
and UO_308 (O_308,N_46982,N_46550);
and UO_309 (O_309,N_49303,N_48176);
xnor UO_310 (O_310,N_46136,N_45938);
or UO_311 (O_311,N_46774,N_48288);
and UO_312 (O_312,N_48039,N_46489);
or UO_313 (O_313,N_48954,N_49610);
xor UO_314 (O_314,N_45406,N_45307);
and UO_315 (O_315,N_49962,N_49553);
nor UO_316 (O_316,N_48688,N_48488);
nor UO_317 (O_317,N_45864,N_47671);
xnor UO_318 (O_318,N_48791,N_47617);
or UO_319 (O_319,N_45357,N_45400);
and UO_320 (O_320,N_45273,N_48144);
and UO_321 (O_321,N_47105,N_47319);
nand UO_322 (O_322,N_48635,N_46976);
nor UO_323 (O_323,N_45678,N_49138);
or UO_324 (O_324,N_48102,N_46098);
and UO_325 (O_325,N_45261,N_49453);
nor UO_326 (O_326,N_45624,N_45093);
and UO_327 (O_327,N_46300,N_48543);
or UO_328 (O_328,N_46668,N_49998);
or UO_329 (O_329,N_48972,N_49832);
nor UO_330 (O_330,N_45736,N_46490);
or UO_331 (O_331,N_45742,N_48261);
nor UO_332 (O_332,N_49575,N_49607);
xor UO_333 (O_333,N_49019,N_48699);
nor UO_334 (O_334,N_48734,N_45176);
or UO_335 (O_335,N_45011,N_45395);
nor UO_336 (O_336,N_48025,N_46327);
xnor UO_337 (O_337,N_49892,N_48470);
xnor UO_338 (O_338,N_48497,N_47495);
or UO_339 (O_339,N_49175,N_49713);
and UO_340 (O_340,N_46811,N_48564);
and UO_341 (O_341,N_46714,N_46004);
xor UO_342 (O_342,N_46875,N_48641);
xnor UO_343 (O_343,N_48760,N_48487);
nand UO_344 (O_344,N_47644,N_47060);
nand UO_345 (O_345,N_47795,N_45841);
xor UO_346 (O_346,N_46124,N_46058);
and UO_347 (O_347,N_48640,N_46709);
nor UO_348 (O_348,N_49880,N_45385);
nand UO_349 (O_349,N_45062,N_49197);
nor UO_350 (O_350,N_45849,N_48519);
nor UO_351 (O_351,N_47307,N_46930);
or UO_352 (O_352,N_49857,N_49876);
xor UO_353 (O_353,N_48296,N_46390);
and UO_354 (O_354,N_45706,N_45569);
nand UO_355 (O_355,N_45459,N_45913);
nor UO_356 (O_356,N_47464,N_47653);
nand UO_357 (O_357,N_47454,N_46180);
nor UO_358 (O_358,N_48711,N_46801);
xnor UO_359 (O_359,N_47629,N_47925);
or UO_360 (O_360,N_46226,N_48006);
nor UO_361 (O_361,N_45496,N_46776);
xnor UO_362 (O_362,N_48354,N_46105);
nor UO_363 (O_363,N_47961,N_46254);
xnor UO_364 (O_364,N_48234,N_49001);
or UO_365 (O_365,N_45305,N_49420);
nor UO_366 (O_366,N_48626,N_48617);
xor UO_367 (O_367,N_46227,N_49509);
or UO_368 (O_368,N_47416,N_49240);
and UO_369 (O_369,N_45972,N_49347);
or UO_370 (O_370,N_45415,N_48273);
nand UO_371 (O_371,N_48980,N_49181);
nand UO_372 (O_372,N_45656,N_47713);
and UO_373 (O_373,N_47959,N_47506);
or UO_374 (O_374,N_45198,N_47696);
xor UO_375 (O_375,N_48850,N_48380);
and UO_376 (O_376,N_47011,N_48755);
nor UO_377 (O_377,N_48205,N_49446);
nand UO_378 (O_378,N_49045,N_48177);
and UO_379 (O_379,N_45945,N_47426);
nand UO_380 (O_380,N_46060,N_48611);
and UO_381 (O_381,N_47342,N_48398);
nand UO_382 (O_382,N_45903,N_45409);
nand UO_383 (O_383,N_47786,N_45719);
nor UO_384 (O_384,N_48561,N_49054);
and UO_385 (O_385,N_45431,N_45291);
nand UO_386 (O_386,N_46526,N_46572);
nand UO_387 (O_387,N_47245,N_48431);
xor UO_388 (O_388,N_48271,N_49289);
nor UO_389 (O_389,N_48299,N_46672);
xnor UO_390 (O_390,N_49033,N_49648);
and UO_391 (O_391,N_49738,N_48362);
or UO_392 (O_392,N_49047,N_45922);
xnor UO_393 (O_393,N_47332,N_46411);
nand UO_394 (O_394,N_48179,N_47746);
xnor UO_395 (O_395,N_45657,N_45184);
xor UO_396 (O_396,N_45545,N_45366);
nor UO_397 (O_397,N_47433,N_45028);
and UO_398 (O_398,N_46018,N_47799);
nor UO_399 (O_399,N_48893,N_49606);
and UO_400 (O_400,N_49505,N_46114);
nand UO_401 (O_401,N_49765,N_48579);
and UO_402 (O_402,N_45652,N_49792);
or UO_403 (O_403,N_46232,N_49873);
nor UO_404 (O_404,N_48324,N_46671);
nand UO_405 (O_405,N_49914,N_48977);
or UO_406 (O_406,N_45684,N_45422);
or UO_407 (O_407,N_49199,N_48565);
nand UO_408 (O_408,N_47510,N_46804);
nor UO_409 (O_409,N_45550,N_47747);
or UO_410 (O_410,N_45585,N_46981);
xnor UO_411 (O_411,N_45073,N_46093);
nand UO_412 (O_412,N_48769,N_46659);
nor UO_413 (O_413,N_46581,N_46219);
xnor UO_414 (O_414,N_48349,N_49890);
and UO_415 (O_415,N_46003,N_49722);
or UO_416 (O_416,N_45616,N_49928);
xnor UO_417 (O_417,N_45003,N_49797);
and UO_418 (O_418,N_45768,N_46535);
xor UO_419 (O_419,N_48333,N_49815);
nor UO_420 (O_420,N_45423,N_45925);
xor UO_421 (O_421,N_46951,N_47796);
nand UO_422 (O_422,N_46142,N_49419);
xor UO_423 (O_423,N_49384,N_48851);
or UO_424 (O_424,N_45118,N_46309);
and UO_425 (O_425,N_47286,N_48766);
xnor UO_426 (O_426,N_47546,N_47181);
and UO_427 (O_427,N_47640,N_45158);
xnor UO_428 (O_428,N_49624,N_46638);
nand UO_429 (O_429,N_49547,N_47344);
nand UO_430 (O_430,N_48817,N_47624);
and UO_431 (O_431,N_45765,N_49094);
or UO_432 (O_432,N_49059,N_49496);
or UO_433 (O_433,N_47605,N_46100);
nand UO_434 (O_434,N_46991,N_47079);
nor UO_435 (O_435,N_49260,N_49236);
nor UO_436 (O_436,N_49445,N_47117);
or UO_437 (O_437,N_49954,N_49602);
xor UO_438 (O_438,N_47164,N_45734);
nand UO_439 (O_439,N_49634,N_48326);
xnor UO_440 (O_440,N_45112,N_48831);
and UO_441 (O_441,N_46615,N_49435);
or UO_442 (O_442,N_48668,N_49081);
xor UO_443 (O_443,N_49562,N_49424);
nor UO_444 (O_444,N_46944,N_46270);
and UO_445 (O_445,N_49948,N_49110);
nor UO_446 (O_446,N_46858,N_46786);
or UO_447 (O_447,N_45523,N_48278);
and UO_448 (O_448,N_47979,N_49000);
nor UO_449 (O_449,N_45601,N_48862);
xor UO_450 (O_450,N_47531,N_46771);
xor UO_451 (O_451,N_47544,N_46474);
xor UO_452 (O_452,N_47378,N_49935);
and UO_453 (O_453,N_48841,N_49357);
xor UO_454 (O_454,N_46820,N_47923);
and UO_455 (O_455,N_48592,N_49824);
and UO_456 (O_456,N_45789,N_46194);
or UO_457 (O_457,N_48282,N_49255);
nor UO_458 (O_458,N_47360,N_46592);
or UO_459 (O_459,N_47649,N_45477);
xor UO_460 (O_460,N_46294,N_46200);
or UO_461 (O_461,N_48857,N_45049);
nand UO_462 (O_462,N_49292,N_47016);
and UO_463 (O_463,N_47666,N_45119);
and UO_464 (O_464,N_47226,N_49055);
and UO_465 (O_465,N_49895,N_47398);
xnor UO_466 (O_466,N_45069,N_49346);
xor UO_467 (O_467,N_49991,N_49769);
nor UO_468 (O_468,N_48979,N_46293);
or UO_469 (O_469,N_45452,N_47932);
nor UO_470 (O_470,N_49363,N_45166);
xnor UO_471 (O_471,N_46836,N_45480);
and UO_472 (O_472,N_45006,N_46873);
and UO_473 (O_473,N_49084,N_49743);
or UO_474 (O_474,N_47738,N_46385);
nor UO_475 (O_475,N_49030,N_48818);
xor UO_476 (O_476,N_46459,N_47545);
and UO_477 (O_477,N_47614,N_48531);
xor UO_478 (O_478,N_46157,N_47623);
or UO_479 (O_479,N_48489,N_47651);
and UO_480 (O_480,N_49655,N_46039);
or UO_481 (O_481,N_47445,N_48939);
or UO_482 (O_482,N_46637,N_45790);
and UO_483 (O_483,N_49608,N_45912);
or UO_484 (O_484,N_49708,N_47478);
nand UO_485 (O_485,N_49391,N_47777);
nor UO_486 (O_486,N_48061,N_48390);
xnor UO_487 (O_487,N_47114,N_46123);
or UO_488 (O_488,N_47424,N_48810);
and UO_489 (O_489,N_47482,N_47870);
nor UO_490 (O_490,N_48169,N_46111);
or UO_491 (O_491,N_46422,N_48786);
nand UO_492 (O_492,N_48891,N_45732);
xnor UO_493 (O_493,N_45337,N_49702);
nand UO_494 (O_494,N_46049,N_45023);
xnor UO_495 (O_495,N_47442,N_48887);
or UO_496 (O_496,N_48528,N_46880);
nand UO_497 (O_497,N_46384,N_47414);
xor UO_498 (O_498,N_46777,N_45941);
and UO_499 (O_499,N_49480,N_46896);
xor UO_500 (O_500,N_49697,N_46380);
and UO_501 (O_501,N_49894,N_49261);
and UO_502 (O_502,N_46570,N_49159);
nor UO_503 (O_503,N_48262,N_47185);
nand UO_504 (O_504,N_49801,N_46282);
and UO_505 (O_505,N_46351,N_47231);
nand UO_506 (O_506,N_47588,N_46445);
or UO_507 (O_507,N_49461,N_48490);
and UO_508 (O_508,N_45429,N_49560);
nand UO_509 (O_509,N_45239,N_45370);
nor UO_510 (O_510,N_48174,N_48925);
xnor UO_511 (O_511,N_48745,N_49126);
nor UO_512 (O_512,N_49443,N_46980);
or UO_513 (O_513,N_48127,N_48439);
nor UO_514 (O_514,N_48546,N_45666);
nor UO_515 (O_515,N_48801,N_45867);
or UO_516 (O_516,N_46383,N_46567);
xnor UO_517 (O_517,N_47712,N_47382);
nor UO_518 (O_518,N_48042,N_48189);
xnor UO_519 (O_519,N_49432,N_46085);
and UO_520 (O_520,N_45321,N_45380);
nor UO_521 (O_521,N_46633,N_47264);
or UO_522 (O_522,N_47618,N_46995);
and UO_523 (O_523,N_45227,N_49654);
or UO_524 (O_524,N_48357,N_47299);
xnor UO_525 (O_525,N_49671,N_48967);
nor UO_526 (O_526,N_49112,N_47405);
or UO_527 (O_527,N_49320,N_47201);
nand UO_528 (O_528,N_48442,N_49850);
or UO_529 (O_529,N_49353,N_49211);
nor UO_530 (O_530,N_49636,N_46767);
nand UO_531 (O_531,N_47560,N_46106);
and UO_532 (O_532,N_47167,N_46794);
or UO_533 (O_533,N_47583,N_46275);
nand UO_534 (O_534,N_46584,N_47917);
or UO_535 (O_535,N_49448,N_46466);
nand UO_536 (O_536,N_45361,N_49851);
nor UO_537 (O_537,N_45362,N_47293);
nor UO_538 (O_538,N_49487,N_48767);
or UO_539 (O_539,N_46301,N_45157);
and UO_540 (O_540,N_48436,N_47688);
nor UO_541 (O_541,N_49525,N_46904);
or UO_542 (O_542,N_46887,N_46362);
xnor UO_543 (O_543,N_45460,N_46149);
or UO_544 (O_544,N_48573,N_49037);
nand UO_545 (O_545,N_48539,N_45478);
and UO_546 (O_546,N_47635,N_48630);
nor UO_547 (O_547,N_45677,N_47981);
nand UO_548 (O_548,N_48676,N_48860);
nand UO_549 (O_549,N_49684,N_46096);
nand UO_550 (O_550,N_46392,N_49013);
nand UO_551 (O_551,N_45990,N_45196);
and UO_552 (O_552,N_47243,N_45644);
nor UO_553 (O_553,N_46224,N_45091);
nand UO_554 (O_554,N_47250,N_46248);
nand UO_555 (O_555,N_47960,N_47928);
or UO_556 (O_556,N_46652,N_48508);
or UO_557 (O_557,N_47620,N_48913);
nand UO_558 (O_558,N_46525,N_49041);
nand UO_559 (O_559,N_47000,N_48569);
nor UO_560 (O_560,N_46235,N_47776);
nor UO_561 (O_561,N_48807,N_48057);
nor UO_562 (O_562,N_46505,N_48447);
or UO_563 (O_563,N_46907,N_47826);
and UO_564 (O_564,N_49978,N_46834);
and UO_565 (O_565,N_48066,N_48429);
and UO_566 (O_566,N_49343,N_47335);
xor UO_567 (O_567,N_47408,N_49248);
xor UO_568 (O_568,N_47337,N_48392);
or UO_569 (O_569,N_46070,N_45309);
nand UO_570 (O_570,N_49568,N_47867);
xnor UO_571 (O_571,N_47711,N_46281);
and UO_572 (O_572,N_45136,N_46073);
xor UO_573 (O_573,N_46233,N_48772);
nor UO_574 (O_574,N_49896,N_45365);
xor UO_575 (O_575,N_45332,N_49745);
nor UO_576 (O_576,N_47728,N_48133);
and UO_577 (O_577,N_46736,N_47968);
or UO_578 (O_578,N_46756,N_46437);
or UO_579 (O_579,N_47736,N_48502);
and UO_580 (O_580,N_47341,N_48196);
nor UO_581 (O_581,N_46969,N_46996);
nand UO_582 (O_582,N_45581,N_45575);
xor UO_583 (O_583,N_45764,N_47377);
or UO_584 (O_584,N_47994,N_48215);
nand UO_585 (O_585,N_45618,N_46175);
nor UO_586 (O_586,N_48335,N_47333);
nand UO_587 (O_587,N_45975,N_49116);
or UO_588 (O_588,N_49355,N_46439);
or UO_589 (O_589,N_45663,N_48775);
and UO_590 (O_590,N_46205,N_45214);
and UO_591 (O_591,N_49328,N_47300);
xnor UO_592 (O_592,N_47349,N_45186);
nor UO_593 (O_593,N_45504,N_47275);
nor UO_594 (O_594,N_47732,N_49049);
and UO_595 (O_595,N_49483,N_49155);
or UO_596 (O_596,N_48212,N_47374);
and UO_597 (O_597,N_45560,N_49096);
or UO_598 (O_598,N_48155,N_49349);
or UO_599 (O_599,N_49115,N_46261);
nand UO_600 (O_600,N_46236,N_48474);
and UO_601 (O_601,N_45448,N_48846);
nand UO_602 (O_602,N_46312,N_49586);
xnor UO_603 (O_603,N_47475,N_47180);
and UO_604 (O_604,N_48784,N_48963);
nand UO_605 (O_605,N_45132,N_48735);
and UO_606 (O_606,N_46623,N_48415);
nand UO_607 (O_607,N_49867,N_46122);
or UO_608 (O_608,N_46130,N_47458);
or UO_609 (O_609,N_46375,N_48405);
and UO_610 (O_610,N_49887,N_47082);
and UO_611 (O_611,N_46582,N_48370);
or UO_612 (O_612,N_47490,N_46322);
nand UO_613 (O_613,N_45424,N_49474);
nor UO_614 (O_614,N_46324,N_48359);
nand UO_615 (O_615,N_45032,N_49158);
xnor UO_616 (O_616,N_48616,N_47566);
or UO_617 (O_617,N_48233,N_46278);
or UO_618 (O_618,N_48572,N_45194);
xnor UO_619 (O_619,N_47107,N_46292);
nor UO_620 (O_620,N_47480,N_47026);
xor UO_621 (O_621,N_46746,N_47717);
and UO_622 (O_622,N_45279,N_46782);
nor UO_623 (O_623,N_49556,N_46650);
nand UO_624 (O_624,N_45347,N_45479);
or UO_625 (O_625,N_45100,N_47784);
or UO_626 (O_626,N_47190,N_47946);
and UO_627 (O_627,N_47296,N_46593);
and UO_628 (O_628,N_46165,N_47368);
and UO_629 (O_629,N_45189,N_47200);
nor UO_630 (O_630,N_48496,N_49167);
nor UO_631 (O_631,N_45682,N_49053);
xnor UO_632 (O_632,N_48293,N_48917);
nor UO_633 (O_633,N_45943,N_49078);
xor UO_634 (O_634,N_47238,N_45787);
nor UO_635 (O_635,N_47843,N_46670);
nor UO_636 (O_636,N_48833,N_46022);
nand UO_637 (O_637,N_45009,N_46162);
or UO_638 (O_638,N_45179,N_49130);
xnor UO_639 (O_639,N_49536,N_47450);
and UO_640 (O_640,N_49027,N_48768);
nor UO_641 (O_641,N_46420,N_49390);
or UO_642 (O_642,N_45304,N_48441);
xnor UO_643 (O_643,N_45507,N_48435);
xnor UO_644 (O_644,N_48973,N_46654);
xnor UO_645 (O_645,N_47155,N_45457);
nand UO_646 (O_646,N_49511,N_47730);
nand UO_647 (O_647,N_47757,N_49596);
or UO_648 (O_648,N_49559,N_47785);
nor UO_649 (O_649,N_45082,N_47965);
and UO_650 (O_650,N_49982,N_46288);
nand UO_651 (O_651,N_47033,N_47045);
xor UO_652 (O_652,N_49280,N_45296);
and UO_653 (O_653,N_45510,N_47865);
or UO_654 (O_654,N_47557,N_48389);
or UO_655 (O_655,N_45092,N_45255);
nand UO_656 (O_656,N_48842,N_45329);
xnor UO_657 (O_657,N_48328,N_48660);
nor UO_658 (O_658,N_46790,N_48899);
nor UO_659 (O_659,N_47389,N_47315);
xor UO_660 (O_660,N_48535,N_48654);
and UO_661 (O_661,N_47638,N_49603);
nor UO_662 (O_662,N_45113,N_46078);
nand UO_663 (O_663,N_48107,N_46796);
nand UO_664 (O_664,N_45427,N_47993);
or UO_665 (O_665,N_48088,N_49604);
xnor UO_666 (O_666,N_49495,N_48247);
nor UO_667 (O_667,N_47385,N_48249);
and UO_668 (O_668,N_47423,N_49295);
xor UO_669 (O_669,N_49905,N_45414);
nand UO_670 (O_670,N_45839,N_49829);
nor UO_671 (O_671,N_47555,N_45489);
nor UO_672 (O_672,N_49118,N_45000);
nor UO_673 (O_673,N_48753,N_49760);
xnor UO_674 (O_674,N_49091,N_49062);
nand UO_675 (O_675,N_48938,N_48725);
nand UO_676 (O_676,N_48619,N_49729);
nor UO_677 (O_677,N_45952,N_47830);
and UO_678 (O_678,N_47985,N_48346);
nand UO_679 (O_679,N_49965,N_48316);
nor UO_680 (O_680,N_45634,N_46464);
xor UO_681 (O_681,N_47686,N_46852);
nor UO_682 (O_682,N_46960,N_48412);
or UO_683 (O_683,N_47343,N_48424);
and UO_684 (O_684,N_48756,N_47077);
or UO_685 (O_685,N_46908,N_49380);
nor UO_686 (O_686,N_48732,N_47948);
xnor UO_687 (O_687,N_47876,N_48192);
xnor UO_688 (O_688,N_48780,N_48175);
nand UO_689 (O_689,N_47310,N_48055);
xor UO_690 (O_690,N_48200,N_49541);
nor UO_691 (O_691,N_45936,N_46475);
nand UO_692 (O_692,N_45906,N_45873);
and UO_693 (O_693,N_45643,N_48075);
nor UO_694 (O_694,N_47999,N_49400);
nand UO_695 (O_695,N_46762,N_48030);
xnor UO_696 (O_696,N_48432,N_48047);
nor UO_697 (O_697,N_49964,N_45065);
nand UO_698 (O_698,N_46011,N_46406);
and UO_699 (O_699,N_48473,N_45253);
xnor UO_700 (O_700,N_47103,N_47846);
xor UO_701 (O_701,N_48751,N_45763);
nor UO_702 (O_702,N_49309,N_49189);
xor UO_703 (O_703,N_48008,N_49847);
or UO_704 (O_704,N_48149,N_48897);
nand UO_705 (O_705,N_46803,N_48353);
or UO_706 (O_706,N_47684,N_45193);
and UO_707 (O_707,N_48504,N_49938);
nand UO_708 (O_708,N_49827,N_46494);
or UO_709 (O_709,N_45201,N_47483);
nor UO_710 (O_710,N_47248,N_48907);
and UO_711 (O_711,N_47809,N_46516);
xnor UO_712 (O_712,N_47133,N_48560);
or UO_713 (O_713,N_47207,N_47896);
xor UO_714 (O_714,N_46829,N_49848);
nor UO_715 (O_715,N_45835,N_45609);
or UO_716 (O_716,N_46528,N_47473);
and UO_717 (O_717,N_48253,N_47030);
and UO_718 (O_718,N_46843,N_46050);
xnor UO_719 (O_719,N_46757,N_47570);
xnor UO_720 (O_720,N_48461,N_45600);
and UO_721 (O_721,N_49592,N_49593);
xnor UO_722 (O_722,N_47236,N_47607);
nand UO_723 (O_723,N_49339,N_45980);
or UO_724 (O_724,N_46075,N_48924);
nand UO_725 (O_725,N_49061,N_47756);
or UO_726 (O_726,N_45024,N_49725);
xnor UO_727 (O_727,N_45451,N_46876);
and UO_728 (O_728,N_46627,N_47710);
xnor UO_729 (O_729,N_46617,N_47119);
or UO_730 (O_730,N_45853,N_47675);
and UO_731 (O_731,N_47068,N_49348);
xnor UO_732 (O_732,N_45971,N_48507);
or UO_733 (O_733,N_49579,N_49600);
and UO_734 (O_734,N_45940,N_46765);
and UO_735 (O_735,N_47139,N_48092);
nand UO_736 (O_736,N_46611,N_47670);
xnor UO_737 (O_737,N_45120,N_47577);
nand UO_738 (O_738,N_47322,N_47611);
and UO_739 (O_739,N_47367,N_45780);
nor UO_740 (O_740,N_45192,N_49361);
or UO_741 (O_741,N_45513,N_49637);
xnor UO_742 (O_742,N_47807,N_48300);
nor UO_743 (O_743,N_48675,N_46241);
xor UO_744 (O_744,N_45883,N_49073);
nand UO_745 (O_745,N_46588,N_45818);
and UO_746 (O_746,N_46044,N_47409);
xor UO_747 (O_747,N_45374,N_48124);
xor UO_748 (O_748,N_45658,N_46543);
or UO_749 (O_749,N_45711,N_47749);
xor UO_750 (O_750,N_46812,N_47436);
xor UO_751 (O_751,N_47612,N_49243);
nor UO_752 (O_752,N_45636,N_45741);
nand UO_753 (O_753,N_47631,N_45359);
xor UO_754 (O_754,N_49150,N_46573);
nand UO_755 (O_755,N_48779,N_47864);
xnor UO_756 (O_756,N_48274,N_48032);
and UO_757 (O_757,N_49783,N_49003);
and UO_758 (O_758,N_49538,N_49961);
nand UO_759 (O_759,N_48994,N_46493);
xnor UO_760 (O_760,N_49106,N_47143);
nor UO_761 (O_761,N_46562,N_49264);
or UO_762 (O_762,N_48285,N_46542);
nand UO_763 (O_763,N_45603,N_45203);
nor UO_764 (O_764,N_46993,N_47006);
xor UO_765 (O_765,N_48073,N_45340);
nor UO_766 (O_766,N_49809,N_48403);
nand UO_767 (O_767,N_47875,N_48658);
nand UO_768 (O_768,N_48077,N_45556);
xnor UO_769 (O_769,N_46632,N_47639);
xnor UO_770 (O_770,N_46088,N_49234);
nand UO_771 (O_771,N_46643,N_47553);
and UO_772 (O_772,N_46214,N_46828);
xor UO_773 (O_773,N_45476,N_49235);
nor UO_774 (O_774,N_49058,N_46127);
nor UO_775 (O_775,N_48182,N_47941);
nor UO_776 (O_776,N_49622,N_46849);
nor UO_777 (O_777,N_47768,N_49028);
and UO_778 (O_778,N_48059,N_48534);
xnor UO_779 (O_779,N_47149,N_47497);
and UO_780 (O_780,N_45498,N_48648);
xor UO_781 (O_781,N_48339,N_47116);
nor UO_782 (O_782,N_49752,N_49316);
nor UO_783 (O_783,N_48513,N_47345);
and UO_784 (O_784,N_45760,N_45673);
nor UO_785 (O_785,N_48084,N_48048);
xor UO_786 (O_786,N_46221,N_49063);
nor UO_787 (O_787,N_45957,N_49257);
and UO_788 (O_788,N_45628,N_48758);
or UO_789 (O_789,N_47004,N_48873);
nand UO_790 (O_790,N_48762,N_45889);
nor UO_791 (O_791,N_46922,N_49955);
or UO_792 (O_792,N_48421,N_46704);
xor UO_793 (O_793,N_47973,N_48020);
and UO_794 (O_794,N_46713,N_49529);
or UO_795 (O_795,N_47358,N_46144);
nand UO_796 (O_796,N_49156,N_45271);
nor UO_797 (O_797,N_49383,N_45891);
xor UO_798 (O_798,N_47668,N_49698);
nand UO_799 (O_799,N_47444,N_49317);
or UO_800 (O_800,N_48582,N_47466);
nor UO_801 (O_801,N_45164,N_46191);
and UO_802 (O_802,N_47324,N_48794);
or UO_803 (O_803,N_47285,N_47814);
xor UO_804 (O_804,N_48885,N_49222);
nor UO_805 (O_805,N_47679,N_45831);
nor UO_806 (O_806,N_45858,N_47914);
nand UO_807 (O_807,N_49712,N_49151);
nand UO_808 (O_808,N_45375,N_49886);
and UO_809 (O_809,N_47278,N_48337);
nand UO_810 (O_810,N_47214,N_46318);
xor UO_811 (O_811,N_45539,N_48605);
nor UO_812 (O_812,N_48167,N_49666);
and UO_813 (O_813,N_46036,N_45602);
nand UO_814 (O_814,N_47910,N_46616);
nor UO_815 (O_815,N_47558,N_48608);
and UO_816 (O_816,N_49653,N_46984);
and UO_817 (O_817,N_48722,N_48081);
or UO_818 (O_818,N_46872,N_48566);
xnor UO_819 (O_819,N_45475,N_46139);
or UO_820 (O_820,N_47655,N_49757);
or UO_821 (O_821,N_49182,N_49837);
xor UO_822 (O_822,N_48718,N_49917);
nor UO_823 (O_823,N_48639,N_48209);
nand UO_824 (O_824,N_46846,N_45247);
and UO_825 (O_825,N_49803,N_46363);
and UO_826 (O_826,N_49051,N_48245);
xor UO_827 (O_827,N_47693,N_49439);
and UO_828 (O_828,N_45294,N_46359);
xor UO_829 (O_829,N_48128,N_46314);
or UO_830 (O_830,N_49044,N_49052);
nand UO_831 (O_831,N_48724,N_46167);
nand UO_832 (O_832,N_45468,N_46835);
or UO_833 (O_833,N_49974,N_46321);
nand UO_834 (O_834,N_46196,N_47326);
nand UO_835 (O_835,N_45907,N_46785);
nand UO_836 (O_836,N_47604,N_47145);
nand UO_837 (O_837,N_46798,N_46721);
xnor UO_838 (O_838,N_49229,N_47842);
or UO_839 (O_839,N_47800,N_45774);
xnor UO_840 (O_840,N_45017,N_47752);
or UO_841 (O_841,N_48856,N_47989);
xnor UO_842 (O_842,N_46262,N_49922);
and UO_843 (O_843,N_47372,N_45074);
xor UO_844 (O_844,N_46566,N_46808);
xnor UO_845 (O_845,N_49526,N_48905);
and UO_846 (O_846,N_46759,N_47891);
nand UO_847 (O_847,N_45199,N_46682);
or UO_848 (O_848,N_49701,N_47494);
and UO_849 (O_849,N_48458,N_49644);
and UO_850 (O_850,N_48239,N_46805);
nor UO_851 (O_851,N_45486,N_47208);
xor UO_852 (O_852,N_46077,N_49069);
nor UO_853 (O_853,N_48284,N_46116);
and UO_854 (O_854,N_46407,N_47859);
nor UO_855 (O_855,N_46575,N_49969);
nor UO_856 (O_856,N_45610,N_45554);
or UO_857 (O_857,N_45868,N_46741);
xnor UO_858 (O_858,N_46972,N_47964);
and UO_859 (O_859,N_45455,N_46962);
or UO_860 (O_860,N_45998,N_49498);
xor UO_861 (O_861,N_46500,N_49093);
or UO_862 (O_862,N_45735,N_47147);
or UO_863 (O_863,N_46900,N_46883);
and UO_864 (O_864,N_49987,N_47256);
or UO_865 (O_865,N_49941,N_45029);
xor UO_866 (O_866,N_49976,N_45984);
and UO_867 (O_867,N_45981,N_46674);
nand UO_868 (O_868,N_49034,N_48792);
or UO_869 (O_869,N_45254,N_45583);
xnor UO_870 (O_870,N_45783,N_49494);
nand UO_871 (O_871,N_48908,N_49311);
nor UO_872 (O_872,N_45037,N_49825);
nand UO_873 (O_873,N_45680,N_45620);
or UO_874 (O_874,N_46104,N_49736);
nor UO_875 (O_875,N_49885,N_47070);
and UO_876 (O_876,N_47916,N_48694);
nand UO_877 (O_877,N_45116,N_46949);
nand UO_878 (O_878,N_48719,N_48523);
or UO_879 (O_879,N_49520,N_49319);
nor UO_880 (O_880,N_45520,N_48898);
nor UO_881 (O_881,N_47525,N_46429);
and UO_882 (O_882,N_48098,N_49609);
or UO_883 (O_883,N_47513,N_47035);
xor UO_884 (O_884,N_47449,N_47443);
and UO_885 (O_885,N_45621,N_49821);
nor UO_886 (O_886,N_48119,N_45167);
or UO_887 (O_887,N_45315,N_49137);
or UO_888 (O_888,N_49213,N_47403);
nor UO_889 (O_889,N_47313,N_45163);
xor UO_890 (O_890,N_49335,N_46886);
nand UO_891 (O_891,N_49187,N_46642);
and UO_892 (O_892,N_45067,N_49784);
nand UO_893 (O_893,N_48304,N_46990);
nand UO_894 (O_894,N_45722,N_49265);
and UO_895 (O_895,N_45646,N_48140);
xnor UO_896 (O_896,N_45535,N_48759);
nand UO_897 (O_897,N_45561,N_45335);
or UO_898 (O_898,N_49877,N_45894);
or UO_899 (O_899,N_47957,N_49578);
and UO_900 (O_900,N_45525,N_45521);
nand UO_901 (O_901,N_45408,N_47126);
nor UO_902 (O_902,N_47905,N_45135);
nand UO_903 (O_903,N_46048,N_47417);
nor UO_904 (O_904,N_48312,N_46590);
or UO_905 (O_905,N_46992,N_47130);
xnor UO_906 (O_906,N_47517,N_49148);
nor UO_907 (O_907,N_48404,N_45001);
xor UO_908 (O_908,N_45829,N_46306);
and UO_909 (O_909,N_47972,N_45961);
nand UO_910 (O_910,N_49709,N_45383);
and UO_911 (O_911,N_47890,N_45467);
and UO_912 (O_912,N_45979,N_45617);
and UO_913 (O_913,N_47211,N_47018);
xnor UO_914 (O_914,N_49992,N_48702);
and UO_915 (O_915,N_48797,N_48526);
or UO_916 (O_916,N_45350,N_49903);
xnor UO_917 (O_917,N_49109,N_48363);
or UO_918 (O_918,N_49679,N_47400);
xor UO_919 (O_919,N_49178,N_46692);
nor UO_920 (O_920,N_46778,N_46173);
xor UO_921 (O_921,N_47847,N_47755);
nand UO_922 (O_922,N_47177,N_48576);
nand UO_923 (O_923,N_47779,N_48911);
xor UO_924 (O_924,N_46448,N_45855);
nor UO_925 (O_925,N_46515,N_46008);
or UO_926 (O_926,N_46212,N_46103);
nor UO_927 (O_927,N_46848,N_48715);
and UO_928 (O_928,N_46517,N_47721);
xor UO_929 (O_929,N_47551,N_45932);
nor UO_930 (O_930,N_48610,N_48618);
and UO_931 (O_931,N_46462,N_46783);
nand UO_932 (O_932,N_49129,N_49281);
xor UO_933 (O_933,N_45150,N_46183);
or UO_934 (O_934,N_49614,N_49372);
nor UO_935 (O_935,N_48665,N_45773);
xor UO_936 (O_936,N_47573,N_47660);
or UO_937 (O_937,N_49715,N_47295);
nand UO_938 (O_938,N_48114,N_48739);
and UO_939 (O_939,N_46460,N_47154);
xor UO_940 (O_940,N_49623,N_46354);
or UO_941 (O_941,N_48777,N_48692);
and UO_942 (O_942,N_49804,N_45436);
or UO_943 (O_943,N_48024,N_48321);
nand UO_944 (O_944,N_46857,N_47025);
xor UO_945 (O_945,N_48580,N_47901);
and UO_946 (O_946,N_45027,N_46307);
and UO_947 (O_947,N_49676,N_49855);
nor UO_948 (O_948,N_46046,N_48667);
or UO_949 (O_949,N_47239,N_48820);
and UO_950 (O_950,N_48997,N_45269);
and UO_951 (O_951,N_46864,N_47550);
and UO_952 (O_952,N_46159,N_48647);
or UO_953 (O_953,N_49007,N_45755);
nor UO_954 (O_954,N_47839,N_49669);
and UO_955 (O_955,N_45825,N_46237);
or UO_956 (O_956,N_48930,N_48947);
and UO_957 (O_957,N_45097,N_48877);
xor UO_958 (O_958,N_48691,N_47895);
nor UO_959 (O_959,N_45784,N_49002);
nor UO_960 (O_960,N_45041,N_47406);
nand UO_961 (O_961,N_46057,N_47390);
nand UO_962 (O_962,N_46014,N_48916);
and UO_963 (O_963,N_46198,N_46108);
and UO_964 (O_964,N_49819,N_49734);
and UO_965 (O_965,N_45660,N_45899);
nor UO_966 (O_966,N_48260,N_49362);
nor UO_967 (O_967,N_48015,N_45083);
nor UO_968 (O_968,N_47708,N_46387);
nor UO_969 (O_969,N_48700,N_48920);
or UO_970 (O_970,N_45517,N_45140);
and UO_971 (O_971,N_48110,N_46476);
nor UO_972 (O_972,N_45445,N_46936);
nand UO_973 (O_973,N_48879,N_46140);
or UO_974 (O_974,N_49470,N_48420);
nor UO_975 (O_975,N_49066,N_45497);
nor UO_976 (O_976,N_45172,N_49533);
nand UO_977 (O_977,N_45342,N_48085);
nor UO_978 (O_978,N_48393,N_47931);
nor UO_979 (O_979,N_46389,N_47944);
nor UO_980 (O_980,N_46626,N_47547);
xnor UO_981 (O_981,N_49287,N_45072);
nand UO_982 (O_982,N_47233,N_46701);
and UO_983 (O_983,N_46533,N_49780);
or UO_984 (O_984,N_48465,N_46443);
or UO_985 (O_985,N_47954,N_46895);
nand UO_986 (O_986,N_49050,N_48463);
nor UO_987 (O_987,N_46814,N_49377);
and UO_988 (O_988,N_45444,N_46987);
xor UO_989 (O_989,N_45363,N_46657);
nor UO_990 (O_990,N_47571,N_49694);
xnor UO_991 (O_991,N_49100,N_45518);
or UO_992 (O_992,N_46491,N_45553);
nand UO_993 (O_993,N_47192,N_47459);
and UO_994 (O_994,N_46552,N_45668);
nor UO_995 (O_995,N_48238,N_45756);
nor UO_996 (O_996,N_47009,N_47727);
nor UO_997 (O_997,N_49183,N_46915);
nor UO_998 (O_998,N_47672,N_47298);
nor UO_999 (O_999,N_49796,N_45519);
nor UO_1000 (O_1000,N_48301,N_46421);
nand UO_1001 (O_1001,N_46304,N_48062);
nand UO_1002 (O_1002,N_49421,N_46230);
nor UO_1003 (O_1003,N_45078,N_47907);
nand UO_1004 (O_1004,N_47987,N_46574);
nand UO_1005 (O_1005,N_49312,N_45056);
or UO_1006 (O_1006,N_47761,N_46512);
or UO_1007 (O_1007,N_45578,N_45978);
nor UO_1008 (O_1008,N_45863,N_49761);
nor UO_1009 (O_1009,N_45746,N_49558);
nand UO_1010 (O_1010,N_48500,N_45372);
or UO_1011 (O_1011,N_47142,N_48147);
nor UO_1012 (O_1012,N_47828,N_46330);
and UO_1013 (O_1013,N_49023,N_48656);
nor UO_1014 (O_1014,N_47125,N_46520);
and UO_1015 (O_1015,N_49274,N_46217);
or UO_1016 (O_1016,N_46513,N_46530);
nand UO_1017 (O_1017,N_47743,N_46740);
xor UO_1018 (O_1018,N_49626,N_48331);
nor UO_1019 (O_1019,N_47581,N_49331);
xnor UO_1020 (O_1020,N_46402,N_46974);
xnor UO_1021 (O_1021,N_47165,N_46583);
nand UO_1022 (O_1022,N_46986,N_45999);
xnor UO_1023 (O_1023,N_48629,N_47855);
nand UO_1024 (O_1024,N_48235,N_48680);
nand UO_1025 (O_1025,N_48153,N_45744);
or UO_1026 (O_1026,N_49450,N_45447);
and UO_1027 (O_1027,N_47539,N_49515);
nor UO_1028 (O_1028,N_49633,N_45759);
and UO_1029 (O_1029,N_49618,N_46587);
nand UO_1030 (O_1030,N_47002,N_47760);
nor UO_1031 (O_1031,N_46597,N_46935);
nor UO_1032 (O_1032,N_48843,N_47230);
nor UO_1033 (O_1033,N_45729,N_49368);
or UO_1034 (O_1034,N_47818,N_46368);
or UO_1035 (O_1035,N_46636,N_48536);
xnor UO_1036 (O_1036,N_48430,N_47578);
xnor UO_1037 (O_1037,N_49465,N_46603);
nand UO_1038 (O_1038,N_46666,N_49645);
nor UO_1039 (O_1039,N_49871,N_49022);
or UO_1040 (O_1040,N_49408,N_46403);
and UO_1041 (O_1041,N_48250,N_46347);
xor UO_1042 (O_1042,N_47595,N_47718);
or UO_1043 (O_1043,N_48950,N_45953);
xor UO_1044 (O_1044,N_45230,N_49889);
or UO_1045 (O_1045,N_46607,N_47146);
nand UO_1046 (O_1046,N_49703,N_49010);
nor UO_1047 (O_1047,N_46366,N_48872);
and UO_1048 (O_1048,N_46807,N_45942);
or UO_1049 (O_1049,N_48575,N_46928);
xnor UO_1050 (O_1050,N_48051,N_48584);
xor UO_1051 (O_1051,N_45094,N_46870);
and UO_1052 (O_1052,N_49228,N_49029);
and UO_1053 (O_1053,N_47469,N_48449);
or UO_1054 (O_1054,N_46279,N_49413);
nand UO_1055 (O_1055,N_47270,N_48427);
nor UO_1056 (O_1056,N_45881,N_49650);
and UO_1057 (O_1057,N_47535,N_47437);
nor UO_1058 (O_1058,N_46898,N_46580);
xnor UO_1059 (O_1059,N_48416,N_49539);
xnor UO_1060 (O_1060,N_48340,N_49661);
nand UO_1061 (O_1061,N_46316,N_49334);
xor UO_1062 (O_1062,N_49594,N_46172);
nand UO_1063 (O_1063,N_47922,N_46725);
nand UO_1064 (O_1064,N_45134,N_47399);
or UO_1065 (O_1065,N_46501,N_49923);
xor UO_1066 (O_1066,N_47943,N_48834);
and UO_1067 (O_1067,N_46877,N_45397);
or UO_1068 (O_1068,N_46035,N_48701);
nor UO_1069 (O_1069,N_48219,N_46040);
nand UO_1070 (O_1070,N_48981,N_47512);
and UO_1071 (O_1071,N_47911,N_46817);
nor UO_1072 (O_1072,N_47351,N_45669);
or UO_1073 (O_1073,N_49830,N_48336);
and UO_1074 (O_1074,N_46748,N_45168);
nor UO_1075 (O_1075,N_47056,N_48381);
nand UO_1076 (O_1076,N_47522,N_46350);
and UO_1077 (O_1077,N_49530,N_45443);
nor UO_1078 (O_1078,N_48134,N_45994);
and UO_1079 (O_1079,N_49221,N_45804);
and UO_1080 (O_1080,N_45376,N_49931);
or UO_1081 (O_1081,N_46916,N_49076);
nand UO_1082 (O_1082,N_45384,N_49425);
or UO_1083 (O_1083,N_47702,N_47884);
nand UO_1084 (O_1084,N_49227,N_49367);
nor UO_1085 (O_1085,N_46856,N_46884);
or UO_1086 (O_1086,N_46357,N_45597);
xor UO_1087 (O_1087,N_46253,N_49111);
and UO_1088 (O_1088,N_45893,N_46888);
and UO_1089 (O_1089,N_47701,N_48373);
and UO_1090 (O_1090,N_46185,N_49774);
xnor UO_1091 (O_1091,N_47312,N_45339);
or UO_1092 (O_1092,N_49947,N_49437);
or UO_1093 (O_1093,N_49071,N_47184);
and UO_1094 (O_1094,N_47392,N_47457);
and UO_1095 (O_1095,N_47013,N_48636);
xor UO_1096 (O_1096,N_49735,N_49401);
nor UO_1097 (O_1097,N_47225,N_47569);
xor UO_1098 (O_1098,N_48096,N_48937);
nand UO_1099 (O_1099,N_48542,N_46446);
or UO_1100 (O_1100,N_47027,N_46201);
nor UO_1101 (O_1101,N_48599,N_49043);
xor UO_1102 (O_1102,N_47020,N_45897);
or UO_1103 (O_1103,N_47418,N_48208);
and UO_1104 (O_1104,N_46145,N_46053);
or UO_1105 (O_1105,N_45010,N_46662);
or UO_1106 (O_1106,N_47279,N_46026);
nand UO_1107 (O_1107,N_49278,N_45540);
nand UO_1108 (O_1108,N_47519,N_47862);
xor UO_1109 (O_1109,N_47793,N_49298);
xor UO_1110 (O_1110,N_45586,N_48974);
or UO_1111 (O_1111,N_45824,N_49351);
and UO_1112 (O_1112,N_49233,N_48604);
nand UO_1113 (O_1113,N_45404,N_45958);
nor UO_1114 (O_1114,N_45563,N_48091);
xor UO_1115 (O_1115,N_46563,N_49168);
xor UO_1116 (O_1116,N_47281,N_49924);
or UO_1117 (O_1117,N_48750,N_47441);
nor UO_1118 (O_1118,N_49933,N_46334);
and UO_1119 (O_1119,N_49621,N_46109);
and UO_1120 (O_1120,N_45161,N_47081);
and UO_1121 (O_1121,N_46063,N_47034);
and UO_1122 (O_1122,N_47415,N_48764);
nand UO_1123 (O_1123,N_46625,N_48737);
nor UO_1124 (O_1124,N_49566,N_49336);
nand UO_1125 (O_1125,N_47040,N_46791);
nand UO_1126 (O_1126,N_48007,N_48023);
nor UO_1127 (O_1127,N_46939,N_46356);
xnor UO_1128 (O_1128,N_47032,N_48187);
xnor UO_1129 (O_1129,N_48964,N_45187);
and UO_1130 (O_1130,N_47869,N_45224);
nand UO_1131 (O_1131,N_45441,N_49569);
and UO_1132 (O_1132,N_48517,N_45288);
or UO_1133 (O_1133,N_49212,N_48368);
nor UO_1134 (O_1134,N_49506,N_45025);
nor UO_1135 (O_1135,N_48103,N_49285);
nand UO_1136 (O_1136,N_46731,N_46074);
and UO_1137 (O_1137,N_47568,N_45509);
nor UO_1138 (O_1138,N_48854,N_48789);
and UO_1139 (O_1139,N_45014,N_45814);
xor UO_1140 (O_1140,N_47219,N_47072);
nor UO_1141 (O_1141,N_48400,N_49389);
xnor UO_1142 (O_1142,N_45847,N_45728);
nand UO_1143 (O_1143,N_48154,N_49060);
nand UO_1144 (O_1144,N_48492,N_46686);
xor UO_1145 (O_1145,N_45612,N_48240);
or UO_1146 (O_1146,N_45524,N_46690);
nand UO_1147 (O_1147,N_47481,N_47501);
or UO_1148 (O_1148,N_45641,N_46071);
nor UO_1149 (O_1149,N_47217,N_46793);
and UO_1150 (O_1150,N_47704,N_48145);
nand UO_1151 (O_1151,N_49932,N_46768);
and UO_1152 (O_1152,N_47942,N_48193);
or UO_1153 (O_1153,N_49843,N_48910);
and UO_1154 (O_1154,N_48163,N_49844);
nand UO_1155 (O_1155,N_47363,N_49036);
nand UO_1156 (O_1156,N_45712,N_48391);
xnor UO_1157 (O_1157,N_48562,N_46199);
nor UO_1158 (O_1158,N_49454,N_49772);
or UO_1159 (O_1159,N_48886,N_48227);
and UO_1160 (O_1160,N_48295,N_47823);
xor UO_1161 (O_1161,N_47446,N_48411);
xor UO_1162 (O_1162,N_47063,N_47825);
or UO_1163 (O_1163,N_48704,N_47735);
nand UO_1164 (O_1164,N_48355,N_45373);
or UO_1165 (O_1165,N_48723,N_48514);
nand UO_1166 (O_1166,N_49731,N_46822);
and UO_1167 (O_1167,N_47852,N_46737);
xor UO_1168 (O_1168,N_47090,N_45830);
and UO_1169 (O_1169,N_46107,N_46072);
nand UO_1170 (O_1170,N_46879,N_49891);
nand UO_1171 (O_1171,N_49460,N_46188);
nor UO_1172 (O_1172,N_47232,N_48845);
nand UO_1173 (O_1173,N_46197,N_45900);
nor UO_1174 (O_1174,N_47259,N_48976);
xnor UO_1175 (O_1175,N_47904,N_46634);
nor UO_1176 (O_1176,N_47067,N_47194);
nor UO_1177 (O_1177,N_47945,N_45921);
and UO_1178 (O_1178,N_46641,N_46685);
nand UO_1179 (O_1179,N_48556,N_48011);
or UO_1180 (O_1180,N_48385,N_46728);
nand UO_1181 (O_1181,N_45031,N_47058);
and UO_1182 (O_1182,N_48827,N_46609);
nand UO_1183 (O_1183,N_47247,N_48946);
and UO_1184 (O_1184,N_45022,N_49249);
and UO_1185 (O_1185,N_49215,N_49601);
nor UO_1186 (O_1186,N_45160,N_46576);
and UO_1187 (O_1187,N_49291,N_47518);
xnor UO_1188 (O_1188,N_45508,N_45589);
nand UO_1189 (O_1189,N_45579,N_48933);
nor UO_1190 (O_1190,N_49639,N_49459);
and UO_1191 (O_1191,N_46398,N_45593);
and UO_1192 (O_1192,N_45068,N_47966);
and UO_1193 (O_1193,N_46859,N_47476);
xnor UO_1194 (O_1194,N_47492,N_48889);
nor UO_1195 (O_1195,N_49216,N_49392);
nand UO_1196 (O_1196,N_47792,N_46220);
or UO_1197 (O_1197,N_48793,N_49527);
xnor UO_1198 (O_1198,N_47306,N_46150);
nand UO_1199 (O_1199,N_49176,N_47148);
and UO_1200 (O_1200,N_49620,N_49719);
nor UO_1201 (O_1201,N_46985,N_48310);
and UO_1202 (O_1202,N_47806,N_47816);
or UO_1203 (O_1203,N_49299,N_46128);
xor UO_1204 (O_1204,N_48945,N_48720);
and UO_1205 (O_1205,N_45674,N_49294);
xnor UO_1206 (O_1206,N_45268,N_48999);
nand UO_1207 (O_1207,N_47305,N_47432);
and UO_1208 (O_1208,N_48251,N_47783);
xor UO_1209 (O_1209,N_48018,N_46177);
and UO_1210 (O_1210,N_47676,N_49219);
or UO_1211 (O_1211,N_45927,N_48679);
and UO_1212 (O_1212,N_47734,N_48131);
xor UO_1213 (O_1213,N_47958,N_47339);
or UO_1214 (O_1214,N_45218,N_48137);
nand UO_1215 (O_1215,N_47909,N_48364);
or UO_1216 (O_1216,N_45779,N_46606);
nand UO_1217 (O_1217,N_46602,N_47098);
nand UO_1218 (O_1218,N_48053,N_48010);
and UO_1219 (O_1219,N_48294,N_48382);
and UO_1220 (O_1220,N_45946,N_45733);
nand UO_1221 (O_1221,N_45501,N_45638);
nor UO_1222 (O_1222,N_49681,N_45221);
and UO_1223 (O_1223,N_45039,N_45075);
nand UO_1224 (O_1224,N_45442,N_46349);
or UO_1225 (O_1225,N_45869,N_45407);
nand UO_1226 (O_1226,N_49997,N_45472);
nor UO_1227 (O_1227,N_48269,N_46019);
nor UO_1228 (O_1228,N_45183,N_45822);
or UO_1229 (O_1229,N_49356,N_47594);
nor UO_1230 (O_1230,N_48870,N_48736);
and UO_1231 (O_1231,N_48281,N_47658);
nor UO_1232 (O_1232,N_46206,N_48303);
or UO_1233 (O_1233,N_45250,N_45976);
xnor UO_1234 (O_1234,N_47769,N_46381);
or UO_1235 (O_1235,N_45147,N_49133);
xnor UO_1236 (O_1236,N_48892,N_45259);
or UO_1237 (O_1237,N_48970,N_49990);
nand UO_1238 (O_1238,N_45012,N_45792);
nor UO_1239 (O_1239,N_45285,N_48591);
nor UO_1240 (O_1240,N_48774,N_46983);
xnor UO_1241 (O_1241,N_46352,N_48409);
or UO_1242 (O_1242,N_47274,N_47401);
and UO_1243 (O_1243,N_46942,N_47930);
xnor UO_1244 (O_1244,N_49861,N_47950);
and UO_1245 (O_1245,N_47836,N_47161);
or UO_1246 (O_1246,N_45596,N_49157);
or UO_1247 (O_1247,N_45085,N_46353);
xor UO_1248 (O_1248,N_45861,N_46578);
or UO_1249 (O_1249,N_48731,N_47970);
nand UO_1250 (O_1250,N_47854,N_45471);
nand UO_1251 (O_1251,N_47361,N_45951);
and UO_1252 (O_1252,N_45738,N_49564);
nor UO_1253 (O_1253,N_45226,N_46323);
xor UO_1254 (O_1254,N_48948,N_46917);
or UO_1255 (O_1255,N_49297,N_49310);
and UO_1256 (O_1256,N_45697,N_48822);
nor UO_1257 (O_1257,N_45267,N_45785);
nor UO_1258 (O_1258,N_48089,N_47938);
nor UO_1259 (O_1259,N_48631,N_47304);
xor UO_1260 (O_1260,N_46396,N_48213);
and UO_1261 (O_1261,N_49838,N_49476);
nor UO_1262 (O_1262,N_48164,N_48044);
and UO_1263 (O_1263,N_46545,N_45299);
or UO_1264 (O_1264,N_49705,N_47782);
and UO_1265 (O_1265,N_45870,N_48847);
nand UO_1266 (O_1266,N_46059,N_46102);
nand UO_1267 (O_1267,N_46579,N_49841);
or UO_1268 (O_1268,N_48798,N_49271);
nand UO_1269 (O_1269,N_47838,N_45788);
or UO_1270 (O_1270,N_47967,N_49101);
nor UO_1271 (O_1271,N_47866,N_48796);
nor UO_1272 (O_1272,N_49411,N_49659);
xor UO_1273 (O_1273,N_49975,N_46425);
or UO_1274 (O_1274,N_48246,N_46325);
or UO_1275 (O_1275,N_45880,N_47564);
and UO_1276 (O_1276,N_49374,N_47533);
nand UO_1277 (O_1277,N_45997,N_49225);
or UO_1278 (O_1278,N_46015,N_47043);
nor UO_1279 (O_1279,N_47726,N_49402);
nand UO_1280 (O_1280,N_47813,N_49581);
nand UO_1281 (O_1281,N_45613,N_49089);
xor UO_1282 (O_1282,N_48265,N_46541);
nand UO_1283 (O_1283,N_47277,N_49365);
and UO_1284 (O_1284,N_47302,N_46537);
or UO_1285 (O_1285,N_48318,N_49849);
and UO_1286 (O_1286,N_47291,N_45059);
nor UO_1287 (O_1287,N_49359,N_47832);
nor UO_1288 (O_1288,N_46927,N_46267);
nor UO_1289 (O_1289,N_47402,N_46478);
nand UO_1290 (O_1290,N_46940,N_48050);
nor UO_1291 (O_1291,N_45054,N_46296);
xor UO_1292 (O_1292,N_45349,N_49364);
or UO_1293 (O_1293,N_45426,N_46937);
and UO_1294 (O_1294,N_47992,N_46640);
or UO_1295 (O_1295,N_49412,N_46115);
nor UO_1296 (O_1296,N_46064,N_45277);
and UO_1297 (O_1297,N_47129,N_48986);
and UO_1298 (O_1298,N_47331,N_45004);
nor UO_1299 (O_1299,N_49160,N_45794);
nand UO_1300 (O_1300,N_46287,N_46415);
xnor UO_1301 (O_1301,N_45799,N_45145);
or UO_1302 (O_1302,N_48252,N_46269);
or UO_1303 (O_1303,N_46376,N_47391);
xor UO_1304 (O_1304,N_45959,N_47790);
nand UO_1305 (O_1305,N_47085,N_47858);
nand UO_1306 (O_1306,N_47168,N_46299);
xor UO_1307 (O_1307,N_45207,N_45456);
xor UO_1308 (O_1308,N_45178,N_45862);
nor UO_1309 (O_1309,N_45910,N_48837);
nor UO_1310 (O_1310,N_45432,N_48317);
and UO_1311 (O_1311,N_46006,N_48129);
xnor UO_1312 (O_1312,N_48306,N_48971);
or UO_1313 (O_1313,N_45750,N_47837);
xor UO_1314 (O_1314,N_45064,N_47576);
nand UO_1315 (O_1315,N_49748,N_46335);
and UO_1316 (O_1316,N_47128,N_45985);
nand UO_1317 (O_1317,N_46258,N_48869);
nand UO_1318 (O_1318,N_48890,N_47050);
xor UO_1319 (O_1319,N_49721,N_49723);
and UO_1320 (O_1320,N_46470,N_45848);
xor UO_1321 (O_1321,N_47404,N_47739);
nand UO_1322 (O_1322,N_46331,N_47681);
or UO_1323 (O_1323,N_46789,N_45470);
nor UO_1324 (O_1324,N_46339,N_47650);
xnor UO_1325 (O_1325,N_45956,N_47724);
nand UO_1326 (O_1326,N_45141,N_46830);
nor UO_1327 (O_1327,N_48342,N_49259);
nor UO_1328 (O_1328,N_47975,N_49146);
xnor UO_1329 (O_1329,N_45892,N_49095);
and UO_1330 (O_1330,N_49918,N_49239);
or UO_1331 (O_1331,N_48748,N_47562);
nor UO_1332 (O_1332,N_46693,N_45036);
nand UO_1333 (O_1333,N_49959,N_48866);
or UO_1334 (O_1334,N_46110,N_47074);
and UO_1335 (O_1335,N_46065,N_47811);
xnor UO_1336 (O_1336,N_45217,N_49737);
xor UO_1337 (O_1337,N_45567,N_49032);
xnor UO_1338 (O_1338,N_49683,N_46496);
nor UO_1339 (O_1339,N_46414,N_46409);
or UO_1340 (O_1340,N_48378,N_47220);
nor UO_1341 (O_1341,N_48438,N_48683);
and UO_1342 (O_1342,N_48478,N_49806);
or UO_1343 (O_1343,N_47527,N_45222);
nor UO_1344 (O_1344,N_45466,N_46499);
and UO_1345 (O_1345,N_45811,N_45740);
nand UO_1346 (O_1346,N_47889,N_49968);
and UO_1347 (O_1347,N_46751,N_45411);
and UO_1348 (O_1348,N_47366,N_46484);
nor UO_1349 (O_1349,N_49649,N_48957);
nand UO_1350 (O_1350,N_45627,N_48672);
or UO_1351 (O_1351,N_47561,N_45303);
nor UO_1352 (O_1352,N_46595,N_49724);
nor UO_1353 (O_1353,N_46559,N_47575);
xnor UO_1354 (O_1354,N_48983,N_46034);
and UO_1355 (O_1355,N_45969,N_46101);
or UO_1356 (O_1356,N_45924,N_48923);
or UO_1357 (O_1357,N_45367,N_45866);
nand UO_1358 (O_1358,N_46030,N_48190);
or UO_1359 (O_1359,N_47952,N_45850);
xnor UO_1360 (O_1360,N_48646,N_49519);
nand UO_1361 (O_1361,N_45705,N_45696);
and UO_1362 (O_1362,N_48703,N_49388);
nor UO_1363 (O_1363,N_46899,N_46379);
nand UO_1364 (O_1364,N_48067,N_47112);
nand UO_1365 (O_1365,N_47173,N_49919);
and UO_1366 (O_1366,N_46477,N_48922);
and UO_1367 (O_1367,N_48965,N_49727);
xnor UO_1368 (O_1368,N_46056,N_45387);
xnor UO_1369 (O_1369,N_48350,N_47144);
xnor UO_1370 (O_1370,N_49305,N_47271);
nor UO_1371 (O_1371,N_49125,N_45313);
xor UO_1372 (O_1372,N_49989,N_48072);
and UO_1373 (O_1373,N_46372,N_45234);
xor UO_1374 (O_1374,N_45718,N_48828);
xnor UO_1375 (O_1375,N_49279,N_47835);
and UO_1376 (O_1376,N_45197,N_45125);
nor UO_1377 (O_1377,N_48268,N_47781);
nor UO_1378 (O_1378,N_45611,N_46433);
and UO_1379 (O_1379,N_49246,N_47395);
xnor UO_1380 (O_1380,N_47524,N_45782);
nor UO_1381 (O_1381,N_45156,N_49673);
or UO_1382 (O_1382,N_48998,N_48674);
xnor UO_1383 (O_1383,N_47186,N_49141);
xnor UO_1384 (O_1384,N_49449,N_49144);
and UO_1385 (O_1385,N_48408,N_45328);
or UO_1386 (O_1386,N_47630,N_48122);
xnor UO_1387 (O_1387,N_45693,N_45699);
nand UO_1388 (O_1388,N_49399,N_47589);
nand UO_1389 (O_1389,N_47269,N_46447);
nand UO_1390 (O_1390,N_45096,N_45195);
or UO_1391 (O_1391,N_48689,N_49136);
xor UO_1392 (O_1392,N_47682,N_46473);
or UO_1393 (O_1393,N_46561,N_45614);
nor UO_1394 (O_1394,N_45402,N_47253);
or UO_1395 (O_1395,N_45727,N_45983);
xnor UO_1396 (O_1396,N_48586,N_48369);
nand UO_1397 (O_1397,N_45534,N_48019);
nor UO_1398 (O_1398,N_47051,N_48505);
or UO_1399 (O_1399,N_49619,N_45559);
nor UO_1400 (O_1400,N_46399,N_47172);
nor UO_1401 (O_1401,N_46881,N_49184);
or UO_1402 (O_1402,N_47489,N_45300);
nor UO_1403 (O_1403,N_49875,N_48402);
and UO_1404 (O_1404,N_49660,N_48852);
and UO_1405 (O_1405,N_49188,N_48941);
and UO_1406 (O_1406,N_45420,N_47266);
and UO_1407 (O_1407,N_45937,N_46245);
or UO_1408 (O_1408,N_46508,N_46806);
xor UO_1409 (O_1409,N_47062,N_47096);
or UO_1410 (O_1410,N_46837,N_49333);
nor UO_1411 (O_1411,N_48896,N_46320);
nand UO_1412 (O_1412,N_46338,N_49910);
xor UO_1413 (O_1413,N_49805,N_47764);
xnor UO_1414 (O_1414,N_49270,N_45594);
nor UO_1415 (O_1415,N_49417,N_45151);
nor UO_1416 (O_1416,N_45512,N_46539);
xnor UO_1417 (O_1417,N_49397,N_46706);
xnor UO_1418 (O_1418,N_49782,N_46630);
and UO_1419 (O_1419,N_47218,N_46256);
xor UO_1420 (O_1420,N_48621,N_49395);
nor UO_1421 (O_1421,N_45104,N_46823);
or UO_1422 (O_1422,N_46868,N_48472);
nand UO_1423 (O_1423,N_48747,N_49977);
and UO_1424 (O_1424,N_45566,N_45801);
nand UO_1425 (O_1425,N_46675,N_49004);
and UO_1426 (O_1426,N_47936,N_47241);
or UO_1427 (O_1427,N_49926,N_49856);
nand UO_1428 (O_1428,N_48138,N_48141);
nand UO_1429 (O_1429,N_45791,N_45964);
xor UO_1430 (O_1430,N_45101,N_49817);
and UO_1431 (O_1431,N_48829,N_49242);
and UO_1432 (O_1432,N_45177,N_45483);
and UO_1433 (O_1433,N_49456,N_48076);
xnor UO_1434 (O_1434,N_45772,N_49678);
or UO_1435 (O_1435,N_48555,N_47052);
xnor UO_1436 (O_1436,N_45348,N_49516);
nor UO_1437 (O_1437,N_49406,N_49366);
and UO_1438 (O_1438,N_48229,N_46506);
xor UO_1439 (O_1439,N_46084,N_48308);
xor UO_1440 (O_1440,N_48778,N_49241);
and UO_1441 (O_1441,N_45576,N_48105);
and UO_1442 (O_1442,N_47872,N_46718);
xnor UO_1443 (O_1443,N_46810,N_49971);
xor UO_1444 (O_1444,N_46242,N_49327);
nand UO_1445 (O_1445,N_47120,N_45911);
nand UO_1446 (O_1446,N_48550,N_49852);
nor UO_1447 (O_1447,N_48160,N_49726);
nand UO_1448 (O_1448,N_45966,N_48501);
nand UO_1449 (O_1449,N_47801,N_47685);
and UO_1450 (O_1450,N_49360,N_46865);
nand UO_1451 (O_1451,N_49513,N_46699);
nor UO_1452 (O_1452,N_45797,N_48445);
nor UO_1453 (O_1453,N_45516,N_46956);
and UO_1454 (O_1454,N_47812,N_49882);
nand UO_1455 (O_1455,N_47157,N_49067);
and UO_1456 (O_1456,N_49981,N_46773);
nor UO_1457 (O_1457,N_46298,N_45793);
or UO_1458 (O_1458,N_48237,N_46374);
nand UO_1459 (O_1459,N_45967,N_48311);
and UO_1460 (O_1460,N_46727,N_48770);
and UO_1461 (O_1461,N_48031,N_48993);
nand UO_1462 (O_1462,N_47703,N_49866);
xnor UO_1463 (O_1463,N_47608,N_49643);
and UO_1464 (O_1464,N_45745,N_47822);
xnor UO_1465 (O_1465,N_47488,N_48884);
xnor UO_1466 (O_1466,N_46954,N_48763);
or UO_1467 (O_1467,N_49481,N_48188);
or UO_1468 (O_1468,N_49570,N_45020);
xnor UO_1469 (O_1469,N_49787,N_46678);
xnor UO_1470 (O_1470,N_47092,N_45716);
or UO_1471 (O_1471,N_46028,N_46405);
and UO_1472 (O_1472,N_45358,N_45515);
nor UO_1473 (O_1473,N_45502,N_45703);
nor UO_1474 (O_1474,N_49398,N_48374);
nand UO_1475 (O_1475,N_49378,N_49031);
or UO_1476 (O_1476,N_45608,N_45159);
and UO_1477 (O_1477,N_47523,N_45421);
nor UO_1478 (O_1478,N_49508,N_48726);
xor UO_1479 (O_1479,N_45918,N_48068);
and UO_1480 (O_1480,N_45410,N_47246);
or UO_1481 (O_1481,N_45871,N_48214);
or UO_1482 (O_1482,N_46418,N_47598);
nor UO_1483 (O_1483,N_47548,N_48776);
nor UO_1484 (O_1484,N_47881,N_47824);
and UO_1485 (O_1485,N_48666,N_47290);
or UO_1486 (O_1486,N_46094,N_49455);
or UO_1487 (O_1487,N_45686,N_48943);
and UO_1488 (O_1488,N_47780,N_45208);
xnor UO_1489 (O_1489,N_46624,N_45413);
xnor UO_1490 (O_1490,N_48457,N_47606);
nor UO_1491 (O_1491,N_46081,N_45185);
or UO_1492 (O_1492,N_45137,N_48944);
xor UO_1493 (O_1493,N_45692,N_48548);
xnor UO_1494 (O_1494,N_45577,N_46069);
nor UO_1495 (O_1495,N_47537,N_47244);
xnor UO_1496 (O_1496,N_45670,N_49452);
and UO_1497 (O_1497,N_47508,N_49056);
and UO_1498 (O_1498,N_48113,N_49469);
nand UO_1499 (O_1499,N_49177,N_49064);
nand UO_1500 (O_1500,N_45331,N_48371);
nor UO_1501 (O_1501,N_45352,N_46938);
nor UO_1502 (O_1502,N_45105,N_49252);
or UO_1503 (O_1503,N_45538,N_46340);
or UO_1504 (O_1504,N_49433,N_46492);
nor UO_1505 (O_1505,N_47330,N_47108);
nand UO_1506 (O_1506,N_49379,N_49430);
nand UO_1507 (O_1507,N_46079,N_47939);
xnor UO_1508 (O_1508,N_45562,N_49224);
xnor UO_1509 (O_1509,N_46739,N_48026);
and UO_1510 (O_1510,N_49699,N_45607);
and UO_1511 (O_1511,N_47520,N_45048);
and UO_1512 (O_1512,N_45739,N_45191);
nand UO_1513 (O_1513,N_48395,N_45914);
or UO_1514 (O_1514,N_47935,N_45572);
xor UO_1515 (O_1515,N_49493,N_45490);
xnor UO_1516 (O_1516,N_47309,N_45263);
xnor UO_1517 (O_1517,N_45388,N_46431);
nor UO_1518 (O_1518,N_45810,N_49046);
or UO_1519 (O_1519,N_45220,N_49685);
nand UO_1520 (O_1520,N_45872,N_47502);
or UO_1521 (O_1521,N_48453,N_45661);
or UO_1522 (O_1522,N_49382,N_45121);
or UO_1523 (O_1523,N_49099,N_49635);
and UO_1524 (O_1524,N_45654,N_49258);
nand UO_1525 (O_1525,N_47053,N_47327);
nand UO_1526 (O_1526,N_45803,N_46067);
nor UO_1527 (O_1527,N_49501,N_47744);
or UO_1528 (O_1528,N_46032,N_47356);
and UO_1529 (O_1529,N_47170,N_49080);
and UO_1530 (O_1530,N_47440,N_45418);
nor UO_1531 (O_1531,N_49718,N_46775);
nand UO_1532 (O_1532,N_45241,N_49908);
xor UO_1533 (O_1533,N_47325,N_49338);
nor UO_1534 (O_1534,N_45131,N_48733);
or UO_1535 (O_1535,N_48094,N_46978);
and UO_1536 (O_1536,N_47493,N_48338);
nor UO_1537 (O_1537,N_48651,N_46733);
nor UO_1538 (O_1538,N_46277,N_49595);
and UO_1539 (O_1539,N_47075,N_45344);
xor UO_1540 (O_1540,N_48223,N_49521);
and UO_1541 (O_1541,N_45381,N_46160);
or UO_1542 (O_1542,N_48606,N_45672);
or UO_1543 (O_1543,N_49009,N_49717);
nor UO_1544 (O_1544,N_47528,N_47373);
or UO_1545 (O_1545,N_47821,N_49139);
and UO_1546 (O_1546,N_49532,N_46061);
nor UO_1547 (O_1547,N_45045,N_48949);
nor UO_1548 (O_1548,N_46955,N_48365);
and UO_1549 (O_1549,N_48713,N_47240);
or UO_1550 (O_1550,N_46166,N_47988);
xnor UO_1551 (O_1551,N_45625,N_46781);
nor UO_1552 (O_1552,N_46920,N_48045);
or UO_1553 (O_1553,N_46156,N_46042);
and UO_1554 (O_1554,N_48126,N_48347);
and UO_1555 (O_1555,N_49117,N_47061);
nor UO_1556 (O_1556,N_47632,N_48815);
or UO_1557 (O_1557,N_45808,N_49662);
and UO_1558 (O_1558,N_49276,N_46719);
xor UO_1559 (O_1559,N_46885,N_47927);
nor UO_1560 (O_1560,N_49766,N_49563);
nand UO_1561 (O_1561,N_46729,N_45832);
nor UO_1562 (O_1562,N_46342,N_48975);
and UO_1563 (O_1563,N_45318,N_49528);
or UO_1564 (O_1564,N_46152,N_48132);
nand UO_1565 (O_1565,N_45171,N_48987);
xor UO_1566 (O_1566,N_46440,N_48583);
nor UO_1567 (O_1567,N_47664,N_47788);
nand UO_1568 (O_1568,N_47099,N_46555);
nand UO_1569 (O_1569,N_45827,N_46163);
and UO_1570 (O_1570,N_46428,N_45995);
or UO_1571 (O_1571,N_45820,N_48225);
or UO_1572 (O_1572,N_49522,N_45805);
and UO_1573 (O_1573,N_46271,N_45047);
nor UO_1574 (O_1574,N_48554,N_48623);
or UO_1575 (O_1575,N_49934,N_45645);
or UO_1576 (O_1576,N_48313,N_48509);
or UO_1577 (O_1577,N_48628,N_49492);
nand UO_1578 (O_1578,N_46143,N_45635);
nor UO_1579 (O_1579,N_48824,N_45974);
and UO_1580 (O_1580,N_47636,N_46012);
nand UO_1581 (O_1581,N_46204,N_47314);
and UO_1582 (O_1582,N_49196,N_49739);
or UO_1583 (O_1583,N_48684,N_48642);
and UO_1584 (O_1584,N_47585,N_46824);
or UO_1585 (O_1585,N_46819,N_47288);
xnor UO_1586 (O_1586,N_45710,N_45662);
or UO_1587 (O_1587,N_47831,N_48956);
nor UO_1588 (O_1588,N_49741,N_48574);
xnor UO_1589 (O_1589,N_46747,N_49214);
and UO_1590 (O_1590,N_46131,N_47487);
nand UO_1591 (O_1591,N_46469,N_49232);
xnor UO_1592 (O_1592,N_49535,N_46598);
and UO_1593 (O_1593,N_46558,N_47767);
xor UO_1594 (O_1594,N_46712,N_49665);
nor UO_1595 (O_1595,N_49174,N_45919);
xnor UO_1596 (O_1596,N_49108,N_48655);
or UO_1597 (O_1597,N_47912,N_48657);
nor UO_1598 (O_1598,N_46442,N_47448);
nor UO_1599 (O_1599,N_47329,N_48989);
and UO_1600 (O_1600,N_45778,N_45016);
and UO_1601 (O_1601,N_45675,N_48181);
and UO_1602 (O_1602,N_47175,N_47980);
xnor UO_1603 (O_1603,N_48942,N_45679);
or UO_1604 (O_1604,N_49580,N_48241);
nor UO_1605 (O_1605,N_49057,N_46037);
nand UO_1606 (O_1606,N_46758,N_48883);
xnor UO_1607 (O_1607,N_46005,N_47775);
nor UO_1608 (O_1608,N_46827,N_45463);
nand UO_1609 (O_1609,N_49696,N_49154);
xnor UO_1610 (O_1610,N_49416,N_45629);
or UO_1611 (O_1611,N_46818,N_45040);
or UO_1612 (O_1612,N_49789,N_46832);
or UO_1613 (O_1613,N_46272,N_45107);
and UO_1614 (O_1614,N_47627,N_45061);
and UO_1615 (O_1615,N_49195,N_49956);
nand UO_1616 (O_1616,N_49277,N_47465);
xnor UO_1617 (O_1617,N_47737,N_46216);
or UO_1618 (O_1618,N_49300,N_48377);
nor UO_1619 (O_1619,N_49440,N_45043);
nand UO_1620 (O_1620,N_48046,N_48279);
and UO_1621 (O_1621,N_46676,N_45726);
xnor UO_1622 (O_1622,N_47622,N_46273);
nand UO_1623 (O_1623,N_49826,N_49198);
xor UO_1624 (O_1624,N_45333,N_49901);
or UO_1625 (O_1625,N_49647,N_45743);
nor UO_1626 (O_1626,N_47407,N_46082);
xnor UO_1627 (O_1627,N_48859,N_47132);
or UO_1628 (O_1628,N_48481,N_49200);
xnor UO_1629 (O_1629,N_47978,N_47413);
nand UO_1630 (O_1630,N_45386,N_47150);
nand UO_1631 (O_1631,N_45143,N_46129);
nand UO_1632 (O_1632,N_47234,N_49488);
xor UO_1633 (O_1633,N_49906,N_49549);
and UO_1634 (O_1634,N_49920,N_48000);
or UO_1635 (O_1635,N_49878,N_46863);
or UO_1636 (O_1636,N_45492,N_47516);
or UO_1637 (O_1637,N_45308,N_47036);
and UO_1638 (O_1638,N_47648,N_49011);
xor UO_1639 (O_1639,N_49776,N_47284);
nor UO_1640 (O_1640,N_46055,N_49810);
and UO_1641 (O_1641,N_45879,N_49085);
nand UO_1642 (O_1642,N_47393,N_45886);
or UO_1643 (O_1643,N_47420,N_48332);
or UO_1644 (O_1644,N_46882,N_47646);
or UO_1645 (O_1645,N_48624,N_49958);
and UO_1646 (O_1646,N_47453,N_47104);
and UO_1647 (O_1647,N_47976,N_49191);
nand UO_1648 (O_1648,N_46591,N_48880);
nor UO_1649 (O_1649,N_49306,N_45844);
and UO_1650 (O_1650,N_48399,N_46538);
or UO_1651 (O_1651,N_49807,N_47163);
nor UO_1652 (O_1652,N_47249,N_47151);
nor UO_1653 (O_1653,N_48204,N_48211);
xnor UO_1654 (O_1654,N_48525,N_48958);
nor UO_1655 (O_1655,N_47174,N_48522);
and UO_1656 (O_1656,N_48620,N_46229);
nand UO_1657 (O_1657,N_46941,N_47977);
nor UO_1658 (O_1658,N_47829,N_47592);
xnor UO_1659 (O_1659,N_48836,N_48738);
or UO_1660 (O_1660,N_48609,N_45664);
or UO_1661 (O_1661,N_48414,N_45558);
nor UO_1662 (O_1662,N_47751,N_49984);
xnor UO_1663 (O_1663,N_45260,N_45401);
nor UO_1664 (O_1664,N_49967,N_46742);
or UO_1665 (O_1665,N_46441,N_49210);
or UO_1666 (O_1666,N_49854,N_46735);
and UO_1667 (O_1667,N_49203,N_45640);
nand UO_1668 (O_1668,N_45631,N_47514);
or UO_1669 (O_1669,N_48510,N_46369);
or UO_1670 (O_1670,N_45274,N_48036);
xor UO_1671 (O_1671,N_46210,N_48021);
xor UO_1672 (O_1672,N_49473,N_49534);
nand UO_1673 (O_1673,N_46451,N_47301);
xnor UO_1674 (O_1674,N_48305,N_49695);
nand UO_1675 (O_1675,N_46839,N_47396);
xnor UO_1676 (O_1676,N_47308,N_48607);
or UO_1677 (O_1677,N_47071,N_47123);
or UO_1678 (O_1678,N_48255,N_49006);
nand UO_1679 (O_1679,N_48248,N_47102);
or UO_1680 (O_1680,N_46722,N_47882);
nand UO_1681 (O_1681,N_48034,N_45543);
and UO_1682 (O_1682,N_48345,N_48275);
xnor UO_1683 (O_1683,N_48121,N_46619);
and UO_1684 (O_1684,N_45252,N_46840);
nand UO_1685 (O_1685,N_48054,N_46404);
xnor UO_1686 (O_1686,N_48002,N_49204);
and UO_1687 (O_1687,N_48111,N_49710);
nor UO_1688 (O_1688,N_49785,N_45720);
and UO_1689 (O_1689,N_45278,N_48095);
and UO_1690 (O_1690,N_46989,N_46847);
xnor UO_1691 (O_1691,N_45346,N_48637);
nand UO_1692 (O_1692,N_45021,N_49750);
nand UO_1693 (O_1693,N_48835,N_45890);
and UO_1694 (O_1694,N_45454,N_46594);
nand UO_1695 (O_1695,N_47365,N_46787);
nand UO_1696 (O_1696,N_49491,N_48049);
nand UO_1697 (O_1697,N_48360,N_47628);
xnor UO_1698 (O_1698,N_47559,N_49759);
nor UO_1699 (O_1699,N_45671,N_46502);
and UO_1700 (O_1700,N_48743,N_49677);
and UO_1701 (O_1701,N_45412,N_47316);
or UO_1702 (O_1702,N_49250,N_46952);
or UO_1703 (O_1703,N_45438,N_48104);
xor UO_1704 (O_1704,N_47714,N_48224);
and UO_1705 (O_1705,N_49444,N_47222);
xnor UO_1706 (O_1706,N_47178,N_48471);
xor UO_1707 (O_1707,N_45127,N_46266);
nand UO_1708 (O_1708,N_45070,N_49065);
or UO_1709 (O_1709,N_45748,N_45493);
xor UO_1710 (O_1710,N_45465,N_45117);
nand UO_1711 (O_1711,N_45464,N_48650);
nor UO_1712 (O_1712,N_45537,N_45484);
xnor UO_1713 (O_1713,N_45338,N_49087);
and UO_1714 (O_1714,N_47228,N_47122);
xnor UO_1715 (O_1715,N_47212,N_47715);
xnor UO_1716 (O_1716,N_45084,N_48687);
nand UO_1717 (O_1717,N_45325,N_45947);
nand UO_1718 (O_1718,N_48511,N_45633);
and UO_1719 (O_1719,N_48570,N_46076);
and UO_1720 (O_1720,N_49670,N_46866);
or UO_1721 (O_1721,N_46921,N_46371);
xnor UO_1722 (O_1722,N_48013,N_45902);
nand UO_1723 (O_1723,N_49088,N_48460);
or UO_1724 (O_1724,N_47819,N_47634);
and UO_1725 (O_1725,N_47877,N_48118);
nor UO_1726 (O_1726,N_49779,N_46038);
or UO_1727 (O_1727,N_48372,N_46531);
nor UO_1728 (O_1728,N_47530,N_45968);
nor UO_1729 (O_1729,N_46906,N_48936);
nor UO_1730 (O_1730,N_45311,N_48454);
nand UO_1731 (O_1731,N_47998,N_47262);
nor UO_1732 (O_1732,N_46091,N_48855);
nor UO_1733 (O_1733,N_49762,N_49711);
nor UO_1734 (O_1734,N_49518,N_49552);
nor UO_1735 (O_1735,N_46395,N_46449);
or UO_1736 (O_1736,N_48557,N_45130);
or UO_1737 (O_1737,N_45928,N_45213);
nor UO_1738 (O_1738,N_46119,N_48348);
nor UO_1739 (O_1739,N_47328,N_46544);
nand UO_1740 (O_1740,N_48161,N_49486);
nor UO_1741 (O_1741,N_45816,N_49940);
nand UO_1742 (O_1742,N_45209,N_46027);
and UO_1743 (O_1743,N_45532,N_45154);
xnor UO_1744 (O_1744,N_46158,N_49823);
and UO_1745 (O_1745,N_47541,N_46784);
nand UO_1746 (O_1746,N_46302,N_45955);
or UO_1747 (O_1747,N_45753,N_48645);
nor UO_1748 (O_1748,N_48266,N_46313);
nor UO_1749 (O_1749,N_47059,N_49231);
and UO_1750 (O_1750,N_46481,N_47410);
nor UO_1751 (O_1751,N_46010,N_49689);
nor UO_1752 (O_1752,N_47883,N_48437);
xor UO_1753 (O_1753,N_45954,N_49646);
nand UO_1754 (O_1754,N_46651,N_48978);
nor UO_1755 (O_1755,N_45681,N_46933);
nand UO_1756 (O_1756,N_45905,N_45702);
nand UO_1757 (O_1757,N_49381,N_45364);
nor UO_1758 (O_1758,N_47731,N_47580);
nand UO_1759 (O_1759,N_47376,N_47659);
xor UO_1760 (O_1760,N_48952,N_47695);
or UO_1761 (O_1761,N_46148,N_45175);
nand UO_1762 (O_1762,N_48515,N_46257);
or UO_1763 (O_1763,N_47064,N_46181);
nand UO_1764 (O_1764,N_46664,N_49512);
nand UO_1765 (O_1765,N_48440,N_49747);
xnor UO_1766 (O_1766,N_49672,N_45651);
nand UO_1767 (O_1767,N_46707,N_49812);
xor UO_1768 (O_1768,N_45111,N_49939);
and UO_1769 (O_1769,N_45933,N_49613);
nor UO_1770 (O_1770,N_47956,N_49165);
nand UO_1771 (O_1771,N_47140,N_47657);
nand UO_1772 (O_1772,N_49616,N_48407);
or UO_1773 (O_1773,N_48109,N_49489);
xnor UO_1774 (O_1774,N_48386,N_47613);
xor UO_1775 (O_1775,N_45319,N_49083);
nand UO_1776 (O_1776,N_45327,N_46423);
or UO_1777 (O_1777,N_46208,N_47861);
or UO_1778 (O_1778,N_49755,N_46315);
and UO_1779 (O_1779,N_48875,N_49912);
or UO_1780 (O_1780,N_45229,N_49396);
nand UO_1781 (O_1781,N_49746,N_49546);
or UO_1782 (O_1782,N_46310,N_47770);
or UO_1783 (O_1783,N_45474,N_46291);
nand UO_1784 (O_1784,N_47224,N_49853);
xor UO_1785 (O_1785,N_49079,N_48895);
nand UO_1786 (O_1786,N_46176,N_48139);
nand UO_1787 (O_1787,N_45876,N_46426);
nor UO_1788 (O_1788,N_49720,N_48038);
xor UO_1789 (O_1789,N_47947,N_46171);
nand UO_1790 (O_1790,N_47827,N_47949);
or UO_1791 (O_1791,N_48484,N_49898);
xor UO_1792 (O_1792,N_48558,N_45162);
or UO_1793 (O_1793,N_46223,N_47915);
or UO_1794 (O_1794,N_45152,N_47690);
and UO_1795 (O_1795,N_47455,N_46305);
xor UO_1796 (O_1796,N_49966,N_45223);
nand UO_1797 (O_1797,N_48330,N_48825);
or UO_1798 (O_1798,N_45626,N_45817);
nor UO_1799 (O_1799,N_47874,N_47538);
or UO_1800 (O_1800,N_46147,N_49943);
and UO_1801 (O_1801,N_48966,N_48578);
or UO_1802 (O_1802,N_49288,N_47532);
xnor UO_1803 (O_1803,N_48995,N_47460);
and UO_1804 (O_1804,N_48996,N_46519);
xor UO_1805 (O_1805,N_47024,N_49332);
xor UO_1806 (O_1806,N_49957,N_46931);
nand UO_1807 (O_1807,N_45777,N_49897);
nand UO_1808 (O_1808,N_47209,N_48961);
nor UO_1809 (O_1809,N_46417,N_49591);
xor UO_1810 (O_1810,N_46903,N_46401);
nand UO_1811 (O_1811,N_48028,N_45836);
nor UO_1812 (O_1812,N_45246,N_48795);
nor UO_1813 (O_1813,N_48541,N_48686);
nor UO_1814 (O_1814,N_46687,N_45992);
and UO_1815 (O_1815,N_48467,N_45499);
xnor UO_1816 (O_1816,N_48678,N_49082);
xor UO_1817 (O_1817,N_48434,N_46068);
or UO_1818 (O_1818,N_46020,N_48448);
or UO_1819 (O_1819,N_48914,N_46203);
nor UO_1820 (O_1820,N_46135,N_48951);
nand UO_1821 (O_1821,N_47834,N_47388);
or UO_1822 (O_1822,N_46914,N_49344);
nor UO_1823 (O_1823,N_47029,N_47109);
nand UO_1824 (O_1824,N_45316,N_46860);
nor UO_1825 (O_1825,N_47265,N_45398);
nand UO_1826 (O_1826,N_45584,N_47203);
or UO_1827 (O_1827,N_46629,N_47127);
nor UO_1828 (O_1828,N_48276,N_45190);
nand UO_1829 (O_1829,N_46943,N_46355);
xor UO_1830 (O_1830,N_48397,N_47046);
or UO_1831 (O_1831,N_48136,N_48881);
nand UO_1832 (O_1832,N_48503,N_46452);
nand UO_1833 (O_1833,N_47197,N_49571);
nand UO_1834 (O_1834,N_49035,N_48712);
and UO_1835 (O_1835,N_47853,N_48571);
and UO_1836 (O_1836,N_47820,N_47906);
xnor UO_1837 (O_1837,N_46815,N_49631);
nor UO_1838 (O_1838,N_48516,N_45877);
and UO_1839 (O_1839,N_49268,N_49074);
or UO_1840 (O_1840,N_47470,N_46599);
and UO_1841 (O_1841,N_49951,N_45295);
or UO_1842 (O_1842,N_46618,N_45389);
and UO_1843 (O_1843,N_49272,N_45055);
nor UO_1844 (O_1844,N_46694,N_46264);
xnor UO_1845 (O_1845,N_49714,N_46002);
or UO_1846 (O_1846,N_49462,N_48953);
nor UO_1847 (O_1847,N_47903,N_45302);
or UO_1848 (O_1848,N_48874,N_49561);
or UO_1849 (O_1849,N_49005,N_46295);
or UO_1850 (O_1850,N_45506,N_45721);
and UO_1851 (O_1851,N_45648,N_45761);
xnor UO_1852 (O_1852,N_45371,N_48257);
nor UO_1853 (O_1853,N_46097,N_48805);
nor UO_1854 (O_1854,N_47336,N_47491);
and UO_1855 (O_1855,N_46514,N_45887);
nor UO_1856 (O_1856,N_49716,N_47091);
and UO_1857 (O_1857,N_45619,N_49840);
xor UO_1858 (O_1858,N_46001,N_48717);
xnor UO_1859 (O_1859,N_47069,N_47748);
or UO_1860 (O_1860,N_47350,N_46647);
nor UO_1861 (O_1861,N_46628,N_47810);
xnor UO_1862 (O_1862,N_45649,N_45211);
nand UO_1863 (O_1863,N_46800,N_45687);
nor UO_1864 (O_1864,N_46416,N_48446);
nand UO_1865 (O_1865,N_45403,N_45355);
nor UO_1866 (O_1866,N_48480,N_48819);
nor UO_1867 (O_1867,N_47003,N_48530);
nand UO_1868 (O_1868,N_48387,N_45482);
xnor UO_1869 (O_1869,N_47740,N_46795);
or UO_1870 (O_1870,N_47073,N_47745);
and UO_1871 (O_1871,N_49617,N_46045);
xnor UO_1872 (O_1872,N_48540,N_48292);
nor UO_1873 (O_1873,N_49244,N_46463);
or UO_1874 (O_1874,N_47353,N_48063);
nand UO_1875 (O_1875,N_47563,N_46412);
nor UO_1876 (O_1876,N_45846,N_46138);
and UO_1877 (O_1877,N_45552,N_46648);
nand UO_1878 (O_1878,N_47242,N_45709);
and UO_1879 (O_1879,N_48811,N_47880);
xor UO_1880 (O_1880,N_49641,N_45182);
xor UO_1881 (O_1881,N_46303,N_48876);
nand UO_1882 (O_1882,N_49668,N_47894);
or UO_1883 (O_1883,N_48012,N_49909);
nand UO_1884 (O_1884,N_49834,N_49767);
and UO_1885 (O_1885,N_49072,N_49457);
nand UO_1886 (O_1886,N_49134,N_46605);
and UO_1887 (O_1887,N_46479,N_48721);
and UO_1888 (O_1888,N_46021,N_48148);
xor UO_1889 (O_1889,N_48614,N_47346);
nor UO_1890 (O_1890,N_47434,N_46182);
nor UO_1891 (O_1891,N_48921,N_49858);
nand UO_1892 (O_1892,N_46265,N_48186);
nor UO_1893 (O_1893,N_45587,N_49742);
nand UO_1894 (O_1894,N_45588,N_46710);
and UO_1895 (O_1895,N_46926,N_49925);
and UO_1896 (O_1896,N_45860,N_47136);
and UO_1897 (O_1897,N_48919,N_47833);
nor UO_1898 (O_1898,N_48499,N_46297);
or UO_1899 (O_1899,N_48696,N_46488);
nor UO_1900 (O_1900,N_47375,N_46534);
and UO_1901 (O_1901,N_48198,N_45991);
nand UO_1902 (O_1902,N_47692,N_49322);
nor UO_1903 (O_1903,N_45973,N_48083);
and UO_1904 (O_1904,N_47986,N_49263);
or UO_1905 (O_1905,N_47955,N_46286);
nand UO_1906 (O_1906,N_48100,N_47014);
nand UO_1907 (O_1907,N_45244,N_47131);
and UO_1908 (O_1908,N_49340,N_47600);
nor UO_1909 (O_1909,N_45865,N_47135);
xor UO_1910 (O_1910,N_47041,N_46134);
or UO_1911 (O_1911,N_45237,N_45058);
nand UO_1912 (O_1912,N_45821,N_49707);
xor UO_1913 (O_1913,N_45930,N_49077);
or UO_1914 (O_1914,N_46153,N_48638);
nand UO_1915 (O_1915,N_46024,N_48201);
or UO_1916 (O_1916,N_49822,N_45574);
or UO_1917 (O_1917,N_45700,N_45008);
nor UO_1918 (O_1918,N_46083,N_49350);
xnor UO_1919 (O_1919,N_45842,N_45769);
or UO_1920 (O_1920,N_49068,N_49778);
xnor UO_1921 (O_1921,N_48894,N_49768);
nand UO_1922 (O_1922,N_46947,N_47995);
and UO_1923 (O_1923,N_46507,N_45806);
and UO_1924 (O_1924,N_47759,N_49025);
or UO_1925 (O_1925,N_47699,N_46743);
xnor UO_1926 (O_1926,N_47572,N_47479);
or UO_1927 (O_1927,N_46644,N_49615);
xor UO_1928 (O_1928,N_49038,N_46724);
or UO_1929 (O_1929,N_45356,N_45330);
xnor UO_1930 (O_1930,N_48106,N_45165);
nand UO_1931 (O_1931,N_49986,N_49143);
xnor UO_1932 (O_1932,N_46726,N_48384);
or UO_1933 (O_1933,N_47673,N_46816);
and UO_1934 (O_1934,N_45290,N_45293);
and UO_1935 (O_1935,N_49020,N_48475);
nor UO_1936 (O_1936,N_49123,N_46763);
and UO_1937 (O_1937,N_49017,N_46168);
or UO_1938 (O_1938,N_47815,N_46041);
nor UO_1939 (O_1939,N_48027,N_48289);
xor UO_1940 (O_1940,N_45215,N_48685);
nor UO_1941 (O_1941,N_45103,N_45840);
and UO_1942 (O_1942,N_46730,N_49652);
and UO_1943 (O_1943,N_48361,N_49410);
and UO_1944 (O_1944,N_48157,N_48915);
or UO_1945 (O_1945,N_45689,N_47355);
and UO_1946 (O_1946,N_46234,N_47565);
nand UO_1947 (O_1947,N_45345,N_45833);
or UO_1948 (O_1948,N_47106,N_48590);
or UO_1949 (O_1949,N_45007,N_46125);
xor UO_1950 (O_1950,N_47590,N_47983);
xnor UO_1951 (O_1951,N_45885,N_49386);
xnor UO_1952 (O_1952,N_45276,N_47940);
nor UO_1953 (O_1953,N_46716,N_48159);
nand UO_1954 (O_1954,N_48017,N_46311);
or UO_1955 (O_1955,N_46099,N_45245);
xor UO_1956 (O_1956,N_45802,N_46890);
nor UO_1957 (O_1957,N_45694,N_49960);
or UO_1958 (O_1958,N_46434,N_46117);
and UO_1959 (O_1959,N_48327,N_47472);
nand UO_1960 (O_1960,N_49544,N_47196);
nand UO_1961 (O_1961,N_45210,N_46377);
or UO_1962 (O_1962,N_49135,N_45109);
nand UO_1963 (O_1963,N_47762,N_46621);
nor UO_1964 (O_1964,N_47031,N_48156);
nor UO_1965 (O_1965,N_49164,N_49337);
nand UO_1966 (O_1966,N_49730,N_47153);
nand UO_1967 (O_1967,N_46684,N_45360);
nor UO_1968 (O_1968,N_49691,N_46080);
and UO_1969 (O_1969,N_47503,N_47179);
nor UO_1970 (O_1970,N_48388,N_45035);
and UO_1971 (O_1971,N_46821,N_45149);
nand UO_1972 (O_1972,N_47609,N_47615);
nor UO_1973 (O_1973,N_49479,N_49700);
nand UO_1974 (O_1974,N_45033,N_46750);
and UO_1975 (O_1975,N_47803,N_46052);
or UO_1976 (O_1976,N_45249,N_45377);
or UO_1977 (O_1977,N_48693,N_46994);
and UO_1978 (O_1978,N_45265,N_46660);
nand UO_1979 (O_1979,N_48826,N_46346);
nor UO_1980 (O_1980,N_46430,N_48984);
and UO_1981 (O_1981,N_47268,N_46946);
nor UO_1982 (O_1982,N_45888,N_45548);
xnor UO_1983 (O_1983,N_49993,N_47089);
nor UO_1984 (O_1984,N_48433,N_45916);
or UO_1985 (O_1985,N_45591,N_49428);
and UO_1986 (O_1986,N_46472,N_46971);
and UO_1987 (O_1987,N_49119,N_49415);
and UO_1988 (O_1988,N_48485,N_45153);
xnor UO_1989 (O_1989,N_49574,N_47362);
and UO_1990 (O_1990,N_49814,N_47556);
nor UO_1991 (O_1991,N_49458,N_46319);
nor UO_1992 (O_1992,N_48086,N_49472);
and UO_1993 (O_1993,N_49576,N_46653);
xor UO_1994 (O_1994,N_45378,N_49587);
nand UO_1995 (O_1995,N_46554,N_47974);
nand UO_1996 (O_1996,N_46170,N_46391);
or UO_1997 (O_1997,N_48418,N_48498);
xor UO_1998 (O_1998,N_47619,N_45106);
xnor UO_1999 (O_1999,N_45115,N_47521);
nand UO_2000 (O_2000,N_45770,N_46189);
xor UO_2001 (O_2001,N_48217,N_47431);
or UO_2002 (O_2002,N_45257,N_46169);
nand UO_2003 (O_2003,N_46400,N_46280);
nor UO_2004 (O_2004,N_46934,N_46336);
xor UO_2005 (O_2005,N_48844,N_46161);
nor UO_2006 (O_2006,N_47805,N_46174);
or UO_2007 (O_2007,N_45233,N_46861);
nand UO_2008 (O_2008,N_47536,N_49122);
or UO_2009 (O_2009,N_49687,N_47202);
xor UO_2010 (O_2010,N_47311,N_49658);
and UO_2011 (O_2011,N_46373,N_48191);
or UO_2012 (O_2012,N_45993,N_45758);
nor UO_2013 (O_2013,N_49972,N_49545);
nand UO_2014 (O_2014,N_46975,N_45248);
nor UO_2015 (O_2015,N_46179,N_47189);
xnor UO_2016 (O_2016,N_46874,N_46703);
and UO_2017 (O_2017,N_46797,N_47379);
xor UO_2018 (O_2018,N_48183,N_46667);
nor UO_2019 (O_2019,N_47621,N_45495);
and UO_2020 (O_2020,N_47439,N_45767);
or UO_2021 (O_2021,N_48315,N_46086);
and UO_2022 (O_2022,N_45256,N_45564);
or UO_2023 (O_2023,N_48452,N_46249);
or UO_2024 (O_2024,N_48982,N_47500);
and UO_2025 (O_2025,N_45086,N_45270);
nand UO_2026 (O_2026,N_46826,N_48533);
xnor UO_2027 (O_2027,N_47534,N_45754);
or UO_2028 (O_2028,N_49423,N_48060);
and UO_2029 (O_2029,N_48158,N_47549);
nand UO_2030 (O_2030,N_47213,N_49253);
nor UO_2031 (O_2031,N_48422,N_47037);
or UO_2032 (O_2032,N_47542,N_45188);
nand UO_2033 (O_2033,N_48037,N_45949);
and UO_2034 (O_2034,N_45044,N_45730);
xor UO_2035 (O_2035,N_47591,N_46932);
nor UO_2036 (O_2036,N_47817,N_46285);
nor UO_2037 (O_2037,N_48901,N_46878);
nor UO_2038 (O_2038,N_47042,N_49008);
xor UO_2039 (O_2039,N_48243,N_47645);
nand UO_2040 (O_2040,N_46540,N_47996);
nor UO_2041 (O_2041,N_45565,N_48858);
nand UO_2042 (O_2042,N_48286,N_46770);
nand UO_2043 (O_2043,N_49098,N_47383);
or UO_2044 (O_2044,N_47095,N_47065);
nor UO_2045 (O_2045,N_46222,N_49429);
nor UO_2046 (O_2046,N_46966,N_45314);
nand UO_2047 (O_2047,N_46967,N_45280);
xor UO_2048 (O_2048,N_47772,N_49120);
xor UO_2049 (O_2049,N_46510,N_45717);
nor UO_2050 (O_2050,N_48627,N_47430);
and UO_2051 (O_2051,N_46631,N_45724);
xnor UO_2052 (O_2052,N_46013,N_47260);
nand UO_2053 (O_2053,N_49952,N_47888);
nand UO_2054 (O_2054,N_49371,N_46178);
or UO_2055 (O_2055,N_45570,N_48486);
or UO_2056 (O_2056,N_46964,N_45630);
nand UO_2057 (O_2057,N_46867,N_45368);
xnor UO_2058 (O_2058,N_46924,N_48888);
or UO_2059 (O_2059,N_45181,N_47633);
nand UO_2060 (O_2060,N_48746,N_47719);
and UO_2061 (O_2061,N_47134,N_48058);
xor UO_2062 (O_2062,N_46016,N_47110);
or UO_2063 (O_2063,N_45731,N_47720);
xnor UO_2064 (O_2064,N_45845,N_49145);
nand UO_2065 (O_2065,N_48236,N_47652);
and UO_2066 (O_2066,N_48969,N_47427);
nand UO_2067 (O_2067,N_49342,N_48287);
and UO_2068 (O_2068,N_48785,N_48871);
or UO_2069 (O_2069,N_46838,N_49510);
and UO_2070 (O_2070,N_48162,N_48375);
nand UO_2071 (O_2071,N_49567,N_47352);
xnor UO_2072 (O_2072,N_46897,N_47038);
nand UO_2073 (O_2073,N_46043,N_48142);
nor UO_2074 (O_2074,N_47272,N_49808);
and UO_2075 (O_2075,N_49555,N_48545);
nand UO_2076 (O_2076,N_47171,N_46854);
or UO_2077 (O_2077,N_47282,N_48230);
nand UO_2078 (O_2078,N_49642,N_47716);
or UO_2079 (O_2079,N_48469,N_47380);
xor UO_2080 (O_2080,N_45099,N_45019);
xor UO_2081 (O_2081,N_49842,N_48291);
or UO_2082 (O_2082,N_46284,N_47066);
and UO_2083 (O_2083,N_46753,N_47498);
or UO_2084 (O_2084,N_49484,N_46344);
or UO_2085 (O_2085,N_47044,N_45243);
and UO_2086 (O_2086,N_48444,N_48813);
nor UO_2087 (O_2087,N_46141,N_49185);
nand UO_2088 (O_2088,N_48529,N_48865);
or UO_2089 (O_2089,N_47540,N_49863);
or UO_2090 (O_2090,N_49879,N_45571);
nand UO_2091 (O_2091,N_47221,N_49341);
and UO_2092 (O_2092,N_47991,N_49431);
or UO_2093 (O_2093,N_48781,N_46799);
nand UO_2094 (O_2094,N_47364,N_48652);
nor UO_2095 (O_2095,N_45275,N_47484);
xor UO_2096 (O_2096,N_46689,N_45963);
nand UO_2097 (O_2097,N_47216,N_49426);
and UO_2098 (O_2098,N_46663,N_48568);
or UO_2099 (O_2099,N_48644,N_49321);
xor UO_2100 (O_2100,N_47297,N_45110);
nor UO_2101 (O_2101,N_45854,N_45708);
and UO_2102 (O_2102,N_48080,N_46388);
nor UO_2103 (O_2103,N_48479,N_46308);
nand UO_2104 (O_2104,N_49307,N_49874);
and UO_2105 (O_2105,N_46889,N_48009);
nor UO_2106 (O_2106,N_47176,N_45251);
nand UO_2107 (O_2107,N_45812,N_47137);
or UO_2108 (O_2108,N_46536,N_48625);
or UO_2109 (O_2109,N_46979,N_46365);
and UO_2110 (O_2110,N_49153,N_45087);
nand UO_2111 (O_2111,N_47229,N_47507);
nor UO_2112 (O_2112,N_46697,N_46669);
or UO_2113 (O_2113,N_46195,N_49302);
nand UO_2114 (O_2114,N_45379,N_49674);
nand UO_2115 (O_2115,N_46764,N_46051);
and UO_2116 (O_2116,N_45301,N_46910);
nand UO_2117 (O_2117,N_46871,N_47191);
nor UO_2118 (O_2118,N_49864,N_46250);
xnor UO_2119 (O_2119,N_48544,N_45659);
nor UO_2120 (O_2120,N_47257,N_46546);
nand UO_2121 (O_2121,N_49995,N_45228);
nor UO_2122 (O_2122,N_46193,N_48343);
nand UO_2123 (O_2123,N_46483,N_49016);
and UO_2124 (O_2124,N_49131,N_48056);
xnor UO_2125 (O_2125,N_46977,N_49500);
xnor UO_2126 (O_2126,N_49326,N_48552);
xnor UO_2127 (O_2127,N_46688,N_45970);
nor UO_2128 (O_2128,N_48932,N_45298);
and UO_2129 (O_2129,N_48456,N_45901);
and UO_2130 (O_2130,N_49014,N_47586);
xor UO_2131 (O_2131,N_48078,N_47048);
xnor UO_2132 (O_2132,N_45698,N_45052);
nor UO_2133 (O_2133,N_46851,N_48757);
xor UO_2134 (O_2134,N_45514,N_48527);
and UO_2135 (O_2135,N_45042,N_47860);
xnor UO_2136 (O_2136,N_49811,N_45297);
nor UO_2137 (O_2137,N_45205,N_48661);
and UO_2138 (O_2138,N_46919,N_47080);
nand UO_2139 (O_2139,N_47900,N_49860);
xnor UO_2140 (O_2140,N_48587,N_48171);
nand UO_2141 (O_2141,N_45437,N_49026);
xor UO_2142 (O_2142,N_45169,N_49942);
nand UO_2143 (O_2143,N_49358,N_47680);
nand UO_2144 (O_2144,N_48800,N_46901);
xnor UO_2145 (O_2145,N_48232,N_49590);
nor UO_2146 (O_2146,N_47267,N_45098);
nor UO_2147 (O_2147,N_49354,N_47753);
nand UO_2148 (O_2148,N_47773,N_48740);
nor UO_2149 (O_2149,N_47892,N_45180);
nand UO_2150 (O_2150,N_45737,N_45449);
and UO_2151 (O_2151,N_47252,N_47963);
nor UO_2152 (O_2152,N_49949,N_46894);
and UO_2153 (O_2153,N_49282,N_48906);
xor UO_2154 (O_2154,N_48074,N_46239);
xnor UO_2155 (O_2155,N_48710,N_47411);
and UO_2156 (O_2156,N_49161,N_46645);
or UO_2157 (O_2157,N_49638,N_46792);
nand UO_2158 (O_2158,N_48356,N_48968);
and UO_2159 (O_2159,N_47215,N_45430);
or UO_2160 (O_2160,N_46009,N_47678);
nand UO_2161 (O_2161,N_48483,N_49180);
nor UO_2162 (O_2162,N_48551,N_48297);
and UO_2163 (O_2163,N_47771,N_46231);
nand UO_2164 (O_2164,N_49477,N_49209);
nor UO_2165 (O_2165,N_49170,N_47338);
xnor UO_2166 (O_2166,N_45002,N_48366);
or UO_2167 (O_2167,N_46614,N_48065);
nand UO_2168 (O_2168,N_47879,N_49688);
or UO_2169 (O_2169,N_45987,N_47750);
or UO_2170 (O_2170,N_47709,N_48520);
and UO_2171 (O_2171,N_48754,N_49786);
and UO_2172 (O_2172,N_49040,N_45063);
nor UO_2173 (O_2173,N_46532,N_49275);
and UO_2174 (O_2174,N_48744,N_45287);
nor UO_2175 (O_2175,N_47094,N_45977);
xor UO_2176 (O_2176,N_48991,N_45231);
nand UO_2177 (O_2177,N_47159,N_49680);
nor UO_2178 (O_2178,N_47021,N_45034);
nor UO_2179 (O_2179,N_47850,N_49202);
nor UO_2180 (O_2180,N_47097,N_48839);
xor UO_2181 (O_2181,N_49039,N_45511);
xor UO_2182 (O_2182,N_47237,N_48087);
nor UO_2183 (O_2183,N_49682,N_47665);
xnor UO_2184 (O_2184,N_48613,N_45416);
nor UO_2185 (O_2185,N_48790,N_49451);
and UO_2186 (O_2186,N_48451,N_46209);
nor UO_2187 (O_2187,N_45077,N_46092);
or UO_2188 (O_2188,N_47371,N_49409);
nand UO_2189 (O_2189,N_45667,N_49706);
nand UO_2190 (O_2190,N_49517,N_45272);
and UO_2191 (O_2191,N_48585,N_48329);
nor UO_2192 (O_2192,N_49086,N_48112);
nor UO_2193 (O_2193,N_49387,N_47047);
or UO_2194 (O_2194,N_45417,N_45549);
or UO_2195 (O_2195,N_48325,N_46317);
and UO_2196 (O_2196,N_49405,N_47115);
nand UO_2197 (O_2197,N_46087,N_48955);
or UO_2198 (O_2198,N_46639,N_47318);
or UO_2199 (O_2199,N_48071,N_46522);
and UO_2200 (O_2200,N_46923,N_48864);
xnor UO_2201 (O_2201,N_49632,N_48615);
xnor UO_2202 (O_2202,N_46965,N_48632);
and UO_2203 (O_2203,N_46419,N_48210);
xnor UO_2204 (O_2204,N_49835,N_49254);
nor UO_2205 (O_2205,N_48594,N_49754);
or UO_2206 (O_2206,N_46909,N_47334);
nor UO_2207 (O_2207,N_48787,N_47019);
xnor UO_2208 (O_2208,N_47435,N_48298);
nand UO_2209 (O_2209,N_46033,N_49828);
or UO_2210 (O_2210,N_46062,N_45200);
or UO_2211 (O_2211,N_45931,N_49927);
nor UO_2212 (O_2212,N_47456,N_47868);
xor UO_2213 (O_2213,N_48459,N_48682);
or UO_2214 (O_2214,N_48927,N_48603);
nor UO_2215 (O_2215,N_46893,N_45807);
or UO_2216 (O_2216,N_49531,N_47984);
or UO_2217 (O_2217,N_46754,N_47258);
or UO_2218 (O_2218,N_46000,N_46408);
or UO_2219 (O_2219,N_47169,N_47597);
nor UO_2220 (O_2220,N_47463,N_47797);
nand UO_2221 (O_2221,N_45066,N_47669);
nand UO_2222 (O_2222,N_49667,N_47422);
nand UO_2223 (O_2223,N_48254,N_49385);
xor UO_2224 (O_2224,N_46090,N_47255);
or UO_2225 (O_2225,N_48494,N_46732);
nor UO_2226 (O_2226,N_47499,N_45647);
and UO_2227 (O_2227,N_48926,N_45122);
nand UO_2228 (O_2228,N_46186,N_48878);
and UO_2229 (O_2229,N_48450,N_46259);
or UO_2230 (O_2230,N_46950,N_45599);
and UO_2231 (O_2231,N_45809,N_45124);
xor UO_2232 (O_2232,N_48992,N_48838);
and UO_2233 (O_2233,N_48812,N_46151);
xor UO_2234 (O_2234,N_49764,N_49788);
nand UO_2235 (O_2235,N_45856,N_48323);
or UO_2236 (O_2236,N_49418,N_47951);
or UO_2237 (O_2237,N_49201,N_49921);
xor UO_2238 (O_2238,N_49630,N_47017);
and UO_2239 (O_2239,N_47347,N_48166);
nor UO_2240 (O_2240,N_45353,N_46348);
or UO_2241 (O_2241,N_46424,N_46495);
xor UO_2242 (O_2242,N_49376,N_49758);
xor UO_2243 (O_2243,N_48902,N_45139);
and UO_2244 (O_2244,N_47587,N_45148);
or UO_2245 (O_2245,N_47138,N_45435);
or UO_2246 (O_2246,N_45939,N_47320);
xnor UO_2247 (O_2247,N_47899,N_46228);
and UO_2248 (O_2248,N_47582,N_46557);
nor UO_2249 (O_2249,N_47384,N_46696);
nand UO_2250 (O_2250,N_45123,N_48302);
nor UO_2251 (O_2251,N_49092,N_45898);
or UO_2252 (O_2252,N_49625,N_49543);
or UO_2253 (O_2253,N_46604,N_46715);
nor UO_2254 (O_2254,N_49205,N_46202);
nand UO_2255 (O_2255,N_46487,N_47674);
nor UO_2256 (O_2256,N_46970,N_45695);
xor UO_2257 (O_2257,N_46953,N_47084);
xnor UO_2258 (O_2258,N_48677,N_48116);
and UO_2259 (O_2259,N_48035,N_47778);
or UO_2260 (O_2260,N_46453,N_48596);
nand UO_2261 (O_2261,N_46382,N_46957);
nand UO_2262 (O_2262,N_45128,N_45341);
xnor UO_2263 (O_2263,N_47610,N_49537);
nor UO_2264 (O_2264,N_47554,N_47857);
and UO_2265 (O_2265,N_47280,N_48476);
nor UO_2266 (O_2266,N_45284,N_46225);
and UO_2267 (O_2267,N_45473,N_49599);
nor UO_2268 (O_2268,N_46529,N_49963);
nor UO_2269 (O_2269,N_45202,N_47078);
xnor UO_2270 (O_2270,N_49149,N_48506);
nand UO_2271 (O_2271,N_46497,N_46358);
nor UO_2272 (O_2272,N_49813,N_49893);
nand UO_2273 (O_2273,N_46600,N_45458);
xor UO_2274 (O_2274,N_46622,N_47007);
nand UO_2275 (O_2275,N_49818,N_45874);
nor UO_2276 (O_2276,N_48681,N_46251);
nand UO_2277 (O_2277,N_48079,N_47844);
nand UO_2278 (O_2278,N_49245,N_47158);
and UO_2279 (O_2279,N_48928,N_45582);
nand UO_2280 (O_2280,N_45826,N_46370);
or UO_2281 (O_2281,N_49313,N_46482);
nor UO_2282 (O_2282,N_45965,N_49179);
xnor UO_2283 (O_2283,N_45155,N_47198);
nor UO_2284 (O_2284,N_48130,N_45500);
xnor UO_2285 (O_2285,N_47093,N_47647);
or UO_2286 (O_2286,N_49773,N_46047);
and UO_2287 (O_2287,N_48263,N_46341);
nor UO_2288 (O_2288,N_47283,N_47637);
xnor UO_2289 (O_2289,N_45306,N_47804);
nand UO_2290 (O_2290,N_47182,N_46361);
or UO_2291 (O_2291,N_47289,N_49105);
nor UO_2292 (O_2292,N_47010,N_49284);
and UO_2293 (O_2293,N_45568,N_47897);
or UO_2294 (O_2294,N_48004,N_47990);
or UO_2295 (O_2295,N_46973,N_46779);
nor UO_2296 (O_2296,N_45884,N_49021);
and UO_2297 (O_2297,N_47425,N_45852);
or UO_2298 (O_2298,N_47913,N_48314);
xnor UO_2299 (O_2299,N_48867,N_47039);
or UO_2300 (O_2300,N_49114,N_47235);
nand UO_2301 (O_2301,N_49507,N_48202);
nand UO_2302 (O_2302,N_48264,N_48940);
nand UO_2303 (O_2303,N_47496,N_46095);
xor UO_2304 (O_2304,N_49911,N_49777);
and UO_2305 (O_2305,N_49597,N_47471);
or UO_2306 (O_2306,N_49888,N_46680);
nor UO_2307 (O_2307,N_48803,N_46456);
nor UO_2308 (O_2308,N_49304,N_45771);
nor UO_2309 (O_2309,N_46635,N_47015);
nor UO_2310 (O_2310,N_48730,N_46268);
nand UO_2311 (O_2311,N_46154,N_47849);
and UO_2312 (O_2312,N_45225,N_48988);
or UO_2313 (O_2313,N_45138,N_45015);
and UO_2314 (O_2314,N_45450,N_46337);
and UO_2315 (O_2315,N_45544,N_49217);
or UO_2316 (O_2316,N_47774,N_45440);
xnor UO_2317 (O_2317,N_46809,N_47742);
or UO_2318 (O_2318,N_47526,N_45382);
or UO_2319 (O_2319,N_47741,N_46556);
or UO_2320 (O_2320,N_48597,N_47387);
xor UO_2321 (O_2321,N_49907,N_46360);
xnor UO_2322 (O_2322,N_49206,N_46146);
and UO_2323 (O_2323,N_47918,N_49839);
and UO_2324 (O_2324,N_46711,N_48029);
or UO_2325 (O_2325,N_47662,N_45605);
xor UO_2326 (O_2326,N_48307,N_47729);
or UO_2327 (O_2327,N_48863,N_48671);
or UO_2328 (O_2328,N_47763,N_45258);
and UO_2329 (O_2329,N_49163,N_46276);
nor UO_2330 (O_2330,N_49870,N_48117);
xnor UO_2331 (O_2331,N_47898,N_45725);
xnor UO_2332 (O_2332,N_49171,N_46290);
nand UO_2333 (O_2333,N_48320,N_49936);
nor UO_2334 (O_2334,N_46912,N_45026);
xor UO_2335 (O_2335,N_49441,N_48985);
and UO_2336 (O_2336,N_49330,N_46025);
and UO_2337 (O_2337,N_47505,N_45238);
and UO_2338 (O_2338,N_45013,N_46504);
and UO_2339 (O_2339,N_47808,N_46444);
nor UO_2340 (O_2340,N_48518,N_45950);
nor UO_2341 (O_2341,N_47698,N_48043);
and UO_2342 (O_2342,N_46192,N_49352);
nor UO_2343 (O_2343,N_48005,N_48849);
nor UO_2344 (O_2344,N_45050,N_49103);
xor UO_2345 (O_2345,N_47504,N_45323);
and UO_2346 (O_2346,N_46565,N_46112);
xor UO_2347 (O_2347,N_49572,N_45343);
nor UO_2348 (O_2348,N_48277,N_47929);
or UO_2349 (O_2349,N_45354,N_48783);
or UO_2350 (O_2350,N_46717,N_49186);
xnor UO_2351 (O_2351,N_49482,N_46959);
nand UO_2352 (O_2352,N_47276,N_47354);
and UO_2353 (O_2353,N_45173,N_45264);
xnor UO_2354 (O_2354,N_49107,N_46432);
xor UO_2355 (O_2355,N_47691,N_47357);
xor UO_2356 (O_2356,N_49588,N_47841);
nand UO_2357 (O_2357,N_48383,N_46283);
and UO_2358 (O_2358,N_45691,N_47934);
nor UO_2359 (O_2359,N_46029,N_49314);
nand UO_2360 (O_2360,N_49301,N_48419);
xor UO_2361 (O_2361,N_47474,N_48477);
nor UO_2362 (O_2362,N_47076,N_49605);
and UO_2363 (O_2363,N_46486,N_48716);
nor UO_2364 (O_2364,N_48823,N_47924);
and UO_2365 (O_2365,N_47642,N_46661);
nand UO_2366 (O_2366,N_49692,N_47593);
xnor UO_2367 (O_2367,N_47758,N_49247);
nand UO_2368 (O_2368,N_46655,N_49127);
xnor UO_2369 (O_2369,N_49868,N_48221);
xor UO_2370 (O_2370,N_48194,N_47008);
or UO_2371 (O_2371,N_45623,N_49836);
or UO_2372 (O_2372,N_48206,N_48152);
and UO_2373 (O_2373,N_47798,N_46378);
xor UO_2374 (O_2374,N_49899,N_48802);
nand UO_2375 (O_2375,N_45528,N_46187);
xor UO_2376 (O_2376,N_48197,N_46121);
nand UO_2377 (O_2377,N_49230,N_46450);
or UO_2378 (O_2378,N_49514,N_48962);
xor UO_2379 (O_2379,N_48808,N_47303);
nand UO_2380 (O_2380,N_49904,N_47428);
xor UO_2381 (O_2381,N_45399,N_46438);
nor UO_2382 (O_2382,N_46620,N_47603);
nand UO_2383 (O_2383,N_46656,N_49097);
xnor UO_2384 (O_2384,N_48108,N_45491);
nor UO_2385 (O_2385,N_49478,N_47188);
and UO_2386 (O_2386,N_48165,N_46244);
nor UO_2387 (O_2387,N_45505,N_46749);
or UO_2388 (O_2388,N_48589,N_46891);
or UO_2389 (O_2389,N_48064,N_45405);
nor UO_2390 (O_2390,N_48581,N_46089);
nor UO_2391 (O_2391,N_47599,N_46518);
nor UO_2392 (O_2392,N_48934,N_48231);
and UO_2393 (O_2393,N_48664,N_46802);
nand UO_2394 (O_2394,N_46761,N_49612);
and UO_2395 (O_2395,N_45920,N_45526);
and UO_2396 (O_2396,N_48588,N_45439);
or UO_2397 (O_2397,N_45266,N_49542);
nand UO_2398 (O_2398,N_48280,N_47452);
and UO_2399 (O_2399,N_46723,N_46780);
nand UO_2400 (O_2400,N_49345,N_47601);
and UO_2401 (O_2401,N_48014,N_45292);
or UO_2402 (O_2402,N_48547,N_46825);
nand UO_2403 (O_2403,N_46649,N_49979);
nor UO_2404 (O_2404,N_48804,N_45555);
nor UO_2405 (O_2405,N_49192,N_45838);
or UO_2406 (O_2406,N_45546,N_48401);
nor UO_2407 (O_2407,N_47509,N_45322);
or UO_2408 (O_2408,N_46333,N_48195);
nand UO_2409 (O_2409,N_45351,N_48706);
xnor UO_2410 (O_2410,N_47055,N_45800);
nor UO_2411 (O_2411,N_46343,N_45798);
xnor UO_2412 (O_2412,N_47005,N_45434);
and UO_2413 (O_2413,N_49582,N_46745);
nor UO_2414 (O_2414,N_48170,N_49881);
xnor UO_2415 (O_2415,N_48909,N_45310);
or UO_2416 (O_2416,N_47706,N_46999);
and UO_2417 (O_2417,N_48272,N_49208);
and UO_2418 (O_2418,N_48861,N_46454);
and UO_2419 (O_2419,N_47982,N_45707);
or UO_2420 (O_2420,N_48259,N_45935);
and UO_2421 (O_2421,N_49793,N_48662);
nand UO_2422 (O_2422,N_45536,N_48410);
nand UO_2423 (O_2423,N_46435,N_48428);
and UO_2424 (O_2424,N_49290,N_49540);
nor UO_2425 (O_2425,N_47802,N_49147);
nand UO_2426 (O_2426,N_45988,N_48633);
nand UO_2427 (O_2427,N_46328,N_49132);
nand UO_2428 (O_2428,N_47596,N_45102);
xor UO_2429 (O_2429,N_45690,N_49075);
and UO_2430 (O_2430,N_48070,N_47205);
nor UO_2431 (O_2431,N_47261,N_49548);
nor UO_2432 (O_2432,N_46255,N_49024);
xor UO_2433 (O_2433,N_45170,N_46997);
and UO_2434 (O_2434,N_48218,N_46658);
xor UO_2435 (O_2435,N_48367,N_49794);
nor UO_2436 (O_2436,N_47451,N_45336);
and UO_2437 (O_2437,N_45503,N_48082);
xnor UO_2438 (O_2438,N_47794,N_47902);
and UO_2439 (O_2439,N_45960,N_49916);
nand UO_2440 (O_2440,N_49262,N_45655);
nand UO_2441 (O_2441,N_46612,N_45235);
or UO_2442 (O_2442,N_49628,N_48728);
nor UO_2443 (O_2443,N_46503,N_49686);
or UO_2444 (O_2444,N_45038,N_49485);
nor UO_2445 (O_2445,N_48052,N_49744);
nor UO_2446 (O_2446,N_46132,N_49872);
nor UO_2447 (O_2447,N_46679,N_49675);
nor UO_2448 (O_2448,N_49573,N_45882);
and UO_2449 (O_2449,N_48495,N_48258);
or UO_2450 (O_2450,N_48729,N_46760);
or UO_2451 (O_2451,N_48882,N_47124);
nand UO_2452 (O_2452,N_45665,N_47515);
xor UO_2453 (O_2453,N_48379,N_48563);
nor UO_2454 (O_2454,N_49369,N_45595);
and UO_2455 (O_2455,N_47468,N_47971);
xor UO_2456 (O_2456,N_49985,N_46247);
nand UO_2457 (O_2457,N_49937,N_48491);
nor UO_2458 (O_2458,N_49442,N_49152);
nand UO_2459 (O_2459,N_49466,N_47574);
nand UO_2460 (O_2460,N_45751,N_48653);
nor UO_2461 (O_2461,N_49172,N_45762);
xnor UO_2462 (O_2462,N_48376,N_46126);
nand UO_2463 (O_2463,N_47697,N_48707);
and UO_2464 (O_2464,N_48462,N_49733);
nor UO_2465 (O_2465,N_45334,N_45394);
and UO_2466 (O_2466,N_45144,N_49375);
nor UO_2467 (O_2467,N_48830,N_47687);
nor UO_2468 (O_2468,N_49664,N_47584);
or UO_2469 (O_2469,N_45592,N_46925);
or UO_2470 (O_2470,N_49447,N_45289);
and UO_2471 (O_2471,N_47921,N_45216);
or UO_2472 (O_2472,N_45219,N_48394);
nand UO_2473 (O_2473,N_49775,N_46853);
xor UO_2474 (O_2474,N_49598,N_45713);
xnor UO_2475 (O_2475,N_47873,N_45146);
or UO_2476 (O_2476,N_47287,N_46744);
and UO_2477 (O_2477,N_45982,N_49795);
and UO_2478 (O_2478,N_45878,N_46589);
or UO_2479 (O_2479,N_47359,N_49207);
or UO_2480 (O_2480,N_48146,N_45813);
nand UO_2481 (O_2481,N_45747,N_47086);
nand UO_2482 (O_2482,N_49930,N_46918);
or UO_2483 (O_2483,N_46720,N_48267);
or UO_2484 (O_2484,N_47254,N_49015);
and UO_2485 (O_2485,N_48090,N_45081);
and UO_2486 (O_2486,N_49318,N_47162);
and UO_2487 (O_2487,N_48832,N_48033);
nand UO_2488 (O_2488,N_48538,N_46066);
and UO_2489 (O_2489,N_49237,N_49583);
nor UO_2490 (O_2490,N_48309,N_47397);
and UO_2491 (O_2491,N_47223,N_49070);
xor UO_2492 (O_2492,N_47273,N_47919);
or UO_2493 (O_2493,N_45529,N_48567);
nand UO_2494 (O_2494,N_45527,N_48782);
and UO_2495 (O_2495,N_49468,N_46752);
nor UO_2496 (O_2496,N_48659,N_45766);
and UO_2497 (O_2497,N_47953,N_47292);
xor UO_2498 (O_2498,N_48482,N_49656);
xor UO_2499 (O_2499,N_47643,N_45369);
xor UO_2500 (O_2500,N_47132,N_49890);
nor UO_2501 (O_2501,N_48735,N_49296);
nor UO_2502 (O_2502,N_49923,N_48272);
nand UO_2503 (O_2503,N_48109,N_48730);
nor UO_2504 (O_2504,N_45731,N_48059);
and UO_2505 (O_2505,N_47519,N_46299);
and UO_2506 (O_2506,N_49580,N_45479);
xor UO_2507 (O_2507,N_48652,N_46114);
or UO_2508 (O_2508,N_45631,N_47605);
and UO_2509 (O_2509,N_45201,N_49014);
and UO_2510 (O_2510,N_48854,N_47628);
nand UO_2511 (O_2511,N_49320,N_49072);
nand UO_2512 (O_2512,N_47973,N_46496);
xor UO_2513 (O_2513,N_49462,N_48452);
xor UO_2514 (O_2514,N_49934,N_49738);
or UO_2515 (O_2515,N_47070,N_47477);
nand UO_2516 (O_2516,N_49114,N_48107);
nor UO_2517 (O_2517,N_49206,N_47019);
nand UO_2518 (O_2518,N_47694,N_48212);
or UO_2519 (O_2519,N_46758,N_45429);
nand UO_2520 (O_2520,N_46938,N_47187);
nand UO_2521 (O_2521,N_49708,N_45401);
and UO_2522 (O_2522,N_48554,N_47188);
xnor UO_2523 (O_2523,N_49775,N_47361);
or UO_2524 (O_2524,N_47453,N_47072);
xor UO_2525 (O_2525,N_48659,N_48177);
or UO_2526 (O_2526,N_46578,N_45580);
and UO_2527 (O_2527,N_47144,N_47177);
or UO_2528 (O_2528,N_46109,N_45135);
nand UO_2529 (O_2529,N_45562,N_49087);
nand UO_2530 (O_2530,N_48102,N_47583);
and UO_2531 (O_2531,N_47130,N_46646);
and UO_2532 (O_2532,N_49316,N_46384);
and UO_2533 (O_2533,N_48696,N_49116);
nor UO_2534 (O_2534,N_46727,N_48187);
and UO_2535 (O_2535,N_45066,N_47227);
or UO_2536 (O_2536,N_48852,N_47344);
nor UO_2537 (O_2537,N_46762,N_49157);
nor UO_2538 (O_2538,N_48296,N_46479);
nand UO_2539 (O_2539,N_46095,N_45722);
nor UO_2540 (O_2540,N_45579,N_48218);
xor UO_2541 (O_2541,N_46504,N_49744);
nand UO_2542 (O_2542,N_45188,N_46900);
or UO_2543 (O_2543,N_45201,N_45574);
and UO_2544 (O_2544,N_47576,N_46752);
nand UO_2545 (O_2545,N_48068,N_45384);
and UO_2546 (O_2546,N_47625,N_45874);
or UO_2547 (O_2547,N_46360,N_47671);
and UO_2548 (O_2548,N_49477,N_46878);
nor UO_2549 (O_2549,N_48598,N_49553);
or UO_2550 (O_2550,N_47637,N_45537);
nor UO_2551 (O_2551,N_49890,N_49762);
nor UO_2552 (O_2552,N_49026,N_46993);
xor UO_2553 (O_2553,N_46741,N_48804);
and UO_2554 (O_2554,N_49875,N_47794);
nand UO_2555 (O_2555,N_49551,N_47200);
and UO_2556 (O_2556,N_46595,N_46567);
and UO_2557 (O_2557,N_46337,N_46357);
nor UO_2558 (O_2558,N_46604,N_47261);
nor UO_2559 (O_2559,N_48314,N_46574);
or UO_2560 (O_2560,N_45004,N_46335);
nor UO_2561 (O_2561,N_48008,N_49824);
nor UO_2562 (O_2562,N_46559,N_47078);
or UO_2563 (O_2563,N_46534,N_48442);
nand UO_2564 (O_2564,N_49155,N_46719);
and UO_2565 (O_2565,N_49119,N_49742);
and UO_2566 (O_2566,N_48602,N_49380);
and UO_2567 (O_2567,N_48365,N_47168);
and UO_2568 (O_2568,N_46478,N_47104);
and UO_2569 (O_2569,N_45999,N_45317);
or UO_2570 (O_2570,N_49038,N_45505);
and UO_2571 (O_2571,N_49930,N_48515);
nand UO_2572 (O_2572,N_46946,N_46340);
or UO_2573 (O_2573,N_47462,N_49323);
nand UO_2574 (O_2574,N_48246,N_45532);
xnor UO_2575 (O_2575,N_49639,N_46366);
or UO_2576 (O_2576,N_48655,N_48187);
nand UO_2577 (O_2577,N_48745,N_48972);
and UO_2578 (O_2578,N_45056,N_47912);
xor UO_2579 (O_2579,N_45476,N_45920);
or UO_2580 (O_2580,N_46703,N_46292);
nor UO_2581 (O_2581,N_47616,N_45437);
or UO_2582 (O_2582,N_47792,N_45550);
nor UO_2583 (O_2583,N_47761,N_49197);
or UO_2584 (O_2584,N_49329,N_49159);
and UO_2585 (O_2585,N_47785,N_49232);
or UO_2586 (O_2586,N_46549,N_46704);
xor UO_2587 (O_2587,N_46076,N_46844);
or UO_2588 (O_2588,N_45952,N_45690);
nand UO_2589 (O_2589,N_48701,N_49604);
and UO_2590 (O_2590,N_47337,N_47751);
nand UO_2591 (O_2591,N_47370,N_45101);
nor UO_2592 (O_2592,N_48008,N_49117);
xnor UO_2593 (O_2593,N_46075,N_47358);
and UO_2594 (O_2594,N_47643,N_45932);
or UO_2595 (O_2595,N_47331,N_47915);
nor UO_2596 (O_2596,N_47269,N_49224);
and UO_2597 (O_2597,N_46910,N_47780);
or UO_2598 (O_2598,N_49120,N_49715);
xor UO_2599 (O_2599,N_46412,N_45213);
nor UO_2600 (O_2600,N_48886,N_48517);
or UO_2601 (O_2601,N_49897,N_49394);
and UO_2602 (O_2602,N_45797,N_48288);
xnor UO_2603 (O_2603,N_45178,N_48173);
or UO_2604 (O_2604,N_49666,N_47115);
xor UO_2605 (O_2605,N_49463,N_45455);
nand UO_2606 (O_2606,N_47166,N_46882);
nor UO_2607 (O_2607,N_47458,N_48203);
or UO_2608 (O_2608,N_45873,N_46456);
xnor UO_2609 (O_2609,N_48187,N_49286);
nor UO_2610 (O_2610,N_46403,N_49669);
nand UO_2611 (O_2611,N_48742,N_46625);
and UO_2612 (O_2612,N_49336,N_48458);
and UO_2613 (O_2613,N_46470,N_45624);
nor UO_2614 (O_2614,N_47021,N_47593);
nand UO_2615 (O_2615,N_47308,N_46368);
nand UO_2616 (O_2616,N_47928,N_48684);
nand UO_2617 (O_2617,N_48304,N_45179);
and UO_2618 (O_2618,N_49752,N_49108);
and UO_2619 (O_2619,N_45472,N_48916);
nor UO_2620 (O_2620,N_47773,N_45498);
nor UO_2621 (O_2621,N_48907,N_47420);
and UO_2622 (O_2622,N_45583,N_48000);
and UO_2623 (O_2623,N_45372,N_45337);
and UO_2624 (O_2624,N_46504,N_48482);
nor UO_2625 (O_2625,N_49587,N_47550);
xnor UO_2626 (O_2626,N_49774,N_49694);
xnor UO_2627 (O_2627,N_48111,N_46669);
and UO_2628 (O_2628,N_45143,N_47625);
or UO_2629 (O_2629,N_47896,N_47333);
xnor UO_2630 (O_2630,N_49545,N_46080);
xnor UO_2631 (O_2631,N_46326,N_48608);
nand UO_2632 (O_2632,N_48186,N_47206);
nand UO_2633 (O_2633,N_48980,N_46535);
or UO_2634 (O_2634,N_48531,N_49619);
or UO_2635 (O_2635,N_45933,N_46494);
nor UO_2636 (O_2636,N_46202,N_49268);
or UO_2637 (O_2637,N_47165,N_47737);
and UO_2638 (O_2638,N_45708,N_45884);
nor UO_2639 (O_2639,N_49066,N_48582);
and UO_2640 (O_2640,N_45422,N_48833);
xor UO_2641 (O_2641,N_47392,N_45212);
nor UO_2642 (O_2642,N_47193,N_47780);
nand UO_2643 (O_2643,N_46547,N_47998);
and UO_2644 (O_2644,N_48299,N_49948);
nor UO_2645 (O_2645,N_45443,N_46228);
nor UO_2646 (O_2646,N_46829,N_47436);
nand UO_2647 (O_2647,N_46118,N_45784);
nor UO_2648 (O_2648,N_45002,N_49624);
nand UO_2649 (O_2649,N_48874,N_45670);
nand UO_2650 (O_2650,N_48855,N_49541);
nor UO_2651 (O_2651,N_47113,N_47176);
or UO_2652 (O_2652,N_46618,N_49889);
or UO_2653 (O_2653,N_48540,N_47223);
nor UO_2654 (O_2654,N_47028,N_48974);
and UO_2655 (O_2655,N_46214,N_45034);
nand UO_2656 (O_2656,N_49900,N_49407);
xor UO_2657 (O_2657,N_46055,N_45241);
or UO_2658 (O_2658,N_45570,N_49187);
and UO_2659 (O_2659,N_47991,N_45698);
or UO_2660 (O_2660,N_45739,N_46155);
or UO_2661 (O_2661,N_49529,N_46780);
and UO_2662 (O_2662,N_48345,N_46597);
and UO_2663 (O_2663,N_49628,N_46258);
or UO_2664 (O_2664,N_49770,N_47668);
or UO_2665 (O_2665,N_48941,N_48763);
nor UO_2666 (O_2666,N_46799,N_47782);
and UO_2667 (O_2667,N_45104,N_47991);
nor UO_2668 (O_2668,N_48617,N_49926);
xor UO_2669 (O_2669,N_48898,N_49791);
and UO_2670 (O_2670,N_45262,N_48038);
nor UO_2671 (O_2671,N_49469,N_48645);
or UO_2672 (O_2672,N_46737,N_45603);
nor UO_2673 (O_2673,N_47062,N_49545);
nor UO_2674 (O_2674,N_48624,N_47642);
nor UO_2675 (O_2675,N_45138,N_48879);
or UO_2676 (O_2676,N_47980,N_46636);
and UO_2677 (O_2677,N_49739,N_48121);
and UO_2678 (O_2678,N_49735,N_45184);
xnor UO_2679 (O_2679,N_46341,N_46119);
nand UO_2680 (O_2680,N_45145,N_49193);
or UO_2681 (O_2681,N_49696,N_48701);
or UO_2682 (O_2682,N_48974,N_46999);
nor UO_2683 (O_2683,N_47940,N_46542);
nand UO_2684 (O_2684,N_48637,N_49658);
and UO_2685 (O_2685,N_49002,N_49610);
nor UO_2686 (O_2686,N_49345,N_45057);
or UO_2687 (O_2687,N_49014,N_47420);
or UO_2688 (O_2688,N_46756,N_45565);
xnor UO_2689 (O_2689,N_45549,N_48730);
nor UO_2690 (O_2690,N_45123,N_49544);
and UO_2691 (O_2691,N_49737,N_45757);
nand UO_2692 (O_2692,N_47354,N_48797);
xnor UO_2693 (O_2693,N_48860,N_48641);
nor UO_2694 (O_2694,N_45241,N_49417);
or UO_2695 (O_2695,N_45247,N_46823);
xor UO_2696 (O_2696,N_49380,N_47068);
or UO_2697 (O_2697,N_45819,N_49590);
nand UO_2698 (O_2698,N_48634,N_47090);
nor UO_2699 (O_2699,N_49166,N_49179);
nor UO_2700 (O_2700,N_48688,N_48476);
nand UO_2701 (O_2701,N_47365,N_47984);
nor UO_2702 (O_2702,N_45305,N_48350);
nor UO_2703 (O_2703,N_49385,N_48023);
or UO_2704 (O_2704,N_48574,N_48561);
nand UO_2705 (O_2705,N_48043,N_45875);
nand UO_2706 (O_2706,N_47338,N_49514);
or UO_2707 (O_2707,N_45868,N_48340);
nand UO_2708 (O_2708,N_49624,N_49074);
nand UO_2709 (O_2709,N_47029,N_47124);
nand UO_2710 (O_2710,N_48125,N_46383);
or UO_2711 (O_2711,N_48203,N_48841);
nand UO_2712 (O_2712,N_46276,N_45616);
nor UO_2713 (O_2713,N_45806,N_48801);
or UO_2714 (O_2714,N_45819,N_47757);
nand UO_2715 (O_2715,N_49042,N_47973);
and UO_2716 (O_2716,N_49628,N_49944);
or UO_2717 (O_2717,N_48279,N_47069);
nor UO_2718 (O_2718,N_47879,N_49267);
or UO_2719 (O_2719,N_49647,N_48009);
nand UO_2720 (O_2720,N_46805,N_45958);
xnor UO_2721 (O_2721,N_46300,N_49404);
and UO_2722 (O_2722,N_48329,N_47288);
xnor UO_2723 (O_2723,N_47854,N_48662);
nor UO_2724 (O_2724,N_49998,N_49254);
and UO_2725 (O_2725,N_45543,N_45175);
nor UO_2726 (O_2726,N_49116,N_49091);
nand UO_2727 (O_2727,N_46543,N_49296);
or UO_2728 (O_2728,N_48348,N_49495);
or UO_2729 (O_2729,N_47731,N_49357);
xor UO_2730 (O_2730,N_47775,N_49880);
nand UO_2731 (O_2731,N_49013,N_49403);
nor UO_2732 (O_2732,N_47845,N_45675);
nand UO_2733 (O_2733,N_49176,N_48628);
and UO_2734 (O_2734,N_46978,N_49197);
and UO_2735 (O_2735,N_45315,N_46757);
nor UO_2736 (O_2736,N_46738,N_45010);
nand UO_2737 (O_2737,N_45011,N_47714);
xor UO_2738 (O_2738,N_47486,N_48718);
xor UO_2739 (O_2739,N_48415,N_45876);
nand UO_2740 (O_2740,N_48512,N_47791);
xor UO_2741 (O_2741,N_48214,N_46853);
nor UO_2742 (O_2742,N_47444,N_47236);
nand UO_2743 (O_2743,N_47682,N_49591);
xor UO_2744 (O_2744,N_46435,N_47530);
nor UO_2745 (O_2745,N_49096,N_47755);
or UO_2746 (O_2746,N_46790,N_47452);
or UO_2747 (O_2747,N_46797,N_45390);
nand UO_2748 (O_2748,N_45209,N_47402);
or UO_2749 (O_2749,N_45485,N_49719);
nor UO_2750 (O_2750,N_49097,N_46164);
nand UO_2751 (O_2751,N_46696,N_47016);
or UO_2752 (O_2752,N_49645,N_46005);
xnor UO_2753 (O_2753,N_46246,N_48236);
nor UO_2754 (O_2754,N_45317,N_47384);
nand UO_2755 (O_2755,N_47197,N_45844);
xor UO_2756 (O_2756,N_45818,N_46489);
or UO_2757 (O_2757,N_47123,N_48492);
nor UO_2758 (O_2758,N_48461,N_46742);
nand UO_2759 (O_2759,N_47312,N_48571);
and UO_2760 (O_2760,N_49794,N_45228);
nor UO_2761 (O_2761,N_49639,N_49015);
nor UO_2762 (O_2762,N_49661,N_46673);
nand UO_2763 (O_2763,N_47520,N_47584);
xor UO_2764 (O_2764,N_47489,N_48983);
nand UO_2765 (O_2765,N_45545,N_47041);
xor UO_2766 (O_2766,N_47694,N_48869);
nor UO_2767 (O_2767,N_49294,N_46782);
nand UO_2768 (O_2768,N_48521,N_47855);
nor UO_2769 (O_2769,N_45418,N_48614);
or UO_2770 (O_2770,N_49943,N_48302);
xnor UO_2771 (O_2771,N_49477,N_49925);
and UO_2772 (O_2772,N_47449,N_45570);
xor UO_2773 (O_2773,N_48128,N_49939);
or UO_2774 (O_2774,N_47435,N_48282);
and UO_2775 (O_2775,N_47231,N_45661);
or UO_2776 (O_2776,N_49499,N_46991);
xor UO_2777 (O_2777,N_48351,N_46793);
nand UO_2778 (O_2778,N_47442,N_48280);
nand UO_2779 (O_2779,N_47353,N_48414);
and UO_2780 (O_2780,N_47577,N_45592);
and UO_2781 (O_2781,N_45242,N_45623);
or UO_2782 (O_2782,N_49155,N_48995);
and UO_2783 (O_2783,N_48720,N_46586);
and UO_2784 (O_2784,N_47322,N_46203);
xor UO_2785 (O_2785,N_48076,N_47420);
nor UO_2786 (O_2786,N_49109,N_46926);
xnor UO_2787 (O_2787,N_45091,N_48308);
nor UO_2788 (O_2788,N_49421,N_49953);
or UO_2789 (O_2789,N_47126,N_45342);
and UO_2790 (O_2790,N_45504,N_48794);
or UO_2791 (O_2791,N_49482,N_48588);
nand UO_2792 (O_2792,N_49744,N_45180);
nor UO_2793 (O_2793,N_47424,N_48574);
or UO_2794 (O_2794,N_49782,N_45622);
and UO_2795 (O_2795,N_49982,N_45632);
nand UO_2796 (O_2796,N_45762,N_46313);
nor UO_2797 (O_2797,N_49836,N_48195);
nand UO_2798 (O_2798,N_48847,N_46019);
nand UO_2799 (O_2799,N_48339,N_49617);
nor UO_2800 (O_2800,N_46131,N_45560);
or UO_2801 (O_2801,N_49696,N_45153);
or UO_2802 (O_2802,N_46599,N_45306);
xor UO_2803 (O_2803,N_46076,N_47689);
or UO_2804 (O_2804,N_47251,N_46921);
and UO_2805 (O_2805,N_45597,N_49610);
and UO_2806 (O_2806,N_45729,N_48311);
nor UO_2807 (O_2807,N_48961,N_49043);
nand UO_2808 (O_2808,N_48597,N_47111);
nand UO_2809 (O_2809,N_48268,N_47688);
nand UO_2810 (O_2810,N_49656,N_49597);
or UO_2811 (O_2811,N_45098,N_46625);
xor UO_2812 (O_2812,N_46148,N_48572);
nand UO_2813 (O_2813,N_47881,N_49420);
or UO_2814 (O_2814,N_47831,N_46229);
or UO_2815 (O_2815,N_49843,N_48794);
xor UO_2816 (O_2816,N_46996,N_48278);
nand UO_2817 (O_2817,N_45542,N_45523);
nand UO_2818 (O_2818,N_48873,N_49059);
and UO_2819 (O_2819,N_45917,N_48574);
or UO_2820 (O_2820,N_46309,N_49074);
or UO_2821 (O_2821,N_46036,N_48468);
xor UO_2822 (O_2822,N_46790,N_46356);
nand UO_2823 (O_2823,N_46506,N_47268);
xor UO_2824 (O_2824,N_48382,N_47415);
nand UO_2825 (O_2825,N_47128,N_46580);
xor UO_2826 (O_2826,N_45049,N_47138);
xor UO_2827 (O_2827,N_49867,N_49071);
nor UO_2828 (O_2828,N_45907,N_46877);
and UO_2829 (O_2829,N_47524,N_46145);
xor UO_2830 (O_2830,N_49202,N_47630);
nand UO_2831 (O_2831,N_45313,N_46407);
xor UO_2832 (O_2832,N_45587,N_49455);
and UO_2833 (O_2833,N_45676,N_49315);
and UO_2834 (O_2834,N_45596,N_45609);
xnor UO_2835 (O_2835,N_47624,N_47051);
nor UO_2836 (O_2836,N_49341,N_48548);
and UO_2837 (O_2837,N_45447,N_46388);
nand UO_2838 (O_2838,N_46695,N_48091);
and UO_2839 (O_2839,N_49408,N_49597);
and UO_2840 (O_2840,N_46985,N_46339);
nor UO_2841 (O_2841,N_45875,N_48272);
nand UO_2842 (O_2842,N_48995,N_48391);
xnor UO_2843 (O_2843,N_45676,N_48287);
nand UO_2844 (O_2844,N_48527,N_49219);
nand UO_2845 (O_2845,N_47983,N_45820);
xor UO_2846 (O_2846,N_46497,N_49841);
xor UO_2847 (O_2847,N_45940,N_48767);
nand UO_2848 (O_2848,N_49702,N_47079);
xor UO_2849 (O_2849,N_49964,N_49534);
nand UO_2850 (O_2850,N_46665,N_49832);
and UO_2851 (O_2851,N_47475,N_48051);
xor UO_2852 (O_2852,N_49424,N_47799);
nand UO_2853 (O_2853,N_46420,N_46802);
and UO_2854 (O_2854,N_46539,N_46167);
nor UO_2855 (O_2855,N_46917,N_49118);
nand UO_2856 (O_2856,N_45444,N_45635);
xor UO_2857 (O_2857,N_47458,N_46413);
xor UO_2858 (O_2858,N_48080,N_48718);
or UO_2859 (O_2859,N_45485,N_48614);
and UO_2860 (O_2860,N_46224,N_48211);
or UO_2861 (O_2861,N_49718,N_45964);
and UO_2862 (O_2862,N_46120,N_48732);
nand UO_2863 (O_2863,N_48111,N_46141);
or UO_2864 (O_2864,N_45835,N_48471);
or UO_2865 (O_2865,N_46829,N_45468);
or UO_2866 (O_2866,N_46111,N_46553);
and UO_2867 (O_2867,N_47859,N_47137);
and UO_2868 (O_2868,N_48928,N_48255);
nand UO_2869 (O_2869,N_48923,N_45874);
and UO_2870 (O_2870,N_47113,N_45421);
nand UO_2871 (O_2871,N_49353,N_49159);
nor UO_2872 (O_2872,N_47012,N_49751);
nor UO_2873 (O_2873,N_47510,N_46109);
nor UO_2874 (O_2874,N_47810,N_48716);
and UO_2875 (O_2875,N_48808,N_47648);
and UO_2876 (O_2876,N_47551,N_49869);
or UO_2877 (O_2877,N_47570,N_47468);
nor UO_2878 (O_2878,N_49937,N_45711);
or UO_2879 (O_2879,N_45612,N_47374);
and UO_2880 (O_2880,N_46363,N_46237);
nand UO_2881 (O_2881,N_45044,N_49669);
xor UO_2882 (O_2882,N_45467,N_47315);
xnor UO_2883 (O_2883,N_49155,N_48055);
or UO_2884 (O_2884,N_45218,N_48382);
or UO_2885 (O_2885,N_45892,N_48370);
nand UO_2886 (O_2886,N_48086,N_49721);
nor UO_2887 (O_2887,N_45208,N_48387);
nand UO_2888 (O_2888,N_49068,N_45069);
and UO_2889 (O_2889,N_46334,N_46385);
nor UO_2890 (O_2890,N_48069,N_49926);
xor UO_2891 (O_2891,N_48548,N_47242);
xnor UO_2892 (O_2892,N_46405,N_45255);
nor UO_2893 (O_2893,N_49242,N_48338);
or UO_2894 (O_2894,N_45222,N_48788);
nor UO_2895 (O_2895,N_45968,N_49029);
nand UO_2896 (O_2896,N_45355,N_47510);
or UO_2897 (O_2897,N_49564,N_45628);
or UO_2898 (O_2898,N_49436,N_46714);
and UO_2899 (O_2899,N_49637,N_46555);
or UO_2900 (O_2900,N_47010,N_49903);
nand UO_2901 (O_2901,N_46636,N_45030);
nand UO_2902 (O_2902,N_45179,N_49931);
or UO_2903 (O_2903,N_48639,N_47029);
or UO_2904 (O_2904,N_45732,N_47013);
or UO_2905 (O_2905,N_48206,N_48531);
xor UO_2906 (O_2906,N_48710,N_47545);
and UO_2907 (O_2907,N_48044,N_49051);
or UO_2908 (O_2908,N_45738,N_48707);
nor UO_2909 (O_2909,N_45329,N_47685);
xnor UO_2910 (O_2910,N_47098,N_46969);
nor UO_2911 (O_2911,N_46063,N_45879);
nand UO_2912 (O_2912,N_47221,N_46120);
nor UO_2913 (O_2913,N_47258,N_47622);
or UO_2914 (O_2914,N_47456,N_45488);
xnor UO_2915 (O_2915,N_49078,N_46002);
and UO_2916 (O_2916,N_48194,N_49800);
or UO_2917 (O_2917,N_45119,N_46989);
nor UO_2918 (O_2918,N_49522,N_48410);
nand UO_2919 (O_2919,N_45832,N_49788);
or UO_2920 (O_2920,N_46022,N_49189);
nor UO_2921 (O_2921,N_45450,N_48921);
and UO_2922 (O_2922,N_46659,N_46916);
nand UO_2923 (O_2923,N_46402,N_48323);
and UO_2924 (O_2924,N_47285,N_48525);
or UO_2925 (O_2925,N_47006,N_49531);
xnor UO_2926 (O_2926,N_48002,N_49348);
and UO_2927 (O_2927,N_45646,N_46962);
nand UO_2928 (O_2928,N_45131,N_48496);
xor UO_2929 (O_2929,N_48235,N_45577);
xor UO_2930 (O_2930,N_46495,N_45853);
nand UO_2931 (O_2931,N_48099,N_46533);
or UO_2932 (O_2932,N_48380,N_46092);
xor UO_2933 (O_2933,N_47640,N_46408);
nand UO_2934 (O_2934,N_45144,N_45150);
nor UO_2935 (O_2935,N_47676,N_48601);
nand UO_2936 (O_2936,N_45483,N_49023);
and UO_2937 (O_2937,N_48140,N_46883);
nor UO_2938 (O_2938,N_49510,N_47357);
nor UO_2939 (O_2939,N_46638,N_46030);
xor UO_2940 (O_2940,N_47597,N_47438);
nand UO_2941 (O_2941,N_46955,N_45198);
xor UO_2942 (O_2942,N_48861,N_49202);
and UO_2943 (O_2943,N_46979,N_45959);
xor UO_2944 (O_2944,N_46027,N_49222);
nand UO_2945 (O_2945,N_48011,N_45006);
and UO_2946 (O_2946,N_45654,N_47831);
nor UO_2947 (O_2947,N_46850,N_47217);
or UO_2948 (O_2948,N_48408,N_45490);
nor UO_2949 (O_2949,N_49088,N_46095);
nand UO_2950 (O_2950,N_49928,N_48218);
or UO_2951 (O_2951,N_49480,N_48862);
nor UO_2952 (O_2952,N_48731,N_46190);
nand UO_2953 (O_2953,N_46020,N_48043);
and UO_2954 (O_2954,N_45508,N_45354);
nor UO_2955 (O_2955,N_48871,N_46389);
xor UO_2956 (O_2956,N_49007,N_48434);
or UO_2957 (O_2957,N_46373,N_46417);
or UO_2958 (O_2958,N_45931,N_49482);
and UO_2959 (O_2959,N_46083,N_46601);
nand UO_2960 (O_2960,N_47526,N_46469);
and UO_2961 (O_2961,N_45392,N_48661);
nand UO_2962 (O_2962,N_48846,N_49675);
nand UO_2963 (O_2963,N_45459,N_46653);
or UO_2964 (O_2964,N_48672,N_49244);
or UO_2965 (O_2965,N_46736,N_46460);
xor UO_2966 (O_2966,N_47927,N_47294);
nor UO_2967 (O_2967,N_49886,N_46826);
or UO_2968 (O_2968,N_48043,N_47999);
xnor UO_2969 (O_2969,N_45099,N_45755);
and UO_2970 (O_2970,N_49354,N_49739);
nand UO_2971 (O_2971,N_49448,N_49408);
nor UO_2972 (O_2972,N_48053,N_48180);
or UO_2973 (O_2973,N_46997,N_49485);
xnor UO_2974 (O_2974,N_46112,N_48661);
and UO_2975 (O_2975,N_48942,N_46567);
xor UO_2976 (O_2976,N_45676,N_47363);
nor UO_2977 (O_2977,N_48537,N_46578);
and UO_2978 (O_2978,N_46497,N_49060);
nand UO_2979 (O_2979,N_46381,N_47029);
and UO_2980 (O_2980,N_47312,N_45568);
nand UO_2981 (O_2981,N_45751,N_49124);
nand UO_2982 (O_2982,N_48599,N_46245);
or UO_2983 (O_2983,N_48181,N_49698);
or UO_2984 (O_2984,N_47419,N_47539);
xor UO_2985 (O_2985,N_46115,N_47851);
and UO_2986 (O_2986,N_47009,N_45147);
xnor UO_2987 (O_2987,N_48709,N_49838);
nor UO_2988 (O_2988,N_48078,N_49938);
nand UO_2989 (O_2989,N_46618,N_45860);
or UO_2990 (O_2990,N_47111,N_47357);
nand UO_2991 (O_2991,N_46834,N_45111);
and UO_2992 (O_2992,N_49571,N_46739);
or UO_2993 (O_2993,N_45959,N_49202);
nand UO_2994 (O_2994,N_49212,N_48680);
and UO_2995 (O_2995,N_48208,N_49092);
and UO_2996 (O_2996,N_47255,N_49807);
xnor UO_2997 (O_2997,N_47458,N_47896);
nor UO_2998 (O_2998,N_45348,N_45198);
or UO_2999 (O_2999,N_47572,N_49324);
nand UO_3000 (O_3000,N_48050,N_46595);
nand UO_3001 (O_3001,N_45329,N_48904);
nor UO_3002 (O_3002,N_46843,N_46798);
and UO_3003 (O_3003,N_49037,N_45081);
nand UO_3004 (O_3004,N_46054,N_49522);
nor UO_3005 (O_3005,N_45546,N_48758);
nand UO_3006 (O_3006,N_47163,N_45206);
nor UO_3007 (O_3007,N_48692,N_48485);
nand UO_3008 (O_3008,N_49182,N_45459);
and UO_3009 (O_3009,N_47572,N_46195);
or UO_3010 (O_3010,N_45786,N_45708);
nor UO_3011 (O_3011,N_45839,N_45060);
xnor UO_3012 (O_3012,N_48171,N_48459);
and UO_3013 (O_3013,N_45896,N_45234);
xnor UO_3014 (O_3014,N_48775,N_46504);
nor UO_3015 (O_3015,N_48209,N_45290);
or UO_3016 (O_3016,N_45706,N_48498);
xnor UO_3017 (O_3017,N_48912,N_48530);
xor UO_3018 (O_3018,N_49759,N_46002);
nor UO_3019 (O_3019,N_46811,N_49393);
and UO_3020 (O_3020,N_49813,N_47220);
and UO_3021 (O_3021,N_47240,N_49600);
and UO_3022 (O_3022,N_49415,N_45855);
xnor UO_3023 (O_3023,N_48429,N_48910);
xor UO_3024 (O_3024,N_48159,N_49943);
or UO_3025 (O_3025,N_47284,N_47049);
or UO_3026 (O_3026,N_48679,N_49852);
nand UO_3027 (O_3027,N_48199,N_48520);
xor UO_3028 (O_3028,N_47259,N_49187);
and UO_3029 (O_3029,N_45720,N_46240);
and UO_3030 (O_3030,N_49011,N_47296);
and UO_3031 (O_3031,N_46585,N_45619);
and UO_3032 (O_3032,N_45842,N_45429);
nand UO_3033 (O_3033,N_47117,N_46425);
and UO_3034 (O_3034,N_46158,N_45016);
nor UO_3035 (O_3035,N_45180,N_48196);
nor UO_3036 (O_3036,N_45015,N_48671);
xor UO_3037 (O_3037,N_48086,N_46070);
nand UO_3038 (O_3038,N_49241,N_45815);
or UO_3039 (O_3039,N_46607,N_46984);
and UO_3040 (O_3040,N_47733,N_48170);
xor UO_3041 (O_3041,N_45651,N_45357);
xor UO_3042 (O_3042,N_49216,N_46054);
xnor UO_3043 (O_3043,N_46047,N_45439);
nand UO_3044 (O_3044,N_46070,N_49670);
nor UO_3045 (O_3045,N_49770,N_48328);
nand UO_3046 (O_3046,N_49330,N_47664);
xor UO_3047 (O_3047,N_46934,N_48107);
and UO_3048 (O_3048,N_45939,N_46944);
and UO_3049 (O_3049,N_48578,N_47814);
and UO_3050 (O_3050,N_45835,N_49491);
xnor UO_3051 (O_3051,N_48127,N_47056);
or UO_3052 (O_3052,N_48724,N_45726);
and UO_3053 (O_3053,N_46118,N_47313);
nor UO_3054 (O_3054,N_49753,N_49278);
and UO_3055 (O_3055,N_45123,N_49130);
xor UO_3056 (O_3056,N_45290,N_46057);
nand UO_3057 (O_3057,N_45178,N_45080);
nand UO_3058 (O_3058,N_47528,N_47518);
or UO_3059 (O_3059,N_49587,N_48718);
nand UO_3060 (O_3060,N_48195,N_49622);
xnor UO_3061 (O_3061,N_49076,N_45071);
nor UO_3062 (O_3062,N_48999,N_47816);
and UO_3063 (O_3063,N_48013,N_47514);
xor UO_3064 (O_3064,N_45693,N_45973);
or UO_3065 (O_3065,N_49171,N_49851);
nand UO_3066 (O_3066,N_46170,N_48458);
or UO_3067 (O_3067,N_45170,N_45289);
xnor UO_3068 (O_3068,N_46589,N_46117);
nand UO_3069 (O_3069,N_46348,N_48118);
and UO_3070 (O_3070,N_48516,N_45907);
and UO_3071 (O_3071,N_46539,N_48226);
xor UO_3072 (O_3072,N_49124,N_45788);
nor UO_3073 (O_3073,N_45555,N_49985);
and UO_3074 (O_3074,N_46892,N_49898);
nand UO_3075 (O_3075,N_49609,N_46643);
nand UO_3076 (O_3076,N_48067,N_46253);
and UO_3077 (O_3077,N_49094,N_45754);
and UO_3078 (O_3078,N_47341,N_46341);
xnor UO_3079 (O_3079,N_48897,N_45791);
or UO_3080 (O_3080,N_46433,N_45339);
and UO_3081 (O_3081,N_47961,N_49064);
nor UO_3082 (O_3082,N_46732,N_45461);
nor UO_3083 (O_3083,N_49998,N_49156);
or UO_3084 (O_3084,N_46187,N_47732);
and UO_3085 (O_3085,N_46149,N_46979);
nor UO_3086 (O_3086,N_46752,N_46373);
xnor UO_3087 (O_3087,N_47963,N_49461);
or UO_3088 (O_3088,N_47761,N_48461);
or UO_3089 (O_3089,N_45811,N_49541);
and UO_3090 (O_3090,N_47292,N_45505);
or UO_3091 (O_3091,N_49217,N_47670);
xnor UO_3092 (O_3092,N_48968,N_46925);
and UO_3093 (O_3093,N_46119,N_49705);
nor UO_3094 (O_3094,N_49062,N_47309);
nor UO_3095 (O_3095,N_45260,N_45410);
and UO_3096 (O_3096,N_45885,N_46572);
or UO_3097 (O_3097,N_48405,N_46221);
xor UO_3098 (O_3098,N_48561,N_45025);
or UO_3099 (O_3099,N_47738,N_47688);
nor UO_3100 (O_3100,N_47163,N_45760);
and UO_3101 (O_3101,N_46586,N_49253);
or UO_3102 (O_3102,N_45222,N_48437);
nand UO_3103 (O_3103,N_48507,N_45195);
and UO_3104 (O_3104,N_47645,N_48953);
xnor UO_3105 (O_3105,N_47207,N_47210);
nand UO_3106 (O_3106,N_47068,N_47229);
xnor UO_3107 (O_3107,N_47810,N_46231);
or UO_3108 (O_3108,N_47404,N_45915);
nand UO_3109 (O_3109,N_49093,N_48263);
xor UO_3110 (O_3110,N_48263,N_46370);
xnor UO_3111 (O_3111,N_45925,N_46326);
or UO_3112 (O_3112,N_45073,N_47987);
or UO_3113 (O_3113,N_46686,N_48599);
and UO_3114 (O_3114,N_49365,N_49325);
nor UO_3115 (O_3115,N_48356,N_46540);
and UO_3116 (O_3116,N_45925,N_49444);
nor UO_3117 (O_3117,N_45106,N_47495);
nand UO_3118 (O_3118,N_46452,N_45785);
nor UO_3119 (O_3119,N_45566,N_46098);
xor UO_3120 (O_3120,N_46623,N_45860);
nor UO_3121 (O_3121,N_48492,N_48084);
nor UO_3122 (O_3122,N_47260,N_48938);
nor UO_3123 (O_3123,N_48621,N_46380);
nor UO_3124 (O_3124,N_46732,N_45488);
xor UO_3125 (O_3125,N_45309,N_48265);
and UO_3126 (O_3126,N_47057,N_45402);
nor UO_3127 (O_3127,N_48449,N_46051);
xor UO_3128 (O_3128,N_49669,N_49924);
xnor UO_3129 (O_3129,N_49522,N_45786);
nand UO_3130 (O_3130,N_45858,N_49163);
xor UO_3131 (O_3131,N_45279,N_47069);
and UO_3132 (O_3132,N_47723,N_45667);
nand UO_3133 (O_3133,N_48140,N_46945);
or UO_3134 (O_3134,N_49303,N_45205);
and UO_3135 (O_3135,N_47189,N_45522);
or UO_3136 (O_3136,N_48717,N_45773);
nand UO_3137 (O_3137,N_45706,N_49575);
or UO_3138 (O_3138,N_49160,N_48678);
and UO_3139 (O_3139,N_49262,N_45012);
and UO_3140 (O_3140,N_45208,N_49398);
nor UO_3141 (O_3141,N_46293,N_45078);
or UO_3142 (O_3142,N_45790,N_45628);
or UO_3143 (O_3143,N_47395,N_49488);
or UO_3144 (O_3144,N_46142,N_45297);
nor UO_3145 (O_3145,N_47641,N_47845);
and UO_3146 (O_3146,N_46974,N_47196);
nor UO_3147 (O_3147,N_49585,N_48000);
or UO_3148 (O_3148,N_49169,N_48543);
and UO_3149 (O_3149,N_46324,N_48680);
or UO_3150 (O_3150,N_48642,N_45747);
or UO_3151 (O_3151,N_48044,N_46282);
nor UO_3152 (O_3152,N_46773,N_45864);
and UO_3153 (O_3153,N_47603,N_48978);
nor UO_3154 (O_3154,N_47549,N_45940);
xnor UO_3155 (O_3155,N_46170,N_45793);
nand UO_3156 (O_3156,N_46065,N_47306);
or UO_3157 (O_3157,N_47771,N_48899);
or UO_3158 (O_3158,N_46099,N_46982);
nor UO_3159 (O_3159,N_49195,N_45591);
and UO_3160 (O_3160,N_47649,N_46512);
nor UO_3161 (O_3161,N_45681,N_49285);
and UO_3162 (O_3162,N_46306,N_46117);
xnor UO_3163 (O_3163,N_46600,N_46801);
or UO_3164 (O_3164,N_47027,N_49496);
nand UO_3165 (O_3165,N_47282,N_47770);
xnor UO_3166 (O_3166,N_45588,N_46057);
nand UO_3167 (O_3167,N_49071,N_46066);
xnor UO_3168 (O_3168,N_45777,N_48233);
nand UO_3169 (O_3169,N_47326,N_46776);
or UO_3170 (O_3170,N_45292,N_48625);
nand UO_3171 (O_3171,N_45516,N_48493);
nor UO_3172 (O_3172,N_48252,N_47743);
xnor UO_3173 (O_3173,N_49359,N_46128);
xnor UO_3174 (O_3174,N_49108,N_46455);
and UO_3175 (O_3175,N_49871,N_49184);
nor UO_3176 (O_3176,N_45489,N_48997);
and UO_3177 (O_3177,N_47289,N_48267);
and UO_3178 (O_3178,N_47575,N_47885);
nor UO_3179 (O_3179,N_49904,N_47936);
nand UO_3180 (O_3180,N_48002,N_47647);
and UO_3181 (O_3181,N_49615,N_49024);
or UO_3182 (O_3182,N_49468,N_48955);
or UO_3183 (O_3183,N_47358,N_46044);
and UO_3184 (O_3184,N_45550,N_46565);
nor UO_3185 (O_3185,N_48450,N_46003);
and UO_3186 (O_3186,N_45412,N_47985);
or UO_3187 (O_3187,N_47671,N_45270);
xor UO_3188 (O_3188,N_47557,N_49950);
xnor UO_3189 (O_3189,N_46223,N_46715);
and UO_3190 (O_3190,N_49132,N_48497);
or UO_3191 (O_3191,N_49923,N_48715);
nand UO_3192 (O_3192,N_45691,N_45036);
nor UO_3193 (O_3193,N_48450,N_46736);
xnor UO_3194 (O_3194,N_45044,N_46785);
xnor UO_3195 (O_3195,N_47819,N_46321);
xnor UO_3196 (O_3196,N_49908,N_45897);
xnor UO_3197 (O_3197,N_45037,N_45848);
xnor UO_3198 (O_3198,N_48889,N_48028);
nor UO_3199 (O_3199,N_49485,N_48489);
nand UO_3200 (O_3200,N_48298,N_47226);
and UO_3201 (O_3201,N_49973,N_46070);
or UO_3202 (O_3202,N_49124,N_49429);
or UO_3203 (O_3203,N_48353,N_47792);
and UO_3204 (O_3204,N_48258,N_48160);
xnor UO_3205 (O_3205,N_45989,N_46817);
xor UO_3206 (O_3206,N_47988,N_47291);
and UO_3207 (O_3207,N_46716,N_45199);
nor UO_3208 (O_3208,N_47524,N_45319);
nand UO_3209 (O_3209,N_45672,N_45765);
and UO_3210 (O_3210,N_45329,N_48956);
xor UO_3211 (O_3211,N_47781,N_46584);
and UO_3212 (O_3212,N_48460,N_49549);
xor UO_3213 (O_3213,N_45181,N_46480);
xor UO_3214 (O_3214,N_48411,N_47375);
nor UO_3215 (O_3215,N_49596,N_46652);
and UO_3216 (O_3216,N_49772,N_45173);
xnor UO_3217 (O_3217,N_45847,N_46752);
xnor UO_3218 (O_3218,N_45106,N_47094);
nand UO_3219 (O_3219,N_47895,N_46114);
xor UO_3220 (O_3220,N_49563,N_48704);
nor UO_3221 (O_3221,N_47829,N_48660);
nor UO_3222 (O_3222,N_47851,N_45201);
or UO_3223 (O_3223,N_49687,N_45369);
nor UO_3224 (O_3224,N_47310,N_48253);
or UO_3225 (O_3225,N_49446,N_49185);
nor UO_3226 (O_3226,N_45851,N_49084);
nand UO_3227 (O_3227,N_45528,N_48988);
xnor UO_3228 (O_3228,N_47075,N_45467);
nand UO_3229 (O_3229,N_45819,N_46626);
nand UO_3230 (O_3230,N_45380,N_47714);
nor UO_3231 (O_3231,N_46678,N_47318);
nor UO_3232 (O_3232,N_46084,N_49592);
or UO_3233 (O_3233,N_45295,N_46216);
nand UO_3234 (O_3234,N_48987,N_48468);
nand UO_3235 (O_3235,N_46745,N_47202);
nand UO_3236 (O_3236,N_48176,N_46531);
and UO_3237 (O_3237,N_49029,N_46538);
nand UO_3238 (O_3238,N_47195,N_45668);
nand UO_3239 (O_3239,N_46330,N_48231);
nand UO_3240 (O_3240,N_45882,N_46468);
nor UO_3241 (O_3241,N_46971,N_47443);
xnor UO_3242 (O_3242,N_46446,N_48688);
nor UO_3243 (O_3243,N_45506,N_46913);
nand UO_3244 (O_3244,N_47274,N_49306);
nor UO_3245 (O_3245,N_47280,N_47328);
nor UO_3246 (O_3246,N_45015,N_46733);
nand UO_3247 (O_3247,N_49189,N_45499);
or UO_3248 (O_3248,N_47201,N_47323);
nor UO_3249 (O_3249,N_45743,N_48129);
and UO_3250 (O_3250,N_45678,N_45779);
nor UO_3251 (O_3251,N_48927,N_48858);
or UO_3252 (O_3252,N_45003,N_48081);
nand UO_3253 (O_3253,N_47428,N_47714);
and UO_3254 (O_3254,N_47020,N_47351);
nand UO_3255 (O_3255,N_47344,N_46457);
and UO_3256 (O_3256,N_49611,N_45844);
and UO_3257 (O_3257,N_48978,N_49174);
xor UO_3258 (O_3258,N_48651,N_46988);
nor UO_3259 (O_3259,N_49208,N_46038);
nand UO_3260 (O_3260,N_47631,N_47405);
nor UO_3261 (O_3261,N_49127,N_46780);
and UO_3262 (O_3262,N_45899,N_45722);
xnor UO_3263 (O_3263,N_49655,N_49369);
xor UO_3264 (O_3264,N_46465,N_47187);
nand UO_3265 (O_3265,N_47167,N_48380);
and UO_3266 (O_3266,N_45452,N_48577);
xnor UO_3267 (O_3267,N_47446,N_49829);
nand UO_3268 (O_3268,N_48919,N_46165);
xor UO_3269 (O_3269,N_47866,N_49677);
xor UO_3270 (O_3270,N_47913,N_47644);
and UO_3271 (O_3271,N_47081,N_49544);
and UO_3272 (O_3272,N_47031,N_48623);
nor UO_3273 (O_3273,N_48164,N_47903);
or UO_3274 (O_3274,N_46272,N_45286);
nor UO_3275 (O_3275,N_49492,N_46886);
nor UO_3276 (O_3276,N_45610,N_46082);
nor UO_3277 (O_3277,N_47927,N_46679);
nor UO_3278 (O_3278,N_48634,N_47360);
nand UO_3279 (O_3279,N_47913,N_45152);
nand UO_3280 (O_3280,N_46773,N_47199);
xor UO_3281 (O_3281,N_48969,N_49896);
xnor UO_3282 (O_3282,N_48976,N_49594);
xor UO_3283 (O_3283,N_45329,N_47908);
xor UO_3284 (O_3284,N_49146,N_48752);
xor UO_3285 (O_3285,N_47833,N_45060);
nor UO_3286 (O_3286,N_46868,N_49119);
or UO_3287 (O_3287,N_49390,N_48518);
nor UO_3288 (O_3288,N_47076,N_49709);
and UO_3289 (O_3289,N_49063,N_48600);
nor UO_3290 (O_3290,N_48352,N_49152);
nor UO_3291 (O_3291,N_45598,N_48221);
or UO_3292 (O_3292,N_46513,N_49255);
nor UO_3293 (O_3293,N_47570,N_46246);
and UO_3294 (O_3294,N_49796,N_48436);
nor UO_3295 (O_3295,N_48942,N_46572);
xnor UO_3296 (O_3296,N_49798,N_49269);
or UO_3297 (O_3297,N_45634,N_48521);
nand UO_3298 (O_3298,N_47157,N_45960);
xor UO_3299 (O_3299,N_45956,N_46726);
nand UO_3300 (O_3300,N_45681,N_46214);
or UO_3301 (O_3301,N_47301,N_46998);
xnor UO_3302 (O_3302,N_46027,N_46398);
nand UO_3303 (O_3303,N_47120,N_48794);
and UO_3304 (O_3304,N_45738,N_45121);
xnor UO_3305 (O_3305,N_46031,N_49550);
xnor UO_3306 (O_3306,N_45691,N_48878);
nor UO_3307 (O_3307,N_49311,N_47628);
nor UO_3308 (O_3308,N_46056,N_49034);
nor UO_3309 (O_3309,N_49661,N_46474);
and UO_3310 (O_3310,N_49628,N_46325);
xnor UO_3311 (O_3311,N_45925,N_49763);
and UO_3312 (O_3312,N_45151,N_48178);
and UO_3313 (O_3313,N_46855,N_48045);
xor UO_3314 (O_3314,N_45261,N_45303);
xnor UO_3315 (O_3315,N_48773,N_46904);
nand UO_3316 (O_3316,N_47490,N_48971);
and UO_3317 (O_3317,N_46806,N_47678);
or UO_3318 (O_3318,N_45352,N_48197);
xor UO_3319 (O_3319,N_45640,N_48265);
nand UO_3320 (O_3320,N_47909,N_45233);
xnor UO_3321 (O_3321,N_47013,N_46352);
nand UO_3322 (O_3322,N_48886,N_45708);
nor UO_3323 (O_3323,N_46359,N_47143);
nand UO_3324 (O_3324,N_47070,N_47177);
nand UO_3325 (O_3325,N_47922,N_45927);
nor UO_3326 (O_3326,N_47465,N_47133);
and UO_3327 (O_3327,N_46165,N_47701);
nand UO_3328 (O_3328,N_46918,N_45737);
xnor UO_3329 (O_3329,N_46120,N_45202);
or UO_3330 (O_3330,N_49644,N_45671);
or UO_3331 (O_3331,N_45542,N_45192);
nand UO_3332 (O_3332,N_46128,N_49700);
nand UO_3333 (O_3333,N_49821,N_48665);
and UO_3334 (O_3334,N_45754,N_47648);
or UO_3335 (O_3335,N_48594,N_45857);
and UO_3336 (O_3336,N_48478,N_48106);
and UO_3337 (O_3337,N_47933,N_49531);
xor UO_3338 (O_3338,N_48033,N_45993);
or UO_3339 (O_3339,N_49222,N_48123);
or UO_3340 (O_3340,N_48658,N_45421);
xnor UO_3341 (O_3341,N_47119,N_45436);
or UO_3342 (O_3342,N_48168,N_49456);
or UO_3343 (O_3343,N_49815,N_47332);
nand UO_3344 (O_3344,N_45130,N_48563);
nor UO_3345 (O_3345,N_49154,N_46773);
nor UO_3346 (O_3346,N_47352,N_45732);
nand UO_3347 (O_3347,N_47792,N_49665);
nand UO_3348 (O_3348,N_48768,N_49720);
nor UO_3349 (O_3349,N_49053,N_45098);
and UO_3350 (O_3350,N_49090,N_48677);
xor UO_3351 (O_3351,N_47266,N_46424);
xor UO_3352 (O_3352,N_45802,N_48146);
nand UO_3353 (O_3353,N_49380,N_47698);
or UO_3354 (O_3354,N_47826,N_48562);
or UO_3355 (O_3355,N_45079,N_47394);
xor UO_3356 (O_3356,N_45505,N_48589);
or UO_3357 (O_3357,N_46301,N_46753);
and UO_3358 (O_3358,N_47467,N_48730);
and UO_3359 (O_3359,N_49201,N_46867);
xor UO_3360 (O_3360,N_48500,N_45808);
xor UO_3361 (O_3361,N_45854,N_49776);
and UO_3362 (O_3362,N_48986,N_49899);
xnor UO_3363 (O_3363,N_48865,N_48590);
xor UO_3364 (O_3364,N_46182,N_47562);
and UO_3365 (O_3365,N_48733,N_45524);
nor UO_3366 (O_3366,N_46863,N_47460);
and UO_3367 (O_3367,N_47003,N_45282);
and UO_3368 (O_3368,N_46865,N_45547);
and UO_3369 (O_3369,N_48239,N_48046);
nor UO_3370 (O_3370,N_48498,N_46373);
xor UO_3371 (O_3371,N_45320,N_47213);
nor UO_3372 (O_3372,N_46275,N_47725);
xnor UO_3373 (O_3373,N_48901,N_49346);
or UO_3374 (O_3374,N_46025,N_46397);
and UO_3375 (O_3375,N_47471,N_46572);
nand UO_3376 (O_3376,N_45018,N_47663);
and UO_3377 (O_3377,N_47979,N_47428);
and UO_3378 (O_3378,N_49277,N_46717);
nor UO_3379 (O_3379,N_47328,N_48272);
and UO_3380 (O_3380,N_47762,N_46684);
xnor UO_3381 (O_3381,N_45972,N_46655);
nand UO_3382 (O_3382,N_46662,N_48140);
xnor UO_3383 (O_3383,N_47256,N_47212);
or UO_3384 (O_3384,N_49551,N_47263);
and UO_3385 (O_3385,N_47353,N_47307);
nand UO_3386 (O_3386,N_45245,N_45317);
or UO_3387 (O_3387,N_48167,N_49124);
nor UO_3388 (O_3388,N_45318,N_48879);
and UO_3389 (O_3389,N_45975,N_49561);
or UO_3390 (O_3390,N_47128,N_47372);
nor UO_3391 (O_3391,N_49727,N_48503);
or UO_3392 (O_3392,N_47239,N_45979);
or UO_3393 (O_3393,N_45008,N_48273);
nor UO_3394 (O_3394,N_46836,N_48461);
and UO_3395 (O_3395,N_46817,N_48776);
or UO_3396 (O_3396,N_46549,N_46682);
nand UO_3397 (O_3397,N_45070,N_47341);
nand UO_3398 (O_3398,N_49258,N_46593);
nand UO_3399 (O_3399,N_46006,N_49490);
xnor UO_3400 (O_3400,N_45778,N_48670);
and UO_3401 (O_3401,N_49777,N_48568);
or UO_3402 (O_3402,N_49729,N_47278);
nor UO_3403 (O_3403,N_48557,N_48234);
nor UO_3404 (O_3404,N_48213,N_46087);
nand UO_3405 (O_3405,N_47112,N_47548);
nand UO_3406 (O_3406,N_49710,N_45942);
nor UO_3407 (O_3407,N_45204,N_48666);
and UO_3408 (O_3408,N_48922,N_48686);
nor UO_3409 (O_3409,N_48218,N_49816);
nand UO_3410 (O_3410,N_47801,N_49124);
or UO_3411 (O_3411,N_45873,N_49951);
nand UO_3412 (O_3412,N_48775,N_49263);
and UO_3413 (O_3413,N_46125,N_49525);
nor UO_3414 (O_3414,N_45238,N_46994);
and UO_3415 (O_3415,N_46783,N_46881);
nand UO_3416 (O_3416,N_49880,N_46873);
xnor UO_3417 (O_3417,N_45766,N_48786);
xnor UO_3418 (O_3418,N_48521,N_45779);
and UO_3419 (O_3419,N_46056,N_47611);
and UO_3420 (O_3420,N_49101,N_46814);
and UO_3421 (O_3421,N_48173,N_47699);
nand UO_3422 (O_3422,N_48462,N_47087);
and UO_3423 (O_3423,N_49423,N_49359);
and UO_3424 (O_3424,N_48575,N_45499);
xnor UO_3425 (O_3425,N_47543,N_45076);
xnor UO_3426 (O_3426,N_46097,N_48288);
xor UO_3427 (O_3427,N_46007,N_48378);
and UO_3428 (O_3428,N_47324,N_47873);
and UO_3429 (O_3429,N_46728,N_48699);
and UO_3430 (O_3430,N_48950,N_45684);
nand UO_3431 (O_3431,N_45641,N_45110);
or UO_3432 (O_3432,N_45435,N_46322);
nand UO_3433 (O_3433,N_46574,N_45317);
nor UO_3434 (O_3434,N_46374,N_45764);
nand UO_3435 (O_3435,N_48083,N_46537);
nor UO_3436 (O_3436,N_45573,N_47015);
nand UO_3437 (O_3437,N_49029,N_45703);
nor UO_3438 (O_3438,N_48474,N_49081);
and UO_3439 (O_3439,N_48363,N_48704);
nand UO_3440 (O_3440,N_48118,N_48596);
nand UO_3441 (O_3441,N_46219,N_45590);
xnor UO_3442 (O_3442,N_45132,N_45384);
xnor UO_3443 (O_3443,N_46364,N_49343);
or UO_3444 (O_3444,N_45314,N_49223);
xnor UO_3445 (O_3445,N_45731,N_46954);
xor UO_3446 (O_3446,N_48319,N_46049);
and UO_3447 (O_3447,N_47345,N_47971);
or UO_3448 (O_3448,N_46166,N_47905);
nand UO_3449 (O_3449,N_47957,N_48888);
xor UO_3450 (O_3450,N_47808,N_49118);
xor UO_3451 (O_3451,N_48819,N_48013);
and UO_3452 (O_3452,N_48147,N_49676);
nor UO_3453 (O_3453,N_45908,N_47359);
or UO_3454 (O_3454,N_46687,N_47303);
and UO_3455 (O_3455,N_49975,N_46936);
or UO_3456 (O_3456,N_49830,N_49054);
xnor UO_3457 (O_3457,N_46200,N_47061);
nand UO_3458 (O_3458,N_47883,N_48074);
and UO_3459 (O_3459,N_49720,N_49918);
nor UO_3460 (O_3460,N_48822,N_48114);
xnor UO_3461 (O_3461,N_46853,N_48116);
nor UO_3462 (O_3462,N_48884,N_45961);
or UO_3463 (O_3463,N_48993,N_47007);
nor UO_3464 (O_3464,N_45922,N_49962);
and UO_3465 (O_3465,N_45040,N_47934);
nor UO_3466 (O_3466,N_45456,N_49161);
or UO_3467 (O_3467,N_46203,N_47379);
and UO_3468 (O_3468,N_49486,N_45267);
and UO_3469 (O_3469,N_48068,N_49288);
or UO_3470 (O_3470,N_49328,N_45698);
xnor UO_3471 (O_3471,N_48435,N_45158);
nor UO_3472 (O_3472,N_48084,N_49620);
or UO_3473 (O_3473,N_49047,N_49398);
nor UO_3474 (O_3474,N_46606,N_47421);
and UO_3475 (O_3475,N_45177,N_48371);
xor UO_3476 (O_3476,N_46063,N_45141);
nor UO_3477 (O_3477,N_49307,N_46850);
or UO_3478 (O_3478,N_49921,N_48341);
or UO_3479 (O_3479,N_45586,N_49628);
xnor UO_3480 (O_3480,N_47156,N_47114);
nand UO_3481 (O_3481,N_48095,N_45901);
nand UO_3482 (O_3482,N_49342,N_48970);
nor UO_3483 (O_3483,N_49253,N_47033);
xor UO_3484 (O_3484,N_49731,N_46776);
and UO_3485 (O_3485,N_49937,N_47550);
or UO_3486 (O_3486,N_47518,N_49307);
nor UO_3487 (O_3487,N_46344,N_45440);
nor UO_3488 (O_3488,N_48310,N_49996);
nand UO_3489 (O_3489,N_47732,N_47150);
xnor UO_3490 (O_3490,N_46624,N_46747);
nor UO_3491 (O_3491,N_45416,N_45414);
or UO_3492 (O_3492,N_48082,N_49151);
nand UO_3493 (O_3493,N_45351,N_47049);
and UO_3494 (O_3494,N_45531,N_49262);
xor UO_3495 (O_3495,N_49221,N_47923);
nor UO_3496 (O_3496,N_48417,N_45236);
nor UO_3497 (O_3497,N_46448,N_48006);
xor UO_3498 (O_3498,N_45502,N_45705);
and UO_3499 (O_3499,N_49680,N_47871);
nand UO_3500 (O_3500,N_49594,N_47526);
xor UO_3501 (O_3501,N_46161,N_45235);
and UO_3502 (O_3502,N_47973,N_49338);
nor UO_3503 (O_3503,N_47303,N_49696);
nor UO_3504 (O_3504,N_49054,N_49663);
nand UO_3505 (O_3505,N_45340,N_47005);
and UO_3506 (O_3506,N_49392,N_47367);
or UO_3507 (O_3507,N_46414,N_49127);
and UO_3508 (O_3508,N_49889,N_45066);
nand UO_3509 (O_3509,N_49979,N_49061);
and UO_3510 (O_3510,N_45824,N_48959);
and UO_3511 (O_3511,N_47774,N_47231);
nor UO_3512 (O_3512,N_47177,N_49897);
or UO_3513 (O_3513,N_49690,N_49883);
and UO_3514 (O_3514,N_46793,N_47561);
nor UO_3515 (O_3515,N_48403,N_47974);
or UO_3516 (O_3516,N_46756,N_49491);
or UO_3517 (O_3517,N_47373,N_48394);
and UO_3518 (O_3518,N_46851,N_45232);
and UO_3519 (O_3519,N_48289,N_49793);
nand UO_3520 (O_3520,N_46080,N_47328);
nand UO_3521 (O_3521,N_49496,N_48900);
nand UO_3522 (O_3522,N_46504,N_46156);
or UO_3523 (O_3523,N_46376,N_46286);
nand UO_3524 (O_3524,N_47951,N_46384);
and UO_3525 (O_3525,N_46126,N_45130);
and UO_3526 (O_3526,N_49184,N_47215);
or UO_3527 (O_3527,N_47349,N_45759);
and UO_3528 (O_3528,N_45309,N_45209);
xor UO_3529 (O_3529,N_46361,N_46708);
nand UO_3530 (O_3530,N_48545,N_49196);
and UO_3531 (O_3531,N_49237,N_49625);
nand UO_3532 (O_3532,N_49341,N_45106);
or UO_3533 (O_3533,N_49640,N_48765);
nand UO_3534 (O_3534,N_46228,N_46046);
and UO_3535 (O_3535,N_47740,N_48313);
and UO_3536 (O_3536,N_49894,N_47450);
xnor UO_3537 (O_3537,N_45807,N_46928);
nor UO_3538 (O_3538,N_46705,N_48255);
nand UO_3539 (O_3539,N_46897,N_48159);
and UO_3540 (O_3540,N_47016,N_49367);
nand UO_3541 (O_3541,N_45885,N_46614);
xnor UO_3542 (O_3542,N_47326,N_49793);
and UO_3543 (O_3543,N_49395,N_46396);
or UO_3544 (O_3544,N_45881,N_48702);
or UO_3545 (O_3545,N_47761,N_45091);
and UO_3546 (O_3546,N_48564,N_49927);
and UO_3547 (O_3547,N_48456,N_49966);
and UO_3548 (O_3548,N_47982,N_47119);
or UO_3549 (O_3549,N_48993,N_47031);
xor UO_3550 (O_3550,N_47258,N_49020);
nor UO_3551 (O_3551,N_46162,N_48170);
xnor UO_3552 (O_3552,N_47451,N_49796);
nor UO_3553 (O_3553,N_46015,N_46863);
and UO_3554 (O_3554,N_46500,N_47452);
xor UO_3555 (O_3555,N_49694,N_45528);
nand UO_3556 (O_3556,N_47879,N_47339);
xor UO_3557 (O_3557,N_49308,N_48955);
or UO_3558 (O_3558,N_45337,N_45986);
or UO_3559 (O_3559,N_47262,N_47523);
xor UO_3560 (O_3560,N_46160,N_46000);
and UO_3561 (O_3561,N_45716,N_49090);
xor UO_3562 (O_3562,N_49076,N_48801);
xor UO_3563 (O_3563,N_48763,N_47157);
nor UO_3564 (O_3564,N_47710,N_45811);
or UO_3565 (O_3565,N_49073,N_48338);
xor UO_3566 (O_3566,N_45592,N_49399);
and UO_3567 (O_3567,N_49980,N_45636);
nand UO_3568 (O_3568,N_46512,N_47239);
nand UO_3569 (O_3569,N_47876,N_47171);
and UO_3570 (O_3570,N_49256,N_45102);
nor UO_3571 (O_3571,N_45545,N_48610);
nor UO_3572 (O_3572,N_49745,N_47587);
and UO_3573 (O_3573,N_49704,N_49610);
xor UO_3574 (O_3574,N_48210,N_45434);
xnor UO_3575 (O_3575,N_45503,N_48199);
and UO_3576 (O_3576,N_49542,N_47846);
and UO_3577 (O_3577,N_48204,N_45519);
nand UO_3578 (O_3578,N_48736,N_45487);
or UO_3579 (O_3579,N_49302,N_46158);
and UO_3580 (O_3580,N_47709,N_45964);
and UO_3581 (O_3581,N_49912,N_46238);
xnor UO_3582 (O_3582,N_46869,N_49924);
xnor UO_3583 (O_3583,N_47354,N_49989);
xor UO_3584 (O_3584,N_45397,N_48910);
nor UO_3585 (O_3585,N_49073,N_49844);
nand UO_3586 (O_3586,N_47176,N_48041);
nand UO_3587 (O_3587,N_49405,N_49114);
nand UO_3588 (O_3588,N_49007,N_46800);
nor UO_3589 (O_3589,N_47516,N_45292);
and UO_3590 (O_3590,N_48976,N_47374);
nor UO_3591 (O_3591,N_49361,N_46668);
and UO_3592 (O_3592,N_47088,N_47439);
and UO_3593 (O_3593,N_47841,N_48376);
or UO_3594 (O_3594,N_48672,N_46170);
nand UO_3595 (O_3595,N_49420,N_45317);
or UO_3596 (O_3596,N_49398,N_49351);
xnor UO_3597 (O_3597,N_45529,N_45995);
and UO_3598 (O_3598,N_48122,N_46499);
nor UO_3599 (O_3599,N_49687,N_45504);
nand UO_3600 (O_3600,N_45151,N_47088);
nand UO_3601 (O_3601,N_46049,N_46817);
and UO_3602 (O_3602,N_46451,N_45532);
nor UO_3603 (O_3603,N_48010,N_46422);
nand UO_3604 (O_3604,N_49672,N_46651);
xnor UO_3605 (O_3605,N_49587,N_45971);
nand UO_3606 (O_3606,N_48103,N_46301);
or UO_3607 (O_3607,N_49970,N_46810);
and UO_3608 (O_3608,N_49735,N_49594);
xnor UO_3609 (O_3609,N_48843,N_47526);
or UO_3610 (O_3610,N_46558,N_46680);
nand UO_3611 (O_3611,N_46507,N_47230);
xnor UO_3612 (O_3612,N_45589,N_48131);
nor UO_3613 (O_3613,N_45251,N_45135);
xnor UO_3614 (O_3614,N_48832,N_46443);
xor UO_3615 (O_3615,N_45406,N_45213);
nor UO_3616 (O_3616,N_48220,N_47371);
xor UO_3617 (O_3617,N_47615,N_47747);
xor UO_3618 (O_3618,N_46309,N_49257);
nand UO_3619 (O_3619,N_47327,N_45284);
nand UO_3620 (O_3620,N_49450,N_46382);
nand UO_3621 (O_3621,N_46866,N_49649);
nor UO_3622 (O_3622,N_46250,N_46181);
nand UO_3623 (O_3623,N_48073,N_49380);
or UO_3624 (O_3624,N_48680,N_49297);
and UO_3625 (O_3625,N_48097,N_46638);
or UO_3626 (O_3626,N_45759,N_47386);
or UO_3627 (O_3627,N_46003,N_45947);
nand UO_3628 (O_3628,N_45861,N_45258);
xor UO_3629 (O_3629,N_49358,N_48101);
and UO_3630 (O_3630,N_46323,N_49216);
nor UO_3631 (O_3631,N_48284,N_48995);
nor UO_3632 (O_3632,N_49384,N_46585);
or UO_3633 (O_3633,N_48940,N_49956);
nand UO_3634 (O_3634,N_45699,N_49413);
and UO_3635 (O_3635,N_48404,N_47047);
or UO_3636 (O_3636,N_49327,N_45695);
nor UO_3637 (O_3637,N_47627,N_48687);
or UO_3638 (O_3638,N_46711,N_47298);
nand UO_3639 (O_3639,N_47921,N_49064);
and UO_3640 (O_3640,N_49771,N_49310);
and UO_3641 (O_3641,N_48185,N_48900);
or UO_3642 (O_3642,N_45918,N_46087);
nand UO_3643 (O_3643,N_48691,N_49499);
nor UO_3644 (O_3644,N_47886,N_46188);
xor UO_3645 (O_3645,N_49450,N_46658);
nand UO_3646 (O_3646,N_48163,N_48206);
and UO_3647 (O_3647,N_47083,N_48802);
or UO_3648 (O_3648,N_48577,N_45119);
or UO_3649 (O_3649,N_49945,N_48787);
nand UO_3650 (O_3650,N_45765,N_47832);
or UO_3651 (O_3651,N_45400,N_47990);
nand UO_3652 (O_3652,N_47381,N_49956);
xnor UO_3653 (O_3653,N_45016,N_45323);
or UO_3654 (O_3654,N_49393,N_49748);
or UO_3655 (O_3655,N_48113,N_47941);
nand UO_3656 (O_3656,N_48719,N_47150);
and UO_3657 (O_3657,N_49090,N_48632);
and UO_3658 (O_3658,N_46103,N_46403);
xnor UO_3659 (O_3659,N_48986,N_49543);
xnor UO_3660 (O_3660,N_48703,N_45743);
or UO_3661 (O_3661,N_47962,N_48966);
xor UO_3662 (O_3662,N_48690,N_45380);
nor UO_3663 (O_3663,N_48936,N_47107);
or UO_3664 (O_3664,N_48663,N_49300);
or UO_3665 (O_3665,N_45641,N_48363);
nor UO_3666 (O_3666,N_48692,N_47546);
nor UO_3667 (O_3667,N_45187,N_45242);
and UO_3668 (O_3668,N_48901,N_49890);
xnor UO_3669 (O_3669,N_47092,N_45983);
xnor UO_3670 (O_3670,N_47569,N_48398);
nor UO_3671 (O_3671,N_47082,N_46612);
xor UO_3672 (O_3672,N_48434,N_49645);
nand UO_3673 (O_3673,N_47731,N_48812);
xnor UO_3674 (O_3674,N_45893,N_47374);
xor UO_3675 (O_3675,N_49751,N_47499);
nand UO_3676 (O_3676,N_48285,N_49552);
nand UO_3677 (O_3677,N_45090,N_49288);
nand UO_3678 (O_3678,N_49878,N_45633);
and UO_3679 (O_3679,N_46733,N_46992);
and UO_3680 (O_3680,N_45165,N_48548);
and UO_3681 (O_3681,N_46932,N_47740);
and UO_3682 (O_3682,N_48162,N_46825);
or UO_3683 (O_3683,N_47937,N_47801);
xnor UO_3684 (O_3684,N_45964,N_46604);
or UO_3685 (O_3685,N_48132,N_49552);
xnor UO_3686 (O_3686,N_47204,N_49487);
nor UO_3687 (O_3687,N_47780,N_48268);
and UO_3688 (O_3688,N_45796,N_46421);
and UO_3689 (O_3689,N_46404,N_46198);
nor UO_3690 (O_3690,N_48187,N_49419);
and UO_3691 (O_3691,N_45618,N_46780);
xnor UO_3692 (O_3692,N_48939,N_49267);
and UO_3693 (O_3693,N_49559,N_45664);
xnor UO_3694 (O_3694,N_45220,N_48683);
and UO_3695 (O_3695,N_49698,N_48369);
or UO_3696 (O_3696,N_45843,N_46532);
nand UO_3697 (O_3697,N_49653,N_49861);
nor UO_3698 (O_3698,N_49316,N_48328);
xor UO_3699 (O_3699,N_48862,N_46343);
xor UO_3700 (O_3700,N_48636,N_46950);
or UO_3701 (O_3701,N_47155,N_49184);
nor UO_3702 (O_3702,N_47144,N_48235);
xor UO_3703 (O_3703,N_46603,N_48398);
nor UO_3704 (O_3704,N_49613,N_47044);
nor UO_3705 (O_3705,N_49069,N_45304);
or UO_3706 (O_3706,N_49537,N_49000);
and UO_3707 (O_3707,N_45564,N_45636);
xor UO_3708 (O_3708,N_45518,N_45232);
and UO_3709 (O_3709,N_45564,N_45506);
nor UO_3710 (O_3710,N_45020,N_49934);
nand UO_3711 (O_3711,N_48442,N_47781);
nor UO_3712 (O_3712,N_48233,N_45365);
nor UO_3713 (O_3713,N_48888,N_46039);
xor UO_3714 (O_3714,N_47442,N_45411);
or UO_3715 (O_3715,N_49442,N_48209);
nor UO_3716 (O_3716,N_48152,N_47467);
nor UO_3717 (O_3717,N_46574,N_45042);
or UO_3718 (O_3718,N_45043,N_46907);
or UO_3719 (O_3719,N_45464,N_47688);
nand UO_3720 (O_3720,N_46652,N_47778);
and UO_3721 (O_3721,N_46852,N_46976);
xor UO_3722 (O_3722,N_48984,N_45668);
nor UO_3723 (O_3723,N_49606,N_49424);
xor UO_3724 (O_3724,N_47583,N_46857);
nand UO_3725 (O_3725,N_45843,N_49469);
nor UO_3726 (O_3726,N_47147,N_46091);
or UO_3727 (O_3727,N_46319,N_49948);
and UO_3728 (O_3728,N_47134,N_49165);
or UO_3729 (O_3729,N_46152,N_46522);
and UO_3730 (O_3730,N_46036,N_47107);
and UO_3731 (O_3731,N_45119,N_49818);
xnor UO_3732 (O_3732,N_46999,N_47281);
and UO_3733 (O_3733,N_46029,N_48886);
xnor UO_3734 (O_3734,N_46770,N_47291);
nor UO_3735 (O_3735,N_45869,N_46245);
or UO_3736 (O_3736,N_48601,N_45737);
xor UO_3737 (O_3737,N_49305,N_48058);
xnor UO_3738 (O_3738,N_45637,N_48844);
nand UO_3739 (O_3739,N_45878,N_45495);
nand UO_3740 (O_3740,N_45340,N_48315);
and UO_3741 (O_3741,N_48177,N_48063);
nor UO_3742 (O_3742,N_47480,N_45037);
nor UO_3743 (O_3743,N_48531,N_49630);
or UO_3744 (O_3744,N_47680,N_45068);
nor UO_3745 (O_3745,N_48609,N_49925);
nor UO_3746 (O_3746,N_46981,N_48208);
and UO_3747 (O_3747,N_48492,N_48054);
and UO_3748 (O_3748,N_45937,N_48704);
or UO_3749 (O_3749,N_46157,N_48419);
or UO_3750 (O_3750,N_45804,N_47361);
and UO_3751 (O_3751,N_48690,N_49670);
and UO_3752 (O_3752,N_45992,N_49604);
nor UO_3753 (O_3753,N_48863,N_48974);
xor UO_3754 (O_3754,N_45987,N_45399);
and UO_3755 (O_3755,N_45284,N_48328);
nor UO_3756 (O_3756,N_46993,N_47032);
and UO_3757 (O_3757,N_46578,N_48598);
xnor UO_3758 (O_3758,N_48047,N_47747);
or UO_3759 (O_3759,N_48705,N_45652);
xor UO_3760 (O_3760,N_45881,N_45705);
nand UO_3761 (O_3761,N_46105,N_45432);
and UO_3762 (O_3762,N_48855,N_49807);
nor UO_3763 (O_3763,N_47835,N_45819);
and UO_3764 (O_3764,N_45190,N_47489);
nor UO_3765 (O_3765,N_49216,N_45726);
nand UO_3766 (O_3766,N_48257,N_45003);
or UO_3767 (O_3767,N_46826,N_45979);
or UO_3768 (O_3768,N_48399,N_49636);
and UO_3769 (O_3769,N_47898,N_49072);
nor UO_3770 (O_3770,N_48410,N_46787);
or UO_3771 (O_3771,N_48827,N_48530);
nor UO_3772 (O_3772,N_48832,N_49299);
and UO_3773 (O_3773,N_46245,N_48211);
nand UO_3774 (O_3774,N_49764,N_45070);
nor UO_3775 (O_3775,N_45853,N_45483);
or UO_3776 (O_3776,N_47473,N_49014);
and UO_3777 (O_3777,N_46075,N_45389);
or UO_3778 (O_3778,N_47790,N_49791);
nand UO_3779 (O_3779,N_49698,N_45985);
and UO_3780 (O_3780,N_48885,N_46585);
nand UO_3781 (O_3781,N_47296,N_47997);
nor UO_3782 (O_3782,N_46684,N_46978);
nor UO_3783 (O_3783,N_49637,N_47921);
or UO_3784 (O_3784,N_49520,N_49142);
and UO_3785 (O_3785,N_48317,N_46418);
nor UO_3786 (O_3786,N_46590,N_48334);
nand UO_3787 (O_3787,N_46171,N_49213);
xor UO_3788 (O_3788,N_49566,N_48068);
nand UO_3789 (O_3789,N_46761,N_48192);
nand UO_3790 (O_3790,N_47718,N_45155);
xnor UO_3791 (O_3791,N_49987,N_48026);
nand UO_3792 (O_3792,N_45636,N_48997);
nand UO_3793 (O_3793,N_47480,N_45875);
or UO_3794 (O_3794,N_47696,N_46962);
nor UO_3795 (O_3795,N_48345,N_49740);
or UO_3796 (O_3796,N_49911,N_47419);
and UO_3797 (O_3797,N_48375,N_45612);
or UO_3798 (O_3798,N_45398,N_46451);
or UO_3799 (O_3799,N_47170,N_48028);
or UO_3800 (O_3800,N_45586,N_45172);
xor UO_3801 (O_3801,N_47600,N_45070);
and UO_3802 (O_3802,N_48360,N_49249);
or UO_3803 (O_3803,N_49504,N_46931);
nand UO_3804 (O_3804,N_48617,N_49302);
xor UO_3805 (O_3805,N_47503,N_46254);
or UO_3806 (O_3806,N_47913,N_45999);
xor UO_3807 (O_3807,N_49845,N_48984);
xor UO_3808 (O_3808,N_46210,N_49402);
nand UO_3809 (O_3809,N_49840,N_49557);
xor UO_3810 (O_3810,N_49620,N_49964);
and UO_3811 (O_3811,N_47956,N_47233);
nand UO_3812 (O_3812,N_49254,N_49674);
xor UO_3813 (O_3813,N_45401,N_49950);
or UO_3814 (O_3814,N_47498,N_45645);
or UO_3815 (O_3815,N_46376,N_48333);
xor UO_3816 (O_3816,N_47328,N_45538);
nand UO_3817 (O_3817,N_49999,N_46836);
nor UO_3818 (O_3818,N_49630,N_48271);
and UO_3819 (O_3819,N_45265,N_45869);
xnor UO_3820 (O_3820,N_45035,N_47893);
and UO_3821 (O_3821,N_49659,N_48850);
and UO_3822 (O_3822,N_47208,N_48064);
xor UO_3823 (O_3823,N_48524,N_47184);
or UO_3824 (O_3824,N_48220,N_45706);
or UO_3825 (O_3825,N_47527,N_49747);
nor UO_3826 (O_3826,N_47912,N_47692);
or UO_3827 (O_3827,N_49622,N_46210);
xnor UO_3828 (O_3828,N_49213,N_47274);
xor UO_3829 (O_3829,N_45986,N_48337);
or UO_3830 (O_3830,N_47885,N_47027);
xor UO_3831 (O_3831,N_47893,N_47799);
and UO_3832 (O_3832,N_48468,N_46972);
or UO_3833 (O_3833,N_45240,N_48575);
and UO_3834 (O_3834,N_48265,N_48147);
nand UO_3835 (O_3835,N_48316,N_45656);
xnor UO_3836 (O_3836,N_45918,N_48453);
nand UO_3837 (O_3837,N_46828,N_47299);
xnor UO_3838 (O_3838,N_49423,N_45276);
or UO_3839 (O_3839,N_49042,N_47339);
xnor UO_3840 (O_3840,N_45744,N_46067);
or UO_3841 (O_3841,N_49707,N_48297);
and UO_3842 (O_3842,N_48115,N_47439);
xor UO_3843 (O_3843,N_46381,N_48729);
xnor UO_3844 (O_3844,N_45104,N_45959);
xnor UO_3845 (O_3845,N_48129,N_49651);
xnor UO_3846 (O_3846,N_47077,N_47862);
xnor UO_3847 (O_3847,N_47445,N_46018);
nand UO_3848 (O_3848,N_46047,N_49790);
or UO_3849 (O_3849,N_47450,N_47819);
nand UO_3850 (O_3850,N_46747,N_49346);
nand UO_3851 (O_3851,N_45303,N_45256);
xor UO_3852 (O_3852,N_46576,N_46417);
and UO_3853 (O_3853,N_45649,N_46247);
nand UO_3854 (O_3854,N_47776,N_49771);
xor UO_3855 (O_3855,N_45861,N_45004);
nand UO_3856 (O_3856,N_47440,N_46921);
nor UO_3857 (O_3857,N_46880,N_49985);
or UO_3858 (O_3858,N_45049,N_49242);
nor UO_3859 (O_3859,N_49049,N_46824);
xor UO_3860 (O_3860,N_46419,N_47417);
nor UO_3861 (O_3861,N_45399,N_45574);
nand UO_3862 (O_3862,N_47986,N_47326);
and UO_3863 (O_3863,N_47963,N_46762);
nor UO_3864 (O_3864,N_47188,N_49316);
nor UO_3865 (O_3865,N_49842,N_49957);
or UO_3866 (O_3866,N_45113,N_46217);
nand UO_3867 (O_3867,N_49986,N_46047);
and UO_3868 (O_3868,N_48186,N_45714);
nor UO_3869 (O_3869,N_46460,N_49110);
xnor UO_3870 (O_3870,N_49224,N_48008);
nand UO_3871 (O_3871,N_46719,N_49109);
xnor UO_3872 (O_3872,N_46062,N_49866);
xnor UO_3873 (O_3873,N_49024,N_47257);
or UO_3874 (O_3874,N_46214,N_45165);
xnor UO_3875 (O_3875,N_47014,N_46338);
nor UO_3876 (O_3876,N_46760,N_48366);
or UO_3877 (O_3877,N_45476,N_47626);
nor UO_3878 (O_3878,N_49912,N_45695);
and UO_3879 (O_3879,N_45575,N_45246);
and UO_3880 (O_3880,N_49713,N_49455);
xor UO_3881 (O_3881,N_47376,N_48686);
xnor UO_3882 (O_3882,N_49511,N_47735);
or UO_3883 (O_3883,N_45435,N_45082);
or UO_3884 (O_3884,N_45591,N_46122);
or UO_3885 (O_3885,N_49927,N_49667);
xnor UO_3886 (O_3886,N_45517,N_46318);
nor UO_3887 (O_3887,N_46010,N_47816);
nand UO_3888 (O_3888,N_46030,N_48479);
or UO_3889 (O_3889,N_47104,N_48859);
or UO_3890 (O_3890,N_46838,N_49142);
and UO_3891 (O_3891,N_47251,N_45031);
nor UO_3892 (O_3892,N_47781,N_45491);
xnor UO_3893 (O_3893,N_49063,N_45049);
xnor UO_3894 (O_3894,N_49453,N_48066);
nand UO_3895 (O_3895,N_49016,N_47457);
and UO_3896 (O_3896,N_46314,N_46748);
or UO_3897 (O_3897,N_49954,N_46166);
nand UO_3898 (O_3898,N_49114,N_46102);
or UO_3899 (O_3899,N_48727,N_47528);
nand UO_3900 (O_3900,N_49376,N_47355);
nand UO_3901 (O_3901,N_47705,N_46971);
and UO_3902 (O_3902,N_48406,N_45197);
xor UO_3903 (O_3903,N_45249,N_48402);
nand UO_3904 (O_3904,N_45333,N_48166);
and UO_3905 (O_3905,N_48881,N_46097);
xor UO_3906 (O_3906,N_49932,N_49584);
nor UO_3907 (O_3907,N_49206,N_47551);
or UO_3908 (O_3908,N_47934,N_46177);
xnor UO_3909 (O_3909,N_46458,N_47290);
nor UO_3910 (O_3910,N_49730,N_45757);
or UO_3911 (O_3911,N_45201,N_47445);
nand UO_3912 (O_3912,N_47708,N_46451);
and UO_3913 (O_3913,N_45052,N_45207);
nor UO_3914 (O_3914,N_45987,N_45890);
nor UO_3915 (O_3915,N_46644,N_46139);
or UO_3916 (O_3916,N_47045,N_48527);
nand UO_3917 (O_3917,N_47804,N_48836);
xor UO_3918 (O_3918,N_48454,N_48108);
and UO_3919 (O_3919,N_47756,N_48914);
xnor UO_3920 (O_3920,N_46861,N_46444);
nor UO_3921 (O_3921,N_47874,N_47386);
nor UO_3922 (O_3922,N_49362,N_45036);
nor UO_3923 (O_3923,N_45866,N_49519);
nor UO_3924 (O_3924,N_48517,N_45281);
xor UO_3925 (O_3925,N_45378,N_45305);
xor UO_3926 (O_3926,N_47345,N_48569);
or UO_3927 (O_3927,N_47553,N_47869);
and UO_3928 (O_3928,N_47388,N_45317);
xor UO_3929 (O_3929,N_49413,N_47211);
nand UO_3930 (O_3930,N_47978,N_48399);
nor UO_3931 (O_3931,N_47535,N_47552);
and UO_3932 (O_3932,N_46756,N_48194);
nand UO_3933 (O_3933,N_45369,N_45874);
nor UO_3934 (O_3934,N_45222,N_49421);
nand UO_3935 (O_3935,N_45762,N_48191);
xor UO_3936 (O_3936,N_48798,N_46520);
nand UO_3937 (O_3937,N_47999,N_46216);
or UO_3938 (O_3938,N_46917,N_48665);
and UO_3939 (O_3939,N_45233,N_49415);
nand UO_3940 (O_3940,N_48848,N_48483);
nand UO_3941 (O_3941,N_48749,N_48269);
xnor UO_3942 (O_3942,N_46609,N_48134);
nor UO_3943 (O_3943,N_46808,N_49503);
or UO_3944 (O_3944,N_46898,N_49308);
or UO_3945 (O_3945,N_48099,N_46112);
nand UO_3946 (O_3946,N_46752,N_49306);
and UO_3947 (O_3947,N_49648,N_46524);
xnor UO_3948 (O_3948,N_49182,N_49849);
nor UO_3949 (O_3949,N_49401,N_46751);
or UO_3950 (O_3950,N_46300,N_49062);
or UO_3951 (O_3951,N_47458,N_48555);
or UO_3952 (O_3952,N_49213,N_48260);
xor UO_3953 (O_3953,N_46412,N_49527);
or UO_3954 (O_3954,N_46458,N_47591);
nor UO_3955 (O_3955,N_46465,N_48515);
xnor UO_3956 (O_3956,N_47391,N_45945);
and UO_3957 (O_3957,N_46680,N_47469);
and UO_3958 (O_3958,N_46376,N_48380);
xor UO_3959 (O_3959,N_45744,N_46989);
or UO_3960 (O_3960,N_48846,N_47056);
or UO_3961 (O_3961,N_48715,N_47189);
and UO_3962 (O_3962,N_45785,N_48735);
xnor UO_3963 (O_3963,N_49179,N_48461);
and UO_3964 (O_3964,N_48931,N_46378);
nor UO_3965 (O_3965,N_47211,N_45112);
xor UO_3966 (O_3966,N_48284,N_45807);
or UO_3967 (O_3967,N_45279,N_45612);
xnor UO_3968 (O_3968,N_48635,N_48923);
or UO_3969 (O_3969,N_49928,N_48198);
xnor UO_3970 (O_3970,N_46251,N_48290);
and UO_3971 (O_3971,N_45294,N_45241);
nand UO_3972 (O_3972,N_45285,N_48746);
nor UO_3973 (O_3973,N_48997,N_47489);
or UO_3974 (O_3974,N_49336,N_45405);
nand UO_3975 (O_3975,N_46507,N_46023);
and UO_3976 (O_3976,N_46176,N_45903);
and UO_3977 (O_3977,N_48549,N_48670);
and UO_3978 (O_3978,N_46063,N_48728);
nor UO_3979 (O_3979,N_47666,N_48078);
xor UO_3980 (O_3980,N_49095,N_45984);
xor UO_3981 (O_3981,N_47216,N_46087);
nand UO_3982 (O_3982,N_47573,N_49678);
or UO_3983 (O_3983,N_49174,N_48039);
or UO_3984 (O_3984,N_45278,N_47634);
xnor UO_3985 (O_3985,N_46557,N_47589);
or UO_3986 (O_3986,N_49526,N_47013);
or UO_3987 (O_3987,N_47743,N_46602);
xor UO_3988 (O_3988,N_47196,N_49460);
nor UO_3989 (O_3989,N_49369,N_45878);
nand UO_3990 (O_3990,N_49959,N_48049);
xnor UO_3991 (O_3991,N_45544,N_46727);
or UO_3992 (O_3992,N_48990,N_48350);
nand UO_3993 (O_3993,N_48470,N_48130);
xnor UO_3994 (O_3994,N_45682,N_47771);
nand UO_3995 (O_3995,N_45116,N_45055);
xor UO_3996 (O_3996,N_45762,N_47456);
and UO_3997 (O_3997,N_49116,N_49954);
nor UO_3998 (O_3998,N_47533,N_49452);
nand UO_3999 (O_3999,N_49198,N_46692);
xnor UO_4000 (O_4000,N_49950,N_45688);
nand UO_4001 (O_4001,N_47505,N_49436);
nand UO_4002 (O_4002,N_45926,N_49959);
xnor UO_4003 (O_4003,N_49186,N_49905);
or UO_4004 (O_4004,N_47077,N_46731);
and UO_4005 (O_4005,N_47395,N_49046);
or UO_4006 (O_4006,N_47837,N_45899);
nor UO_4007 (O_4007,N_45845,N_49148);
nor UO_4008 (O_4008,N_45110,N_48412);
nand UO_4009 (O_4009,N_49811,N_45531);
or UO_4010 (O_4010,N_48395,N_45075);
nand UO_4011 (O_4011,N_46685,N_47602);
and UO_4012 (O_4012,N_48046,N_46734);
or UO_4013 (O_4013,N_46194,N_46608);
xnor UO_4014 (O_4014,N_48822,N_46601);
and UO_4015 (O_4015,N_48049,N_46483);
nand UO_4016 (O_4016,N_49801,N_48134);
and UO_4017 (O_4017,N_47192,N_46687);
xor UO_4018 (O_4018,N_47050,N_45648);
nor UO_4019 (O_4019,N_45251,N_46285);
and UO_4020 (O_4020,N_45492,N_47268);
and UO_4021 (O_4021,N_46709,N_45995);
or UO_4022 (O_4022,N_48392,N_48047);
nand UO_4023 (O_4023,N_46011,N_46910);
nor UO_4024 (O_4024,N_48543,N_49075);
xnor UO_4025 (O_4025,N_45161,N_45592);
and UO_4026 (O_4026,N_46119,N_48463);
xnor UO_4027 (O_4027,N_48927,N_46180);
nand UO_4028 (O_4028,N_46064,N_47393);
nor UO_4029 (O_4029,N_47259,N_48743);
or UO_4030 (O_4030,N_46427,N_46887);
and UO_4031 (O_4031,N_48634,N_45468);
nand UO_4032 (O_4032,N_45486,N_47236);
and UO_4033 (O_4033,N_48119,N_45773);
nand UO_4034 (O_4034,N_45060,N_48214);
or UO_4035 (O_4035,N_46264,N_45652);
or UO_4036 (O_4036,N_45416,N_49526);
nand UO_4037 (O_4037,N_45199,N_47169);
xor UO_4038 (O_4038,N_48574,N_49803);
nand UO_4039 (O_4039,N_49359,N_47633);
or UO_4040 (O_4040,N_48734,N_47841);
nand UO_4041 (O_4041,N_48787,N_49763);
xnor UO_4042 (O_4042,N_45855,N_48306);
nor UO_4043 (O_4043,N_46377,N_48006);
or UO_4044 (O_4044,N_49090,N_45180);
nor UO_4045 (O_4045,N_46162,N_48573);
or UO_4046 (O_4046,N_48680,N_49331);
xor UO_4047 (O_4047,N_46578,N_49929);
and UO_4048 (O_4048,N_48038,N_45158);
nor UO_4049 (O_4049,N_49352,N_49143);
nor UO_4050 (O_4050,N_49165,N_45542);
nor UO_4051 (O_4051,N_46218,N_45413);
xnor UO_4052 (O_4052,N_48483,N_48442);
xnor UO_4053 (O_4053,N_45730,N_46162);
nor UO_4054 (O_4054,N_49302,N_45810);
and UO_4055 (O_4055,N_45857,N_46336);
nor UO_4056 (O_4056,N_48178,N_49537);
xor UO_4057 (O_4057,N_48579,N_45836);
nand UO_4058 (O_4058,N_45023,N_45389);
and UO_4059 (O_4059,N_45736,N_45038);
xor UO_4060 (O_4060,N_45247,N_47313);
nand UO_4061 (O_4061,N_47060,N_48637);
or UO_4062 (O_4062,N_46050,N_46375);
or UO_4063 (O_4063,N_47382,N_45434);
nor UO_4064 (O_4064,N_47493,N_48429);
and UO_4065 (O_4065,N_45987,N_49242);
nand UO_4066 (O_4066,N_46356,N_49778);
and UO_4067 (O_4067,N_49026,N_45093);
or UO_4068 (O_4068,N_49426,N_49831);
nor UO_4069 (O_4069,N_46007,N_46639);
nor UO_4070 (O_4070,N_46592,N_49528);
and UO_4071 (O_4071,N_48042,N_46382);
or UO_4072 (O_4072,N_48738,N_47292);
and UO_4073 (O_4073,N_49345,N_48582);
and UO_4074 (O_4074,N_47542,N_48651);
xor UO_4075 (O_4075,N_45661,N_49535);
or UO_4076 (O_4076,N_47250,N_46236);
or UO_4077 (O_4077,N_49965,N_48798);
nand UO_4078 (O_4078,N_45246,N_49759);
or UO_4079 (O_4079,N_47666,N_45940);
and UO_4080 (O_4080,N_47344,N_46969);
xor UO_4081 (O_4081,N_45655,N_48915);
nand UO_4082 (O_4082,N_45037,N_49814);
or UO_4083 (O_4083,N_49273,N_45566);
nor UO_4084 (O_4084,N_49679,N_46846);
xnor UO_4085 (O_4085,N_48144,N_46769);
or UO_4086 (O_4086,N_49533,N_46774);
xnor UO_4087 (O_4087,N_46562,N_49237);
or UO_4088 (O_4088,N_47427,N_47511);
or UO_4089 (O_4089,N_48872,N_46313);
and UO_4090 (O_4090,N_47524,N_49044);
or UO_4091 (O_4091,N_48021,N_49794);
nand UO_4092 (O_4092,N_45247,N_47489);
nor UO_4093 (O_4093,N_48103,N_46743);
nor UO_4094 (O_4094,N_47740,N_49691);
xor UO_4095 (O_4095,N_48160,N_45598);
and UO_4096 (O_4096,N_47748,N_48605);
xor UO_4097 (O_4097,N_48184,N_48049);
nand UO_4098 (O_4098,N_46493,N_45900);
and UO_4099 (O_4099,N_45358,N_49215);
nor UO_4100 (O_4100,N_45250,N_47762);
and UO_4101 (O_4101,N_49172,N_46906);
nand UO_4102 (O_4102,N_49385,N_48938);
xnor UO_4103 (O_4103,N_47401,N_48600);
or UO_4104 (O_4104,N_49824,N_49248);
xor UO_4105 (O_4105,N_48917,N_45335);
xnor UO_4106 (O_4106,N_47305,N_47846);
or UO_4107 (O_4107,N_46440,N_47840);
or UO_4108 (O_4108,N_46691,N_46080);
and UO_4109 (O_4109,N_45298,N_49997);
nor UO_4110 (O_4110,N_45152,N_45569);
nor UO_4111 (O_4111,N_45063,N_45096);
and UO_4112 (O_4112,N_49767,N_48723);
or UO_4113 (O_4113,N_48447,N_48802);
and UO_4114 (O_4114,N_48284,N_45897);
xnor UO_4115 (O_4115,N_46096,N_48665);
and UO_4116 (O_4116,N_46698,N_46202);
nor UO_4117 (O_4117,N_48975,N_48776);
nand UO_4118 (O_4118,N_47702,N_45890);
nand UO_4119 (O_4119,N_48975,N_48529);
xnor UO_4120 (O_4120,N_46761,N_49362);
and UO_4121 (O_4121,N_47119,N_47270);
and UO_4122 (O_4122,N_49769,N_47621);
nor UO_4123 (O_4123,N_47170,N_47915);
and UO_4124 (O_4124,N_48832,N_48917);
xnor UO_4125 (O_4125,N_49034,N_49127);
and UO_4126 (O_4126,N_45926,N_45346);
or UO_4127 (O_4127,N_47750,N_46296);
nor UO_4128 (O_4128,N_47213,N_48780);
and UO_4129 (O_4129,N_49251,N_48743);
nand UO_4130 (O_4130,N_45622,N_46074);
xnor UO_4131 (O_4131,N_49927,N_48346);
or UO_4132 (O_4132,N_47349,N_46331);
nand UO_4133 (O_4133,N_49538,N_49725);
nand UO_4134 (O_4134,N_47372,N_45059);
nor UO_4135 (O_4135,N_45723,N_48271);
nand UO_4136 (O_4136,N_48814,N_49720);
xor UO_4137 (O_4137,N_45339,N_46611);
and UO_4138 (O_4138,N_47275,N_49085);
nor UO_4139 (O_4139,N_45400,N_45860);
or UO_4140 (O_4140,N_49276,N_49799);
nand UO_4141 (O_4141,N_45381,N_49391);
and UO_4142 (O_4142,N_49175,N_47450);
xor UO_4143 (O_4143,N_47763,N_46450);
and UO_4144 (O_4144,N_46080,N_49505);
xnor UO_4145 (O_4145,N_48254,N_45787);
xor UO_4146 (O_4146,N_47324,N_46017);
nor UO_4147 (O_4147,N_46156,N_47944);
nand UO_4148 (O_4148,N_45513,N_47824);
nand UO_4149 (O_4149,N_48901,N_49375);
and UO_4150 (O_4150,N_49375,N_47977);
nand UO_4151 (O_4151,N_45227,N_46138);
nand UO_4152 (O_4152,N_48233,N_45527);
and UO_4153 (O_4153,N_49106,N_45551);
and UO_4154 (O_4154,N_47283,N_48727);
or UO_4155 (O_4155,N_48704,N_45657);
or UO_4156 (O_4156,N_49042,N_48805);
and UO_4157 (O_4157,N_46145,N_49669);
nor UO_4158 (O_4158,N_48039,N_46326);
or UO_4159 (O_4159,N_47234,N_47876);
xnor UO_4160 (O_4160,N_45807,N_49033);
or UO_4161 (O_4161,N_48833,N_49819);
nor UO_4162 (O_4162,N_48208,N_49705);
and UO_4163 (O_4163,N_47590,N_45682);
nand UO_4164 (O_4164,N_48226,N_45388);
and UO_4165 (O_4165,N_45094,N_49857);
or UO_4166 (O_4166,N_48095,N_47109);
or UO_4167 (O_4167,N_46253,N_48419);
nand UO_4168 (O_4168,N_49262,N_48625);
nand UO_4169 (O_4169,N_49449,N_47828);
and UO_4170 (O_4170,N_46586,N_48395);
nand UO_4171 (O_4171,N_47567,N_45146);
and UO_4172 (O_4172,N_46959,N_46605);
nand UO_4173 (O_4173,N_46850,N_48052);
and UO_4174 (O_4174,N_49148,N_45766);
nor UO_4175 (O_4175,N_47050,N_49305);
and UO_4176 (O_4176,N_49240,N_47511);
nand UO_4177 (O_4177,N_46890,N_46103);
nand UO_4178 (O_4178,N_48965,N_48103);
or UO_4179 (O_4179,N_47697,N_49362);
nand UO_4180 (O_4180,N_47253,N_47836);
nand UO_4181 (O_4181,N_47966,N_49232);
nor UO_4182 (O_4182,N_48640,N_45106);
nor UO_4183 (O_4183,N_45859,N_47335);
and UO_4184 (O_4184,N_45386,N_46383);
and UO_4185 (O_4185,N_45508,N_46680);
and UO_4186 (O_4186,N_48857,N_47403);
nor UO_4187 (O_4187,N_47412,N_49672);
nand UO_4188 (O_4188,N_49423,N_45492);
or UO_4189 (O_4189,N_49320,N_49352);
nor UO_4190 (O_4190,N_48760,N_49827);
or UO_4191 (O_4191,N_46517,N_46806);
xor UO_4192 (O_4192,N_47118,N_46294);
and UO_4193 (O_4193,N_45855,N_46953);
nand UO_4194 (O_4194,N_46365,N_45095);
nand UO_4195 (O_4195,N_49027,N_49704);
nor UO_4196 (O_4196,N_46235,N_45061);
nor UO_4197 (O_4197,N_49517,N_46539);
or UO_4198 (O_4198,N_47388,N_49919);
or UO_4199 (O_4199,N_49857,N_49755);
and UO_4200 (O_4200,N_49686,N_49431);
or UO_4201 (O_4201,N_46173,N_45181);
xnor UO_4202 (O_4202,N_45004,N_47841);
or UO_4203 (O_4203,N_45056,N_47275);
or UO_4204 (O_4204,N_45553,N_46425);
xor UO_4205 (O_4205,N_48549,N_49390);
nor UO_4206 (O_4206,N_47313,N_46226);
or UO_4207 (O_4207,N_46263,N_47569);
nand UO_4208 (O_4208,N_49999,N_48233);
nor UO_4209 (O_4209,N_48431,N_48390);
xor UO_4210 (O_4210,N_46623,N_45438);
and UO_4211 (O_4211,N_46025,N_49907);
or UO_4212 (O_4212,N_48095,N_46157);
nand UO_4213 (O_4213,N_45231,N_45140);
nor UO_4214 (O_4214,N_49538,N_47724);
and UO_4215 (O_4215,N_47155,N_47010);
xnor UO_4216 (O_4216,N_45494,N_46173);
nor UO_4217 (O_4217,N_48745,N_49814);
nor UO_4218 (O_4218,N_48668,N_48874);
xnor UO_4219 (O_4219,N_48424,N_45940);
nor UO_4220 (O_4220,N_47033,N_45845);
nor UO_4221 (O_4221,N_46381,N_49595);
nand UO_4222 (O_4222,N_48027,N_49040);
and UO_4223 (O_4223,N_49206,N_48878);
nand UO_4224 (O_4224,N_49708,N_46105);
xnor UO_4225 (O_4225,N_46615,N_47416);
xnor UO_4226 (O_4226,N_48648,N_47830);
or UO_4227 (O_4227,N_47392,N_46043);
nor UO_4228 (O_4228,N_47247,N_47892);
xnor UO_4229 (O_4229,N_46183,N_48797);
nand UO_4230 (O_4230,N_49467,N_49307);
or UO_4231 (O_4231,N_47093,N_47777);
xor UO_4232 (O_4232,N_46314,N_48812);
xnor UO_4233 (O_4233,N_49330,N_45231);
and UO_4234 (O_4234,N_49519,N_49873);
nor UO_4235 (O_4235,N_45987,N_49438);
or UO_4236 (O_4236,N_49178,N_49268);
nor UO_4237 (O_4237,N_45543,N_48305);
or UO_4238 (O_4238,N_45935,N_49382);
nand UO_4239 (O_4239,N_46475,N_48355);
nand UO_4240 (O_4240,N_45289,N_47516);
and UO_4241 (O_4241,N_45101,N_49534);
nand UO_4242 (O_4242,N_46043,N_45921);
xor UO_4243 (O_4243,N_49340,N_49104);
and UO_4244 (O_4244,N_49311,N_47689);
xor UO_4245 (O_4245,N_49944,N_48141);
nor UO_4246 (O_4246,N_46986,N_48519);
xor UO_4247 (O_4247,N_46946,N_46064);
or UO_4248 (O_4248,N_48091,N_46866);
or UO_4249 (O_4249,N_49677,N_47206);
and UO_4250 (O_4250,N_49762,N_49142);
or UO_4251 (O_4251,N_47088,N_46519);
or UO_4252 (O_4252,N_48477,N_46251);
nand UO_4253 (O_4253,N_48973,N_49394);
nand UO_4254 (O_4254,N_49982,N_45597);
and UO_4255 (O_4255,N_49942,N_45928);
nor UO_4256 (O_4256,N_48225,N_46740);
and UO_4257 (O_4257,N_45517,N_45397);
and UO_4258 (O_4258,N_46117,N_45685);
or UO_4259 (O_4259,N_45580,N_45839);
xor UO_4260 (O_4260,N_48486,N_49568);
or UO_4261 (O_4261,N_47658,N_47177);
and UO_4262 (O_4262,N_45923,N_48799);
xor UO_4263 (O_4263,N_45886,N_46769);
nor UO_4264 (O_4264,N_48585,N_45672);
and UO_4265 (O_4265,N_49049,N_46067);
nor UO_4266 (O_4266,N_49668,N_48445);
xnor UO_4267 (O_4267,N_49095,N_48585);
and UO_4268 (O_4268,N_46167,N_49532);
nand UO_4269 (O_4269,N_45608,N_45517);
nand UO_4270 (O_4270,N_49242,N_46707);
or UO_4271 (O_4271,N_45447,N_46100);
nor UO_4272 (O_4272,N_45820,N_47417);
and UO_4273 (O_4273,N_47166,N_48226);
or UO_4274 (O_4274,N_49576,N_45605);
nand UO_4275 (O_4275,N_46690,N_48528);
nor UO_4276 (O_4276,N_49049,N_48694);
xor UO_4277 (O_4277,N_47205,N_49748);
xnor UO_4278 (O_4278,N_48284,N_45224);
or UO_4279 (O_4279,N_49604,N_46188);
or UO_4280 (O_4280,N_48015,N_46391);
and UO_4281 (O_4281,N_49709,N_47847);
or UO_4282 (O_4282,N_47230,N_45751);
nor UO_4283 (O_4283,N_48517,N_48911);
or UO_4284 (O_4284,N_48977,N_49160);
or UO_4285 (O_4285,N_47883,N_46007);
nor UO_4286 (O_4286,N_47994,N_46058);
or UO_4287 (O_4287,N_49206,N_45038);
or UO_4288 (O_4288,N_47489,N_48333);
nor UO_4289 (O_4289,N_47212,N_47604);
nor UO_4290 (O_4290,N_48232,N_46582);
and UO_4291 (O_4291,N_45643,N_46160);
or UO_4292 (O_4292,N_46365,N_49451);
xor UO_4293 (O_4293,N_49767,N_49694);
or UO_4294 (O_4294,N_45105,N_48264);
xnor UO_4295 (O_4295,N_45422,N_49421);
or UO_4296 (O_4296,N_46116,N_49722);
and UO_4297 (O_4297,N_47773,N_47267);
or UO_4298 (O_4298,N_48257,N_47105);
nand UO_4299 (O_4299,N_47451,N_45611);
and UO_4300 (O_4300,N_45028,N_45316);
or UO_4301 (O_4301,N_46632,N_49367);
nand UO_4302 (O_4302,N_46704,N_45762);
and UO_4303 (O_4303,N_47477,N_49695);
nand UO_4304 (O_4304,N_46831,N_49652);
nor UO_4305 (O_4305,N_47887,N_49318);
nand UO_4306 (O_4306,N_45974,N_47090);
xor UO_4307 (O_4307,N_46813,N_49226);
nor UO_4308 (O_4308,N_47998,N_45532);
xnor UO_4309 (O_4309,N_47766,N_45751);
xnor UO_4310 (O_4310,N_47877,N_46019);
xor UO_4311 (O_4311,N_48806,N_47812);
or UO_4312 (O_4312,N_45073,N_47927);
nand UO_4313 (O_4313,N_45870,N_49289);
xor UO_4314 (O_4314,N_49608,N_46955);
or UO_4315 (O_4315,N_49290,N_46095);
nand UO_4316 (O_4316,N_45968,N_45707);
xnor UO_4317 (O_4317,N_48423,N_48595);
xnor UO_4318 (O_4318,N_47366,N_49484);
or UO_4319 (O_4319,N_47571,N_46362);
or UO_4320 (O_4320,N_49542,N_46053);
nand UO_4321 (O_4321,N_47461,N_49307);
or UO_4322 (O_4322,N_46501,N_46752);
or UO_4323 (O_4323,N_49812,N_49873);
and UO_4324 (O_4324,N_48259,N_48704);
and UO_4325 (O_4325,N_45886,N_46502);
nor UO_4326 (O_4326,N_47356,N_46927);
xor UO_4327 (O_4327,N_47991,N_47841);
nor UO_4328 (O_4328,N_49225,N_45155);
and UO_4329 (O_4329,N_49746,N_49156);
and UO_4330 (O_4330,N_45171,N_45631);
nand UO_4331 (O_4331,N_48028,N_47757);
xnor UO_4332 (O_4332,N_48982,N_49594);
or UO_4333 (O_4333,N_47941,N_49791);
and UO_4334 (O_4334,N_45099,N_45601);
or UO_4335 (O_4335,N_46456,N_49522);
or UO_4336 (O_4336,N_48251,N_46891);
and UO_4337 (O_4337,N_47388,N_46413);
and UO_4338 (O_4338,N_48224,N_47919);
xor UO_4339 (O_4339,N_46765,N_46036);
nand UO_4340 (O_4340,N_48918,N_48674);
nor UO_4341 (O_4341,N_49808,N_47348);
xnor UO_4342 (O_4342,N_48089,N_47287);
nor UO_4343 (O_4343,N_45127,N_49379);
nand UO_4344 (O_4344,N_45898,N_48278);
nand UO_4345 (O_4345,N_47459,N_46471);
nand UO_4346 (O_4346,N_46554,N_47753);
xor UO_4347 (O_4347,N_46422,N_45937);
or UO_4348 (O_4348,N_48733,N_46459);
and UO_4349 (O_4349,N_47756,N_48378);
or UO_4350 (O_4350,N_48590,N_49754);
or UO_4351 (O_4351,N_49734,N_45340);
or UO_4352 (O_4352,N_45225,N_45234);
and UO_4353 (O_4353,N_46156,N_46847);
xnor UO_4354 (O_4354,N_49604,N_49213);
nand UO_4355 (O_4355,N_49267,N_47865);
nor UO_4356 (O_4356,N_48705,N_46351);
or UO_4357 (O_4357,N_48768,N_46035);
nor UO_4358 (O_4358,N_48970,N_48645);
xnor UO_4359 (O_4359,N_46270,N_48699);
and UO_4360 (O_4360,N_48674,N_45075);
or UO_4361 (O_4361,N_46331,N_49927);
nand UO_4362 (O_4362,N_45330,N_47547);
xor UO_4363 (O_4363,N_48908,N_45019);
nand UO_4364 (O_4364,N_45716,N_48375);
nand UO_4365 (O_4365,N_48863,N_48888);
nor UO_4366 (O_4366,N_47668,N_45515);
xnor UO_4367 (O_4367,N_47226,N_49041);
or UO_4368 (O_4368,N_48008,N_45589);
nor UO_4369 (O_4369,N_47697,N_48615);
xnor UO_4370 (O_4370,N_48644,N_45121);
or UO_4371 (O_4371,N_46273,N_45472);
nand UO_4372 (O_4372,N_45461,N_47821);
xor UO_4373 (O_4373,N_46223,N_49750);
and UO_4374 (O_4374,N_47328,N_46458);
nand UO_4375 (O_4375,N_49269,N_45137);
nor UO_4376 (O_4376,N_47949,N_45480);
nand UO_4377 (O_4377,N_49980,N_49995);
nand UO_4378 (O_4378,N_46449,N_45974);
and UO_4379 (O_4379,N_46910,N_45029);
or UO_4380 (O_4380,N_45700,N_45005);
and UO_4381 (O_4381,N_47669,N_48057);
or UO_4382 (O_4382,N_46276,N_46332);
xnor UO_4383 (O_4383,N_49977,N_45746);
xor UO_4384 (O_4384,N_48866,N_48816);
xnor UO_4385 (O_4385,N_48875,N_49939);
xor UO_4386 (O_4386,N_48739,N_47024);
or UO_4387 (O_4387,N_46712,N_48805);
and UO_4388 (O_4388,N_49886,N_45101);
nand UO_4389 (O_4389,N_46941,N_47140);
nor UO_4390 (O_4390,N_47140,N_45604);
nand UO_4391 (O_4391,N_49447,N_49030);
or UO_4392 (O_4392,N_49519,N_47929);
nor UO_4393 (O_4393,N_45824,N_47969);
nand UO_4394 (O_4394,N_45665,N_46758);
or UO_4395 (O_4395,N_49480,N_45883);
nand UO_4396 (O_4396,N_47468,N_45107);
nor UO_4397 (O_4397,N_48456,N_49994);
xor UO_4398 (O_4398,N_45403,N_46325);
nor UO_4399 (O_4399,N_45814,N_48325);
nor UO_4400 (O_4400,N_45481,N_45659);
and UO_4401 (O_4401,N_47371,N_46077);
or UO_4402 (O_4402,N_46046,N_48290);
or UO_4403 (O_4403,N_46262,N_46556);
xor UO_4404 (O_4404,N_48071,N_47262);
and UO_4405 (O_4405,N_45672,N_45994);
and UO_4406 (O_4406,N_46595,N_45754);
or UO_4407 (O_4407,N_45768,N_49803);
xor UO_4408 (O_4408,N_49076,N_49160);
or UO_4409 (O_4409,N_45653,N_49361);
and UO_4410 (O_4410,N_47938,N_46116);
and UO_4411 (O_4411,N_47793,N_48007);
or UO_4412 (O_4412,N_49828,N_45258);
xnor UO_4413 (O_4413,N_49618,N_47632);
or UO_4414 (O_4414,N_48668,N_45403);
or UO_4415 (O_4415,N_47427,N_45016);
or UO_4416 (O_4416,N_46960,N_45053);
and UO_4417 (O_4417,N_47566,N_46877);
nand UO_4418 (O_4418,N_48586,N_47934);
nor UO_4419 (O_4419,N_49583,N_45417);
or UO_4420 (O_4420,N_48309,N_47973);
or UO_4421 (O_4421,N_49289,N_49411);
xor UO_4422 (O_4422,N_45022,N_46276);
nand UO_4423 (O_4423,N_47071,N_46547);
or UO_4424 (O_4424,N_49237,N_46807);
nand UO_4425 (O_4425,N_48188,N_45033);
nand UO_4426 (O_4426,N_46442,N_46783);
xnor UO_4427 (O_4427,N_48118,N_46018);
and UO_4428 (O_4428,N_47776,N_46641);
and UO_4429 (O_4429,N_47118,N_47509);
nand UO_4430 (O_4430,N_48403,N_48435);
and UO_4431 (O_4431,N_49520,N_45079);
xnor UO_4432 (O_4432,N_47121,N_48955);
or UO_4433 (O_4433,N_46729,N_48886);
nand UO_4434 (O_4434,N_49531,N_45093);
or UO_4435 (O_4435,N_45670,N_47277);
nor UO_4436 (O_4436,N_48149,N_47780);
nor UO_4437 (O_4437,N_49506,N_49303);
nor UO_4438 (O_4438,N_48519,N_45649);
nand UO_4439 (O_4439,N_45054,N_48922);
nor UO_4440 (O_4440,N_48873,N_46277);
nor UO_4441 (O_4441,N_48122,N_48681);
nand UO_4442 (O_4442,N_46207,N_46373);
xor UO_4443 (O_4443,N_45863,N_47268);
nand UO_4444 (O_4444,N_47745,N_49376);
xnor UO_4445 (O_4445,N_49912,N_48445);
and UO_4446 (O_4446,N_48427,N_47037);
or UO_4447 (O_4447,N_47350,N_48340);
xor UO_4448 (O_4448,N_46649,N_47534);
nand UO_4449 (O_4449,N_45659,N_47647);
xor UO_4450 (O_4450,N_46635,N_47501);
nand UO_4451 (O_4451,N_47444,N_49858);
xor UO_4452 (O_4452,N_46568,N_46450);
or UO_4453 (O_4453,N_48395,N_45142);
nand UO_4454 (O_4454,N_45630,N_48313);
or UO_4455 (O_4455,N_45234,N_48539);
nor UO_4456 (O_4456,N_47984,N_49548);
or UO_4457 (O_4457,N_46953,N_48023);
xnor UO_4458 (O_4458,N_48927,N_49428);
nor UO_4459 (O_4459,N_45725,N_48562);
and UO_4460 (O_4460,N_47573,N_47710);
nor UO_4461 (O_4461,N_47950,N_46236);
and UO_4462 (O_4462,N_46759,N_47248);
nor UO_4463 (O_4463,N_48725,N_47885);
nor UO_4464 (O_4464,N_49875,N_49388);
and UO_4465 (O_4465,N_45425,N_49512);
and UO_4466 (O_4466,N_45073,N_46059);
xnor UO_4467 (O_4467,N_47934,N_45975);
nor UO_4468 (O_4468,N_48679,N_47789);
nor UO_4469 (O_4469,N_45066,N_45385);
nand UO_4470 (O_4470,N_45409,N_46791);
xor UO_4471 (O_4471,N_45168,N_47165);
xor UO_4472 (O_4472,N_47041,N_46024);
and UO_4473 (O_4473,N_47396,N_49704);
xor UO_4474 (O_4474,N_49698,N_48089);
nor UO_4475 (O_4475,N_48073,N_48686);
nand UO_4476 (O_4476,N_48909,N_46848);
or UO_4477 (O_4477,N_46792,N_45504);
xor UO_4478 (O_4478,N_46438,N_45441);
and UO_4479 (O_4479,N_49444,N_49278);
nor UO_4480 (O_4480,N_46444,N_47048);
and UO_4481 (O_4481,N_47989,N_45196);
and UO_4482 (O_4482,N_47032,N_45644);
nor UO_4483 (O_4483,N_45372,N_47351);
nor UO_4484 (O_4484,N_49279,N_47279);
or UO_4485 (O_4485,N_48124,N_46001);
or UO_4486 (O_4486,N_48420,N_48803);
nand UO_4487 (O_4487,N_45389,N_49703);
nor UO_4488 (O_4488,N_45840,N_45764);
xnor UO_4489 (O_4489,N_47858,N_49612);
nand UO_4490 (O_4490,N_47389,N_49509);
xnor UO_4491 (O_4491,N_47078,N_45237);
nand UO_4492 (O_4492,N_49404,N_46860);
or UO_4493 (O_4493,N_46946,N_49493);
xnor UO_4494 (O_4494,N_49712,N_46557);
or UO_4495 (O_4495,N_47448,N_45669);
or UO_4496 (O_4496,N_49285,N_48595);
xor UO_4497 (O_4497,N_45099,N_45824);
nand UO_4498 (O_4498,N_46154,N_47063);
and UO_4499 (O_4499,N_49247,N_45883);
or UO_4500 (O_4500,N_48893,N_48325);
or UO_4501 (O_4501,N_46268,N_49675);
nand UO_4502 (O_4502,N_46363,N_49811);
and UO_4503 (O_4503,N_45640,N_45831);
or UO_4504 (O_4504,N_46462,N_49162);
nand UO_4505 (O_4505,N_48723,N_48283);
and UO_4506 (O_4506,N_47202,N_49987);
and UO_4507 (O_4507,N_47189,N_49510);
nand UO_4508 (O_4508,N_45041,N_49104);
and UO_4509 (O_4509,N_48382,N_47665);
and UO_4510 (O_4510,N_45384,N_47170);
or UO_4511 (O_4511,N_47301,N_48312);
and UO_4512 (O_4512,N_46586,N_47722);
or UO_4513 (O_4513,N_49643,N_49287);
nor UO_4514 (O_4514,N_46134,N_48524);
xnor UO_4515 (O_4515,N_45728,N_48669);
xnor UO_4516 (O_4516,N_49311,N_45398);
nand UO_4517 (O_4517,N_49547,N_46647);
nor UO_4518 (O_4518,N_45497,N_46413);
xor UO_4519 (O_4519,N_46135,N_48377);
and UO_4520 (O_4520,N_49747,N_45460);
and UO_4521 (O_4521,N_49789,N_48620);
xor UO_4522 (O_4522,N_45686,N_45094);
nor UO_4523 (O_4523,N_49755,N_47892);
and UO_4524 (O_4524,N_45187,N_48571);
or UO_4525 (O_4525,N_45323,N_46701);
nand UO_4526 (O_4526,N_48957,N_47008);
nand UO_4527 (O_4527,N_49302,N_48523);
xnor UO_4528 (O_4528,N_48703,N_47783);
nand UO_4529 (O_4529,N_48356,N_45789);
nor UO_4530 (O_4530,N_48409,N_47313);
or UO_4531 (O_4531,N_49414,N_48137);
and UO_4532 (O_4532,N_49625,N_49274);
nor UO_4533 (O_4533,N_49834,N_49333);
nand UO_4534 (O_4534,N_46035,N_49823);
nand UO_4535 (O_4535,N_49289,N_49408);
xor UO_4536 (O_4536,N_45396,N_48712);
nand UO_4537 (O_4537,N_45116,N_45577);
and UO_4538 (O_4538,N_49399,N_45093);
xor UO_4539 (O_4539,N_46799,N_47517);
xor UO_4540 (O_4540,N_49204,N_46683);
xnor UO_4541 (O_4541,N_46737,N_47046);
nor UO_4542 (O_4542,N_45798,N_46495);
nor UO_4543 (O_4543,N_45069,N_49203);
nor UO_4544 (O_4544,N_45399,N_46209);
nand UO_4545 (O_4545,N_48659,N_48989);
xnor UO_4546 (O_4546,N_46720,N_47368);
nor UO_4547 (O_4547,N_45783,N_47254);
xor UO_4548 (O_4548,N_48562,N_49381);
nand UO_4549 (O_4549,N_47221,N_47338);
or UO_4550 (O_4550,N_46271,N_48251);
or UO_4551 (O_4551,N_49607,N_48370);
xnor UO_4552 (O_4552,N_46266,N_47359);
xor UO_4553 (O_4553,N_49736,N_45134);
and UO_4554 (O_4554,N_49725,N_47995);
or UO_4555 (O_4555,N_46765,N_49241);
or UO_4556 (O_4556,N_47277,N_46859);
nand UO_4557 (O_4557,N_47625,N_49667);
or UO_4558 (O_4558,N_45448,N_47644);
nor UO_4559 (O_4559,N_46624,N_48175);
nand UO_4560 (O_4560,N_45184,N_48073);
and UO_4561 (O_4561,N_48326,N_47550);
nor UO_4562 (O_4562,N_45194,N_46404);
xnor UO_4563 (O_4563,N_45293,N_49029);
nor UO_4564 (O_4564,N_46495,N_45202);
xor UO_4565 (O_4565,N_46610,N_46376);
xor UO_4566 (O_4566,N_48780,N_48542);
nor UO_4567 (O_4567,N_49038,N_46045);
and UO_4568 (O_4568,N_46844,N_49285);
nor UO_4569 (O_4569,N_45947,N_49834);
xnor UO_4570 (O_4570,N_49687,N_49614);
xnor UO_4571 (O_4571,N_46332,N_46028);
or UO_4572 (O_4572,N_46632,N_47604);
or UO_4573 (O_4573,N_48374,N_46037);
nor UO_4574 (O_4574,N_47900,N_49443);
xor UO_4575 (O_4575,N_47769,N_47580);
xor UO_4576 (O_4576,N_46948,N_46393);
and UO_4577 (O_4577,N_49498,N_45270);
or UO_4578 (O_4578,N_49373,N_46160);
nor UO_4579 (O_4579,N_46234,N_47340);
xnor UO_4580 (O_4580,N_49035,N_48158);
nand UO_4581 (O_4581,N_48218,N_47879);
nand UO_4582 (O_4582,N_46844,N_45667);
xnor UO_4583 (O_4583,N_47060,N_49498);
nand UO_4584 (O_4584,N_49907,N_46621);
nor UO_4585 (O_4585,N_49660,N_46292);
nor UO_4586 (O_4586,N_47775,N_47410);
nand UO_4587 (O_4587,N_47911,N_49098);
nor UO_4588 (O_4588,N_45369,N_49643);
or UO_4589 (O_4589,N_45128,N_47728);
nor UO_4590 (O_4590,N_48738,N_45318);
and UO_4591 (O_4591,N_45741,N_49600);
or UO_4592 (O_4592,N_45654,N_46846);
nor UO_4593 (O_4593,N_47528,N_46813);
and UO_4594 (O_4594,N_47323,N_47229);
and UO_4595 (O_4595,N_47994,N_46484);
nor UO_4596 (O_4596,N_49724,N_46357);
xnor UO_4597 (O_4597,N_45979,N_45283);
nand UO_4598 (O_4598,N_46479,N_45566);
nand UO_4599 (O_4599,N_46012,N_46086);
xnor UO_4600 (O_4600,N_49912,N_48910);
or UO_4601 (O_4601,N_46369,N_45051);
or UO_4602 (O_4602,N_45495,N_46535);
nand UO_4603 (O_4603,N_46507,N_48825);
or UO_4604 (O_4604,N_49869,N_49257);
nand UO_4605 (O_4605,N_48205,N_48605);
nor UO_4606 (O_4606,N_47114,N_45547);
nor UO_4607 (O_4607,N_48931,N_46794);
or UO_4608 (O_4608,N_47402,N_46226);
xnor UO_4609 (O_4609,N_48963,N_47007);
and UO_4610 (O_4610,N_45709,N_47301);
or UO_4611 (O_4611,N_47654,N_47748);
nand UO_4612 (O_4612,N_47717,N_45728);
xor UO_4613 (O_4613,N_48421,N_48127);
and UO_4614 (O_4614,N_47310,N_48628);
nand UO_4615 (O_4615,N_49852,N_45790);
and UO_4616 (O_4616,N_46185,N_46765);
or UO_4617 (O_4617,N_45123,N_49966);
xnor UO_4618 (O_4618,N_47347,N_46279);
xor UO_4619 (O_4619,N_46131,N_48646);
nor UO_4620 (O_4620,N_48163,N_45734);
or UO_4621 (O_4621,N_45957,N_48850);
and UO_4622 (O_4622,N_49717,N_49815);
nor UO_4623 (O_4623,N_46478,N_45132);
xnor UO_4624 (O_4624,N_46231,N_49567);
or UO_4625 (O_4625,N_49469,N_48028);
nor UO_4626 (O_4626,N_45233,N_47333);
and UO_4627 (O_4627,N_47935,N_49543);
nor UO_4628 (O_4628,N_48981,N_45211);
and UO_4629 (O_4629,N_48503,N_45357);
or UO_4630 (O_4630,N_47910,N_46463);
nand UO_4631 (O_4631,N_47960,N_49968);
xor UO_4632 (O_4632,N_46533,N_47855);
and UO_4633 (O_4633,N_47522,N_48462);
nand UO_4634 (O_4634,N_49759,N_47280);
nand UO_4635 (O_4635,N_46661,N_45333);
and UO_4636 (O_4636,N_47112,N_47984);
or UO_4637 (O_4637,N_49662,N_45330);
nand UO_4638 (O_4638,N_47532,N_47602);
or UO_4639 (O_4639,N_46797,N_49952);
nor UO_4640 (O_4640,N_47737,N_48571);
nor UO_4641 (O_4641,N_46950,N_49114);
or UO_4642 (O_4642,N_49491,N_45233);
nand UO_4643 (O_4643,N_49839,N_49439);
and UO_4644 (O_4644,N_46643,N_49382);
nor UO_4645 (O_4645,N_46846,N_45926);
nand UO_4646 (O_4646,N_45496,N_46097);
and UO_4647 (O_4647,N_45649,N_45986);
nand UO_4648 (O_4648,N_48194,N_45428);
xor UO_4649 (O_4649,N_49963,N_48342);
or UO_4650 (O_4650,N_47757,N_47107);
nor UO_4651 (O_4651,N_46427,N_48613);
xor UO_4652 (O_4652,N_46457,N_49331);
xnor UO_4653 (O_4653,N_47238,N_49600);
nand UO_4654 (O_4654,N_47371,N_47663);
or UO_4655 (O_4655,N_45599,N_46976);
or UO_4656 (O_4656,N_46655,N_48197);
or UO_4657 (O_4657,N_45854,N_47899);
nor UO_4658 (O_4658,N_49962,N_49162);
or UO_4659 (O_4659,N_48969,N_49717);
and UO_4660 (O_4660,N_47812,N_46353);
or UO_4661 (O_4661,N_47442,N_45886);
nor UO_4662 (O_4662,N_49944,N_45751);
xnor UO_4663 (O_4663,N_48325,N_45309);
and UO_4664 (O_4664,N_48578,N_45767);
xnor UO_4665 (O_4665,N_47662,N_46386);
nor UO_4666 (O_4666,N_49794,N_46134);
xnor UO_4667 (O_4667,N_49197,N_48985);
and UO_4668 (O_4668,N_46886,N_46744);
nor UO_4669 (O_4669,N_49667,N_45058);
and UO_4670 (O_4670,N_46168,N_46290);
and UO_4671 (O_4671,N_45585,N_46696);
and UO_4672 (O_4672,N_49246,N_49836);
or UO_4673 (O_4673,N_49379,N_45568);
nand UO_4674 (O_4674,N_49428,N_46320);
and UO_4675 (O_4675,N_47132,N_45514);
xnor UO_4676 (O_4676,N_49655,N_48032);
nor UO_4677 (O_4677,N_45263,N_45402);
and UO_4678 (O_4678,N_47904,N_48902);
nor UO_4679 (O_4679,N_49646,N_45885);
and UO_4680 (O_4680,N_49485,N_49272);
nor UO_4681 (O_4681,N_46324,N_48517);
nor UO_4682 (O_4682,N_48512,N_47152);
nor UO_4683 (O_4683,N_48022,N_48657);
and UO_4684 (O_4684,N_46702,N_47418);
and UO_4685 (O_4685,N_49170,N_48232);
or UO_4686 (O_4686,N_45276,N_48945);
xnor UO_4687 (O_4687,N_48150,N_46314);
or UO_4688 (O_4688,N_48675,N_47849);
and UO_4689 (O_4689,N_45635,N_47011);
xnor UO_4690 (O_4690,N_46607,N_46374);
nor UO_4691 (O_4691,N_49015,N_48163);
nand UO_4692 (O_4692,N_49617,N_47496);
or UO_4693 (O_4693,N_46073,N_46049);
and UO_4694 (O_4694,N_46250,N_49222);
nand UO_4695 (O_4695,N_49082,N_45707);
or UO_4696 (O_4696,N_46143,N_49507);
nand UO_4697 (O_4697,N_45420,N_45729);
nand UO_4698 (O_4698,N_46319,N_49789);
xor UO_4699 (O_4699,N_46064,N_45352);
xnor UO_4700 (O_4700,N_49417,N_49525);
or UO_4701 (O_4701,N_49958,N_46715);
xnor UO_4702 (O_4702,N_47079,N_46554);
xnor UO_4703 (O_4703,N_49044,N_49739);
xnor UO_4704 (O_4704,N_45503,N_45479);
or UO_4705 (O_4705,N_49336,N_45994);
or UO_4706 (O_4706,N_48676,N_46448);
or UO_4707 (O_4707,N_49387,N_49674);
nand UO_4708 (O_4708,N_48126,N_45255);
nand UO_4709 (O_4709,N_49535,N_45089);
or UO_4710 (O_4710,N_49687,N_45567);
xor UO_4711 (O_4711,N_45246,N_46775);
and UO_4712 (O_4712,N_45492,N_48836);
nor UO_4713 (O_4713,N_47424,N_47266);
xnor UO_4714 (O_4714,N_47813,N_45217);
nor UO_4715 (O_4715,N_45916,N_46017);
or UO_4716 (O_4716,N_47678,N_45995);
nand UO_4717 (O_4717,N_46002,N_45538);
or UO_4718 (O_4718,N_49393,N_48537);
nand UO_4719 (O_4719,N_47829,N_45317);
or UO_4720 (O_4720,N_46572,N_49902);
nor UO_4721 (O_4721,N_49339,N_49345);
xor UO_4722 (O_4722,N_49145,N_48220);
nor UO_4723 (O_4723,N_49623,N_48869);
nand UO_4724 (O_4724,N_45636,N_48246);
nor UO_4725 (O_4725,N_45713,N_49842);
and UO_4726 (O_4726,N_47044,N_48840);
nand UO_4727 (O_4727,N_46449,N_48996);
nor UO_4728 (O_4728,N_49729,N_45395);
and UO_4729 (O_4729,N_46946,N_46268);
xor UO_4730 (O_4730,N_45443,N_46203);
or UO_4731 (O_4731,N_45107,N_48944);
nor UO_4732 (O_4732,N_45129,N_46409);
xor UO_4733 (O_4733,N_47619,N_45362);
and UO_4734 (O_4734,N_46593,N_49485);
and UO_4735 (O_4735,N_47230,N_49079);
nand UO_4736 (O_4736,N_45414,N_46532);
nand UO_4737 (O_4737,N_46626,N_46201);
nand UO_4738 (O_4738,N_46091,N_45227);
or UO_4739 (O_4739,N_46853,N_48616);
nand UO_4740 (O_4740,N_46871,N_45317);
xnor UO_4741 (O_4741,N_45102,N_46586);
xor UO_4742 (O_4742,N_45108,N_47114);
and UO_4743 (O_4743,N_48416,N_46811);
and UO_4744 (O_4744,N_47435,N_48103);
xor UO_4745 (O_4745,N_47163,N_48158);
nand UO_4746 (O_4746,N_48654,N_45582);
nor UO_4747 (O_4747,N_49022,N_45693);
nor UO_4748 (O_4748,N_46673,N_48833);
xor UO_4749 (O_4749,N_48311,N_45694);
nand UO_4750 (O_4750,N_45290,N_45395);
or UO_4751 (O_4751,N_45035,N_49407);
nand UO_4752 (O_4752,N_48403,N_47317);
xor UO_4753 (O_4753,N_49352,N_45406);
or UO_4754 (O_4754,N_49372,N_45798);
nor UO_4755 (O_4755,N_49452,N_46220);
nor UO_4756 (O_4756,N_48471,N_48076);
and UO_4757 (O_4757,N_47140,N_48820);
xor UO_4758 (O_4758,N_48667,N_45503);
xnor UO_4759 (O_4759,N_45310,N_46161);
xnor UO_4760 (O_4760,N_45011,N_48695);
nor UO_4761 (O_4761,N_46567,N_48203);
xnor UO_4762 (O_4762,N_46124,N_46096);
or UO_4763 (O_4763,N_45925,N_46072);
xor UO_4764 (O_4764,N_49619,N_48756);
xnor UO_4765 (O_4765,N_48550,N_48677);
nand UO_4766 (O_4766,N_46936,N_47676);
nor UO_4767 (O_4767,N_49014,N_46643);
or UO_4768 (O_4768,N_48266,N_46375);
or UO_4769 (O_4769,N_45164,N_47944);
or UO_4770 (O_4770,N_45922,N_48729);
or UO_4771 (O_4771,N_47392,N_46244);
nand UO_4772 (O_4772,N_45893,N_46049);
nor UO_4773 (O_4773,N_47304,N_47843);
nor UO_4774 (O_4774,N_47767,N_45206);
or UO_4775 (O_4775,N_45800,N_49917);
xnor UO_4776 (O_4776,N_46149,N_49646);
or UO_4777 (O_4777,N_48807,N_48873);
and UO_4778 (O_4778,N_46342,N_45714);
or UO_4779 (O_4779,N_46967,N_46213);
xor UO_4780 (O_4780,N_46401,N_46742);
nor UO_4781 (O_4781,N_47374,N_47115);
nand UO_4782 (O_4782,N_49289,N_45126);
nand UO_4783 (O_4783,N_47747,N_47689);
and UO_4784 (O_4784,N_47140,N_48731);
and UO_4785 (O_4785,N_46000,N_47599);
nor UO_4786 (O_4786,N_49181,N_45090);
or UO_4787 (O_4787,N_46171,N_48644);
xnor UO_4788 (O_4788,N_46378,N_46466);
and UO_4789 (O_4789,N_47487,N_48416);
or UO_4790 (O_4790,N_45906,N_46996);
nor UO_4791 (O_4791,N_49707,N_46494);
or UO_4792 (O_4792,N_46800,N_46534);
or UO_4793 (O_4793,N_48418,N_45903);
or UO_4794 (O_4794,N_45896,N_45652);
nor UO_4795 (O_4795,N_49100,N_45053);
nand UO_4796 (O_4796,N_49927,N_49326);
nor UO_4797 (O_4797,N_48485,N_45892);
and UO_4798 (O_4798,N_47835,N_45143);
nand UO_4799 (O_4799,N_46549,N_48538);
xor UO_4800 (O_4800,N_46227,N_49452);
or UO_4801 (O_4801,N_46796,N_46497);
nor UO_4802 (O_4802,N_45678,N_47191);
or UO_4803 (O_4803,N_47897,N_45637);
or UO_4804 (O_4804,N_48847,N_48810);
nand UO_4805 (O_4805,N_45148,N_48259);
nor UO_4806 (O_4806,N_45213,N_45591);
or UO_4807 (O_4807,N_45787,N_48101);
and UO_4808 (O_4808,N_49278,N_47014);
xor UO_4809 (O_4809,N_49690,N_45024);
xor UO_4810 (O_4810,N_48074,N_49870);
xor UO_4811 (O_4811,N_49017,N_48109);
nand UO_4812 (O_4812,N_48117,N_47094);
xnor UO_4813 (O_4813,N_47395,N_48119);
xor UO_4814 (O_4814,N_49421,N_48137);
and UO_4815 (O_4815,N_46990,N_46424);
and UO_4816 (O_4816,N_46389,N_46870);
xor UO_4817 (O_4817,N_48271,N_45776);
and UO_4818 (O_4818,N_48746,N_46038);
nor UO_4819 (O_4819,N_49801,N_47317);
nand UO_4820 (O_4820,N_46548,N_45970);
and UO_4821 (O_4821,N_45708,N_47724);
xnor UO_4822 (O_4822,N_47134,N_45828);
nand UO_4823 (O_4823,N_47450,N_47955);
xor UO_4824 (O_4824,N_49153,N_45728);
or UO_4825 (O_4825,N_46726,N_48847);
nor UO_4826 (O_4826,N_49915,N_48939);
and UO_4827 (O_4827,N_49519,N_47268);
or UO_4828 (O_4828,N_48168,N_48245);
or UO_4829 (O_4829,N_46087,N_49078);
nor UO_4830 (O_4830,N_49322,N_45662);
nand UO_4831 (O_4831,N_48349,N_46874);
and UO_4832 (O_4832,N_47260,N_48812);
nand UO_4833 (O_4833,N_45565,N_45100);
or UO_4834 (O_4834,N_45971,N_46369);
and UO_4835 (O_4835,N_48238,N_49387);
xnor UO_4836 (O_4836,N_48188,N_45432);
or UO_4837 (O_4837,N_45245,N_46962);
or UO_4838 (O_4838,N_45459,N_48582);
or UO_4839 (O_4839,N_49494,N_47800);
nand UO_4840 (O_4840,N_47147,N_46935);
or UO_4841 (O_4841,N_48273,N_49595);
or UO_4842 (O_4842,N_45586,N_49026);
and UO_4843 (O_4843,N_45029,N_49889);
xnor UO_4844 (O_4844,N_49606,N_49741);
nand UO_4845 (O_4845,N_46751,N_46240);
and UO_4846 (O_4846,N_45217,N_45553);
xor UO_4847 (O_4847,N_46259,N_49644);
or UO_4848 (O_4848,N_49757,N_49432);
nand UO_4849 (O_4849,N_48094,N_45600);
nand UO_4850 (O_4850,N_45133,N_47772);
xnor UO_4851 (O_4851,N_46130,N_45847);
and UO_4852 (O_4852,N_47613,N_49004);
nand UO_4853 (O_4853,N_49448,N_49281);
or UO_4854 (O_4854,N_47003,N_49750);
nand UO_4855 (O_4855,N_49597,N_49149);
xor UO_4856 (O_4856,N_45905,N_48713);
and UO_4857 (O_4857,N_48130,N_48878);
xor UO_4858 (O_4858,N_47487,N_45645);
or UO_4859 (O_4859,N_45025,N_47488);
xnor UO_4860 (O_4860,N_45061,N_45262);
nand UO_4861 (O_4861,N_47937,N_48412);
xnor UO_4862 (O_4862,N_45579,N_48726);
nor UO_4863 (O_4863,N_47278,N_45065);
nor UO_4864 (O_4864,N_46733,N_48849);
nand UO_4865 (O_4865,N_49901,N_47106);
xor UO_4866 (O_4866,N_49752,N_47593);
nor UO_4867 (O_4867,N_47680,N_47080);
xor UO_4868 (O_4868,N_48655,N_46218);
or UO_4869 (O_4869,N_45467,N_48938);
nand UO_4870 (O_4870,N_45394,N_46900);
or UO_4871 (O_4871,N_48811,N_45174);
or UO_4872 (O_4872,N_45094,N_48135);
or UO_4873 (O_4873,N_49751,N_49060);
nand UO_4874 (O_4874,N_48829,N_47251);
nand UO_4875 (O_4875,N_46343,N_47011);
or UO_4876 (O_4876,N_49966,N_48166);
nor UO_4877 (O_4877,N_45614,N_48886);
nor UO_4878 (O_4878,N_49070,N_45570);
or UO_4879 (O_4879,N_48709,N_45039);
and UO_4880 (O_4880,N_48957,N_48749);
nand UO_4881 (O_4881,N_49551,N_45311);
xnor UO_4882 (O_4882,N_49093,N_46610);
nand UO_4883 (O_4883,N_48899,N_47532);
nor UO_4884 (O_4884,N_46622,N_49035);
xnor UO_4885 (O_4885,N_47977,N_45925);
nand UO_4886 (O_4886,N_45263,N_47171);
xor UO_4887 (O_4887,N_45016,N_46862);
and UO_4888 (O_4888,N_46378,N_47803);
or UO_4889 (O_4889,N_48721,N_49533);
nor UO_4890 (O_4890,N_49067,N_48474);
nand UO_4891 (O_4891,N_46350,N_49755);
xnor UO_4892 (O_4892,N_48873,N_48944);
nor UO_4893 (O_4893,N_47946,N_45827);
nor UO_4894 (O_4894,N_49898,N_48159);
or UO_4895 (O_4895,N_49476,N_46130);
or UO_4896 (O_4896,N_47154,N_45310);
and UO_4897 (O_4897,N_47970,N_49429);
and UO_4898 (O_4898,N_47505,N_48032);
or UO_4899 (O_4899,N_47897,N_47944);
nand UO_4900 (O_4900,N_46249,N_46699);
xnor UO_4901 (O_4901,N_46397,N_47357);
or UO_4902 (O_4902,N_49330,N_45634);
and UO_4903 (O_4903,N_46747,N_49141);
and UO_4904 (O_4904,N_48685,N_48329);
nand UO_4905 (O_4905,N_45680,N_47019);
xnor UO_4906 (O_4906,N_49063,N_48381);
nor UO_4907 (O_4907,N_46820,N_46473);
and UO_4908 (O_4908,N_49163,N_47845);
or UO_4909 (O_4909,N_49157,N_45488);
and UO_4910 (O_4910,N_46266,N_46627);
nand UO_4911 (O_4911,N_47390,N_47954);
or UO_4912 (O_4912,N_46782,N_47949);
or UO_4913 (O_4913,N_49828,N_46252);
xor UO_4914 (O_4914,N_49680,N_49068);
or UO_4915 (O_4915,N_49094,N_48294);
xor UO_4916 (O_4916,N_49595,N_47684);
or UO_4917 (O_4917,N_45365,N_47824);
or UO_4918 (O_4918,N_46105,N_45062);
or UO_4919 (O_4919,N_48112,N_47567);
nand UO_4920 (O_4920,N_48726,N_47088);
or UO_4921 (O_4921,N_45617,N_46859);
xor UO_4922 (O_4922,N_45351,N_47861);
nand UO_4923 (O_4923,N_48869,N_48573);
xnor UO_4924 (O_4924,N_45286,N_46121);
nor UO_4925 (O_4925,N_47742,N_49403);
or UO_4926 (O_4926,N_48175,N_48974);
nor UO_4927 (O_4927,N_46773,N_45056);
and UO_4928 (O_4928,N_46626,N_45388);
or UO_4929 (O_4929,N_46696,N_48221);
or UO_4930 (O_4930,N_46982,N_46100);
nor UO_4931 (O_4931,N_48952,N_49030);
xor UO_4932 (O_4932,N_45128,N_46336);
nor UO_4933 (O_4933,N_45110,N_48801);
nand UO_4934 (O_4934,N_48998,N_49325);
xor UO_4935 (O_4935,N_48851,N_46648);
nand UO_4936 (O_4936,N_49037,N_45023);
xor UO_4937 (O_4937,N_47443,N_48900);
nor UO_4938 (O_4938,N_47474,N_45837);
or UO_4939 (O_4939,N_47684,N_47929);
xnor UO_4940 (O_4940,N_48164,N_46054);
nor UO_4941 (O_4941,N_46259,N_48726);
and UO_4942 (O_4942,N_45182,N_49699);
and UO_4943 (O_4943,N_46977,N_48325);
nand UO_4944 (O_4944,N_48181,N_45541);
and UO_4945 (O_4945,N_45439,N_45795);
xor UO_4946 (O_4946,N_46805,N_49134);
nand UO_4947 (O_4947,N_49359,N_49178);
or UO_4948 (O_4948,N_49082,N_47773);
or UO_4949 (O_4949,N_49123,N_46969);
nand UO_4950 (O_4950,N_48917,N_45145);
or UO_4951 (O_4951,N_45902,N_47854);
and UO_4952 (O_4952,N_47805,N_46917);
and UO_4953 (O_4953,N_47285,N_47645);
or UO_4954 (O_4954,N_45267,N_45027);
nand UO_4955 (O_4955,N_49948,N_48313);
and UO_4956 (O_4956,N_49127,N_47922);
xor UO_4957 (O_4957,N_45939,N_45797);
nor UO_4958 (O_4958,N_47580,N_45369);
nand UO_4959 (O_4959,N_47200,N_48782);
nor UO_4960 (O_4960,N_46328,N_49544);
xor UO_4961 (O_4961,N_49914,N_49671);
or UO_4962 (O_4962,N_47582,N_47541);
nor UO_4963 (O_4963,N_46216,N_46990);
nor UO_4964 (O_4964,N_47290,N_48259);
nor UO_4965 (O_4965,N_47602,N_46114);
and UO_4966 (O_4966,N_45115,N_49087);
nand UO_4967 (O_4967,N_45345,N_45402);
and UO_4968 (O_4968,N_45141,N_46887);
or UO_4969 (O_4969,N_45925,N_45006);
and UO_4970 (O_4970,N_46132,N_46323);
xnor UO_4971 (O_4971,N_48994,N_48467);
nand UO_4972 (O_4972,N_46783,N_48338);
xnor UO_4973 (O_4973,N_49933,N_48672);
or UO_4974 (O_4974,N_48678,N_49716);
and UO_4975 (O_4975,N_49090,N_46743);
or UO_4976 (O_4976,N_48826,N_47300);
nand UO_4977 (O_4977,N_46684,N_47229);
nor UO_4978 (O_4978,N_49911,N_46532);
xnor UO_4979 (O_4979,N_46709,N_47473);
nor UO_4980 (O_4980,N_48319,N_49098);
xor UO_4981 (O_4981,N_48054,N_48703);
or UO_4982 (O_4982,N_45055,N_48377);
nand UO_4983 (O_4983,N_46078,N_48231);
or UO_4984 (O_4984,N_45103,N_49917);
xnor UO_4985 (O_4985,N_47983,N_45510);
and UO_4986 (O_4986,N_49547,N_49200);
or UO_4987 (O_4987,N_47191,N_46706);
or UO_4988 (O_4988,N_47369,N_45221);
xor UO_4989 (O_4989,N_46803,N_45746);
xor UO_4990 (O_4990,N_47255,N_46058);
xor UO_4991 (O_4991,N_46260,N_49309);
xor UO_4992 (O_4992,N_49845,N_49095);
and UO_4993 (O_4993,N_48878,N_48186);
nor UO_4994 (O_4994,N_46329,N_47189);
nand UO_4995 (O_4995,N_45156,N_47137);
and UO_4996 (O_4996,N_47932,N_46592);
or UO_4997 (O_4997,N_49740,N_45124);
xor UO_4998 (O_4998,N_46355,N_49505);
xnor UO_4999 (O_4999,N_48467,N_48937);
endmodule