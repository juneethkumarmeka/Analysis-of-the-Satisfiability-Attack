module basic_500_3000_500_50_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_343,In_243);
or U1 (N_1,In_380,In_13);
nor U2 (N_2,In_262,In_184);
and U3 (N_3,In_374,In_132);
and U4 (N_4,In_62,In_319);
nand U5 (N_5,In_362,In_269);
or U6 (N_6,In_457,In_142);
nand U7 (N_7,In_229,In_417);
and U8 (N_8,In_321,In_8);
nor U9 (N_9,In_30,In_279);
nand U10 (N_10,In_353,In_146);
nor U11 (N_11,In_356,In_10);
nor U12 (N_12,In_18,In_348);
nor U13 (N_13,In_139,In_340);
and U14 (N_14,In_401,In_33);
nor U15 (N_15,In_301,In_94);
xor U16 (N_16,In_28,In_241);
and U17 (N_17,In_67,In_347);
nor U18 (N_18,In_332,In_434);
and U19 (N_19,In_224,In_100);
nor U20 (N_20,In_267,In_22);
or U21 (N_21,In_496,In_144);
nand U22 (N_22,In_64,In_75);
or U23 (N_23,In_447,In_494);
or U24 (N_24,In_1,In_44);
nand U25 (N_25,In_463,In_412);
or U26 (N_26,In_225,In_15);
or U27 (N_27,In_237,In_289);
nor U28 (N_28,In_394,In_349);
nor U29 (N_29,In_242,In_85);
xnor U30 (N_30,In_248,In_69);
nor U31 (N_31,In_315,In_440);
nand U32 (N_32,In_140,In_57);
nor U33 (N_33,In_247,In_71);
nor U34 (N_34,In_82,In_129);
or U35 (N_35,In_35,In_369);
or U36 (N_36,In_125,In_351);
nor U37 (N_37,In_192,In_120);
and U38 (N_38,In_367,In_209);
and U39 (N_39,In_395,In_421);
and U40 (N_40,In_471,In_212);
and U41 (N_41,In_83,In_190);
or U42 (N_42,In_154,In_105);
or U43 (N_43,In_24,In_424);
nand U44 (N_44,In_177,In_450);
or U45 (N_45,In_387,In_404);
or U46 (N_46,In_406,In_264);
nand U47 (N_47,In_66,In_413);
and U48 (N_48,In_26,In_165);
nor U49 (N_49,In_381,In_271);
xnor U50 (N_50,In_290,In_300);
nor U51 (N_51,In_286,In_98);
nor U52 (N_52,In_377,In_163);
and U53 (N_53,In_388,In_200);
and U54 (N_54,In_27,In_160);
and U55 (N_55,In_275,In_400);
or U56 (N_56,In_446,In_256);
nand U57 (N_57,In_164,In_432);
nor U58 (N_58,In_152,In_458);
and U59 (N_59,In_95,In_442);
nor U60 (N_60,In_285,In_341);
or U61 (N_61,In_390,In_73);
or U62 (N_62,In_255,In_115);
or U63 (N_63,In_123,N_21);
or U64 (N_64,N_33,In_488);
or U65 (N_65,N_10,In_182);
nor U66 (N_66,In_304,In_445);
and U67 (N_67,In_203,In_430);
or U68 (N_68,N_18,In_183);
nor U69 (N_69,In_202,In_478);
nor U70 (N_70,In_408,In_378);
and U71 (N_71,In_309,In_364);
or U72 (N_72,In_342,In_169);
and U73 (N_73,In_52,N_56);
nand U74 (N_74,In_86,In_119);
nand U75 (N_75,In_368,In_195);
nand U76 (N_76,N_7,In_17);
and U77 (N_77,In_174,In_19);
and U78 (N_78,In_330,In_466);
nor U79 (N_79,In_234,In_138);
nor U80 (N_80,In_205,N_57);
and U81 (N_81,In_425,N_29);
or U82 (N_82,In_124,In_423);
nand U83 (N_83,In_477,In_467);
and U84 (N_84,In_4,In_322);
nand U85 (N_85,In_436,In_312);
nor U86 (N_86,In_37,In_486);
nand U87 (N_87,In_7,In_5);
nand U88 (N_88,In_439,In_173);
and U89 (N_89,In_136,In_253);
nand U90 (N_90,In_396,N_19);
and U91 (N_91,In_270,In_431);
nor U92 (N_92,In_150,In_335);
nor U93 (N_93,In_110,In_426);
nor U94 (N_94,N_4,N_38);
or U95 (N_95,In_462,In_298);
and U96 (N_96,In_282,In_272);
and U97 (N_97,In_51,In_371);
nand U98 (N_98,In_422,In_379);
and U99 (N_99,In_61,N_44);
nand U100 (N_100,In_295,In_53);
or U101 (N_101,In_366,In_46);
nand U102 (N_102,In_460,In_157);
and U103 (N_103,In_280,In_42);
nand U104 (N_104,In_102,In_104);
or U105 (N_105,In_25,In_170);
or U106 (N_106,In_187,In_38);
nor U107 (N_107,N_49,N_39);
and U108 (N_108,In_411,N_17);
nand U109 (N_109,In_418,N_16);
and U110 (N_110,In_331,In_178);
and U111 (N_111,In_313,In_435);
and U112 (N_112,In_360,In_108);
nor U113 (N_113,In_88,N_12);
or U114 (N_114,In_16,In_148);
nand U115 (N_115,N_8,In_161);
nor U116 (N_116,In_84,In_410);
xor U117 (N_117,In_245,In_441);
or U118 (N_118,In_97,N_55);
or U119 (N_119,In_481,N_15);
and U120 (N_120,In_333,N_63);
nand U121 (N_121,In_68,In_427);
nand U122 (N_122,N_92,In_128);
and U123 (N_123,N_109,In_48);
and U124 (N_124,N_94,In_45);
nor U125 (N_125,In_11,In_116);
or U126 (N_126,In_327,In_236);
nand U127 (N_127,In_420,In_111);
nor U128 (N_128,N_118,In_409);
and U129 (N_129,In_240,In_386);
nand U130 (N_130,N_74,In_393);
nand U131 (N_131,N_28,In_199);
nand U132 (N_132,In_489,In_249);
and U133 (N_133,N_27,In_59);
and U134 (N_134,In_109,N_45);
nand U135 (N_135,N_34,N_52);
or U136 (N_136,In_106,N_96);
nand U137 (N_137,In_311,In_172);
and U138 (N_138,N_3,In_168);
and U139 (N_139,N_51,In_107);
nand U140 (N_140,In_399,N_5);
nand U141 (N_141,In_112,In_323);
nor U142 (N_142,N_59,In_383);
nor U143 (N_143,In_235,In_126);
xnor U144 (N_144,N_11,In_118);
nand U145 (N_145,In_363,In_252);
nor U146 (N_146,In_0,In_87);
nor U147 (N_147,In_449,In_493);
nand U148 (N_148,In_357,In_238);
nand U149 (N_149,N_107,N_85);
nor U150 (N_150,N_106,N_81);
and U151 (N_151,In_302,In_14);
and U152 (N_152,In_263,In_92);
and U153 (N_153,In_254,N_20);
or U154 (N_154,N_91,In_96);
xnor U155 (N_155,In_151,In_438);
nand U156 (N_156,In_257,In_491);
nand U157 (N_157,N_90,In_207);
or U158 (N_158,N_95,N_77);
xor U159 (N_159,In_281,In_41);
nand U160 (N_160,In_153,In_284);
and U161 (N_161,N_0,N_64);
or U162 (N_162,In_188,In_149);
nand U163 (N_163,N_62,In_218);
nand U164 (N_164,In_419,In_29);
and U165 (N_165,In_305,In_266);
or U166 (N_166,In_158,In_497);
nand U167 (N_167,In_310,N_35);
nand U168 (N_168,In_358,In_317);
nor U169 (N_169,N_42,N_58);
nand U170 (N_170,In_337,In_78);
nand U171 (N_171,N_80,In_455);
nor U172 (N_172,N_53,In_359);
nor U173 (N_173,In_246,In_32);
nand U174 (N_174,In_402,In_495);
and U175 (N_175,In_288,In_346);
nor U176 (N_176,In_171,N_43);
nor U177 (N_177,In_329,N_114);
nand U178 (N_178,In_265,N_87);
or U179 (N_179,In_375,N_26);
nor U180 (N_180,N_140,N_160);
nand U181 (N_181,N_65,In_318);
nor U182 (N_182,N_89,N_2);
or U183 (N_183,N_124,In_297);
nor U184 (N_184,In_56,In_376);
nand U185 (N_185,In_370,In_197);
or U186 (N_186,N_79,N_165);
nand U187 (N_187,N_9,N_30);
or U188 (N_188,In_336,N_163);
or U189 (N_189,In_244,N_171);
and U190 (N_190,In_117,N_123);
and U191 (N_191,In_499,In_214);
nor U192 (N_192,In_372,In_415);
nor U193 (N_193,N_76,In_216);
nand U194 (N_194,In_193,In_273);
nor U195 (N_195,In_23,N_61);
nor U196 (N_196,N_69,In_208);
or U197 (N_197,In_155,N_37);
nor U198 (N_198,In_480,N_40);
or U199 (N_199,N_120,In_47);
or U200 (N_200,In_429,In_326);
nand U201 (N_201,In_222,In_454);
or U202 (N_202,In_277,N_88);
and U203 (N_203,In_227,In_80);
nand U204 (N_204,N_46,N_100);
xor U205 (N_205,N_175,N_130);
or U206 (N_206,N_23,In_484);
or U207 (N_207,In_451,N_116);
and U208 (N_208,In_444,In_191);
nor U209 (N_209,In_143,In_127);
nand U210 (N_210,In_186,In_159);
or U211 (N_211,N_177,In_476);
or U212 (N_212,N_99,In_475);
nand U213 (N_213,In_292,In_81);
or U214 (N_214,In_226,N_155);
or U215 (N_215,In_461,In_40);
nand U216 (N_216,In_328,In_93);
and U217 (N_217,In_65,In_141);
nand U218 (N_218,In_433,In_6);
nand U219 (N_219,N_179,N_66);
and U220 (N_220,In_403,N_146);
nor U221 (N_221,In_354,In_180);
nor U222 (N_222,In_479,N_131);
or U223 (N_223,In_334,N_122);
nor U224 (N_224,In_391,In_70);
or U225 (N_225,N_167,N_138);
or U226 (N_226,N_1,In_36);
nand U227 (N_227,In_268,In_133);
nor U228 (N_228,N_141,In_147);
nor U229 (N_229,N_152,N_108);
xnor U230 (N_230,N_31,In_459);
nand U231 (N_231,In_99,N_166);
nand U232 (N_232,In_181,In_355);
nand U233 (N_233,In_145,In_261);
and U234 (N_234,In_350,N_73);
and U235 (N_235,N_143,N_119);
nand U236 (N_236,In_464,N_148);
nor U237 (N_237,In_465,In_55);
nor U238 (N_238,In_338,In_131);
nand U239 (N_239,In_316,In_122);
nand U240 (N_240,N_178,In_114);
nand U241 (N_241,N_224,In_325);
xor U242 (N_242,N_211,N_129);
and U243 (N_243,In_274,In_175);
or U244 (N_244,N_68,In_239);
nor U245 (N_245,In_58,In_384);
nand U246 (N_246,N_67,In_217);
nor U247 (N_247,In_306,N_223);
and U248 (N_248,N_149,In_228);
or U249 (N_249,In_223,N_207);
nand U250 (N_250,In_3,In_89);
and U251 (N_251,In_179,In_166);
or U252 (N_252,In_130,N_101);
or U253 (N_253,N_137,N_125);
or U254 (N_254,N_13,N_219);
and U255 (N_255,N_220,N_72);
or U256 (N_256,In_452,In_2);
and U257 (N_257,N_172,In_385);
or U258 (N_258,In_54,N_198);
or U259 (N_259,In_314,In_20);
and U260 (N_260,N_194,In_291);
nor U261 (N_261,N_126,In_198);
nand U262 (N_262,N_230,N_221);
or U263 (N_263,In_470,In_185);
nor U264 (N_264,N_159,N_164);
nor U265 (N_265,N_193,N_217);
nand U266 (N_266,N_151,N_113);
or U267 (N_267,N_98,N_112);
nand U268 (N_268,N_234,In_414);
or U269 (N_269,N_84,In_162);
nor U270 (N_270,N_227,In_221);
nand U271 (N_271,N_229,In_382);
or U272 (N_272,N_176,In_294);
nand U273 (N_273,In_448,N_218);
nand U274 (N_274,N_182,N_204);
and U275 (N_275,N_97,N_190);
and U276 (N_276,In_39,In_456);
or U277 (N_277,In_296,In_72);
nor U278 (N_278,N_83,N_169);
nor U279 (N_279,In_437,In_219);
nand U280 (N_280,N_54,N_201);
nand U281 (N_281,In_90,In_474);
or U282 (N_282,In_492,N_36);
nand U283 (N_283,In_34,In_339);
and U284 (N_284,N_213,N_226);
and U285 (N_285,In_259,In_283);
nor U286 (N_286,N_41,In_134);
or U287 (N_287,N_233,N_188);
nor U288 (N_288,In_12,N_191);
or U289 (N_289,In_156,In_487);
nor U290 (N_290,N_215,In_91);
or U291 (N_291,In_103,N_174);
nand U292 (N_292,N_104,N_212);
nand U293 (N_293,In_230,In_9);
or U294 (N_294,In_76,N_181);
nand U295 (N_295,In_63,In_49);
xnor U296 (N_296,In_324,In_398);
nor U297 (N_297,In_260,In_167);
nand U298 (N_298,N_110,N_22);
nand U299 (N_299,In_50,N_153);
nand U300 (N_300,N_267,In_201);
and U301 (N_301,N_78,N_214);
nor U302 (N_302,In_21,N_293);
or U303 (N_303,N_195,In_79);
and U304 (N_304,N_144,N_197);
and U305 (N_305,N_298,N_295);
nor U306 (N_306,N_134,N_186);
and U307 (N_307,N_161,N_286);
nand U308 (N_308,In_345,N_262);
and U309 (N_309,N_278,N_290);
nand U310 (N_310,N_71,N_6);
nor U311 (N_311,N_285,In_233);
nor U312 (N_312,In_250,N_277);
xor U313 (N_313,N_264,N_238);
nor U314 (N_314,N_292,N_157);
nand U315 (N_315,In_308,In_352);
nand U316 (N_316,N_206,N_82);
and U317 (N_317,In_60,N_75);
nand U318 (N_318,In_498,N_135);
nor U319 (N_319,In_189,In_344);
or U320 (N_320,N_273,N_192);
nand U321 (N_321,In_407,N_139);
nand U322 (N_322,N_252,N_14);
nand U323 (N_323,N_24,In_392);
and U324 (N_324,N_265,N_200);
and U325 (N_325,N_296,N_136);
and U326 (N_326,N_283,N_111);
nand U327 (N_327,N_173,N_25);
or U328 (N_328,N_271,N_121);
nand U329 (N_329,N_168,In_373);
or U330 (N_330,N_103,N_102);
nor U331 (N_331,In_258,In_31);
or U332 (N_332,N_47,N_269);
nand U333 (N_333,N_245,N_258);
and U334 (N_334,N_261,N_281);
or U335 (N_335,N_239,N_115);
or U336 (N_336,In_472,N_133);
nand U337 (N_337,N_196,N_127);
nor U338 (N_338,N_259,N_249);
and U339 (N_339,N_170,In_428);
or U340 (N_340,N_232,In_135);
or U341 (N_341,In_210,N_70);
and U342 (N_342,In_278,N_244);
and U343 (N_343,In_137,In_77);
nand U344 (N_344,N_142,N_253);
and U345 (N_345,In_361,N_299);
nand U346 (N_346,N_86,In_485);
or U347 (N_347,In_113,In_405);
nand U348 (N_348,In_299,In_397);
or U349 (N_349,N_251,In_121);
nor U350 (N_350,N_246,In_206);
or U351 (N_351,N_50,In_211);
nor U352 (N_352,N_272,N_93);
nor U353 (N_353,N_257,N_154);
or U354 (N_354,N_202,In_482);
nor U355 (N_355,In_176,In_473);
and U356 (N_356,In_232,N_240);
and U357 (N_357,N_270,In_416);
and U358 (N_358,In_453,N_189);
and U359 (N_359,In_196,In_443);
nand U360 (N_360,N_248,N_336);
or U361 (N_361,N_305,In_215);
and U362 (N_362,N_289,N_355);
nor U363 (N_363,N_294,N_250);
nand U364 (N_364,N_288,N_158);
nand U365 (N_365,N_353,N_222);
and U366 (N_366,In_276,N_274);
nor U367 (N_367,In_389,N_242);
nor U368 (N_368,In_101,N_310);
and U369 (N_369,N_335,In_307);
nor U370 (N_370,N_333,N_337);
or U371 (N_371,N_128,N_302);
or U372 (N_372,N_216,N_260);
or U373 (N_373,N_352,In_365);
and U374 (N_374,N_325,N_280);
nor U375 (N_375,N_328,N_60);
and U376 (N_376,N_275,N_351);
and U377 (N_377,N_301,N_330);
nor U378 (N_378,N_350,N_237);
and U379 (N_379,N_48,N_236);
and U380 (N_380,N_318,N_340);
nand U381 (N_381,N_324,N_331);
or U382 (N_382,N_334,In_320);
nor U383 (N_383,In_231,N_346);
nor U384 (N_384,N_311,N_282);
and U385 (N_385,N_156,In_287);
nand U386 (N_386,N_205,In_469);
nor U387 (N_387,N_147,N_326);
or U388 (N_388,In_483,In_194);
nor U389 (N_389,N_309,N_354);
or U390 (N_390,N_344,N_183);
nand U391 (N_391,N_210,N_150);
and U392 (N_392,N_279,N_341);
nor U393 (N_393,N_321,In_468);
nor U394 (N_394,N_185,N_268);
nand U395 (N_395,N_358,N_162);
nand U396 (N_396,N_348,In_213);
or U397 (N_397,N_357,In_303);
nand U398 (N_398,N_105,N_291);
or U399 (N_399,In_220,N_316);
and U400 (N_400,N_132,N_332);
or U401 (N_401,N_312,N_199);
or U402 (N_402,In_251,N_247);
nor U403 (N_403,N_208,N_225);
or U404 (N_404,N_319,N_209);
or U405 (N_405,N_349,N_359);
and U406 (N_406,N_329,In_293);
and U407 (N_407,N_117,N_254);
nor U408 (N_408,N_339,N_184);
nand U409 (N_409,N_356,N_180);
nor U410 (N_410,N_263,N_306);
and U411 (N_411,N_203,N_266);
or U412 (N_412,N_313,N_145);
nor U413 (N_413,N_297,In_204);
nand U414 (N_414,N_276,N_300);
and U415 (N_415,N_315,N_32);
or U416 (N_416,N_342,N_322);
nand U417 (N_417,N_228,N_255);
nor U418 (N_418,N_303,N_304);
nor U419 (N_419,N_343,N_307);
and U420 (N_420,N_394,N_241);
or U421 (N_421,N_404,N_320);
and U422 (N_422,N_410,N_243);
and U423 (N_423,N_380,N_395);
nand U424 (N_424,N_397,N_398);
or U425 (N_425,N_389,N_363);
nand U426 (N_426,N_338,N_408);
nand U427 (N_427,N_347,N_374);
or U428 (N_428,N_407,N_235);
or U429 (N_429,N_376,N_368);
and U430 (N_430,N_317,N_370);
and U431 (N_431,N_366,N_287);
or U432 (N_432,N_393,N_409);
or U433 (N_433,N_412,N_365);
and U434 (N_434,N_417,N_369);
or U435 (N_435,N_401,In_43);
nor U436 (N_436,N_411,N_345);
and U437 (N_437,N_381,N_378);
and U438 (N_438,N_323,N_327);
or U439 (N_439,N_364,N_403);
or U440 (N_440,N_387,N_388);
nand U441 (N_441,N_231,N_386);
nand U442 (N_442,N_390,N_383);
nand U443 (N_443,N_379,N_377);
nor U444 (N_444,N_413,N_362);
nor U445 (N_445,N_382,N_284);
nor U446 (N_446,N_399,N_187);
or U447 (N_447,N_406,In_74);
nor U448 (N_448,N_414,N_308);
nand U449 (N_449,N_416,N_402);
nor U450 (N_450,N_360,N_367);
nor U451 (N_451,N_385,N_415);
or U452 (N_452,N_375,N_405);
and U453 (N_453,N_384,N_391);
xnor U454 (N_454,N_256,N_400);
nor U455 (N_455,N_392,N_419);
nor U456 (N_456,N_314,N_396);
nor U457 (N_457,N_371,N_372);
and U458 (N_458,In_490,N_361);
nor U459 (N_459,N_418,N_373);
nand U460 (N_460,N_375,N_393);
or U461 (N_461,In_43,N_345);
and U462 (N_462,N_410,N_370);
nand U463 (N_463,N_383,N_361);
nor U464 (N_464,N_405,N_397);
nand U465 (N_465,N_397,N_287);
nand U466 (N_466,N_388,N_371);
nand U467 (N_467,N_385,N_317);
nand U468 (N_468,N_384,N_381);
nor U469 (N_469,N_327,N_361);
and U470 (N_470,N_383,N_347);
nor U471 (N_471,N_415,N_417);
nor U472 (N_472,N_366,N_368);
nor U473 (N_473,N_373,N_365);
or U474 (N_474,N_371,N_404);
and U475 (N_475,N_416,N_381);
nand U476 (N_476,N_376,N_414);
or U477 (N_477,N_400,N_347);
and U478 (N_478,N_409,N_401);
and U479 (N_479,N_362,N_368);
nand U480 (N_480,N_424,N_478);
nor U481 (N_481,N_433,N_451);
nor U482 (N_482,N_423,N_466);
nor U483 (N_483,N_438,N_459);
or U484 (N_484,N_461,N_469);
and U485 (N_485,N_426,N_452);
xor U486 (N_486,N_464,N_421);
or U487 (N_487,N_436,N_434);
or U488 (N_488,N_477,N_471);
nor U489 (N_489,N_457,N_425);
nand U490 (N_490,N_476,N_442);
nor U491 (N_491,N_474,N_462);
and U492 (N_492,N_427,N_467);
xor U493 (N_493,N_479,N_429);
or U494 (N_494,N_439,N_422);
and U495 (N_495,N_454,N_458);
nand U496 (N_496,N_473,N_441);
or U497 (N_497,N_443,N_465);
or U498 (N_498,N_437,N_440);
or U499 (N_499,N_463,N_428);
and U500 (N_500,N_450,N_430);
nor U501 (N_501,N_446,N_449);
xor U502 (N_502,N_468,N_453);
or U503 (N_503,N_447,N_472);
nor U504 (N_504,N_431,N_456);
and U505 (N_505,N_448,N_435);
and U506 (N_506,N_470,N_475);
xor U507 (N_507,N_444,N_455);
nor U508 (N_508,N_420,N_445);
and U509 (N_509,N_432,N_460);
and U510 (N_510,N_429,N_477);
or U511 (N_511,N_476,N_464);
nand U512 (N_512,N_462,N_431);
and U513 (N_513,N_457,N_431);
and U514 (N_514,N_460,N_424);
or U515 (N_515,N_426,N_433);
or U516 (N_516,N_427,N_435);
or U517 (N_517,N_478,N_451);
nor U518 (N_518,N_455,N_420);
or U519 (N_519,N_474,N_459);
and U520 (N_520,N_447,N_458);
and U521 (N_521,N_453,N_467);
nor U522 (N_522,N_473,N_422);
nand U523 (N_523,N_442,N_440);
nor U524 (N_524,N_434,N_459);
and U525 (N_525,N_471,N_427);
nor U526 (N_526,N_445,N_478);
nor U527 (N_527,N_473,N_435);
or U528 (N_528,N_479,N_445);
nor U529 (N_529,N_464,N_449);
nand U530 (N_530,N_471,N_428);
and U531 (N_531,N_477,N_444);
nand U532 (N_532,N_452,N_467);
nand U533 (N_533,N_421,N_447);
nand U534 (N_534,N_437,N_433);
or U535 (N_535,N_468,N_459);
and U536 (N_536,N_458,N_461);
or U537 (N_537,N_433,N_475);
or U538 (N_538,N_431,N_464);
or U539 (N_539,N_467,N_438);
or U540 (N_540,N_507,N_518);
and U541 (N_541,N_484,N_482);
and U542 (N_542,N_488,N_539);
nand U543 (N_543,N_516,N_521);
nor U544 (N_544,N_520,N_494);
nand U545 (N_545,N_490,N_514);
nor U546 (N_546,N_525,N_501);
nand U547 (N_547,N_503,N_505);
nand U548 (N_548,N_531,N_529);
nand U549 (N_549,N_530,N_495);
or U550 (N_550,N_536,N_496);
nor U551 (N_551,N_491,N_486);
nor U552 (N_552,N_526,N_533);
nor U553 (N_553,N_500,N_510);
and U554 (N_554,N_522,N_492);
nand U555 (N_555,N_535,N_538);
and U556 (N_556,N_537,N_480);
nor U557 (N_557,N_512,N_524);
nor U558 (N_558,N_497,N_489);
nand U559 (N_559,N_504,N_517);
and U560 (N_560,N_487,N_508);
nand U561 (N_561,N_532,N_523);
and U562 (N_562,N_499,N_498);
or U563 (N_563,N_481,N_485);
and U564 (N_564,N_493,N_506);
and U565 (N_565,N_511,N_534);
nor U566 (N_566,N_502,N_519);
and U567 (N_567,N_509,N_513);
or U568 (N_568,N_527,N_483);
nand U569 (N_569,N_515,N_528);
and U570 (N_570,N_503,N_533);
nand U571 (N_571,N_510,N_486);
and U572 (N_572,N_533,N_481);
nor U573 (N_573,N_484,N_500);
or U574 (N_574,N_510,N_509);
or U575 (N_575,N_526,N_480);
or U576 (N_576,N_532,N_521);
and U577 (N_577,N_528,N_485);
nand U578 (N_578,N_527,N_510);
and U579 (N_579,N_487,N_537);
or U580 (N_580,N_489,N_491);
and U581 (N_581,N_493,N_481);
or U582 (N_582,N_497,N_505);
and U583 (N_583,N_513,N_481);
and U584 (N_584,N_494,N_539);
nor U585 (N_585,N_495,N_481);
or U586 (N_586,N_518,N_537);
nor U587 (N_587,N_503,N_537);
and U588 (N_588,N_490,N_506);
nand U589 (N_589,N_534,N_514);
nand U590 (N_590,N_492,N_528);
and U591 (N_591,N_493,N_482);
and U592 (N_592,N_505,N_525);
or U593 (N_593,N_491,N_519);
nand U594 (N_594,N_491,N_528);
or U595 (N_595,N_485,N_508);
xnor U596 (N_596,N_482,N_507);
and U597 (N_597,N_519,N_513);
nor U598 (N_598,N_488,N_521);
nor U599 (N_599,N_530,N_482);
nand U600 (N_600,N_573,N_581);
and U601 (N_601,N_583,N_585);
nand U602 (N_602,N_556,N_580);
or U603 (N_603,N_560,N_592);
and U604 (N_604,N_582,N_595);
nor U605 (N_605,N_551,N_568);
and U606 (N_606,N_578,N_594);
nor U607 (N_607,N_579,N_549);
and U608 (N_608,N_547,N_542);
or U609 (N_609,N_562,N_575);
xor U610 (N_610,N_548,N_561);
and U611 (N_611,N_543,N_596);
and U612 (N_612,N_599,N_558);
and U613 (N_613,N_591,N_555);
or U614 (N_614,N_572,N_552);
and U615 (N_615,N_545,N_593);
and U616 (N_616,N_584,N_571);
or U617 (N_617,N_565,N_588);
or U618 (N_618,N_597,N_589);
nand U619 (N_619,N_563,N_557);
nor U620 (N_620,N_586,N_577);
or U621 (N_621,N_564,N_559);
nand U622 (N_622,N_587,N_598);
and U623 (N_623,N_553,N_541);
or U624 (N_624,N_576,N_544);
nand U625 (N_625,N_567,N_554);
nand U626 (N_626,N_570,N_550);
and U627 (N_627,N_590,N_574);
or U628 (N_628,N_566,N_569);
or U629 (N_629,N_540,N_546);
nand U630 (N_630,N_573,N_541);
and U631 (N_631,N_554,N_587);
nand U632 (N_632,N_544,N_556);
nand U633 (N_633,N_585,N_598);
nand U634 (N_634,N_560,N_565);
and U635 (N_635,N_587,N_589);
or U636 (N_636,N_599,N_594);
and U637 (N_637,N_572,N_554);
and U638 (N_638,N_550,N_593);
nor U639 (N_639,N_586,N_592);
or U640 (N_640,N_577,N_545);
or U641 (N_641,N_595,N_587);
or U642 (N_642,N_594,N_591);
nand U643 (N_643,N_596,N_579);
or U644 (N_644,N_564,N_552);
nand U645 (N_645,N_579,N_562);
nor U646 (N_646,N_557,N_580);
and U647 (N_647,N_545,N_595);
or U648 (N_648,N_583,N_548);
nand U649 (N_649,N_584,N_556);
nor U650 (N_650,N_597,N_592);
or U651 (N_651,N_569,N_565);
or U652 (N_652,N_572,N_578);
and U653 (N_653,N_581,N_565);
nor U654 (N_654,N_591,N_552);
and U655 (N_655,N_573,N_586);
nor U656 (N_656,N_582,N_558);
or U657 (N_657,N_597,N_576);
nor U658 (N_658,N_543,N_593);
nor U659 (N_659,N_574,N_576);
and U660 (N_660,N_640,N_659);
nor U661 (N_661,N_651,N_646);
or U662 (N_662,N_639,N_653);
and U663 (N_663,N_610,N_626);
or U664 (N_664,N_657,N_631);
nor U665 (N_665,N_635,N_645);
nand U666 (N_666,N_642,N_654);
nor U667 (N_667,N_618,N_602);
or U668 (N_668,N_605,N_603);
nor U669 (N_669,N_630,N_628);
and U670 (N_670,N_607,N_611);
nor U671 (N_671,N_612,N_617);
or U672 (N_672,N_634,N_623);
nand U673 (N_673,N_627,N_606);
and U674 (N_674,N_656,N_632);
xnor U675 (N_675,N_644,N_600);
or U676 (N_676,N_629,N_624);
and U677 (N_677,N_609,N_608);
nor U678 (N_678,N_619,N_625);
and U679 (N_679,N_649,N_614);
nor U680 (N_680,N_647,N_621);
nor U681 (N_681,N_650,N_641);
nand U682 (N_682,N_620,N_648);
nand U683 (N_683,N_616,N_613);
and U684 (N_684,N_633,N_637);
nand U685 (N_685,N_601,N_652);
nand U686 (N_686,N_622,N_636);
nand U687 (N_687,N_655,N_643);
and U688 (N_688,N_658,N_604);
and U689 (N_689,N_638,N_615);
nand U690 (N_690,N_642,N_648);
or U691 (N_691,N_638,N_658);
nand U692 (N_692,N_651,N_653);
nor U693 (N_693,N_643,N_652);
nand U694 (N_694,N_644,N_623);
or U695 (N_695,N_621,N_649);
nand U696 (N_696,N_654,N_659);
nor U697 (N_697,N_612,N_620);
nand U698 (N_698,N_659,N_617);
and U699 (N_699,N_625,N_604);
or U700 (N_700,N_633,N_649);
nor U701 (N_701,N_648,N_604);
or U702 (N_702,N_621,N_637);
nor U703 (N_703,N_633,N_636);
nor U704 (N_704,N_643,N_617);
nand U705 (N_705,N_659,N_626);
and U706 (N_706,N_650,N_653);
nand U707 (N_707,N_610,N_609);
and U708 (N_708,N_617,N_623);
nand U709 (N_709,N_657,N_609);
and U710 (N_710,N_608,N_636);
or U711 (N_711,N_627,N_622);
nor U712 (N_712,N_605,N_656);
nand U713 (N_713,N_629,N_627);
nor U714 (N_714,N_617,N_656);
nor U715 (N_715,N_607,N_623);
and U716 (N_716,N_621,N_642);
nand U717 (N_717,N_658,N_619);
or U718 (N_718,N_608,N_658);
and U719 (N_719,N_618,N_637);
nor U720 (N_720,N_689,N_698);
nand U721 (N_721,N_661,N_693);
or U722 (N_722,N_673,N_660);
or U723 (N_723,N_664,N_670);
nand U724 (N_724,N_697,N_712);
or U725 (N_725,N_678,N_667);
nor U726 (N_726,N_703,N_690);
and U727 (N_727,N_692,N_686);
or U728 (N_728,N_714,N_717);
and U729 (N_729,N_700,N_696);
or U730 (N_730,N_676,N_668);
and U731 (N_731,N_707,N_671);
nor U732 (N_732,N_680,N_688);
and U733 (N_733,N_665,N_682);
and U734 (N_734,N_701,N_695);
nor U735 (N_735,N_669,N_685);
or U736 (N_736,N_716,N_677);
nand U737 (N_737,N_706,N_702);
and U738 (N_738,N_675,N_705);
nand U739 (N_739,N_683,N_713);
nand U740 (N_740,N_718,N_709);
nand U741 (N_741,N_662,N_708);
or U742 (N_742,N_694,N_687);
nand U743 (N_743,N_674,N_663);
or U744 (N_744,N_672,N_711);
and U745 (N_745,N_681,N_715);
xor U746 (N_746,N_666,N_684);
or U747 (N_747,N_710,N_679);
or U748 (N_748,N_691,N_699);
or U749 (N_749,N_719,N_704);
and U750 (N_750,N_698,N_660);
and U751 (N_751,N_666,N_711);
nand U752 (N_752,N_676,N_700);
or U753 (N_753,N_677,N_713);
xor U754 (N_754,N_671,N_705);
and U755 (N_755,N_695,N_665);
or U756 (N_756,N_715,N_672);
or U757 (N_757,N_692,N_688);
nor U758 (N_758,N_709,N_694);
nor U759 (N_759,N_663,N_667);
and U760 (N_760,N_667,N_705);
or U761 (N_761,N_686,N_711);
and U762 (N_762,N_660,N_686);
xnor U763 (N_763,N_662,N_717);
and U764 (N_764,N_717,N_686);
and U765 (N_765,N_676,N_716);
nor U766 (N_766,N_710,N_675);
or U767 (N_767,N_665,N_672);
and U768 (N_768,N_661,N_668);
nand U769 (N_769,N_710,N_682);
nor U770 (N_770,N_686,N_706);
nand U771 (N_771,N_681,N_701);
nor U772 (N_772,N_699,N_680);
or U773 (N_773,N_691,N_673);
and U774 (N_774,N_660,N_696);
nand U775 (N_775,N_711,N_695);
nor U776 (N_776,N_666,N_716);
nor U777 (N_777,N_675,N_668);
nand U778 (N_778,N_703,N_684);
nor U779 (N_779,N_705,N_666);
nor U780 (N_780,N_765,N_767);
and U781 (N_781,N_739,N_770);
or U782 (N_782,N_731,N_752);
and U783 (N_783,N_775,N_742);
or U784 (N_784,N_776,N_757);
nand U785 (N_785,N_773,N_753);
nor U786 (N_786,N_729,N_728);
and U787 (N_787,N_762,N_732);
nand U788 (N_788,N_744,N_763);
and U789 (N_789,N_745,N_725);
nor U790 (N_790,N_721,N_758);
or U791 (N_791,N_774,N_751);
nand U792 (N_792,N_730,N_756);
or U793 (N_793,N_748,N_736);
or U794 (N_794,N_766,N_754);
or U795 (N_795,N_734,N_771);
nand U796 (N_796,N_755,N_759);
and U797 (N_797,N_747,N_768);
and U798 (N_798,N_746,N_769);
and U799 (N_799,N_778,N_733);
nor U800 (N_800,N_740,N_722);
nor U801 (N_801,N_743,N_779);
or U802 (N_802,N_727,N_724);
nand U803 (N_803,N_741,N_761);
and U804 (N_804,N_737,N_738);
and U805 (N_805,N_760,N_726);
nand U806 (N_806,N_749,N_720);
nor U807 (N_807,N_772,N_764);
and U808 (N_808,N_777,N_723);
and U809 (N_809,N_735,N_750);
nand U810 (N_810,N_762,N_730);
nor U811 (N_811,N_739,N_740);
and U812 (N_812,N_723,N_778);
or U813 (N_813,N_726,N_763);
and U814 (N_814,N_773,N_730);
nor U815 (N_815,N_756,N_746);
or U816 (N_816,N_722,N_746);
nand U817 (N_817,N_720,N_740);
or U818 (N_818,N_776,N_742);
nand U819 (N_819,N_772,N_760);
nand U820 (N_820,N_736,N_720);
and U821 (N_821,N_768,N_722);
nand U822 (N_822,N_750,N_731);
nand U823 (N_823,N_751,N_741);
and U824 (N_824,N_734,N_746);
nand U825 (N_825,N_762,N_775);
nor U826 (N_826,N_758,N_748);
nand U827 (N_827,N_771,N_738);
nand U828 (N_828,N_774,N_750);
and U829 (N_829,N_740,N_732);
nand U830 (N_830,N_751,N_736);
nand U831 (N_831,N_774,N_776);
nor U832 (N_832,N_724,N_757);
nor U833 (N_833,N_732,N_757);
and U834 (N_834,N_729,N_771);
nand U835 (N_835,N_765,N_741);
nand U836 (N_836,N_770,N_724);
nor U837 (N_837,N_735,N_744);
nor U838 (N_838,N_761,N_768);
and U839 (N_839,N_744,N_751);
nand U840 (N_840,N_817,N_826);
nor U841 (N_841,N_808,N_796);
nand U842 (N_842,N_787,N_837);
nand U843 (N_843,N_824,N_815);
nand U844 (N_844,N_802,N_828);
and U845 (N_845,N_806,N_827);
or U846 (N_846,N_816,N_795);
nor U847 (N_847,N_780,N_812);
nand U848 (N_848,N_794,N_798);
nand U849 (N_849,N_805,N_789);
or U850 (N_850,N_797,N_801);
nand U851 (N_851,N_781,N_810);
or U852 (N_852,N_804,N_807);
and U853 (N_853,N_790,N_822);
or U854 (N_854,N_831,N_835);
or U855 (N_855,N_793,N_836);
or U856 (N_856,N_811,N_791);
nor U857 (N_857,N_820,N_799);
or U858 (N_858,N_829,N_809);
nand U859 (N_859,N_818,N_792);
nor U860 (N_860,N_823,N_821);
nand U861 (N_861,N_832,N_785);
nor U862 (N_862,N_825,N_783);
nand U863 (N_863,N_830,N_800);
nor U864 (N_864,N_819,N_813);
nand U865 (N_865,N_838,N_784);
or U866 (N_866,N_834,N_839);
nand U867 (N_867,N_833,N_782);
or U868 (N_868,N_788,N_814);
or U869 (N_869,N_786,N_803);
and U870 (N_870,N_801,N_800);
nand U871 (N_871,N_828,N_796);
nor U872 (N_872,N_791,N_780);
or U873 (N_873,N_824,N_836);
or U874 (N_874,N_788,N_780);
or U875 (N_875,N_801,N_822);
nand U876 (N_876,N_826,N_829);
and U877 (N_877,N_791,N_825);
nor U878 (N_878,N_788,N_820);
nand U879 (N_879,N_790,N_833);
and U880 (N_880,N_784,N_821);
or U881 (N_881,N_797,N_825);
and U882 (N_882,N_830,N_799);
nand U883 (N_883,N_814,N_780);
nor U884 (N_884,N_835,N_827);
nand U885 (N_885,N_819,N_790);
and U886 (N_886,N_815,N_806);
nand U887 (N_887,N_825,N_805);
or U888 (N_888,N_810,N_791);
nor U889 (N_889,N_821,N_792);
nor U890 (N_890,N_837,N_816);
nor U891 (N_891,N_822,N_783);
or U892 (N_892,N_839,N_805);
nand U893 (N_893,N_789,N_784);
and U894 (N_894,N_808,N_816);
nor U895 (N_895,N_808,N_804);
and U896 (N_896,N_825,N_794);
nand U897 (N_897,N_813,N_833);
or U898 (N_898,N_839,N_799);
or U899 (N_899,N_794,N_831);
nor U900 (N_900,N_880,N_875);
and U901 (N_901,N_888,N_855);
nand U902 (N_902,N_897,N_863);
and U903 (N_903,N_898,N_850);
or U904 (N_904,N_858,N_865);
nor U905 (N_905,N_853,N_879);
and U906 (N_906,N_859,N_852);
nand U907 (N_907,N_877,N_894);
nand U908 (N_908,N_889,N_890);
nor U909 (N_909,N_868,N_848);
or U910 (N_910,N_886,N_861);
nand U911 (N_911,N_895,N_862);
xnor U912 (N_912,N_843,N_869);
nand U913 (N_913,N_882,N_878);
nor U914 (N_914,N_857,N_871);
or U915 (N_915,N_842,N_892);
nand U916 (N_916,N_899,N_840);
nor U917 (N_917,N_866,N_856);
nor U918 (N_918,N_872,N_845);
nand U919 (N_919,N_893,N_884);
or U920 (N_920,N_864,N_883);
or U921 (N_921,N_881,N_860);
nor U922 (N_922,N_851,N_867);
nor U923 (N_923,N_846,N_849);
or U924 (N_924,N_847,N_885);
nand U925 (N_925,N_844,N_887);
nand U926 (N_926,N_874,N_896);
or U927 (N_927,N_873,N_891);
nand U928 (N_928,N_854,N_876);
or U929 (N_929,N_870,N_841);
or U930 (N_930,N_897,N_885);
and U931 (N_931,N_889,N_884);
and U932 (N_932,N_894,N_843);
nand U933 (N_933,N_890,N_864);
and U934 (N_934,N_894,N_898);
or U935 (N_935,N_897,N_867);
and U936 (N_936,N_858,N_855);
or U937 (N_937,N_840,N_875);
nor U938 (N_938,N_871,N_886);
nand U939 (N_939,N_852,N_892);
xor U940 (N_940,N_845,N_864);
and U941 (N_941,N_878,N_860);
nor U942 (N_942,N_859,N_885);
nand U943 (N_943,N_868,N_846);
xnor U944 (N_944,N_869,N_867);
nand U945 (N_945,N_863,N_865);
xnor U946 (N_946,N_875,N_898);
or U947 (N_947,N_889,N_868);
nand U948 (N_948,N_899,N_848);
or U949 (N_949,N_873,N_878);
and U950 (N_950,N_899,N_844);
or U951 (N_951,N_871,N_891);
nor U952 (N_952,N_875,N_876);
nand U953 (N_953,N_882,N_858);
or U954 (N_954,N_874,N_877);
or U955 (N_955,N_877,N_840);
nor U956 (N_956,N_845,N_841);
and U957 (N_957,N_857,N_848);
or U958 (N_958,N_896,N_856);
nand U959 (N_959,N_849,N_871);
and U960 (N_960,N_928,N_938);
or U961 (N_961,N_937,N_907);
and U962 (N_962,N_900,N_910);
and U963 (N_963,N_918,N_911);
nand U964 (N_964,N_926,N_916);
or U965 (N_965,N_944,N_950);
nand U966 (N_966,N_955,N_951);
nand U967 (N_967,N_925,N_901);
nor U968 (N_968,N_946,N_953);
nand U969 (N_969,N_936,N_917);
or U970 (N_970,N_905,N_932);
nor U971 (N_971,N_920,N_903);
nand U972 (N_972,N_941,N_913);
xnor U973 (N_973,N_908,N_919);
nand U974 (N_974,N_942,N_949);
and U975 (N_975,N_939,N_902);
nand U976 (N_976,N_958,N_906);
or U977 (N_977,N_915,N_929);
and U978 (N_978,N_947,N_959);
nor U979 (N_979,N_914,N_940);
and U980 (N_980,N_943,N_935);
nor U981 (N_981,N_952,N_945);
or U982 (N_982,N_948,N_957);
nor U983 (N_983,N_927,N_923);
or U984 (N_984,N_912,N_921);
nor U985 (N_985,N_922,N_909);
nand U986 (N_986,N_924,N_931);
or U987 (N_987,N_956,N_930);
or U988 (N_988,N_933,N_954);
or U989 (N_989,N_904,N_934);
nor U990 (N_990,N_915,N_950);
or U991 (N_991,N_919,N_958);
or U992 (N_992,N_946,N_923);
nand U993 (N_993,N_923,N_913);
and U994 (N_994,N_900,N_925);
or U995 (N_995,N_929,N_921);
or U996 (N_996,N_908,N_907);
nor U997 (N_997,N_927,N_926);
or U998 (N_998,N_932,N_950);
nor U999 (N_999,N_936,N_943);
and U1000 (N_1000,N_937,N_915);
or U1001 (N_1001,N_901,N_956);
or U1002 (N_1002,N_959,N_917);
and U1003 (N_1003,N_925,N_916);
or U1004 (N_1004,N_912,N_946);
nand U1005 (N_1005,N_909,N_917);
and U1006 (N_1006,N_930,N_946);
and U1007 (N_1007,N_933,N_920);
nor U1008 (N_1008,N_916,N_946);
or U1009 (N_1009,N_940,N_941);
xnor U1010 (N_1010,N_952,N_914);
or U1011 (N_1011,N_934,N_919);
and U1012 (N_1012,N_956,N_920);
nor U1013 (N_1013,N_912,N_925);
and U1014 (N_1014,N_941,N_922);
and U1015 (N_1015,N_917,N_951);
nand U1016 (N_1016,N_911,N_954);
or U1017 (N_1017,N_949,N_919);
nand U1018 (N_1018,N_912,N_913);
nor U1019 (N_1019,N_935,N_929);
and U1020 (N_1020,N_986,N_970);
nand U1021 (N_1021,N_989,N_995);
or U1022 (N_1022,N_1009,N_963);
nand U1023 (N_1023,N_994,N_981);
or U1024 (N_1024,N_1018,N_1002);
nor U1025 (N_1025,N_1011,N_1000);
nor U1026 (N_1026,N_979,N_964);
and U1027 (N_1027,N_975,N_977);
and U1028 (N_1028,N_1003,N_982);
nand U1029 (N_1029,N_1014,N_961);
nor U1030 (N_1030,N_983,N_972);
nand U1031 (N_1031,N_1015,N_973);
or U1032 (N_1032,N_998,N_1008);
or U1033 (N_1033,N_969,N_978);
or U1034 (N_1034,N_968,N_993);
or U1035 (N_1035,N_1017,N_990);
and U1036 (N_1036,N_991,N_985);
nand U1037 (N_1037,N_1006,N_1019);
or U1038 (N_1038,N_1001,N_996);
and U1039 (N_1039,N_984,N_992);
nor U1040 (N_1040,N_976,N_1004);
nand U1041 (N_1041,N_999,N_1010);
and U1042 (N_1042,N_971,N_966);
nor U1043 (N_1043,N_997,N_1005);
or U1044 (N_1044,N_967,N_988);
and U1045 (N_1045,N_980,N_960);
nand U1046 (N_1046,N_965,N_962);
or U1047 (N_1047,N_1007,N_987);
nand U1048 (N_1048,N_974,N_1012);
or U1049 (N_1049,N_1016,N_1013);
or U1050 (N_1050,N_964,N_972);
and U1051 (N_1051,N_1016,N_964);
nand U1052 (N_1052,N_961,N_991);
nand U1053 (N_1053,N_1006,N_1015);
nor U1054 (N_1054,N_993,N_1003);
or U1055 (N_1055,N_968,N_1016);
and U1056 (N_1056,N_1008,N_1011);
nand U1057 (N_1057,N_976,N_962);
or U1058 (N_1058,N_1009,N_1014);
nor U1059 (N_1059,N_988,N_964);
or U1060 (N_1060,N_1011,N_987);
or U1061 (N_1061,N_997,N_1002);
nor U1062 (N_1062,N_961,N_1008);
or U1063 (N_1063,N_980,N_985);
or U1064 (N_1064,N_980,N_990);
and U1065 (N_1065,N_1008,N_1014);
or U1066 (N_1066,N_1014,N_1002);
and U1067 (N_1067,N_981,N_1009);
or U1068 (N_1068,N_970,N_1001);
and U1069 (N_1069,N_971,N_992);
or U1070 (N_1070,N_995,N_974);
and U1071 (N_1071,N_969,N_995);
or U1072 (N_1072,N_986,N_985);
xnor U1073 (N_1073,N_974,N_1009);
or U1074 (N_1074,N_991,N_987);
nand U1075 (N_1075,N_1019,N_986);
nor U1076 (N_1076,N_1008,N_1007);
and U1077 (N_1077,N_996,N_998);
xor U1078 (N_1078,N_968,N_971);
and U1079 (N_1079,N_1001,N_1019);
nor U1080 (N_1080,N_1030,N_1025);
and U1081 (N_1081,N_1053,N_1034);
nand U1082 (N_1082,N_1075,N_1065);
or U1083 (N_1083,N_1070,N_1049);
nor U1084 (N_1084,N_1046,N_1074);
nand U1085 (N_1085,N_1039,N_1033);
nor U1086 (N_1086,N_1052,N_1045);
nand U1087 (N_1087,N_1069,N_1040);
nand U1088 (N_1088,N_1077,N_1071);
nor U1089 (N_1089,N_1051,N_1044);
nand U1090 (N_1090,N_1056,N_1062);
and U1091 (N_1091,N_1041,N_1035);
or U1092 (N_1092,N_1037,N_1050);
nor U1093 (N_1093,N_1031,N_1054);
nand U1094 (N_1094,N_1060,N_1068);
and U1095 (N_1095,N_1020,N_1027);
nor U1096 (N_1096,N_1024,N_1032);
and U1097 (N_1097,N_1022,N_1067);
and U1098 (N_1098,N_1048,N_1073);
or U1099 (N_1099,N_1047,N_1076);
nor U1100 (N_1100,N_1028,N_1072);
xor U1101 (N_1101,N_1021,N_1058);
nor U1102 (N_1102,N_1042,N_1079);
nor U1103 (N_1103,N_1066,N_1023);
nand U1104 (N_1104,N_1064,N_1055);
or U1105 (N_1105,N_1057,N_1029);
nand U1106 (N_1106,N_1078,N_1038);
nor U1107 (N_1107,N_1036,N_1061);
nor U1108 (N_1108,N_1026,N_1043);
nand U1109 (N_1109,N_1063,N_1059);
nor U1110 (N_1110,N_1048,N_1049);
nand U1111 (N_1111,N_1059,N_1042);
or U1112 (N_1112,N_1025,N_1034);
nand U1113 (N_1113,N_1066,N_1041);
nor U1114 (N_1114,N_1026,N_1063);
nand U1115 (N_1115,N_1023,N_1048);
or U1116 (N_1116,N_1057,N_1050);
and U1117 (N_1117,N_1046,N_1054);
xnor U1118 (N_1118,N_1032,N_1029);
nand U1119 (N_1119,N_1054,N_1034);
nand U1120 (N_1120,N_1054,N_1035);
nor U1121 (N_1121,N_1021,N_1069);
nor U1122 (N_1122,N_1062,N_1060);
nand U1123 (N_1123,N_1058,N_1040);
nor U1124 (N_1124,N_1034,N_1023);
or U1125 (N_1125,N_1079,N_1075);
nor U1126 (N_1126,N_1031,N_1045);
nor U1127 (N_1127,N_1028,N_1043);
or U1128 (N_1128,N_1050,N_1030);
nand U1129 (N_1129,N_1051,N_1025);
and U1130 (N_1130,N_1039,N_1045);
and U1131 (N_1131,N_1037,N_1056);
nor U1132 (N_1132,N_1022,N_1043);
nand U1133 (N_1133,N_1048,N_1054);
nand U1134 (N_1134,N_1056,N_1066);
or U1135 (N_1135,N_1020,N_1074);
nor U1136 (N_1136,N_1053,N_1024);
nand U1137 (N_1137,N_1036,N_1064);
nor U1138 (N_1138,N_1045,N_1047);
nor U1139 (N_1139,N_1065,N_1052);
or U1140 (N_1140,N_1119,N_1089);
or U1141 (N_1141,N_1103,N_1087);
and U1142 (N_1142,N_1113,N_1106);
nor U1143 (N_1143,N_1122,N_1099);
and U1144 (N_1144,N_1133,N_1090);
or U1145 (N_1145,N_1081,N_1125);
nor U1146 (N_1146,N_1083,N_1129);
nor U1147 (N_1147,N_1084,N_1127);
nor U1148 (N_1148,N_1093,N_1112);
nor U1149 (N_1149,N_1086,N_1091);
nor U1150 (N_1150,N_1094,N_1139);
nor U1151 (N_1151,N_1105,N_1130);
nor U1152 (N_1152,N_1097,N_1088);
nor U1153 (N_1153,N_1114,N_1138);
and U1154 (N_1154,N_1124,N_1116);
and U1155 (N_1155,N_1137,N_1100);
or U1156 (N_1156,N_1132,N_1115);
nor U1157 (N_1157,N_1110,N_1102);
nor U1158 (N_1158,N_1098,N_1111);
nor U1159 (N_1159,N_1082,N_1134);
and U1160 (N_1160,N_1123,N_1085);
nand U1161 (N_1161,N_1092,N_1109);
nand U1162 (N_1162,N_1104,N_1095);
nand U1163 (N_1163,N_1117,N_1136);
nor U1164 (N_1164,N_1128,N_1120);
nand U1165 (N_1165,N_1135,N_1108);
and U1166 (N_1166,N_1101,N_1107);
nand U1167 (N_1167,N_1080,N_1096);
nand U1168 (N_1168,N_1126,N_1118);
and U1169 (N_1169,N_1121,N_1131);
and U1170 (N_1170,N_1121,N_1096);
nor U1171 (N_1171,N_1115,N_1102);
nand U1172 (N_1172,N_1118,N_1100);
nand U1173 (N_1173,N_1123,N_1090);
and U1174 (N_1174,N_1117,N_1111);
xor U1175 (N_1175,N_1121,N_1138);
nor U1176 (N_1176,N_1103,N_1120);
and U1177 (N_1177,N_1086,N_1111);
nand U1178 (N_1178,N_1139,N_1096);
or U1179 (N_1179,N_1096,N_1125);
or U1180 (N_1180,N_1084,N_1080);
or U1181 (N_1181,N_1115,N_1113);
nor U1182 (N_1182,N_1135,N_1087);
nand U1183 (N_1183,N_1129,N_1089);
nor U1184 (N_1184,N_1130,N_1102);
nor U1185 (N_1185,N_1088,N_1129);
or U1186 (N_1186,N_1113,N_1130);
nand U1187 (N_1187,N_1103,N_1116);
nand U1188 (N_1188,N_1119,N_1088);
and U1189 (N_1189,N_1101,N_1125);
and U1190 (N_1190,N_1118,N_1121);
and U1191 (N_1191,N_1108,N_1122);
and U1192 (N_1192,N_1084,N_1120);
and U1193 (N_1193,N_1112,N_1119);
and U1194 (N_1194,N_1131,N_1106);
nand U1195 (N_1195,N_1118,N_1138);
or U1196 (N_1196,N_1099,N_1125);
nand U1197 (N_1197,N_1119,N_1117);
nor U1198 (N_1198,N_1129,N_1116);
nand U1199 (N_1199,N_1082,N_1083);
and U1200 (N_1200,N_1144,N_1154);
nor U1201 (N_1201,N_1148,N_1169);
or U1202 (N_1202,N_1150,N_1195);
nand U1203 (N_1203,N_1185,N_1153);
nor U1204 (N_1204,N_1149,N_1189);
nor U1205 (N_1205,N_1165,N_1171);
nor U1206 (N_1206,N_1199,N_1188);
and U1207 (N_1207,N_1147,N_1177);
nand U1208 (N_1208,N_1160,N_1190);
nor U1209 (N_1209,N_1196,N_1151);
or U1210 (N_1210,N_1198,N_1155);
nor U1211 (N_1211,N_1193,N_1146);
nor U1212 (N_1212,N_1173,N_1164);
nor U1213 (N_1213,N_1163,N_1186);
and U1214 (N_1214,N_1162,N_1176);
and U1215 (N_1215,N_1187,N_1178);
and U1216 (N_1216,N_1180,N_1157);
nor U1217 (N_1217,N_1182,N_1166);
and U1218 (N_1218,N_1194,N_1140);
nand U1219 (N_1219,N_1191,N_1159);
or U1220 (N_1220,N_1141,N_1183);
xor U1221 (N_1221,N_1181,N_1168);
nor U1222 (N_1222,N_1156,N_1152);
nand U1223 (N_1223,N_1192,N_1161);
and U1224 (N_1224,N_1158,N_1143);
or U1225 (N_1225,N_1184,N_1142);
nand U1226 (N_1226,N_1197,N_1175);
nand U1227 (N_1227,N_1170,N_1174);
nand U1228 (N_1228,N_1167,N_1179);
nand U1229 (N_1229,N_1145,N_1172);
xnor U1230 (N_1230,N_1167,N_1183);
xor U1231 (N_1231,N_1142,N_1154);
nor U1232 (N_1232,N_1168,N_1175);
nand U1233 (N_1233,N_1194,N_1164);
or U1234 (N_1234,N_1192,N_1191);
and U1235 (N_1235,N_1179,N_1175);
nor U1236 (N_1236,N_1193,N_1195);
nor U1237 (N_1237,N_1161,N_1176);
nor U1238 (N_1238,N_1190,N_1192);
nor U1239 (N_1239,N_1162,N_1193);
nor U1240 (N_1240,N_1191,N_1167);
or U1241 (N_1241,N_1140,N_1147);
or U1242 (N_1242,N_1173,N_1156);
and U1243 (N_1243,N_1158,N_1178);
nor U1244 (N_1244,N_1158,N_1187);
and U1245 (N_1245,N_1182,N_1152);
and U1246 (N_1246,N_1196,N_1169);
or U1247 (N_1247,N_1198,N_1177);
nand U1248 (N_1248,N_1141,N_1173);
nor U1249 (N_1249,N_1183,N_1176);
nand U1250 (N_1250,N_1155,N_1145);
and U1251 (N_1251,N_1182,N_1159);
nor U1252 (N_1252,N_1178,N_1162);
or U1253 (N_1253,N_1144,N_1147);
or U1254 (N_1254,N_1174,N_1179);
and U1255 (N_1255,N_1180,N_1166);
or U1256 (N_1256,N_1141,N_1177);
nor U1257 (N_1257,N_1173,N_1143);
or U1258 (N_1258,N_1188,N_1148);
and U1259 (N_1259,N_1156,N_1170);
nand U1260 (N_1260,N_1221,N_1203);
nor U1261 (N_1261,N_1250,N_1223);
nor U1262 (N_1262,N_1207,N_1219);
nand U1263 (N_1263,N_1234,N_1226);
and U1264 (N_1264,N_1204,N_1247);
or U1265 (N_1265,N_1236,N_1227);
nand U1266 (N_1266,N_1241,N_1256);
or U1267 (N_1267,N_1254,N_1249);
nand U1268 (N_1268,N_1217,N_1215);
nand U1269 (N_1269,N_1228,N_1252);
or U1270 (N_1270,N_1239,N_1202);
or U1271 (N_1271,N_1240,N_1231);
or U1272 (N_1272,N_1230,N_1206);
nor U1273 (N_1273,N_1222,N_1211);
or U1274 (N_1274,N_1232,N_1208);
nand U1275 (N_1275,N_1224,N_1200);
or U1276 (N_1276,N_1253,N_1244);
nand U1277 (N_1277,N_1235,N_1248);
or U1278 (N_1278,N_1213,N_1229);
and U1279 (N_1279,N_1251,N_1259);
and U1280 (N_1280,N_1212,N_1258);
nand U1281 (N_1281,N_1237,N_1225);
or U1282 (N_1282,N_1216,N_1214);
nor U1283 (N_1283,N_1238,N_1257);
or U1284 (N_1284,N_1243,N_1246);
or U1285 (N_1285,N_1210,N_1255);
nor U1286 (N_1286,N_1220,N_1218);
or U1287 (N_1287,N_1205,N_1201);
and U1288 (N_1288,N_1209,N_1242);
nor U1289 (N_1289,N_1233,N_1245);
and U1290 (N_1290,N_1251,N_1201);
and U1291 (N_1291,N_1217,N_1203);
nor U1292 (N_1292,N_1247,N_1248);
and U1293 (N_1293,N_1212,N_1234);
nand U1294 (N_1294,N_1250,N_1214);
nand U1295 (N_1295,N_1250,N_1203);
and U1296 (N_1296,N_1217,N_1208);
or U1297 (N_1297,N_1247,N_1210);
nand U1298 (N_1298,N_1247,N_1202);
or U1299 (N_1299,N_1245,N_1250);
xnor U1300 (N_1300,N_1225,N_1247);
and U1301 (N_1301,N_1218,N_1224);
nor U1302 (N_1302,N_1201,N_1243);
or U1303 (N_1303,N_1205,N_1212);
nor U1304 (N_1304,N_1210,N_1219);
or U1305 (N_1305,N_1238,N_1226);
or U1306 (N_1306,N_1227,N_1259);
and U1307 (N_1307,N_1237,N_1240);
and U1308 (N_1308,N_1250,N_1222);
and U1309 (N_1309,N_1219,N_1258);
and U1310 (N_1310,N_1202,N_1227);
or U1311 (N_1311,N_1258,N_1253);
nand U1312 (N_1312,N_1249,N_1257);
or U1313 (N_1313,N_1254,N_1237);
nor U1314 (N_1314,N_1243,N_1206);
or U1315 (N_1315,N_1212,N_1225);
or U1316 (N_1316,N_1219,N_1227);
nand U1317 (N_1317,N_1233,N_1200);
nor U1318 (N_1318,N_1226,N_1251);
or U1319 (N_1319,N_1247,N_1222);
nor U1320 (N_1320,N_1288,N_1267);
nor U1321 (N_1321,N_1294,N_1316);
nand U1322 (N_1322,N_1278,N_1309);
nor U1323 (N_1323,N_1300,N_1308);
or U1324 (N_1324,N_1313,N_1295);
nand U1325 (N_1325,N_1264,N_1274);
and U1326 (N_1326,N_1293,N_1270);
or U1327 (N_1327,N_1284,N_1265);
nand U1328 (N_1328,N_1272,N_1289);
or U1329 (N_1329,N_1310,N_1318);
and U1330 (N_1330,N_1297,N_1273);
nand U1331 (N_1331,N_1305,N_1291);
and U1332 (N_1332,N_1290,N_1282);
nor U1333 (N_1333,N_1299,N_1268);
or U1334 (N_1334,N_1266,N_1319);
nand U1335 (N_1335,N_1261,N_1315);
or U1336 (N_1336,N_1280,N_1303);
nand U1337 (N_1337,N_1285,N_1307);
nand U1338 (N_1338,N_1302,N_1260);
and U1339 (N_1339,N_1311,N_1269);
nand U1340 (N_1340,N_1281,N_1304);
and U1341 (N_1341,N_1262,N_1271);
and U1342 (N_1342,N_1275,N_1277);
and U1343 (N_1343,N_1306,N_1279);
and U1344 (N_1344,N_1314,N_1317);
nor U1345 (N_1345,N_1263,N_1301);
or U1346 (N_1346,N_1296,N_1286);
or U1347 (N_1347,N_1298,N_1276);
nand U1348 (N_1348,N_1283,N_1287);
and U1349 (N_1349,N_1312,N_1292);
and U1350 (N_1350,N_1262,N_1299);
nand U1351 (N_1351,N_1271,N_1317);
nand U1352 (N_1352,N_1274,N_1313);
nor U1353 (N_1353,N_1314,N_1307);
or U1354 (N_1354,N_1284,N_1313);
nand U1355 (N_1355,N_1316,N_1296);
nand U1356 (N_1356,N_1273,N_1311);
or U1357 (N_1357,N_1284,N_1303);
nand U1358 (N_1358,N_1262,N_1297);
and U1359 (N_1359,N_1277,N_1265);
or U1360 (N_1360,N_1283,N_1292);
nand U1361 (N_1361,N_1314,N_1294);
nand U1362 (N_1362,N_1276,N_1284);
nor U1363 (N_1363,N_1264,N_1291);
or U1364 (N_1364,N_1281,N_1264);
nor U1365 (N_1365,N_1292,N_1265);
nor U1366 (N_1366,N_1296,N_1295);
nand U1367 (N_1367,N_1319,N_1315);
and U1368 (N_1368,N_1316,N_1283);
nand U1369 (N_1369,N_1317,N_1303);
nor U1370 (N_1370,N_1301,N_1291);
and U1371 (N_1371,N_1273,N_1310);
or U1372 (N_1372,N_1282,N_1275);
nor U1373 (N_1373,N_1319,N_1269);
or U1374 (N_1374,N_1274,N_1295);
and U1375 (N_1375,N_1298,N_1309);
nand U1376 (N_1376,N_1317,N_1297);
nand U1377 (N_1377,N_1316,N_1309);
nor U1378 (N_1378,N_1262,N_1296);
nor U1379 (N_1379,N_1264,N_1293);
nor U1380 (N_1380,N_1367,N_1373);
or U1381 (N_1381,N_1349,N_1331);
or U1382 (N_1382,N_1358,N_1326);
or U1383 (N_1383,N_1347,N_1370);
or U1384 (N_1384,N_1359,N_1372);
or U1385 (N_1385,N_1352,N_1353);
or U1386 (N_1386,N_1375,N_1337);
and U1387 (N_1387,N_1356,N_1341);
nand U1388 (N_1388,N_1344,N_1335);
nand U1389 (N_1389,N_1369,N_1350);
and U1390 (N_1390,N_1325,N_1364);
or U1391 (N_1391,N_1379,N_1323);
nand U1392 (N_1392,N_1357,N_1321);
and U1393 (N_1393,N_1376,N_1366);
nand U1394 (N_1394,N_1361,N_1354);
nor U1395 (N_1395,N_1332,N_1322);
nand U1396 (N_1396,N_1328,N_1346);
and U1397 (N_1397,N_1345,N_1342);
nand U1398 (N_1398,N_1324,N_1371);
nor U1399 (N_1399,N_1333,N_1338);
nand U1400 (N_1400,N_1368,N_1327);
and U1401 (N_1401,N_1336,N_1320);
nor U1402 (N_1402,N_1330,N_1363);
nand U1403 (N_1403,N_1374,N_1348);
nand U1404 (N_1404,N_1360,N_1334);
nand U1405 (N_1405,N_1365,N_1329);
nand U1406 (N_1406,N_1339,N_1362);
nor U1407 (N_1407,N_1378,N_1355);
nand U1408 (N_1408,N_1377,N_1343);
and U1409 (N_1409,N_1340,N_1351);
and U1410 (N_1410,N_1377,N_1327);
nor U1411 (N_1411,N_1358,N_1332);
nand U1412 (N_1412,N_1379,N_1334);
nand U1413 (N_1413,N_1360,N_1324);
nand U1414 (N_1414,N_1325,N_1323);
nand U1415 (N_1415,N_1360,N_1342);
nand U1416 (N_1416,N_1327,N_1332);
nand U1417 (N_1417,N_1366,N_1363);
or U1418 (N_1418,N_1342,N_1329);
nand U1419 (N_1419,N_1358,N_1379);
and U1420 (N_1420,N_1341,N_1350);
nor U1421 (N_1421,N_1361,N_1333);
nand U1422 (N_1422,N_1375,N_1373);
and U1423 (N_1423,N_1329,N_1341);
or U1424 (N_1424,N_1373,N_1371);
nand U1425 (N_1425,N_1365,N_1349);
or U1426 (N_1426,N_1325,N_1376);
or U1427 (N_1427,N_1350,N_1347);
nand U1428 (N_1428,N_1376,N_1350);
nor U1429 (N_1429,N_1332,N_1323);
nor U1430 (N_1430,N_1368,N_1324);
or U1431 (N_1431,N_1343,N_1328);
or U1432 (N_1432,N_1325,N_1373);
or U1433 (N_1433,N_1356,N_1357);
or U1434 (N_1434,N_1326,N_1338);
nand U1435 (N_1435,N_1369,N_1372);
or U1436 (N_1436,N_1353,N_1367);
nor U1437 (N_1437,N_1342,N_1363);
or U1438 (N_1438,N_1338,N_1331);
nand U1439 (N_1439,N_1325,N_1379);
or U1440 (N_1440,N_1393,N_1382);
nand U1441 (N_1441,N_1403,N_1408);
or U1442 (N_1442,N_1428,N_1426);
and U1443 (N_1443,N_1402,N_1389);
and U1444 (N_1444,N_1400,N_1385);
nor U1445 (N_1445,N_1419,N_1406);
nor U1446 (N_1446,N_1388,N_1409);
nand U1447 (N_1447,N_1436,N_1390);
or U1448 (N_1448,N_1430,N_1407);
or U1449 (N_1449,N_1438,N_1399);
nor U1450 (N_1450,N_1412,N_1422);
or U1451 (N_1451,N_1417,N_1414);
nand U1452 (N_1452,N_1424,N_1401);
nand U1453 (N_1453,N_1386,N_1384);
nand U1454 (N_1454,N_1395,N_1387);
or U1455 (N_1455,N_1420,N_1432);
nor U1456 (N_1456,N_1433,N_1429);
or U1457 (N_1457,N_1413,N_1397);
or U1458 (N_1458,N_1394,N_1435);
nand U1459 (N_1459,N_1425,N_1380);
nand U1460 (N_1460,N_1415,N_1437);
nand U1461 (N_1461,N_1405,N_1416);
nor U1462 (N_1462,N_1391,N_1381);
and U1463 (N_1463,N_1404,N_1411);
nor U1464 (N_1464,N_1383,N_1396);
and U1465 (N_1465,N_1427,N_1398);
or U1466 (N_1466,N_1418,N_1410);
nand U1467 (N_1467,N_1392,N_1434);
or U1468 (N_1468,N_1421,N_1423);
nor U1469 (N_1469,N_1439,N_1431);
nand U1470 (N_1470,N_1421,N_1436);
and U1471 (N_1471,N_1384,N_1416);
and U1472 (N_1472,N_1381,N_1410);
nor U1473 (N_1473,N_1383,N_1380);
xnor U1474 (N_1474,N_1411,N_1403);
or U1475 (N_1475,N_1381,N_1412);
and U1476 (N_1476,N_1392,N_1439);
and U1477 (N_1477,N_1431,N_1408);
or U1478 (N_1478,N_1405,N_1435);
nand U1479 (N_1479,N_1437,N_1391);
nor U1480 (N_1480,N_1400,N_1423);
nor U1481 (N_1481,N_1397,N_1405);
and U1482 (N_1482,N_1390,N_1420);
nand U1483 (N_1483,N_1439,N_1398);
or U1484 (N_1484,N_1438,N_1420);
nor U1485 (N_1485,N_1425,N_1434);
and U1486 (N_1486,N_1401,N_1393);
and U1487 (N_1487,N_1422,N_1424);
nor U1488 (N_1488,N_1417,N_1392);
nand U1489 (N_1489,N_1428,N_1424);
nor U1490 (N_1490,N_1430,N_1403);
nand U1491 (N_1491,N_1415,N_1436);
or U1492 (N_1492,N_1417,N_1410);
nand U1493 (N_1493,N_1401,N_1403);
or U1494 (N_1494,N_1388,N_1390);
and U1495 (N_1495,N_1382,N_1387);
nor U1496 (N_1496,N_1382,N_1403);
nand U1497 (N_1497,N_1436,N_1427);
or U1498 (N_1498,N_1437,N_1432);
nand U1499 (N_1499,N_1426,N_1401);
or U1500 (N_1500,N_1456,N_1459);
nand U1501 (N_1501,N_1478,N_1442);
and U1502 (N_1502,N_1461,N_1482);
nor U1503 (N_1503,N_1443,N_1492);
and U1504 (N_1504,N_1495,N_1441);
or U1505 (N_1505,N_1448,N_1468);
or U1506 (N_1506,N_1489,N_1490);
nand U1507 (N_1507,N_1472,N_1455);
nor U1508 (N_1508,N_1485,N_1446);
nor U1509 (N_1509,N_1470,N_1498);
or U1510 (N_1510,N_1479,N_1451);
nand U1511 (N_1511,N_1449,N_1462);
nor U1512 (N_1512,N_1471,N_1477);
and U1513 (N_1513,N_1487,N_1474);
or U1514 (N_1514,N_1499,N_1496);
and U1515 (N_1515,N_1453,N_1466);
or U1516 (N_1516,N_1486,N_1491);
nand U1517 (N_1517,N_1463,N_1494);
nand U1518 (N_1518,N_1497,N_1484);
nand U1519 (N_1519,N_1444,N_1458);
nand U1520 (N_1520,N_1488,N_1452);
and U1521 (N_1521,N_1476,N_1450);
or U1522 (N_1522,N_1440,N_1454);
or U1523 (N_1523,N_1483,N_1460);
nor U1524 (N_1524,N_1493,N_1447);
or U1525 (N_1525,N_1481,N_1465);
nand U1526 (N_1526,N_1480,N_1457);
nand U1527 (N_1527,N_1473,N_1467);
or U1528 (N_1528,N_1464,N_1475);
nand U1529 (N_1529,N_1445,N_1469);
nand U1530 (N_1530,N_1445,N_1467);
nor U1531 (N_1531,N_1460,N_1473);
nand U1532 (N_1532,N_1445,N_1493);
and U1533 (N_1533,N_1452,N_1471);
nand U1534 (N_1534,N_1449,N_1461);
nor U1535 (N_1535,N_1444,N_1464);
nor U1536 (N_1536,N_1450,N_1451);
nor U1537 (N_1537,N_1484,N_1494);
and U1538 (N_1538,N_1495,N_1489);
and U1539 (N_1539,N_1493,N_1485);
nand U1540 (N_1540,N_1459,N_1479);
or U1541 (N_1541,N_1444,N_1492);
nand U1542 (N_1542,N_1468,N_1469);
and U1543 (N_1543,N_1477,N_1450);
nor U1544 (N_1544,N_1470,N_1474);
nand U1545 (N_1545,N_1450,N_1471);
nor U1546 (N_1546,N_1474,N_1486);
or U1547 (N_1547,N_1447,N_1492);
and U1548 (N_1548,N_1472,N_1440);
nor U1549 (N_1549,N_1485,N_1499);
nand U1550 (N_1550,N_1460,N_1496);
nand U1551 (N_1551,N_1446,N_1467);
nand U1552 (N_1552,N_1487,N_1470);
nand U1553 (N_1553,N_1467,N_1447);
and U1554 (N_1554,N_1480,N_1460);
nand U1555 (N_1555,N_1498,N_1471);
and U1556 (N_1556,N_1446,N_1451);
nor U1557 (N_1557,N_1456,N_1479);
nor U1558 (N_1558,N_1493,N_1488);
nand U1559 (N_1559,N_1464,N_1474);
or U1560 (N_1560,N_1520,N_1525);
or U1561 (N_1561,N_1553,N_1508);
and U1562 (N_1562,N_1555,N_1557);
nor U1563 (N_1563,N_1511,N_1544);
nand U1564 (N_1564,N_1552,N_1517);
nor U1565 (N_1565,N_1521,N_1545);
nand U1566 (N_1566,N_1534,N_1539);
and U1567 (N_1567,N_1542,N_1506);
nand U1568 (N_1568,N_1527,N_1523);
or U1569 (N_1569,N_1548,N_1526);
nand U1570 (N_1570,N_1541,N_1522);
or U1571 (N_1571,N_1533,N_1547);
nand U1572 (N_1572,N_1514,N_1510);
nand U1573 (N_1573,N_1524,N_1537);
nand U1574 (N_1574,N_1500,N_1513);
and U1575 (N_1575,N_1531,N_1504);
nand U1576 (N_1576,N_1543,N_1558);
xnor U1577 (N_1577,N_1505,N_1529);
and U1578 (N_1578,N_1530,N_1551);
nand U1579 (N_1579,N_1556,N_1518);
nor U1580 (N_1580,N_1519,N_1501);
nor U1581 (N_1581,N_1503,N_1540);
nor U1582 (N_1582,N_1546,N_1549);
nand U1583 (N_1583,N_1532,N_1509);
nor U1584 (N_1584,N_1535,N_1538);
nor U1585 (N_1585,N_1559,N_1512);
or U1586 (N_1586,N_1550,N_1502);
nand U1587 (N_1587,N_1516,N_1507);
or U1588 (N_1588,N_1515,N_1528);
nor U1589 (N_1589,N_1536,N_1554);
and U1590 (N_1590,N_1503,N_1505);
or U1591 (N_1591,N_1535,N_1521);
or U1592 (N_1592,N_1502,N_1554);
or U1593 (N_1593,N_1525,N_1556);
and U1594 (N_1594,N_1522,N_1503);
or U1595 (N_1595,N_1522,N_1531);
or U1596 (N_1596,N_1553,N_1543);
and U1597 (N_1597,N_1503,N_1527);
or U1598 (N_1598,N_1525,N_1524);
nor U1599 (N_1599,N_1505,N_1524);
or U1600 (N_1600,N_1523,N_1504);
nor U1601 (N_1601,N_1540,N_1555);
or U1602 (N_1602,N_1523,N_1518);
nor U1603 (N_1603,N_1505,N_1556);
and U1604 (N_1604,N_1537,N_1545);
and U1605 (N_1605,N_1555,N_1536);
and U1606 (N_1606,N_1525,N_1502);
or U1607 (N_1607,N_1536,N_1516);
and U1608 (N_1608,N_1523,N_1537);
nand U1609 (N_1609,N_1500,N_1550);
xor U1610 (N_1610,N_1512,N_1551);
nor U1611 (N_1611,N_1540,N_1510);
and U1612 (N_1612,N_1514,N_1521);
nand U1613 (N_1613,N_1532,N_1527);
and U1614 (N_1614,N_1544,N_1539);
and U1615 (N_1615,N_1524,N_1558);
and U1616 (N_1616,N_1537,N_1559);
and U1617 (N_1617,N_1556,N_1547);
nor U1618 (N_1618,N_1543,N_1507);
nand U1619 (N_1619,N_1534,N_1557);
or U1620 (N_1620,N_1601,N_1605);
nand U1621 (N_1621,N_1580,N_1600);
nand U1622 (N_1622,N_1581,N_1566);
nand U1623 (N_1623,N_1613,N_1596);
or U1624 (N_1624,N_1571,N_1602);
nor U1625 (N_1625,N_1563,N_1597);
and U1626 (N_1626,N_1574,N_1599);
and U1627 (N_1627,N_1603,N_1591);
and U1628 (N_1628,N_1585,N_1573);
or U1629 (N_1629,N_1565,N_1611);
or U1630 (N_1630,N_1577,N_1575);
and U1631 (N_1631,N_1586,N_1572);
nor U1632 (N_1632,N_1576,N_1562);
nand U1633 (N_1633,N_1560,N_1590);
nand U1634 (N_1634,N_1612,N_1589);
nor U1635 (N_1635,N_1608,N_1568);
nand U1636 (N_1636,N_1616,N_1593);
and U1637 (N_1637,N_1588,N_1598);
nand U1638 (N_1638,N_1564,N_1583);
or U1639 (N_1639,N_1578,N_1609);
nor U1640 (N_1640,N_1561,N_1569);
nor U1641 (N_1641,N_1618,N_1619);
nand U1642 (N_1642,N_1587,N_1604);
xor U1643 (N_1643,N_1594,N_1615);
nand U1644 (N_1644,N_1617,N_1579);
and U1645 (N_1645,N_1592,N_1607);
and U1646 (N_1646,N_1567,N_1582);
and U1647 (N_1647,N_1606,N_1610);
nand U1648 (N_1648,N_1584,N_1595);
and U1649 (N_1649,N_1614,N_1570);
nor U1650 (N_1650,N_1584,N_1587);
or U1651 (N_1651,N_1584,N_1570);
nand U1652 (N_1652,N_1594,N_1579);
and U1653 (N_1653,N_1618,N_1562);
or U1654 (N_1654,N_1610,N_1589);
nand U1655 (N_1655,N_1585,N_1616);
and U1656 (N_1656,N_1577,N_1562);
or U1657 (N_1657,N_1583,N_1577);
or U1658 (N_1658,N_1607,N_1614);
and U1659 (N_1659,N_1617,N_1589);
or U1660 (N_1660,N_1565,N_1570);
nand U1661 (N_1661,N_1582,N_1618);
nand U1662 (N_1662,N_1592,N_1563);
and U1663 (N_1663,N_1603,N_1562);
or U1664 (N_1664,N_1593,N_1579);
or U1665 (N_1665,N_1613,N_1577);
or U1666 (N_1666,N_1604,N_1598);
nor U1667 (N_1667,N_1605,N_1572);
or U1668 (N_1668,N_1563,N_1561);
nand U1669 (N_1669,N_1581,N_1569);
and U1670 (N_1670,N_1601,N_1575);
or U1671 (N_1671,N_1603,N_1608);
and U1672 (N_1672,N_1583,N_1578);
nand U1673 (N_1673,N_1599,N_1592);
and U1674 (N_1674,N_1592,N_1584);
or U1675 (N_1675,N_1605,N_1568);
and U1676 (N_1676,N_1611,N_1598);
nor U1677 (N_1677,N_1598,N_1583);
nor U1678 (N_1678,N_1611,N_1566);
nor U1679 (N_1679,N_1610,N_1609);
nor U1680 (N_1680,N_1653,N_1627);
or U1681 (N_1681,N_1665,N_1661);
nor U1682 (N_1682,N_1655,N_1654);
nand U1683 (N_1683,N_1649,N_1624);
nor U1684 (N_1684,N_1671,N_1648);
and U1685 (N_1685,N_1658,N_1643);
and U1686 (N_1686,N_1650,N_1668);
nand U1687 (N_1687,N_1638,N_1621);
nand U1688 (N_1688,N_1647,N_1676);
and U1689 (N_1689,N_1652,N_1645);
nand U1690 (N_1690,N_1677,N_1679);
and U1691 (N_1691,N_1626,N_1620);
or U1692 (N_1692,N_1660,N_1666);
nand U1693 (N_1693,N_1630,N_1635);
nand U1694 (N_1694,N_1644,N_1623);
and U1695 (N_1695,N_1669,N_1642);
nor U1696 (N_1696,N_1639,N_1659);
nand U1697 (N_1697,N_1641,N_1633);
and U1698 (N_1698,N_1646,N_1656);
nor U1699 (N_1699,N_1663,N_1625);
or U1700 (N_1700,N_1678,N_1622);
and U1701 (N_1701,N_1640,N_1629);
or U1702 (N_1702,N_1673,N_1631);
or U1703 (N_1703,N_1628,N_1636);
or U1704 (N_1704,N_1651,N_1637);
and U1705 (N_1705,N_1634,N_1667);
nand U1706 (N_1706,N_1632,N_1657);
and U1707 (N_1707,N_1670,N_1664);
or U1708 (N_1708,N_1675,N_1674);
and U1709 (N_1709,N_1662,N_1672);
nor U1710 (N_1710,N_1648,N_1629);
nor U1711 (N_1711,N_1626,N_1655);
nor U1712 (N_1712,N_1627,N_1666);
nand U1713 (N_1713,N_1669,N_1676);
and U1714 (N_1714,N_1645,N_1636);
nor U1715 (N_1715,N_1665,N_1668);
and U1716 (N_1716,N_1637,N_1669);
nor U1717 (N_1717,N_1638,N_1630);
nand U1718 (N_1718,N_1652,N_1677);
and U1719 (N_1719,N_1660,N_1670);
nor U1720 (N_1720,N_1678,N_1638);
and U1721 (N_1721,N_1628,N_1626);
or U1722 (N_1722,N_1621,N_1622);
nand U1723 (N_1723,N_1669,N_1624);
or U1724 (N_1724,N_1642,N_1645);
or U1725 (N_1725,N_1671,N_1643);
or U1726 (N_1726,N_1675,N_1665);
or U1727 (N_1727,N_1676,N_1662);
nor U1728 (N_1728,N_1675,N_1649);
nand U1729 (N_1729,N_1660,N_1659);
nand U1730 (N_1730,N_1626,N_1634);
nand U1731 (N_1731,N_1665,N_1625);
nor U1732 (N_1732,N_1663,N_1627);
or U1733 (N_1733,N_1645,N_1630);
nor U1734 (N_1734,N_1676,N_1625);
or U1735 (N_1735,N_1649,N_1633);
or U1736 (N_1736,N_1654,N_1635);
and U1737 (N_1737,N_1634,N_1657);
and U1738 (N_1738,N_1675,N_1667);
or U1739 (N_1739,N_1641,N_1624);
nand U1740 (N_1740,N_1725,N_1737);
nor U1741 (N_1741,N_1731,N_1712);
and U1742 (N_1742,N_1710,N_1701);
nor U1743 (N_1743,N_1684,N_1717);
nand U1744 (N_1744,N_1708,N_1735);
or U1745 (N_1745,N_1723,N_1682);
nand U1746 (N_1746,N_1702,N_1730);
nand U1747 (N_1747,N_1729,N_1700);
nor U1748 (N_1748,N_1722,N_1706);
nand U1749 (N_1749,N_1709,N_1715);
and U1750 (N_1750,N_1685,N_1719);
or U1751 (N_1751,N_1698,N_1724);
xor U1752 (N_1752,N_1694,N_1697);
nor U1753 (N_1753,N_1705,N_1681);
and U1754 (N_1754,N_1707,N_1732);
nor U1755 (N_1755,N_1695,N_1728);
and U1756 (N_1756,N_1716,N_1683);
nand U1757 (N_1757,N_1690,N_1711);
and U1758 (N_1758,N_1680,N_1721);
nand U1759 (N_1759,N_1738,N_1696);
or U1760 (N_1760,N_1691,N_1688);
nor U1761 (N_1761,N_1704,N_1699);
nand U1762 (N_1762,N_1692,N_1686);
nor U1763 (N_1763,N_1733,N_1693);
and U1764 (N_1764,N_1727,N_1736);
nor U1765 (N_1765,N_1689,N_1720);
and U1766 (N_1766,N_1726,N_1739);
and U1767 (N_1767,N_1714,N_1703);
nor U1768 (N_1768,N_1713,N_1687);
nand U1769 (N_1769,N_1718,N_1734);
or U1770 (N_1770,N_1688,N_1708);
nor U1771 (N_1771,N_1723,N_1716);
nand U1772 (N_1772,N_1736,N_1703);
or U1773 (N_1773,N_1713,N_1699);
nand U1774 (N_1774,N_1690,N_1705);
or U1775 (N_1775,N_1706,N_1693);
or U1776 (N_1776,N_1689,N_1732);
and U1777 (N_1777,N_1706,N_1737);
nor U1778 (N_1778,N_1698,N_1702);
or U1779 (N_1779,N_1698,N_1731);
nor U1780 (N_1780,N_1724,N_1733);
nand U1781 (N_1781,N_1695,N_1713);
or U1782 (N_1782,N_1708,N_1723);
or U1783 (N_1783,N_1731,N_1728);
xor U1784 (N_1784,N_1724,N_1709);
and U1785 (N_1785,N_1683,N_1696);
nand U1786 (N_1786,N_1687,N_1691);
nand U1787 (N_1787,N_1723,N_1712);
or U1788 (N_1788,N_1689,N_1723);
nand U1789 (N_1789,N_1724,N_1708);
and U1790 (N_1790,N_1687,N_1726);
nor U1791 (N_1791,N_1722,N_1705);
and U1792 (N_1792,N_1730,N_1690);
nand U1793 (N_1793,N_1713,N_1688);
nand U1794 (N_1794,N_1731,N_1696);
and U1795 (N_1795,N_1719,N_1714);
or U1796 (N_1796,N_1709,N_1704);
or U1797 (N_1797,N_1706,N_1681);
nand U1798 (N_1798,N_1685,N_1695);
or U1799 (N_1799,N_1726,N_1722);
nand U1800 (N_1800,N_1775,N_1751);
or U1801 (N_1801,N_1772,N_1766);
and U1802 (N_1802,N_1770,N_1793);
nor U1803 (N_1803,N_1782,N_1758);
nand U1804 (N_1804,N_1745,N_1746);
xor U1805 (N_1805,N_1774,N_1750);
nand U1806 (N_1806,N_1794,N_1767);
or U1807 (N_1807,N_1743,N_1762);
or U1808 (N_1808,N_1779,N_1796);
and U1809 (N_1809,N_1777,N_1753);
nand U1810 (N_1810,N_1754,N_1756);
nor U1811 (N_1811,N_1761,N_1744);
nor U1812 (N_1812,N_1781,N_1778);
or U1813 (N_1813,N_1760,N_1747);
nand U1814 (N_1814,N_1780,N_1769);
nand U1815 (N_1815,N_1757,N_1786);
or U1816 (N_1816,N_1749,N_1768);
nor U1817 (N_1817,N_1773,N_1787);
and U1818 (N_1818,N_1752,N_1759);
or U1819 (N_1819,N_1790,N_1797);
nor U1820 (N_1820,N_1798,N_1792);
nor U1821 (N_1821,N_1789,N_1742);
nand U1822 (N_1822,N_1799,N_1755);
nand U1823 (N_1823,N_1741,N_1791);
nor U1824 (N_1824,N_1763,N_1748);
nand U1825 (N_1825,N_1783,N_1795);
nand U1826 (N_1826,N_1776,N_1740);
nand U1827 (N_1827,N_1788,N_1771);
and U1828 (N_1828,N_1764,N_1784);
nand U1829 (N_1829,N_1765,N_1785);
nor U1830 (N_1830,N_1748,N_1791);
or U1831 (N_1831,N_1773,N_1772);
nor U1832 (N_1832,N_1767,N_1748);
or U1833 (N_1833,N_1774,N_1779);
or U1834 (N_1834,N_1748,N_1783);
and U1835 (N_1835,N_1772,N_1748);
nand U1836 (N_1836,N_1791,N_1788);
nand U1837 (N_1837,N_1760,N_1741);
nand U1838 (N_1838,N_1742,N_1766);
or U1839 (N_1839,N_1797,N_1767);
nor U1840 (N_1840,N_1778,N_1786);
nor U1841 (N_1841,N_1772,N_1741);
nor U1842 (N_1842,N_1768,N_1792);
or U1843 (N_1843,N_1776,N_1757);
and U1844 (N_1844,N_1770,N_1769);
nor U1845 (N_1845,N_1768,N_1772);
and U1846 (N_1846,N_1792,N_1787);
nor U1847 (N_1847,N_1744,N_1743);
nand U1848 (N_1848,N_1798,N_1757);
or U1849 (N_1849,N_1752,N_1742);
and U1850 (N_1850,N_1780,N_1772);
and U1851 (N_1851,N_1777,N_1791);
nand U1852 (N_1852,N_1760,N_1793);
or U1853 (N_1853,N_1785,N_1793);
nor U1854 (N_1854,N_1792,N_1746);
or U1855 (N_1855,N_1786,N_1792);
nand U1856 (N_1856,N_1768,N_1752);
and U1857 (N_1857,N_1743,N_1740);
and U1858 (N_1858,N_1741,N_1781);
nor U1859 (N_1859,N_1795,N_1788);
nand U1860 (N_1860,N_1850,N_1838);
and U1861 (N_1861,N_1818,N_1847);
and U1862 (N_1862,N_1851,N_1812);
or U1863 (N_1863,N_1811,N_1805);
or U1864 (N_1864,N_1841,N_1854);
nor U1865 (N_1865,N_1857,N_1848);
nand U1866 (N_1866,N_1833,N_1837);
nor U1867 (N_1867,N_1843,N_1813);
or U1868 (N_1868,N_1802,N_1806);
nand U1869 (N_1869,N_1803,N_1824);
nand U1870 (N_1870,N_1817,N_1821);
or U1871 (N_1871,N_1820,N_1822);
and U1872 (N_1872,N_1836,N_1800);
or U1873 (N_1873,N_1830,N_1825);
and U1874 (N_1874,N_1829,N_1809);
nand U1875 (N_1875,N_1858,N_1859);
nor U1876 (N_1876,N_1846,N_1807);
nor U1877 (N_1877,N_1834,N_1855);
nand U1878 (N_1878,N_1845,N_1853);
or U1879 (N_1879,N_1842,N_1828);
and U1880 (N_1880,N_1835,N_1815);
or U1881 (N_1881,N_1856,N_1844);
and U1882 (N_1882,N_1827,N_1826);
nor U1883 (N_1883,N_1831,N_1816);
nand U1884 (N_1884,N_1810,N_1852);
nor U1885 (N_1885,N_1832,N_1804);
nor U1886 (N_1886,N_1808,N_1814);
nor U1887 (N_1887,N_1823,N_1840);
or U1888 (N_1888,N_1849,N_1819);
nand U1889 (N_1889,N_1839,N_1801);
nor U1890 (N_1890,N_1822,N_1805);
and U1891 (N_1891,N_1842,N_1830);
nor U1892 (N_1892,N_1856,N_1842);
or U1893 (N_1893,N_1826,N_1848);
or U1894 (N_1894,N_1831,N_1815);
nand U1895 (N_1895,N_1806,N_1836);
or U1896 (N_1896,N_1836,N_1804);
nand U1897 (N_1897,N_1819,N_1814);
nor U1898 (N_1898,N_1850,N_1802);
nor U1899 (N_1899,N_1839,N_1847);
and U1900 (N_1900,N_1806,N_1835);
nor U1901 (N_1901,N_1806,N_1831);
and U1902 (N_1902,N_1832,N_1825);
or U1903 (N_1903,N_1830,N_1852);
nand U1904 (N_1904,N_1827,N_1855);
or U1905 (N_1905,N_1843,N_1859);
or U1906 (N_1906,N_1856,N_1823);
nand U1907 (N_1907,N_1802,N_1836);
nand U1908 (N_1908,N_1857,N_1850);
or U1909 (N_1909,N_1844,N_1800);
nand U1910 (N_1910,N_1832,N_1803);
or U1911 (N_1911,N_1842,N_1841);
and U1912 (N_1912,N_1840,N_1813);
or U1913 (N_1913,N_1853,N_1857);
nand U1914 (N_1914,N_1835,N_1832);
nor U1915 (N_1915,N_1806,N_1843);
nor U1916 (N_1916,N_1818,N_1821);
or U1917 (N_1917,N_1848,N_1805);
and U1918 (N_1918,N_1835,N_1854);
or U1919 (N_1919,N_1834,N_1824);
or U1920 (N_1920,N_1876,N_1906);
nand U1921 (N_1921,N_1910,N_1889);
or U1922 (N_1922,N_1900,N_1918);
nand U1923 (N_1923,N_1885,N_1916);
nor U1924 (N_1924,N_1899,N_1898);
nor U1925 (N_1925,N_1877,N_1911);
and U1926 (N_1926,N_1873,N_1867);
nor U1927 (N_1927,N_1888,N_1871);
or U1928 (N_1928,N_1896,N_1872);
xor U1929 (N_1929,N_1860,N_1866);
or U1930 (N_1930,N_1882,N_1892);
and U1931 (N_1931,N_1903,N_1878);
nand U1932 (N_1932,N_1905,N_1879);
nor U1933 (N_1933,N_1880,N_1890);
or U1934 (N_1934,N_1875,N_1915);
nand U1935 (N_1935,N_1904,N_1907);
and U1936 (N_1936,N_1864,N_1874);
nor U1937 (N_1937,N_1919,N_1901);
or U1938 (N_1938,N_1886,N_1893);
nand U1939 (N_1939,N_1865,N_1913);
and U1940 (N_1940,N_1884,N_1914);
nand U1941 (N_1941,N_1870,N_1891);
and U1942 (N_1942,N_1902,N_1883);
or U1943 (N_1943,N_1887,N_1881);
and U1944 (N_1944,N_1897,N_1908);
or U1945 (N_1945,N_1894,N_1861);
nor U1946 (N_1946,N_1917,N_1912);
and U1947 (N_1947,N_1863,N_1895);
or U1948 (N_1948,N_1869,N_1862);
or U1949 (N_1949,N_1868,N_1909);
nand U1950 (N_1950,N_1913,N_1863);
nor U1951 (N_1951,N_1902,N_1898);
and U1952 (N_1952,N_1883,N_1877);
and U1953 (N_1953,N_1884,N_1904);
nor U1954 (N_1954,N_1882,N_1908);
nor U1955 (N_1955,N_1862,N_1909);
or U1956 (N_1956,N_1908,N_1919);
nand U1957 (N_1957,N_1905,N_1916);
nand U1958 (N_1958,N_1895,N_1878);
or U1959 (N_1959,N_1889,N_1919);
nand U1960 (N_1960,N_1905,N_1887);
nor U1961 (N_1961,N_1896,N_1862);
nor U1962 (N_1962,N_1879,N_1910);
nor U1963 (N_1963,N_1863,N_1910);
nor U1964 (N_1964,N_1891,N_1910);
xnor U1965 (N_1965,N_1870,N_1893);
nand U1966 (N_1966,N_1863,N_1879);
and U1967 (N_1967,N_1883,N_1919);
or U1968 (N_1968,N_1918,N_1893);
nor U1969 (N_1969,N_1876,N_1885);
or U1970 (N_1970,N_1864,N_1900);
nor U1971 (N_1971,N_1895,N_1873);
or U1972 (N_1972,N_1899,N_1901);
and U1973 (N_1973,N_1874,N_1877);
and U1974 (N_1974,N_1894,N_1904);
nor U1975 (N_1975,N_1915,N_1919);
nor U1976 (N_1976,N_1860,N_1905);
nand U1977 (N_1977,N_1876,N_1908);
xnor U1978 (N_1978,N_1869,N_1864);
nand U1979 (N_1979,N_1915,N_1892);
nand U1980 (N_1980,N_1945,N_1964);
nand U1981 (N_1981,N_1950,N_1922);
or U1982 (N_1982,N_1961,N_1973);
nor U1983 (N_1983,N_1966,N_1977);
xnor U1984 (N_1984,N_1942,N_1954);
nand U1985 (N_1985,N_1970,N_1946);
nor U1986 (N_1986,N_1928,N_1941);
nor U1987 (N_1987,N_1971,N_1960);
or U1988 (N_1988,N_1931,N_1929);
nand U1989 (N_1989,N_1924,N_1920);
or U1990 (N_1990,N_1959,N_1978);
and U1991 (N_1991,N_1965,N_1934);
nor U1992 (N_1992,N_1940,N_1939);
xor U1993 (N_1993,N_1948,N_1962);
and U1994 (N_1994,N_1937,N_1963);
nor U1995 (N_1995,N_1951,N_1925);
nand U1996 (N_1996,N_1975,N_1974);
nor U1997 (N_1997,N_1953,N_1926);
xor U1998 (N_1998,N_1927,N_1923);
xnor U1999 (N_1999,N_1955,N_1932);
or U2000 (N_2000,N_1952,N_1944);
or U2001 (N_2001,N_1935,N_1949);
nand U2002 (N_2002,N_1972,N_1969);
or U2003 (N_2003,N_1947,N_1976);
and U2004 (N_2004,N_1930,N_1968);
nor U2005 (N_2005,N_1979,N_1958);
and U2006 (N_2006,N_1956,N_1938);
nand U2007 (N_2007,N_1921,N_1943);
or U2008 (N_2008,N_1967,N_1957);
nor U2009 (N_2009,N_1936,N_1933);
and U2010 (N_2010,N_1959,N_1956);
and U2011 (N_2011,N_1939,N_1971);
and U2012 (N_2012,N_1977,N_1961);
and U2013 (N_2013,N_1967,N_1979);
nand U2014 (N_2014,N_1945,N_1939);
nor U2015 (N_2015,N_1930,N_1950);
or U2016 (N_2016,N_1924,N_1937);
nor U2017 (N_2017,N_1931,N_1947);
and U2018 (N_2018,N_1967,N_1975);
or U2019 (N_2019,N_1926,N_1923);
nor U2020 (N_2020,N_1964,N_1957);
nor U2021 (N_2021,N_1934,N_1948);
nand U2022 (N_2022,N_1927,N_1922);
or U2023 (N_2023,N_1951,N_1922);
nand U2024 (N_2024,N_1937,N_1945);
nand U2025 (N_2025,N_1942,N_1950);
nor U2026 (N_2026,N_1952,N_1923);
or U2027 (N_2027,N_1967,N_1936);
or U2028 (N_2028,N_1936,N_1970);
or U2029 (N_2029,N_1961,N_1958);
or U2030 (N_2030,N_1937,N_1943);
nor U2031 (N_2031,N_1931,N_1969);
nor U2032 (N_2032,N_1960,N_1977);
nor U2033 (N_2033,N_1969,N_1927);
nor U2034 (N_2034,N_1944,N_1945);
nor U2035 (N_2035,N_1921,N_1949);
and U2036 (N_2036,N_1967,N_1942);
or U2037 (N_2037,N_1962,N_1936);
nor U2038 (N_2038,N_1979,N_1977);
nand U2039 (N_2039,N_1924,N_1965);
or U2040 (N_2040,N_2027,N_1988);
nand U2041 (N_2041,N_2010,N_2034);
nor U2042 (N_2042,N_2015,N_2030);
and U2043 (N_2043,N_2004,N_2000);
nand U2044 (N_2044,N_2038,N_1996);
and U2045 (N_2045,N_2029,N_1984);
nand U2046 (N_2046,N_1998,N_1990);
nand U2047 (N_2047,N_1997,N_2017);
and U2048 (N_2048,N_2009,N_1991);
nor U2049 (N_2049,N_2023,N_1987);
nand U2050 (N_2050,N_2008,N_2003);
and U2051 (N_2051,N_2037,N_2033);
nor U2052 (N_2052,N_2025,N_1985);
nand U2053 (N_2053,N_2007,N_1999);
nand U2054 (N_2054,N_1995,N_2026);
nand U2055 (N_2055,N_1980,N_2031);
nor U2056 (N_2056,N_2036,N_1981);
nand U2057 (N_2057,N_2018,N_1989);
or U2058 (N_2058,N_2019,N_2016);
nor U2059 (N_2059,N_2002,N_2028);
nand U2060 (N_2060,N_2024,N_1983);
nor U2061 (N_2061,N_1992,N_2039);
or U2062 (N_2062,N_2014,N_2006);
and U2063 (N_2063,N_2022,N_1994);
and U2064 (N_2064,N_2035,N_2020);
and U2065 (N_2065,N_2021,N_2011);
nand U2066 (N_2066,N_2001,N_2005);
nor U2067 (N_2067,N_1993,N_2032);
nor U2068 (N_2068,N_2013,N_1982);
nor U2069 (N_2069,N_2012,N_1986);
nand U2070 (N_2070,N_2001,N_1991);
and U2071 (N_2071,N_2011,N_2028);
and U2072 (N_2072,N_2021,N_2019);
and U2073 (N_2073,N_1982,N_1985);
nand U2074 (N_2074,N_2010,N_2026);
and U2075 (N_2075,N_1994,N_2018);
nand U2076 (N_2076,N_2036,N_2011);
nor U2077 (N_2077,N_2000,N_2024);
and U2078 (N_2078,N_2007,N_2006);
nand U2079 (N_2079,N_1991,N_1986);
nand U2080 (N_2080,N_2006,N_2035);
nand U2081 (N_2081,N_2009,N_1995);
or U2082 (N_2082,N_2008,N_1999);
and U2083 (N_2083,N_2029,N_1991);
or U2084 (N_2084,N_1983,N_2037);
and U2085 (N_2085,N_2000,N_2029);
nor U2086 (N_2086,N_2030,N_2026);
or U2087 (N_2087,N_1984,N_1994);
and U2088 (N_2088,N_1986,N_2020);
and U2089 (N_2089,N_2021,N_2016);
nor U2090 (N_2090,N_2033,N_2027);
or U2091 (N_2091,N_2004,N_1990);
and U2092 (N_2092,N_1994,N_2002);
nor U2093 (N_2093,N_2037,N_2029);
nand U2094 (N_2094,N_1994,N_1983);
and U2095 (N_2095,N_2005,N_2009);
nand U2096 (N_2096,N_2025,N_2014);
nor U2097 (N_2097,N_2034,N_2005);
or U2098 (N_2098,N_2001,N_2021);
or U2099 (N_2099,N_2004,N_2017);
and U2100 (N_2100,N_2055,N_2069);
nor U2101 (N_2101,N_2071,N_2092);
and U2102 (N_2102,N_2046,N_2098);
or U2103 (N_2103,N_2045,N_2057);
and U2104 (N_2104,N_2064,N_2070);
and U2105 (N_2105,N_2050,N_2075);
and U2106 (N_2106,N_2094,N_2084);
or U2107 (N_2107,N_2068,N_2076);
or U2108 (N_2108,N_2072,N_2052);
nand U2109 (N_2109,N_2082,N_2062);
and U2110 (N_2110,N_2051,N_2044);
nand U2111 (N_2111,N_2083,N_2088);
nor U2112 (N_2112,N_2043,N_2079);
nand U2113 (N_2113,N_2065,N_2060);
nor U2114 (N_2114,N_2091,N_2087);
or U2115 (N_2115,N_2056,N_2063);
nand U2116 (N_2116,N_2049,N_2061);
and U2117 (N_2117,N_2080,N_2048);
nand U2118 (N_2118,N_2096,N_2099);
or U2119 (N_2119,N_2089,N_2097);
or U2120 (N_2120,N_2067,N_2042);
or U2121 (N_2121,N_2078,N_2058);
nand U2122 (N_2122,N_2090,N_2059);
and U2123 (N_2123,N_2077,N_2053);
and U2124 (N_2124,N_2040,N_2047);
nand U2125 (N_2125,N_2041,N_2066);
nor U2126 (N_2126,N_2095,N_2093);
nor U2127 (N_2127,N_2086,N_2085);
or U2128 (N_2128,N_2073,N_2054);
or U2129 (N_2129,N_2074,N_2081);
or U2130 (N_2130,N_2073,N_2098);
and U2131 (N_2131,N_2055,N_2064);
and U2132 (N_2132,N_2073,N_2082);
nand U2133 (N_2133,N_2049,N_2040);
or U2134 (N_2134,N_2090,N_2086);
and U2135 (N_2135,N_2064,N_2062);
nand U2136 (N_2136,N_2046,N_2069);
nand U2137 (N_2137,N_2045,N_2054);
and U2138 (N_2138,N_2094,N_2065);
nand U2139 (N_2139,N_2063,N_2048);
nand U2140 (N_2140,N_2067,N_2075);
nor U2141 (N_2141,N_2084,N_2088);
and U2142 (N_2142,N_2043,N_2051);
xnor U2143 (N_2143,N_2062,N_2087);
and U2144 (N_2144,N_2064,N_2052);
nor U2145 (N_2145,N_2080,N_2096);
nor U2146 (N_2146,N_2047,N_2064);
and U2147 (N_2147,N_2071,N_2069);
and U2148 (N_2148,N_2076,N_2070);
nor U2149 (N_2149,N_2077,N_2089);
or U2150 (N_2150,N_2055,N_2058);
nor U2151 (N_2151,N_2041,N_2095);
nor U2152 (N_2152,N_2081,N_2057);
and U2153 (N_2153,N_2072,N_2068);
nand U2154 (N_2154,N_2043,N_2094);
nand U2155 (N_2155,N_2061,N_2073);
nor U2156 (N_2156,N_2072,N_2050);
and U2157 (N_2157,N_2089,N_2047);
nand U2158 (N_2158,N_2085,N_2076);
nor U2159 (N_2159,N_2044,N_2056);
nand U2160 (N_2160,N_2122,N_2100);
nor U2161 (N_2161,N_2101,N_2113);
and U2162 (N_2162,N_2108,N_2128);
nand U2163 (N_2163,N_2156,N_2118);
and U2164 (N_2164,N_2143,N_2149);
nand U2165 (N_2165,N_2102,N_2151);
nor U2166 (N_2166,N_2157,N_2145);
or U2167 (N_2167,N_2130,N_2114);
or U2168 (N_2168,N_2139,N_2159);
or U2169 (N_2169,N_2129,N_2115);
nand U2170 (N_2170,N_2125,N_2110);
or U2171 (N_2171,N_2124,N_2116);
nand U2172 (N_2172,N_2133,N_2137);
nor U2173 (N_2173,N_2105,N_2111);
nand U2174 (N_2174,N_2123,N_2140);
and U2175 (N_2175,N_2150,N_2126);
nor U2176 (N_2176,N_2144,N_2147);
and U2177 (N_2177,N_2136,N_2104);
nor U2178 (N_2178,N_2134,N_2132);
nand U2179 (N_2179,N_2127,N_2142);
or U2180 (N_2180,N_2153,N_2146);
or U2181 (N_2181,N_2155,N_2154);
and U2182 (N_2182,N_2106,N_2107);
nor U2183 (N_2183,N_2109,N_2119);
or U2184 (N_2184,N_2138,N_2131);
nor U2185 (N_2185,N_2121,N_2120);
nor U2186 (N_2186,N_2148,N_2152);
or U2187 (N_2187,N_2117,N_2112);
nor U2188 (N_2188,N_2158,N_2135);
and U2189 (N_2189,N_2103,N_2141);
nand U2190 (N_2190,N_2112,N_2106);
or U2191 (N_2191,N_2151,N_2129);
nand U2192 (N_2192,N_2116,N_2133);
nand U2193 (N_2193,N_2107,N_2100);
or U2194 (N_2194,N_2157,N_2137);
nand U2195 (N_2195,N_2142,N_2110);
nand U2196 (N_2196,N_2145,N_2112);
or U2197 (N_2197,N_2119,N_2156);
nor U2198 (N_2198,N_2101,N_2127);
or U2199 (N_2199,N_2155,N_2158);
or U2200 (N_2200,N_2127,N_2114);
nand U2201 (N_2201,N_2145,N_2102);
or U2202 (N_2202,N_2134,N_2121);
or U2203 (N_2203,N_2129,N_2139);
or U2204 (N_2204,N_2113,N_2156);
or U2205 (N_2205,N_2133,N_2156);
nand U2206 (N_2206,N_2145,N_2153);
or U2207 (N_2207,N_2129,N_2147);
nor U2208 (N_2208,N_2137,N_2108);
and U2209 (N_2209,N_2128,N_2139);
or U2210 (N_2210,N_2157,N_2127);
or U2211 (N_2211,N_2149,N_2144);
or U2212 (N_2212,N_2129,N_2145);
nand U2213 (N_2213,N_2140,N_2111);
nand U2214 (N_2214,N_2154,N_2128);
or U2215 (N_2215,N_2119,N_2143);
nand U2216 (N_2216,N_2122,N_2133);
and U2217 (N_2217,N_2143,N_2145);
nor U2218 (N_2218,N_2121,N_2109);
nand U2219 (N_2219,N_2101,N_2133);
nand U2220 (N_2220,N_2195,N_2187);
or U2221 (N_2221,N_2215,N_2180);
xor U2222 (N_2222,N_2204,N_2209);
nand U2223 (N_2223,N_2217,N_2190);
nand U2224 (N_2224,N_2202,N_2166);
and U2225 (N_2225,N_2175,N_2201);
nor U2226 (N_2226,N_2206,N_2198);
or U2227 (N_2227,N_2199,N_2218);
and U2228 (N_2228,N_2167,N_2181);
and U2229 (N_2229,N_2210,N_2219);
nand U2230 (N_2230,N_2212,N_2192);
nor U2231 (N_2231,N_2184,N_2205);
nand U2232 (N_2232,N_2168,N_2213);
nand U2233 (N_2233,N_2162,N_2207);
or U2234 (N_2234,N_2188,N_2165);
nand U2235 (N_2235,N_2176,N_2214);
nor U2236 (N_2236,N_2182,N_2185);
nand U2237 (N_2237,N_2203,N_2186);
or U2238 (N_2238,N_2171,N_2208);
nand U2239 (N_2239,N_2163,N_2189);
or U2240 (N_2240,N_2216,N_2160);
nand U2241 (N_2241,N_2169,N_2161);
or U2242 (N_2242,N_2200,N_2172);
nor U2243 (N_2243,N_2183,N_2193);
and U2244 (N_2244,N_2211,N_2179);
nand U2245 (N_2245,N_2194,N_2173);
or U2246 (N_2246,N_2174,N_2170);
or U2247 (N_2247,N_2191,N_2196);
and U2248 (N_2248,N_2197,N_2164);
nand U2249 (N_2249,N_2177,N_2178);
and U2250 (N_2250,N_2175,N_2210);
nor U2251 (N_2251,N_2163,N_2175);
nand U2252 (N_2252,N_2201,N_2161);
and U2253 (N_2253,N_2180,N_2200);
or U2254 (N_2254,N_2202,N_2187);
nor U2255 (N_2255,N_2164,N_2174);
or U2256 (N_2256,N_2163,N_2212);
nand U2257 (N_2257,N_2162,N_2180);
nand U2258 (N_2258,N_2190,N_2167);
nor U2259 (N_2259,N_2215,N_2173);
or U2260 (N_2260,N_2171,N_2209);
or U2261 (N_2261,N_2186,N_2161);
nand U2262 (N_2262,N_2168,N_2204);
nand U2263 (N_2263,N_2204,N_2171);
and U2264 (N_2264,N_2192,N_2194);
nand U2265 (N_2265,N_2212,N_2197);
nand U2266 (N_2266,N_2165,N_2178);
and U2267 (N_2267,N_2213,N_2202);
or U2268 (N_2268,N_2217,N_2169);
nand U2269 (N_2269,N_2160,N_2211);
and U2270 (N_2270,N_2198,N_2212);
nor U2271 (N_2271,N_2212,N_2217);
nand U2272 (N_2272,N_2207,N_2160);
nand U2273 (N_2273,N_2212,N_2176);
nand U2274 (N_2274,N_2172,N_2208);
and U2275 (N_2275,N_2203,N_2180);
or U2276 (N_2276,N_2194,N_2179);
nand U2277 (N_2277,N_2197,N_2170);
nor U2278 (N_2278,N_2205,N_2162);
nand U2279 (N_2279,N_2218,N_2169);
nor U2280 (N_2280,N_2273,N_2266);
and U2281 (N_2281,N_2222,N_2248);
nand U2282 (N_2282,N_2252,N_2240);
nand U2283 (N_2283,N_2267,N_2227);
nand U2284 (N_2284,N_2268,N_2251);
and U2285 (N_2285,N_2228,N_2236);
nand U2286 (N_2286,N_2243,N_2244);
or U2287 (N_2287,N_2261,N_2220);
nor U2288 (N_2288,N_2238,N_2269);
nor U2289 (N_2289,N_2242,N_2250);
or U2290 (N_2290,N_2235,N_2274);
nor U2291 (N_2291,N_2254,N_2270);
nor U2292 (N_2292,N_2279,N_2226);
nor U2293 (N_2293,N_2255,N_2231);
or U2294 (N_2294,N_2271,N_2256);
and U2295 (N_2295,N_2277,N_2265);
nor U2296 (N_2296,N_2246,N_2276);
nor U2297 (N_2297,N_2230,N_2278);
nand U2298 (N_2298,N_2258,N_2232);
or U2299 (N_2299,N_2221,N_2247);
nor U2300 (N_2300,N_2233,N_2262);
nor U2301 (N_2301,N_2241,N_2257);
nand U2302 (N_2302,N_2259,N_2272);
nand U2303 (N_2303,N_2245,N_2264);
xor U2304 (N_2304,N_2263,N_2229);
and U2305 (N_2305,N_2249,N_2225);
and U2306 (N_2306,N_2239,N_2237);
or U2307 (N_2307,N_2224,N_2260);
and U2308 (N_2308,N_2234,N_2253);
nand U2309 (N_2309,N_2223,N_2275);
and U2310 (N_2310,N_2268,N_2241);
or U2311 (N_2311,N_2253,N_2275);
nor U2312 (N_2312,N_2256,N_2253);
and U2313 (N_2313,N_2225,N_2272);
and U2314 (N_2314,N_2270,N_2258);
or U2315 (N_2315,N_2240,N_2278);
and U2316 (N_2316,N_2232,N_2244);
nor U2317 (N_2317,N_2250,N_2276);
xnor U2318 (N_2318,N_2224,N_2239);
nor U2319 (N_2319,N_2263,N_2267);
nor U2320 (N_2320,N_2257,N_2272);
and U2321 (N_2321,N_2244,N_2225);
or U2322 (N_2322,N_2243,N_2279);
or U2323 (N_2323,N_2255,N_2274);
and U2324 (N_2324,N_2260,N_2258);
and U2325 (N_2325,N_2256,N_2230);
nor U2326 (N_2326,N_2234,N_2232);
or U2327 (N_2327,N_2266,N_2229);
nand U2328 (N_2328,N_2275,N_2243);
and U2329 (N_2329,N_2274,N_2260);
nor U2330 (N_2330,N_2247,N_2243);
or U2331 (N_2331,N_2227,N_2260);
nor U2332 (N_2332,N_2266,N_2270);
or U2333 (N_2333,N_2227,N_2276);
or U2334 (N_2334,N_2254,N_2242);
or U2335 (N_2335,N_2263,N_2237);
and U2336 (N_2336,N_2238,N_2259);
and U2337 (N_2337,N_2279,N_2221);
or U2338 (N_2338,N_2265,N_2253);
and U2339 (N_2339,N_2260,N_2246);
nor U2340 (N_2340,N_2307,N_2334);
nor U2341 (N_2341,N_2309,N_2337);
or U2342 (N_2342,N_2315,N_2286);
or U2343 (N_2343,N_2339,N_2308);
nand U2344 (N_2344,N_2293,N_2291);
nor U2345 (N_2345,N_2314,N_2304);
and U2346 (N_2346,N_2284,N_2332);
nand U2347 (N_2347,N_2311,N_2300);
xor U2348 (N_2348,N_2280,N_2325);
or U2349 (N_2349,N_2320,N_2290);
or U2350 (N_2350,N_2316,N_2281);
or U2351 (N_2351,N_2330,N_2287);
nor U2352 (N_2352,N_2305,N_2323);
nor U2353 (N_2353,N_2328,N_2324);
nor U2354 (N_2354,N_2318,N_2317);
and U2355 (N_2355,N_2312,N_2333);
nor U2356 (N_2356,N_2336,N_2306);
nor U2357 (N_2357,N_2322,N_2329);
nor U2358 (N_2358,N_2335,N_2298);
and U2359 (N_2359,N_2288,N_2319);
nor U2360 (N_2360,N_2338,N_2299);
or U2361 (N_2361,N_2296,N_2282);
nand U2362 (N_2362,N_2326,N_2295);
nor U2363 (N_2363,N_2331,N_2289);
nand U2364 (N_2364,N_2310,N_2321);
nor U2365 (N_2365,N_2285,N_2292);
nor U2366 (N_2366,N_2297,N_2327);
and U2367 (N_2367,N_2302,N_2283);
and U2368 (N_2368,N_2313,N_2303);
nor U2369 (N_2369,N_2301,N_2294);
nor U2370 (N_2370,N_2313,N_2282);
or U2371 (N_2371,N_2319,N_2297);
and U2372 (N_2372,N_2313,N_2300);
nand U2373 (N_2373,N_2325,N_2286);
nor U2374 (N_2374,N_2320,N_2323);
xnor U2375 (N_2375,N_2288,N_2295);
or U2376 (N_2376,N_2315,N_2297);
nor U2377 (N_2377,N_2287,N_2305);
nor U2378 (N_2378,N_2295,N_2313);
and U2379 (N_2379,N_2283,N_2327);
nand U2380 (N_2380,N_2314,N_2281);
or U2381 (N_2381,N_2302,N_2308);
or U2382 (N_2382,N_2290,N_2339);
or U2383 (N_2383,N_2306,N_2292);
nor U2384 (N_2384,N_2337,N_2320);
or U2385 (N_2385,N_2311,N_2337);
nor U2386 (N_2386,N_2310,N_2335);
or U2387 (N_2387,N_2285,N_2321);
nand U2388 (N_2388,N_2306,N_2319);
nand U2389 (N_2389,N_2299,N_2306);
or U2390 (N_2390,N_2305,N_2310);
nor U2391 (N_2391,N_2324,N_2296);
or U2392 (N_2392,N_2281,N_2318);
or U2393 (N_2393,N_2324,N_2339);
or U2394 (N_2394,N_2338,N_2297);
and U2395 (N_2395,N_2310,N_2316);
or U2396 (N_2396,N_2300,N_2335);
nand U2397 (N_2397,N_2281,N_2304);
nor U2398 (N_2398,N_2319,N_2321);
and U2399 (N_2399,N_2291,N_2319);
or U2400 (N_2400,N_2371,N_2341);
nand U2401 (N_2401,N_2399,N_2386);
nand U2402 (N_2402,N_2388,N_2354);
or U2403 (N_2403,N_2342,N_2385);
and U2404 (N_2404,N_2396,N_2366);
or U2405 (N_2405,N_2347,N_2383);
or U2406 (N_2406,N_2370,N_2357);
nand U2407 (N_2407,N_2353,N_2346);
or U2408 (N_2408,N_2377,N_2340);
and U2409 (N_2409,N_2373,N_2369);
nor U2410 (N_2410,N_2361,N_2356);
nand U2411 (N_2411,N_2376,N_2344);
nand U2412 (N_2412,N_2363,N_2395);
nor U2413 (N_2413,N_2378,N_2390);
and U2414 (N_2414,N_2393,N_2372);
nor U2415 (N_2415,N_2382,N_2368);
or U2416 (N_2416,N_2345,N_2379);
and U2417 (N_2417,N_2398,N_2389);
and U2418 (N_2418,N_2348,N_2394);
nor U2419 (N_2419,N_2391,N_2381);
nor U2420 (N_2420,N_2397,N_2343);
nand U2421 (N_2421,N_2374,N_2365);
and U2422 (N_2422,N_2384,N_2349);
or U2423 (N_2423,N_2375,N_2359);
or U2424 (N_2424,N_2362,N_2387);
nor U2425 (N_2425,N_2355,N_2352);
nand U2426 (N_2426,N_2351,N_2380);
nand U2427 (N_2427,N_2360,N_2392);
and U2428 (N_2428,N_2350,N_2358);
and U2429 (N_2429,N_2367,N_2364);
xnor U2430 (N_2430,N_2365,N_2352);
and U2431 (N_2431,N_2349,N_2340);
nor U2432 (N_2432,N_2344,N_2359);
or U2433 (N_2433,N_2392,N_2382);
or U2434 (N_2434,N_2354,N_2385);
and U2435 (N_2435,N_2392,N_2389);
and U2436 (N_2436,N_2340,N_2351);
nand U2437 (N_2437,N_2341,N_2399);
nor U2438 (N_2438,N_2381,N_2364);
nor U2439 (N_2439,N_2349,N_2372);
nand U2440 (N_2440,N_2376,N_2355);
nor U2441 (N_2441,N_2390,N_2393);
or U2442 (N_2442,N_2352,N_2353);
or U2443 (N_2443,N_2365,N_2346);
and U2444 (N_2444,N_2376,N_2392);
or U2445 (N_2445,N_2392,N_2365);
nor U2446 (N_2446,N_2353,N_2354);
nand U2447 (N_2447,N_2382,N_2363);
and U2448 (N_2448,N_2393,N_2356);
and U2449 (N_2449,N_2347,N_2349);
nand U2450 (N_2450,N_2394,N_2381);
and U2451 (N_2451,N_2362,N_2371);
nand U2452 (N_2452,N_2380,N_2358);
nand U2453 (N_2453,N_2395,N_2360);
nor U2454 (N_2454,N_2396,N_2378);
nor U2455 (N_2455,N_2392,N_2348);
or U2456 (N_2456,N_2349,N_2367);
nor U2457 (N_2457,N_2345,N_2343);
and U2458 (N_2458,N_2378,N_2372);
and U2459 (N_2459,N_2365,N_2347);
or U2460 (N_2460,N_2405,N_2403);
or U2461 (N_2461,N_2459,N_2411);
or U2462 (N_2462,N_2451,N_2408);
nor U2463 (N_2463,N_2424,N_2418);
or U2464 (N_2464,N_2427,N_2410);
nand U2465 (N_2465,N_2428,N_2401);
and U2466 (N_2466,N_2407,N_2439);
or U2467 (N_2467,N_2448,N_2409);
or U2468 (N_2468,N_2438,N_2443);
nand U2469 (N_2469,N_2414,N_2426);
nand U2470 (N_2470,N_2421,N_2440);
or U2471 (N_2471,N_2400,N_2452);
nor U2472 (N_2472,N_2455,N_2423);
nand U2473 (N_2473,N_2447,N_2442);
and U2474 (N_2474,N_2415,N_2431);
nor U2475 (N_2475,N_2416,N_2433);
or U2476 (N_2476,N_2434,N_2445);
nand U2477 (N_2477,N_2402,N_2422);
nor U2478 (N_2478,N_2404,N_2425);
and U2479 (N_2479,N_2412,N_2449);
and U2480 (N_2480,N_2432,N_2430);
or U2481 (N_2481,N_2444,N_2446);
and U2482 (N_2482,N_2450,N_2429);
or U2483 (N_2483,N_2457,N_2436);
nor U2484 (N_2484,N_2417,N_2441);
or U2485 (N_2485,N_2437,N_2435);
or U2486 (N_2486,N_2453,N_2406);
and U2487 (N_2487,N_2456,N_2454);
and U2488 (N_2488,N_2458,N_2419);
and U2489 (N_2489,N_2420,N_2413);
nor U2490 (N_2490,N_2427,N_2430);
nor U2491 (N_2491,N_2456,N_2443);
or U2492 (N_2492,N_2446,N_2447);
nor U2493 (N_2493,N_2453,N_2422);
nor U2494 (N_2494,N_2432,N_2458);
or U2495 (N_2495,N_2422,N_2448);
nor U2496 (N_2496,N_2401,N_2423);
or U2497 (N_2497,N_2437,N_2423);
nor U2498 (N_2498,N_2431,N_2401);
nor U2499 (N_2499,N_2455,N_2450);
nor U2500 (N_2500,N_2441,N_2432);
nor U2501 (N_2501,N_2420,N_2438);
nand U2502 (N_2502,N_2435,N_2431);
nand U2503 (N_2503,N_2407,N_2421);
nor U2504 (N_2504,N_2401,N_2405);
or U2505 (N_2505,N_2456,N_2403);
or U2506 (N_2506,N_2410,N_2455);
nor U2507 (N_2507,N_2457,N_2424);
or U2508 (N_2508,N_2406,N_2457);
and U2509 (N_2509,N_2441,N_2413);
or U2510 (N_2510,N_2434,N_2401);
or U2511 (N_2511,N_2440,N_2452);
or U2512 (N_2512,N_2443,N_2433);
nor U2513 (N_2513,N_2430,N_2453);
nor U2514 (N_2514,N_2434,N_2431);
nand U2515 (N_2515,N_2433,N_2410);
or U2516 (N_2516,N_2429,N_2423);
or U2517 (N_2517,N_2427,N_2451);
nand U2518 (N_2518,N_2412,N_2402);
nor U2519 (N_2519,N_2457,N_2421);
nand U2520 (N_2520,N_2496,N_2464);
or U2521 (N_2521,N_2506,N_2481);
and U2522 (N_2522,N_2517,N_2482);
nand U2523 (N_2523,N_2507,N_2461);
or U2524 (N_2524,N_2490,N_2492);
or U2525 (N_2525,N_2474,N_2487);
nor U2526 (N_2526,N_2493,N_2484);
nor U2527 (N_2527,N_2472,N_2498);
nand U2528 (N_2528,N_2518,N_2516);
nor U2529 (N_2529,N_2480,N_2502);
or U2530 (N_2530,N_2514,N_2500);
nor U2531 (N_2531,N_2491,N_2477);
nand U2532 (N_2532,N_2489,N_2497);
nor U2533 (N_2533,N_2468,N_2504);
or U2534 (N_2534,N_2488,N_2505);
and U2535 (N_2535,N_2503,N_2478);
nand U2536 (N_2536,N_2467,N_2469);
nor U2537 (N_2537,N_2463,N_2470);
nor U2538 (N_2538,N_2495,N_2509);
nor U2539 (N_2539,N_2519,N_2511);
nor U2540 (N_2540,N_2486,N_2475);
and U2541 (N_2541,N_2510,N_2515);
nand U2542 (N_2542,N_2462,N_2485);
or U2543 (N_2543,N_2471,N_2460);
or U2544 (N_2544,N_2494,N_2512);
nand U2545 (N_2545,N_2473,N_2499);
or U2546 (N_2546,N_2508,N_2483);
and U2547 (N_2547,N_2466,N_2465);
or U2548 (N_2548,N_2513,N_2476);
and U2549 (N_2549,N_2501,N_2479);
or U2550 (N_2550,N_2490,N_2480);
nand U2551 (N_2551,N_2495,N_2499);
nand U2552 (N_2552,N_2490,N_2500);
nor U2553 (N_2553,N_2463,N_2460);
and U2554 (N_2554,N_2501,N_2514);
nand U2555 (N_2555,N_2481,N_2476);
nand U2556 (N_2556,N_2473,N_2477);
and U2557 (N_2557,N_2510,N_2502);
and U2558 (N_2558,N_2516,N_2488);
nand U2559 (N_2559,N_2517,N_2503);
nand U2560 (N_2560,N_2519,N_2485);
or U2561 (N_2561,N_2515,N_2504);
or U2562 (N_2562,N_2479,N_2518);
and U2563 (N_2563,N_2500,N_2508);
or U2564 (N_2564,N_2483,N_2515);
nor U2565 (N_2565,N_2475,N_2479);
and U2566 (N_2566,N_2504,N_2481);
nand U2567 (N_2567,N_2479,N_2466);
nand U2568 (N_2568,N_2518,N_2491);
nor U2569 (N_2569,N_2500,N_2489);
and U2570 (N_2570,N_2510,N_2506);
and U2571 (N_2571,N_2489,N_2510);
or U2572 (N_2572,N_2492,N_2501);
or U2573 (N_2573,N_2497,N_2468);
and U2574 (N_2574,N_2475,N_2465);
nand U2575 (N_2575,N_2510,N_2467);
nand U2576 (N_2576,N_2505,N_2513);
and U2577 (N_2577,N_2484,N_2512);
or U2578 (N_2578,N_2505,N_2464);
nand U2579 (N_2579,N_2508,N_2507);
and U2580 (N_2580,N_2568,N_2558);
and U2581 (N_2581,N_2536,N_2526);
nor U2582 (N_2582,N_2560,N_2578);
nand U2583 (N_2583,N_2566,N_2554);
nor U2584 (N_2584,N_2557,N_2531);
or U2585 (N_2585,N_2547,N_2553);
and U2586 (N_2586,N_2540,N_2532);
nand U2587 (N_2587,N_2535,N_2570);
and U2588 (N_2588,N_2575,N_2572);
or U2589 (N_2589,N_2524,N_2521);
or U2590 (N_2590,N_2574,N_2565);
or U2591 (N_2591,N_2520,N_2556);
nand U2592 (N_2592,N_2528,N_2530);
nor U2593 (N_2593,N_2525,N_2569);
or U2594 (N_2594,N_2523,N_2573);
or U2595 (N_2595,N_2522,N_2539);
nor U2596 (N_2596,N_2563,N_2544);
nor U2597 (N_2597,N_2579,N_2552);
nor U2598 (N_2598,N_2533,N_2541);
or U2599 (N_2599,N_2550,N_2576);
nand U2600 (N_2600,N_2561,N_2546);
nor U2601 (N_2601,N_2543,N_2548);
nand U2602 (N_2602,N_2551,N_2564);
or U2603 (N_2603,N_2534,N_2555);
and U2604 (N_2604,N_2538,N_2545);
and U2605 (N_2605,N_2537,N_2571);
nand U2606 (N_2606,N_2562,N_2577);
nand U2607 (N_2607,N_2549,N_2559);
nand U2608 (N_2608,N_2527,N_2542);
nand U2609 (N_2609,N_2529,N_2567);
and U2610 (N_2610,N_2529,N_2527);
and U2611 (N_2611,N_2554,N_2532);
and U2612 (N_2612,N_2560,N_2564);
nand U2613 (N_2613,N_2530,N_2523);
nor U2614 (N_2614,N_2576,N_2568);
nor U2615 (N_2615,N_2559,N_2529);
nor U2616 (N_2616,N_2520,N_2549);
or U2617 (N_2617,N_2575,N_2564);
and U2618 (N_2618,N_2575,N_2561);
nand U2619 (N_2619,N_2555,N_2526);
nand U2620 (N_2620,N_2521,N_2552);
or U2621 (N_2621,N_2565,N_2528);
and U2622 (N_2622,N_2551,N_2537);
and U2623 (N_2623,N_2552,N_2577);
nor U2624 (N_2624,N_2574,N_2550);
and U2625 (N_2625,N_2541,N_2572);
nand U2626 (N_2626,N_2525,N_2557);
nand U2627 (N_2627,N_2556,N_2576);
or U2628 (N_2628,N_2528,N_2538);
nand U2629 (N_2629,N_2552,N_2526);
and U2630 (N_2630,N_2579,N_2557);
nand U2631 (N_2631,N_2555,N_2543);
or U2632 (N_2632,N_2530,N_2578);
nand U2633 (N_2633,N_2556,N_2560);
nor U2634 (N_2634,N_2535,N_2556);
nand U2635 (N_2635,N_2572,N_2542);
and U2636 (N_2636,N_2550,N_2569);
nor U2637 (N_2637,N_2555,N_2528);
nor U2638 (N_2638,N_2526,N_2537);
or U2639 (N_2639,N_2559,N_2535);
and U2640 (N_2640,N_2639,N_2594);
and U2641 (N_2641,N_2596,N_2632);
and U2642 (N_2642,N_2623,N_2618);
and U2643 (N_2643,N_2582,N_2585);
nor U2644 (N_2644,N_2600,N_2610);
nand U2645 (N_2645,N_2631,N_2634);
or U2646 (N_2646,N_2599,N_2633);
or U2647 (N_2647,N_2628,N_2588);
nor U2648 (N_2648,N_2614,N_2611);
nand U2649 (N_2649,N_2625,N_2580);
and U2650 (N_2650,N_2604,N_2629);
nand U2651 (N_2651,N_2606,N_2638);
nor U2652 (N_2652,N_2613,N_2607);
nand U2653 (N_2653,N_2593,N_2617);
nor U2654 (N_2654,N_2584,N_2619);
nand U2655 (N_2655,N_2598,N_2592);
and U2656 (N_2656,N_2581,N_2602);
nand U2657 (N_2657,N_2624,N_2591);
or U2658 (N_2658,N_2636,N_2587);
nand U2659 (N_2659,N_2609,N_2601);
nor U2660 (N_2660,N_2590,N_2603);
and U2661 (N_2661,N_2616,N_2627);
and U2662 (N_2662,N_2608,N_2589);
nand U2663 (N_2663,N_2637,N_2621);
nor U2664 (N_2664,N_2605,N_2615);
and U2665 (N_2665,N_2635,N_2626);
nand U2666 (N_2666,N_2630,N_2583);
nand U2667 (N_2667,N_2595,N_2620);
nor U2668 (N_2668,N_2586,N_2612);
nand U2669 (N_2669,N_2622,N_2597);
xor U2670 (N_2670,N_2632,N_2589);
and U2671 (N_2671,N_2583,N_2635);
or U2672 (N_2672,N_2582,N_2632);
nand U2673 (N_2673,N_2586,N_2635);
or U2674 (N_2674,N_2637,N_2583);
nor U2675 (N_2675,N_2597,N_2623);
or U2676 (N_2676,N_2614,N_2598);
nor U2677 (N_2677,N_2603,N_2630);
nor U2678 (N_2678,N_2611,N_2595);
or U2679 (N_2679,N_2586,N_2591);
nand U2680 (N_2680,N_2622,N_2593);
or U2681 (N_2681,N_2580,N_2637);
or U2682 (N_2682,N_2623,N_2629);
nor U2683 (N_2683,N_2601,N_2603);
and U2684 (N_2684,N_2612,N_2580);
and U2685 (N_2685,N_2621,N_2639);
nand U2686 (N_2686,N_2608,N_2596);
xor U2687 (N_2687,N_2599,N_2623);
and U2688 (N_2688,N_2611,N_2620);
or U2689 (N_2689,N_2633,N_2596);
or U2690 (N_2690,N_2600,N_2625);
nor U2691 (N_2691,N_2586,N_2632);
nand U2692 (N_2692,N_2616,N_2626);
or U2693 (N_2693,N_2596,N_2601);
or U2694 (N_2694,N_2626,N_2584);
and U2695 (N_2695,N_2612,N_2602);
and U2696 (N_2696,N_2610,N_2586);
and U2697 (N_2697,N_2595,N_2623);
nor U2698 (N_2698,N_2612,N_2601);
and U2699 (N_2699,N_2591,N_2581);
or U2700 (N_2700,N_2698,N_2641);
and U2701 (N_2701,N_2667,N_2672);
nand U2702 (N_2702,N_2687,N_2683);
or U2703 (N_2703,N_2643,N_2642);
nand U2704 (N_2704,N_2671,N_2668);
nand U2705 (N_2705,N_2665,N_2697);
and U2706 (N_2706,N_2658,N_2659);
nor U2707 (N_2707,N_2640,N_2688);
and U2708 (N_2708,N_2645,N_2660);
nor U2709 (N_2709,N_2684,N_2675);
nand U2710 (N_2710,N_2680,N_2666);
nor U2711 (N_2711,N_2670,N_2690);
nor U2712 (N_2712,N_2651,N_2661);
and U2713 (N_2713,N_2646,N_2663);
and U2714 (N_2714,N_2691,N_2699);
nor U2715 (N_2715,N_2694,N_2647);
or U2716 (N_2716,N_2674,N_2662);
nor U2717 (N_2717,N_2676,N_2669);
and U2718 (N_2718,N_2692,N_2673);
nor U2719 (N_2719,N_2677,N_2656);
nor U2720 (N_2720,N_2695,N_2655);
nand U2721 (N_2721,N_2679,N_2681);
or U2722 (N_2722,N_2686,N_2648);
nor U2723 (N_2723,N_2689,N_2657);
and U2724 (N_2724,N_2650,N_2678);
nor U2725 (N_2725,N_2664,N_2693);
or U2726 (N_2726,N_2652,N_2653);
nand U2727 (N_2727,N_2644,N_2682);
nor U2728 (N_2728,N_2696,N_2654);
nand U2729 (N_2729,N_2649,N_2685);
nor U2730 (N_2730,N_2660,N_2666);
xor U2731 (N_2731,N_2651,N_2642);
or U2732 (N_2732,N_2659,N_2666);
nand U2733 (N_2733,N_2671,N_2656);
nand U2734 (N_2734,N_2687,N_2692);
or U2735 (N_2735,N_2645,N_2647);
or U2736 (N_2736,N_2659,N_2683);
or U2737 (N_2737,N_2645,N_2680);
and U2738 (N_2738,N_2683,N_2666);
nand U2739 (N_2739,N_2689,N_2697);
nand U2740 (N_2740,N_2661,N_2688);
nor U2741 (N_2741,N_2658,N_2672);
and U2742 (N_2742,N_2690,N_2692);
nor U2743 (N_2743,N_2665,N_2678);
and U2744 (N_2744,N_2667,N_2656);
nor U2745 (N_2745,N_2664,N_2678);
or U2746 (N_2746,N_2660,N_2678);
nor U2747 (N_2747,N_2642,N_2673);
nand U2748 (N_2748,N_2672,N_2641);
nand U2749 (N_2749,N_2653,N_2656);
and U2750 (N_2750,N_2648,N_2689);
nor U2751 (N_2751,N_2669,N_2678);
nand U2752 (N_2752,N_2666,N_2685);
and U2753 (N_2753,N_2697,N_2640);
nor U2754 (N_2754,N_2670,N_2649);
nor U2755 (N_2755,N_2697,N_2650);
or U2756 (N_2756,N_2642,N_2658);
or U2757 (N_2757,N_2659,N_2696);
and U2758 (N_2758,N_2694,N_2681);
or U2759 (N_2759,N_2690,N_2644);
nand U2760 (N_2760,N_2756,N_2722);
or U2761 (N_2761,N_2736,N_2748);
nor U2762 (N_2762,N_2730,N_2739);
nor U2763 (N_2763,N_2734,N_2711);
nor U2764 (N_2764,N_2731,N_2716);
and U2765 (N_2765,N_2719,N_2751);
nand U2766 (N_2766,N_2754,N_2742);
nand U2767 (N_2767,N_2732,N_2749);
nand U2768 (N_2768,N_2738,N_2704);
nor U2769 (N_2769,N_2728,N_2720);
nor U2770 (N_2770,N_2705,N_2724);
nand U2771 (N_2771,N_2725,N_2709);
nand U2772 (N_2772,N_2712,N_2700);
and U2773 (N_2773,N_2707,N_2721);
nand U2774 (N_2774,N_2717,N_2723);
nor U2775 (N_2775,N_2726,N_2706);
nor U2776 (N_2776,N_2741,N_2713);
nand U2777 (N_2777,N_2757,N_2752);
nor U2778 (N_2778,N_2737,N_2702);
or U2779 (N_2779,N_2744,N_2755);
nand U2780 (N_2780,N_2743,N_2759);
and U2781 (N_2781,N_2729,N_2708);
nand U2782 (N_2782,N_2745,N_2750);
and U2783 (N_2783,N_2715,N_2701);
nand U2784 (N_2784,N_2727,N_2740);
nand U2785 (N_2785,N_2747,N_2710);
or U2786 (N_2786,N_2758,N_2714);
or U2787 (N_2787,N_2703,N_2746);
and U2788 (N_2788,N_2733,N_2718);
and U2789 (N_2789,N_2735,N_2753);
and U2790 (N_2790,N_2741,N_2754);
nor U2791 (N_2791,N_2714,N_2731);
or U2792 (N_2792,N_2706,N_2749);
or U2793 (N_2793,N_2722,N_2748);
and U2794 (N_2794,N_2752,N_2703);
nand U2795 (N_2795,N_2732,N_2737);
and U2796 (N_2796,N_2722,N_2703);
and U2797 (N_2797,N_2718,N_2759);
nor U2798 (N_2798,N_2711,N_2745);
and U2799 (N_2799,N_2713,N_2734);
xor U2800 (N_2800,N_2748,N_2746);
or U2801 (N_2801,N_2726,N_2719);
and U2802 (N_2802,N_2708,N_2740);
or U2803 (N_2803,N_2717,N_2759);
or U2804 (N_2804,N_2714,N_2744);
nor U2805 (N_2805,N_2754,N_2748);
nand U2806 (N_2806,N_2701,N_2740);
nor U2807 (N_2807,N_2741,N_2712);
nand U2808 (N_2808,N_2759,N_2735);
or U2809 (N_2809,N_2715,N_2751);
or U2810 (N_2810,N_2719,N_2734);
nor U2811 (N_2811,N_2740,N_2715);
nor U2812 (N_2812,N_2743,N_2717);
and U2813 (N_2813,N_2701,N_2703);
nor U2814 (N_2814,N_2713,N_2759);
and U2815 (N_2815,N_2741,N_2702);
nand U2816 (N_2816,N_2736,N_2724);
nor U2817 (N_2817,N_2700,N_2725);
and U2818 (N_2818,N_2704,N_2733);
nand U2819 (N_2819,N_2750,N_2710);
and U2820 (N_2820,N_2817,N_2761);
nor U2821 (N_2821,N_2769,N_2778);
and U2822 (N_2822,N_2771,N_2809);
nand U2823 (N_2823,N_2784,N_2819);
nor U2824 (N_2824,N_2779,N_2764);
nor U2825 (N_2825,N_2777,N_2799);
nor U2826 (N_2826,N_2791,N_2788);
nand U2827 (N_2827,N_2770,N_2760);
or U2828 (N_2828,N_2776,N_2785);
or U2829 (N_2829,N_2763,N_2767);
and U2830 (N_2830,N_2803,N_2774);
and U2831 (N_2831,N_2793,N_2786);
and U2832 (N_2832,N_2811,N_2801);
or U2833 (N_2833,N_2762,N_2813);
or U2834 (N_2834,N_2815,N_2816);
nand U2835 (N_2835,N_2798,N_2802);
nand U2836 (N_2836,N_2806,N_2768);
and U2837 (N_2837,N_2782,N_2808);
or U2838 (N_2838,N_2765,N_2787);
nand U2839 (N_2839,N_2804,N_2794);
nor U2840 (N_2840,N_2800,N_2810);
and U2841 (N_2841,N_2807,N_2795);
and U2842 (N_2842,N_2805,N_2772);
nor U2843 (N_2843,N_2814,N_2789);
nor U2844 (N_2844,N_2790,N_2818);
nand U2845 (N_2845,N_2781,N_2783);
or U2846 (N_2846,N_2775,N_2797);
nand U2847 (N_2847,N_2796,N_2766);
nand U2848 (N_2848,N_2780,N_2812);
nand U2849 (N_2849,N_2792,N_2773);
nand U2850 (N_2850,N_2797,N_2787);
xor U2851 (N_2851,N_2793,N_2795);
or U2852 (N_2852,N_2772,N_2788);
nor U2853 (N_2853,N_2768,N_2765);
nand U2854 (N_2854,N_2806,N_2792);
nor U2855 (N_2855,N_2786,N_2819);
and U2856 (N_2856,N_2760,N_2817);
and U2857 (N_2857,N_2808,N_2767);
and U2858 (N_2858,N_2765,N_2796);
nor U2859 (N_2859,N_2774,N_2781);
nand U2860 (N_2860,N_2818,N_2771);
nand U2861 (N_2861,N_2809,N_2761);
and U2862 (N_2862,N_2766,N_2803);
or U2863 (N_2863,N_2767,N_2797);
and U2864 (N_2864,N_2812,N_2808);
nand U2865 (N_2865,N_2776,N_2778);
or U2866 (N_2866,N_2817,N_2800);
nand U2867 (N_2867,N_2816,N_2805);
and U2868 (N_2868,N_2783,N_2769);
and U2869 (N_2869,N_2762,N_2773);
and U2870 (N_2870,N_2808,N_2780);
and U2871 (N_2871,N_2799,N_2776);
or U2872 (N_2872,N_2777,N_2802);
and U2873 (N_2873,N_2817,N_2787);
or U2874 (N_2874,N_2816,N_2786);
nor U2875 (N_2875,N_2765,N_2783);
nand U2876 (N_2876,N_2763,N_2776);
nor U2877 (N_2877,N_2811,N_2808);
and U2878 (N_2878,N_2786,N_2797);
nor U2879 (N_2879,N_2760,N_2805);
nor U2880 (N_2880,N_2867,N_2873);
nor U2881 (N_2881,N_2863,N_2875);
nand U2882 (N_2882,N_2870,N_2838);
or U2883 (N_2883,N_2861,N_2874);
nor U2884 (N_2884,N_2831,N_2840);
or U2885 (N_2885,N_2872,N_2878);
and U2886 (N_2886,N_2842,N_2830);
or U2887 (N_2887,N_2828,N_2858);
or U2888 (N_2888,N_2823,N_2839);
or U2889 (N_2889,N_2827,N_2862);
xor U2890 (N_2890,N_2834,N_2848);
and U2891 (N_2891,N_2869,N_2847);
or U2892 (N_2892,N_2849,N_2829);
nor U2893 (N_2893,N_2859,N_2846);
nand U2894 (N_2894,N_2857,N_2852);
or U2895 (N_2895,N_2876,N_2821);
nand U2896 (N_2896,N_2826,N_2864);
nor U2897 (N_2897,N_2868,N_2856);
and U2898 (N_2898,N_2825,N_2820);
nor U2899 (N_2899,N_2835,N_2854);
or U2900 (N_2900,N_2879,N_2865);
nand U2901 (N_2901,N_2836,N_2851);
and U2902 (N_2902,N_2833,N_2850);
and U2903 (N_2903,N_2822,N_2860);
or U2904 (N_2904,N_2832,N_2877);
or U2905 (N_2905,N_2845,N_2853);
nor U2906 (N_2906,N_2871,N_2855);
nor U2907 (N_2907,N_2837,N_2843);
and U2908 (N_2908,N_2824,N_2844);
and U2909 (N_2909,N_2841,N_2866);
or U2910 (N_2910,N_2862,N_2840);
nand U2911 (N_2911,N_2853,N_2832);
or U2912 (N_2912,N_2872,N_2829);
nand U2913 (N_2913,N_2831,N_2824);
and U2914 (N_2914,N_2857,N_2844);
nand U2915 (N_2915,N_2856,N_2840);
nor U2916 (N_2916,N_2840,N_2869);
nand U2917 (N_2917,N_2870,N_2847);
or U2918 (N_2918,N_2877,N_2825);
nor U2919 (N_2919,N_2829,N_2852);
nor U2920 (N_2920,N_2831,N_2873);
nor U2921 (N_2921,N_2865,N_2827);
and U2922 (N_2922,N_2873,N_2845);
and U2923 (N_2923,N_2831,N_2854);
nor U2924 (N_2924,N_2864,N_2830);
nand U2925 (N_2925,N_2820,N_2878);
nor U2926 (N_2926,N_2874,N_2846);
or U2927 (N_2927,N_2856,N_2850);
and U2928 (N_2928,N_2870,N_2845);
or U2929 (N_2929,N_2830,N_2876);
nand U2930 (N_2930,N_2866,N_2846);
nand U2931 (N_2931,N_2851,N_2840);
or U2932 (N_2932,N_2824,N_2846);
nand U2933 (N_2933,N_2878,N_2853);
nand U2934 (N_2934,N_2870,N_2842);
nand U2935 (N_2935,N_2865,N_2869);
nand U2936 (N_2936,N_2830,N_2851);
or U2937 (N_2937,N_2862,N_2833);
and U2938 (N_2938,N_2853,N_2831);
nand U2939 (N_2939,N_2874,N_2845);
or U2940 (N_2940,N_2903,N_2881);
or U2941 (N_2941,N_2925,N_2927);
and U2942 (N_2942,N_2884,N_2930);
nand U2943 (N_2943,N_2919,N_2911);
nor U2944 (N_2944,N_2923,N_2887);
and U2945 (N_2945,N_2894,N_2916);
or U2946 (N_2946,N_2915,N_2921);
or U2947 (N_2947,N_2934,N_2888);
nor U2948 (N_2948,N_2939,N_2933);
nand U2949 (N_2949,N_2883,N_2924);
or U2950 (N_2950,N_2929,N_2902);
nor U2951 (N_2951,N_2935,N_2886);
or U2952 (N_2952,N_2910,N_2898);
nor U2953 (N_2953,N_2922,N_2892);
or U2954 (N_2954,N_2908,N_2901);
nor U2955 (N_2955,N_2897,N_2900);
nand U2956 (N_2956,N_2913,N_2904);
or U2957 (N_2957,N_2918,N_2936);
or U2958 (N_2958,N_2891,N_2926);
nor U2959 (N_2959,N_2938,N_2906);
nor U2960 (N_2960,N_2920,N_2928);
nor U2961 (N_2961,N_2899,N_2937);
or U2962 (N_2962,N_2885,N_2912);
or U2963 (N_2963,N_2896,N_2932);
or U2964 (N_2964,N_2893,N_2882);
nand U2965 (N_2965,N_2880,N_2889);
and U2966 (N_2966,N_2909,N_2890);
nor U2967 (N_2967,N_2931,N_2914);
or U2968 (N_2968,N_2905,N_2917);
and U2969 (N_2969,N_2895,N_2907);
and U2970 (N_2970,N_2930,N_2883);
nor U2971 (N_2971,N_2918,N_2917);
or U2972 (N_2972,N_2925,N_2913);
and U2973 (N_2973,N_2936,N_2927);
nor U2974 (N_2974,N_2903,N_2915);
or U2975 (N_2975,N_2939,N_2899);
nand U2976 (N_2976,N_2886,N_2919);
and U2977 (N_2977,N_2935,N_2910);
and U2978 (N_2978,N_2933,N_2897);
nor U2979 (N_2979,N_2906,N_2920);
or U2980 (N_2980,N_2929,N_2888);
nand U2981 (N_2981,N_2916,N_2895);
nand U2982 (N_2982,N_2936,N_2898);
and U2983 (N_2983,N_2907,N_2915);
or U2984 (N_2984,N_2922,N_2890);
nand U2985 (N_2985,N_2931,N_2899);
nand U2986 (N_2986,N_2912,N_2906);
nor U2987 (N_2987,N_2901,N_2920);
or U2988 (N_2988,N_2938,N_2939);
or U2989 (N_2989,N_2909,N_2897);
or U2990 (N_2990,N_2920,N_2892);
or U2991 (N_2991,N_2925,N_2901);
and U2992 (N_2992,N_2890,N_2924);
and U2993 (N_2993,N_2895,N_2910);
nand U2994 (N_2994,N_2883,N_2909);
nand U2995 (N_2995,N_2939,N_2890);
nor U2996 (N_2996,N_2903,N_2880);
nor U2997 (N_2997,N_2886,N_2939);
nand U2998 (N_2998,N_2896,N_2890);
and U2999 (N_2999,N_2939,N_2904);
nor UO_0 (O_0,N_2980,N_2971);
nor UO_1 (O_1,N_2992,N_2960);
or UO_2 (O_2,N_2985,N_2998);
and UO_3 (O_3,N_2989,N_2967);
nor UO_4 (O_4,N_2951,N_2946);
and UO_5 (O_5,N_2963,N_2997);
nor UO_6 (O_6,N_2945,N_2990);
and UO_7 (O_7,N_2948,N_2995);
nor UO_8 (O_8,N_2987,N_2962);
and UO_9 (O_9,N_2942,N_2999);
and UO_10 (O_10,N_2981,N_2965);
nor UO_11 (O_11,N_2983,N_2975);
or UO_12 (O_12,N_2968,N_2940);
xnor UO_13 (O_13,N_2972,N_2941);
and UO_14 (O_14,N_2955,N_2961);
or UO_15 (O_15,N_2991,N_2994);
and UO_16 (O_16,N_2986,N_2982);
nor UO_17 (O_17,N_2979,N_2966);
and UO_18 (O_18,N_2953,N_2974);
nand UO_19 (O_19,N_2977,N_2959);
nand UO_20 (O_20,N_2944,N_2952);
and UO_21 (O_21,N_2988,N_2950);
nor UO_22 (O_22,N_2984,N_2969);
or UO_23 (O_23,N_2947,N_2970);
or UO_24 (O_24,N_2949,N_2993);
or UO_25 (O_25,N_2996,N_2978);
and UO_26 (O_26,N_2964,N_2958);
nor UO_27 (O_27,N_2943,N_2973);
nand UO_28 (O_28,N_2957,N_2956);
and UO_29 (O_29,N_2954,N_2976);
and UO_30 (O_30,N_2986,N_2973);
nor UO_31 (O_31,N_2942,N_2980);
nand UO_32 (O_32,N_2963,N_2970);
and UO_33 (O_33,N_2981,N_2953);
nand UO_34 (O_34,N_2953,N_2996);
nand UO_35 (O_35,N_2994,N_2975);
nor UO_36 (O_36,N_2973,N_2951);
or UO_37 (O_37,N_2970,N_2941);
nand UO_38 (O_38,N_2971,N_2957);
nand UO_39 (O_39,N_2982,N_2940);
nand UO_40 (O_40,N_2967,N_2941);
nor UO_41 (O_41,N_2982,N_2995);
nor UO_42 (O_42,N_2940,N_2981);
nand UO_43 (O_43,N_2950,N_2972);
nor UO_44 (O_44,N_2967,N_2950);
or UO_45 (O_45,N_2970,N_2948);
or UO_46 (O_46,N_2955,N_2997);
or UO_47 (O_47,N_2985,N_2962);
nor UO_48 (O_48,N_2951,N_2969);
nand UO_49 (O_49,N_2973,N_2945);
and UO_50 (O_50,N_2976,N_2992);
nand UO_51 (O_51,N_2978,N_2979);
nor UO_52 (O_52,N_2996,N_2956);
nand UO_53 (O_53,N_2975,N_2943);
and UO_54 (O_54,N_2981,N_2980);
nor UO_55 (O_55,N_2989,N_2997);
nor UO_56 (O_56,N_2975,N_2987);
nand UO_57 (O_57,N_2967,N_2953);
or UO_58 (O_58,N_2985,N_2969);
or UO_59 (O_59,N_2986,N_2960);
nand UO_60 (O_60,N_2979,N_2973);
nor UO_61 (O_61,N_2947,N_2943);
nor UO_62 (O_62,N_2943,N_2972);
and UO_63 (O_63,N_2947,N_2964);
nand UO_64 (O_64,N_2964,N_2981);
or UO_65 (O_65,N_2950,N_2983);
nand UO_66 (O_66,N_2970,N_2981);
or UO_67 (O_67,N_2999,N_2956);
nor UO_68 (O_68,N_2947,N_2961);
nand UO_69 (O_69,N_2954,N_2984);
nor UO_70 (O_70,N_2958,N_2981);
nand UO_71 (O_71,N_2973,N_2987);
xnor UO_72 (O_72,N_2953,N_2963);
nand UO_73 (O_73,N_2952,N_2940);
nand UO_74 (O_74,N_2997,N_2992);
and UO_75 (O_75,N_2994,N_2945);
nor UO_76 (O_76,N_2951,N_2964);
or UO_77 (O_77,N_2989,N_2964);
and UO_78 (O_78,N_2981,N_2983);
and UO_79 (O_79,N_2981,N_2996);
or UO_80 (O_80,N_2973,N_2989);
or UO_81 (O_81,N_2970,N_2951);
and UO_82 (O_82,N_2987,N_2992);
and UO_83 (O_83,N_2971,N_2982);
nand UO_84 (O_84,N_2958,N_2976);
and UO_85 (O_85,N_2957,N_2969);
nand UO_86 (O_86,N_2944,N_2950);
and UO_87 (O_87,N_2955,N_2972);
and UO_88 (O_88,N_2990,N_2948);
nand UO_89 (O_89,N_2967,N_2966);
and UO_90 (O_90,N_2962,N_2994);
or UO_91 (O_91,N_2996,N_2955);
nand UO_92 (O_92,N_2992,N_2945);
nand UO_93 (O_93,N_2976,N_2940);
and UO_94 (O_94,N_2999,N_2958);
or UO_95 (O_95,N_2949,N_2957);
nor UO_96 (O_96,N_2980,N_2978);
nor UO_97 (O_97,N_2959,N_2953);
or UO_98 (O_98,N_2943,N_2951);
or UO_99 (O_99,N_2965,N_2974);
nand UO_100 (O_100,N_2976,N_2965);
or UO_101 (O_101,N_2972,N_2971);
nor UO_102 (O_102,N_2969,N_2994);
nor UO_103 (O_103,N_2971,N_2950);
nand UO_104 (O_104,N_2957,N_2959);
and UO_105 (O_105,N_2970,N_2950);
nor UO_106 (O_106,N_2980,N_2989);
nand UO_107 (O_107,N_2974,N_2940);
or UO_108 (O_108,N_2969,N_2989);
and UO_109 (O_109,N_2962,N_2995);
nor UO_110 (O_110,N_2948,N_2999);
or UO_111 (O_111,N_2942,N_2961);
and UO_112 (O_112,N_2975,N_2950);
nor UO_113 (O_113,N_2987,N_2959);
and UO_114 (O_114,N_2981,N_2963);
and UO_115 (O_115,N_2946,N_2981);
or UO_116 (O_116,N_2969,N_2992);
or UO_117 (O_117,N_2964,N_2948);
or UO_118 (O_118,N_2946,N_2993);
and UO_119 (O_119,N_2946,N_2986);
and UO_120 (O_120,N_2942,N_2989);
and UO_121 (O_121,N_2974,N_2946);
or UO_122 (O_122,N_2951,N_2977);
nor UO_123 (O_123,N_2966,N_2941);
nand UO_124 (O_124,N_2998,N_2968);
nand UO_125 (O_125,N_2954,N_2963);
nand UO_126 (O_126,N_2962,N_2998);
nor UO_127 (O_127,N_2969,N_2991);
nand UO_128 (O_128,N_2978,N_2997);
and UO_129 (O_129,N_2952,N_2970);
and UO_130 (O_130,N_2960,N_2967);
or UO_131 (O_131,N_2971,N_2970);
nand UO_132 (O_132,N_2968,N_2985);
nor UO_133 (O_133,N_2951,N_2940);
or UO_134 (O_134,N_2989,N_2957);
and UO_135 (O_135,N_2965,N_2970);
and UO_136 (O_136,N_2948,N_2947);
and UO_137 (O_137,N_2962,N_2966);
or UO_138 (O_138,N_2989,N_2988);
or UO_139 (O_139,N_2958,N_2954);
and UO_140 (O_140,N_2945,N_2947);
nor UO_141 (O_141,N_2974,N_2996);
and UO_142 (O_142,N_2977,N_2952);
nor UO_143 (O_143,N_2940,N_2984);
nor UO_144 (O_144,N_2981,N_2978);
and UO_145 (O_145,N_2988,N_2995);
or UO_146 (O_146,N_2964,N_2987);
nor UO_147 (O_147,N_2942,N_2979);
or UO_148 (O_148,N_2984,N_2949);
and UO_149 (O_149,N_2980,N_2984);
or UO_150 (O_150,N_2963,N_2971);
or UO_151 (O_151,N_2977,N_2954);
nand UO_152 (O_152,N_2961,N_2967);
nand UO_153 (O_153,N_2992,N_2993);
and UO_154 (O_154,N_2955,N_2992);
nand UO_155 (O_155,N_2940,N_2987);
and UO_156 (O_156,N_2954,N_2946);
and UO_157 (O_157,N_2996,N_2994);
nor UO_158 (O_158,N_2965,N_2941);
nor UO_159 (O_159,N_2992,N_2978);
nand UO_160 (O_160,N_2990,N_2988);
and UO_161 (O_161,N_2942,N_2947);
and UO_162 (O_162,N_2987,N_2952);
and UO_163 (O_163,N_2967,N_2963);
or UO_164 (O_164,N_2966,N_2995);
nor UO_165 (O_165,N_2949,N_2942);
nand UO_166 (O_166,N_2978,N_2983);
nor UO_167 (O_167,N_2958,N_2986);
and UO_168 (O_168,N_2989,N_2940);
or UO_169 (O_169,N_2949,N_2996);
nand UO_170 (O_170,N_2986,N_2999);
nand UO_171 (O_171,N_2980,N_2999);
nand UO_172 (O_172,N_2995,N_2945);
or UO_173 (O_173,N_2995,N_2947);
and UO_174 (O_174,N_2948,N_2982);
or UO_175 (O_175,N_2946,N_2994);
or UO_176 (O_176,N_2947,N_2985);
nand UO_177 (O_177,N_2992,N_2965);
and UO_178 (O_178,N_2977,N_2961);
and UO_179 (O_179,N_2953,N_2956);
and UO_180 (O_180,N_2979,N_2941);
nand UO_181 (O_181,N_2986,N_2975);
nand UO_182 (O_182,N_2943,N_2948);
nor UO_183 (O_183,N_2990,N_2961);
or UO_184 (O_184,N_2941,N_2944);
and UO_185 (O_185,N_2943,N_2962);
or UO_186 (O_186,N_2943,N_2989);
nor UO_187 (O_187,N_2984,N_2945);
nand UO_188 (O_188,N_2950,N_2942);
nor UO_189 (O_189,N_2942,N_2983);
or UO_190 (O_190,N_2992,N_2974);
and UO_191 (O_191,N_2979,N_2947);
nand UO_192 (O_192,N_2980,N_2988);
and UO_193 (O_193,N_2956,N_2960);
or UO_194 (O_194,N_2976,N_2993);
and UO_195 (O_195,N_2942,N_2953);
or UO_196 (O_196,N_2998,N_2961);
nand UO_197 (O_197,N_2975,N_2973);
nand UO_198 (O_198,N_2963,N_2994);
or UO_199 (O_199,N_2956,N_2980);
or UO_200 (O_200,N_2972,N_2962);
or UO_201 (O_201,N_2942,N_2996);
nand UO_202 (O_202,N_2995,N_2986);
or UO_203 (O_203,N_2943,N_2965);
nand UO_204 (O_204,N_2970,N_2959);
nand UO_205 (O_205,N_2971,N_2977);
and UO_206 (O_206,N_2953,N_2984);
and UO_207 (O_207,N_2965,N_2996);
and UO_208 (O_208,N_2971,N_2960);
nor UO_209 (O_209,N_2990,N_2952);
nor UO_210 (O_210,N_2949,N_2999);
nand UO_211 (O_211,N_2987,N_2970);
nor UO_212 (O_212,N_2998,N_2977);
or UO_213 (O_213,N_2948,N_2958);
xor UO_214 (O_214,N_2958,N_2975);
and UO_215 (O_215,N_2992,N_2990);
or UO_216 (O_216,N_2991,N_2943);
nor UO_217 (O_217,N_2988,N_2997);
nand UO_218 (O_218,N_2959,N_2941);
nand UO_219 (O_219,N_2950,N_2943);
nand UO_220 (O_220,N_2941,N_2997);
nand UO_221 (O_221,N_2941,N_2978);
or UO_222 (O_222,N_2991,N_2964);
or UO_223 (O_223,N_2964,N_2999);
nor UO_224 (O_224,N_2973,N_2953);
and UO_225 (O_225,N_2964,N_2977);
and UO_226 (O_226,N_2984,N_2970);
and UO_227 (O_227,N_2996,N_2979);
nor UO_228 (O_228,N_2964,N_2953);
nor UO_229 (O_229,N_2990,N_2987);
and UO_230 (O_230,N_2974,N_2971);
and UO_231 (O_231,N_2969,N_2997);
nor UO_232 (O_232,N_2940,N_2945);
and UO_233 (O_233,N_2951,N_2989);
nand UO_234 (O_234,N_2969,N_2954);
and UO_235 (O_235,N_2991,N_2957);
nor UO_236 (O_236,N_2947,N_2988);
and UO_237 (O_237,N_2947,N_2956);
nor UO_238 (O_238,N_2975,N_2944);
or UO_239 (O_239,N_2994,N_2942);
nand UO_240 (O_240,N_2973,N_2959);
or UO_241 (O_241,N_2991,N_2976);
nor UO_242 (O_242,N_2989,N_2945);
and UO_243 (O_243,N_2993,N_2987);
nand UO_244 (O_244,N_2952,N_2972);
and UO_245 (O_245,N_2940,N_2953);
and UO_246 (O_246,N_2942,N_2940);
nand UO_247 (O_247,N_2983,N_2989);
and UO_248 (O_248,N_2949,N_2991);
nor UO_249 (O_249,N_2993,N_2943);
nand UO_250 (O_250,N_2997,N_2950);
or UO_251 (O_251,N_2998,N_2959);
nor UO_252 (O_252,N_2949,N_2977);
xnor UO_253 (O_253,N_2947,N_2955);
nor UO_254 (O_254,N_2979,N_2982);
nand UO_255 (O_255,N_2941,N_2969);
and UO_256 (O_256,N_2943,N_2968);
and UO_257 (O_257,N_2997,N_2970);
nand UO_258 (O_258,N_2954,N_2968);
or UO_259 (O_259,N_2941,N_2983);
or UO_260 (O_260,N_2995,N_2954);
nand UO_261 (O_261,N_2947,N_2949);
nand UO_262 (O_262,N_2990,N_2967);
nor UO_263 (O_263,N_2944,N_2953);
nor UO_264 (O_264,N_2964,N_2993);
nor UO_265 (O_265,N_2977,N_2957);
or UO_266 (O_266,N_2940,N_2941);
nand UO_267 (O_267,N_2977,N_2955);
nand UO_268 (O_268,N_2974,N_2983);
nor UO_269 (O_269,N_2980,N_2979);
nor UO_270 (O_270,N_2985,N_2971);
nor UO_271 (O_271,N_2997,N_2942);
nand UO_272 (O_272,N_2960,N_2982);
or UO_273 (O_273,N_2959,N_2950);
nor UO_274 (O_274,N_2985,N_2944);
nand UO_275 (O_275,N_2972,N_2975);
nor UO_276 (O_276,N_2967,N_2992);
and UO_277 (O_277,N_2999,N_2963);
and UO_278 (O_278,N_2979,N_2965);
nor UO_279 (O_279,N_2966,N_2991);
or UO_280 (O_280,N_2999,N_2955);
and UO_281 (O_281,N_2970,N_2998);
and UO_282 (O_282,N_2946,N_2940);
nand UO_283 (O_283,N_2984,N_2973);
nor UO_284 (O_284,N_2998,N_2954);
or UO_285 (O_285,N_2940,N_2980);
nand UO_286 (O_286,N_2978,N_2942);
nor UO_287 (O_287,N_2965,N_2990);
nand UO_288 (O_288,N_2981,N_2993);
or UO_289 (O_289,N_2956,N_2961);
nor UO_290 (O_290,N_2961,N_2960);
or UO_291 (O_291,N_2978,N_2984);
nand UO_292 (O_292,N_2976,N_2969);
nand UO_293 (O_293,N_2965,N_2946);
nand UO_294 (O_294,N_2979,N_2969);
nor UO_295 (O_295,N_2945,N_2982);
or UO_296 (O_296,N_2968,N_2965);
nand UO_297 (O_297,N_2984,N_2944);
and UO_298 (O_298,N_2984,N_2982);
nor UO_299 (O_299,N_2992,N_2998);
or UO_300 (O_300,N_2977,N_2968);
nand UO_301 (O_301,N_2970,N_2995);
and UO_302 (O_302,N_2969,N_2948);
nor UO_303 (O_303,N_2958,N_2941);
xor UO_304 (O_304,N_2966,N_2977);
nor UO_305 (O_305,N_2952,N_2991);
nand UO_306 (O_306,N_2971,N_2940);
nand UO_307 (O_307,N_2960,N_2944);
nor UO_308 (O_308,N_2946,N_2967);
nor UO_309 (O_309,N_2960,N_2969);
or UO_310 (O_310,N_2969,N_2998);
or UO_311 (O_311,N_2967,N_2975);
or UO_312 (O_312,N_2944,N_2980);
and UO_313 (O_313,N_2943,N_2945);
nor UO_314 (O_314,N_2953,N_2943);
and UO_315 (O_315,N_2958,N_2947);
or UO_316 (O_316,N_2947,N_2971);
or UO_317 (O_317,N_2990,N_2986);
nand UO_318 (O_318,N_2952,N_2988);
and UO_319 (O_319,N_2974,N_2961);
and UO_320 (O_320,N_2949,N_2990);
nand UO_321 (O_321,N_2941,N_2976);
or UO_322 (O_322,N_2995,N_2942);
and UO_323 (O_323,N_2960,N_2952);
nand UO_324 (O_324,N_2979,N_2998);
and UO_325 (O_325,N_2968,N_2982);
nand UO_326 (O_326,N_2954,N_2961);
nand UO_327 (O_327,N_2952,N_2948);
or UO_328 (O_328,N_2945,N_2966);
or UO_329 (O_329,N_2940,N_2955);
nand UO_330 (O_330,N_2948,N_2972);
and UO_331 (O_331,N_2955,N_2998);
nor UO_332 (O_332,N_2979,N_2940);
nor UO_333 (O_333,N_2977,N_2996);
nand UO_334 (O_334,N_2962,N_2971);
nor UO_335 (O_335,N_2947,N_2957);
and UO_336 (O_336,N_2995,N_2978);
and UO_337 (O_337,N_2976,N_2950);
nand UO_338 (O_338,N_2971,N_2994);
nor UO_339 (O_339,N_2980,N_2945);
nor UO_340 (O_340,N_2949,N_2945);
and UO_341 (O_341,N_2950,N_2960);
nand UO_342 (O_342,N_2952,N_2963);
nor UO_343 (O_343,N_2988,N_2998);
and UO_344 (O_344,N_2944,N_2963);
nand UO_345 (O_345,N_2941,N_2962);
and UO_346 (O_346,N_2978,N_2973);
or UO_347 (O_347,N_2968,N_2942);
nor UO_348 (O_348,N_2956,N_2983);
and UO_349 (O_349,N_2986,N_2976);
and UO_350 (O_350,N_2989,N_2959);
and UO_351 (O_351,N_2991,N_2951);
and UO_352 (O_352,N_2986,N_2944);
nand UO_353 (O_353,N_2959,N_2967);
or UO_354 (O_354,N_2973,N_2941);
or UO_355 (O_355,N_2993,N_2967);
or UO_356 (O_356,N_2977,N_2941);
nand UO_357 (O_357,N_2984,N_2999);
nand UO_358 (O_358,N_2974,N_2959);
nor UO_359 (O_359,N_2983,N_2957);
nand UO_360 (O_360,N_2994,N_2965);
and UO_361 (O_361,N_2981,N_2994);
nand UO_362 (O_362,N_2967,N_2986);
or UO_363 (O_363,N_2956,N_2976);
and UO_364 (O_364,N_2956,N_2974);
or UO_365 (O_365,N_2941,N_2982);
and UO_366 (O_366,N_2985,N_2990);
or UO_367 (O_367,N_2951,N_2966);
and UO_368 (O_368,N_2956,N_2958);
or UO_369 (O_369,N_2974,N_2973);
or UO_370 (O_370,N_2991,N_2948);
and UO_371 (O_371,N_2964,N_2967);
or UO_372 (O_372,N_2945,N_2958);
nor UO_373 (O_373,N_2963,N_2958);
nor UO_374 (O_374,N_2994,N_2999);
or UO_375 (O_375,N_2942,N_2970);
and UO_376 (O_376,N_2950,N_2998);
and UO_377 (O_377,N_2973,N_2995);
and UO_378 (O_378,N_2978,N_2967);
and UO_379 (O_379,N_2996,N_2951);
or UO_380 (O_380,N_2959,N_2943);
nand UO_381 (O_381,N_2987,N_2960);
nor UO_382 (O_382,N_2962,N_2999);
or UO_383 (O_383,N_2952,N_2965);
and UO_384 (O_384,N_2956,N_2978);
nand UO_385 (O_385,N_2958,N_2961);
or UO_386 (O_386,N_2976,N_2955);
and UO_387 (O_387,N_2988,N_2978);
nand UO_388 (O_388,N_2989,N_2990);
nor UO_389 (O_389,N_2994,N_2944);
nor UO_390 (O_390,N_2943,N_2966);
and UO_391 (O_391,N_2962,N_2955);
and UO_392 (O_392,N_2959,N_2945);
or UO_393 (O_393,N_2987,N_2963);
nor UO_394 (O_394,N_2979,N_2957);
nor UO_395 (O_395,N_2957,N_2986);
or UO_396 (O_396,N_2993,N_2978);
nand UO_397 (O_397,N_2961,N_2980);
nand UO_398 (O_398,N_2947,N_2960);
nor UO_399 (O_399,N_2976,N_2951);
nand UO_400 (O_400,N_2966,N_2980);
nor UO_401 (O_401,N_2958,N_2989);
or UO_402 (O_402,N_2995,N_2946);
and UO_403 (O_403,N_2942,N_2945);
and UO_404 (O_404,N_2981,N_2995);
and UO_405 (O_405,N_2997,N_2951);
nand UO_406 (O_406,N_2967,N_2948);
and UO_407 (O_407,N_2944,N_2947);
nand UO_408 (O_408,N_2960,N_2973);
and UO_409 (O_409,N_2966,N_2946);
or UO_410 (O_410,N_2940,N_2948);
nor UO_411 (O_411,N_2998,N_2983);
or UO_412 (O_412,N_2971,N_2996);
or UO_413 (O_413,N_2990,N_2968);
nor UO_414 (O_414,N_2981,N_2955);
nor UO_415 (O_415,N_2970,N_2986);
or UO_416 (O_416,N_2981,N_2972);
nor UO_417 (O_417,N_2992,N_2952);
nand UO_418 (O_418,N_2956,N_2991);
and UO_419 (O_419,N_2996,N_2984);
and UO_420 (O_420,N_2947,N_2998);
and UO_421 (O_421,N_2995,N_2977);
nand UO_422 (O_422,N_2994,N_2982);
or UO_423 (O_423,N_2947,N_2981);
or UO_424 (O_424,N_2980,N_2954);
nand UO_425 (O_425,N_2958,N_2972);
nor UO_426 (O_426,N_2991,N_2963);
and UO_427 (O_427,N_2973,N_2993);
and UO_428 (O_428,N_2997,N_2986);
nor UO_429 (O_429,N_2989,N_2984);
or UO_430 (O_430,N_2978,N_2975);
nand UO_431 (O_431,N_2998,N_2973);
or UO_432 (O_432,N_2969,N_2983);
nand UO_433 (O_433,N_2978,N_2999);
nand UO_434 (O_434,N_2942,N_2972);
and UO_435 (O_435,N_2987,N_2941);
nor UO_436 (O_436,N_2944,N_2995);
nand UO_437 (O_437,N_2982,N_2974);
nand UO_438 (O_438,N_2945,N_2970);
nor UO_439 (O_439,N_2999,N_2993);
and UO_440 (O_440,N_2985,N_2961);
or UO_441 (O_441,N_2996,N_2987);
nor UO_442 (O_442,N_2953,N_2995);
and UO_443 (O_443,N_2950,N_2977);
nor UO_444 (O_444,N_2951,N_2986);
nor UO_445 (O_445,N_2982,N_2997);
nor UO_446 (O_446,N_2983,N_2995);
and UO_447 (O_447,N_2978,N_2945);
and UO_448 (O_448,N_2980,N_2959);
and UO_449 (O_449,N_2941,N_2991);
and UO_450 (O_450,N_2968,N_2949);
and UO_451 (O_451,N_2991,N_2959);
nor UO_452 (O_452,N_2974,N_2957);
or UO_453 (O_453,N_2981,N_2974);
and UO_454 (O_454,N_2944,N_2943);
and UO_455 (O_455,N_2953,N_2982);
or UO_456 (O_456,N_2955,N_2982);
nand UO_457 (O_457,N_2975,N_2965);
nor UO_458 (O_458,N_2989,N_2975);
or UO_459 (O_459,N_2974,N_2952);
nor UO_460 (O_460,N_2965,N_2987);
nand UO_461 (O_461,N_2948,N_2979);
and UO_462 (O_462,N_2998,N_2964);
nand UO_463 (O_463,N_2976,N_2984);
nand UO_464 (O_464,N_2946,N_2941);
and UO_465 (O_465,N_2985,N_2953);
nand UO_466 (O_466,N_2994,N_2952);
nor UO_467 (O_467,N_2966,N_2987);
or UO_468 (O_468,N_2943,N_2997);
nor UO_469 (O_469,N_2951,N_2960);
nor UO_470 (O_470,N_2995,N_2949);
nor UO_471 (O_471,N_2984,N_2995);
nand UO_472 (O_472,N_2996,N_2991);
nand UO_473 (O_473,N_2944,N_2992);
or UO_474 (O_474,N_2965,N_2940);
nor UO_475 (O_475,N_2972,N_2965);
nand UO_476 (O_476,N_2971,N_2967);
and UO_477 (O_477,N_2960,N_2972);
nor UO_478 (O_478,N_2960,N_2989);
nor UO_479 (O_479,N_2990,N_2973);
nand UO_480 (O_480,N_2988,N_2973);
nand UO_481 (O_481,N_2971,N_2987);
nand UO_482 (O_482,N_2993,N_2969);
nor UO_483 (O_483,N_2964,N_2975);
nand UO_484 (O_484,N_2976,N_2946);
nor UO_485 (O_485,N_2975,N_2996);
or UO_486 (O_486,N_2996,N_2976);
or UO_487 (O_487,N_2980,N_2992);
or UO_488 (O_488,N_2960,N_2979);
nand UO_489 (O_489,N_2970,N_2977);
nand UO_490 (O_490,N_2969,N_2972);
or UO_491 (O_491,N_2993,N_2985);
and UO_492 (O_492,N_2983,N_2985);
nor UO_493 (O_493,N_2955,N_2965);
and UO_494 (O_494,N_2956,N_2995);
or UO_495 (O_495,N_2966,N_2981);
nand UO_496 (O_496,N_2986,N_2983);
and UO_497 (O_497,N_2941,N_2975);
nand UO_498 (O_498,N_2968,N_2974);
and UO_499 (O_499,N_2974,N_2986);
endmodule