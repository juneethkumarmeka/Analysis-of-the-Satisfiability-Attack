module basic_1500_15000_2000_3_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10032,N_10033,N_10035,N_10037,N_10038,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10050,N_10051,N_10052,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10064,N_10065,N_10067,N_10068,N_10069,N_10071,N_10072,N_10074,N_10075,N_10076,N_10077,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10092,N_10093,N_10094,N_10096,N_10100,N_10101,N_10102,N_10104,N_10106,N_10107,N_10108,N_10109,N_10110,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10129,N_10130,N_10131,N_10132,N_10134,N_10138,N_10139,N_10140,N_10141,N_10144,N_10145,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10173,N_10174,N_10175,N_10177,N_10180,N_10181,N_10183,N_10185,N_10187,N_10188,N_10189,N_10191,N_10192,N_10194,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10207,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10247,N_10248,N_10249,N_10251,N_10252,N_10255,N_10256,N_10257,N_10259,N_10260,N_10261,N_10262,N_10263,N_10265,N_10266,N_10267,N_10268,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10287,N_10288,N_10289,N_10290,N_10291,N_10293,N_10295,N_10296,N_10298,N_10301,N_10302,N_10303,N_10304,N_10305,N_10307,N_10309,N_10310,N_10311,N_10312,N_10313,N_10315,N_10316,N_10317,N_10319,N_10321,N_10322,N_10323,N_10325,N_10326,N_10331,N_10333,N_10335,N_10336,N_10337,N_10339,N_10341,N_10343,N_10344,N_10345,N_10347,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10357,N_10360,N_10362,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10385,N_10386,N_10389,N_10390,N_10391,N_10393,N_10394,N_10395,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10413,N_10415,N_10416,N_10417,N_10418,N_10420,N_10421,N_10422,N_10424,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10436,N_10438,N_10439,N_10441,N_10443,N_10444,N_10445,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10458,N_10460,N_10461,N_10462,N_10465,N_10466,N_10468,N_10469,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10487,N_10488,N_10490,N_10491,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10501,N_10502,N_10504,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10518,N_10520,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10542,N_10543,N_10544,N_10545,N_10546,N_10548,N_10550,N_10551,N_10552,N_10553,N_10555,N_10556,N_10559,N_10560,N_10562,N_10563,N_10564,N_10565,N_10568,N_10570,N_10572,N_10573,N_10574,N_10575,N_10576,N_10578,N_10579,N_10581,N_10582,N_10583,N_10585,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10604,N_10605,N_10607,N_10608,N_10610,N_10611,N_10612,N_10614,N_10616,N_10617,N_10618,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10629,N_10630,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10641,N_10642,N_10645,N_10646,N_10647,N_10648,N_10649,N_10651,N_10652,N_10653,N_10654,N_10656,N_10658,N_10659,N_10661,N_10662,N_10664,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10679,N_10680,N_10682,N_10683,N_10685,N_10686,N_10688,N_10689,N_10690,N_10691,N_10692,N_10694,N_10695,N_10697,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10712,N_10714,N_10715,N_10717,N_10719,N_10720,N_10722,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10743,N_10744,N_10745,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10757,N_10758,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10775,N_10776,N_10777,N_10778,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10788,N_10789,N_10791,N_10792,N_10793,N_10795,N_10797,N_10798,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10807,N_10808,N_10809,N_10810,N_10811,N_10813,N_10814,N_10816,N_10818,N_10820,N_10821,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10842,N_10843,N_10844,N_10845,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10857,N_10858,N_10859,N_10860,N_10861,N_10864,N_10865,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10887,N_10888,N_10892,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10914,N_10915,N_10917,N_10920,N_10921,N_10922,N_10923,N_10926,N_10927,N_10928,N_10929,N_10931,N_10933,N_10938,N_10939,N_10940,N_10941,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10954,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10964,N_10966,N_10967,N_10968,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10979,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10995,N_10996,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11022,N_11023,N_11024,N_11026,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11042,N_11043,N_11044,N_11045,N_11046,N_11049,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11065,N_11067,N_11068,N_11069,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11086,N_11087,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11097,N_11098,N_11099,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11123,N_11124,N_11125,N_11128,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11147,N_11148,N_11149,N_11151,N_11152,N_11153,N_11154,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11190,N_11191,N_11192,N_11193,N_11195,N_11196,N_11198,N_11199,N_11200,N_11201,N_11203,N_11204,N_11206,N_11210,N_11211,N_11212,N_11213,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11224,N_11225,N_11226,N_11227,N_11229,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11281,N_11283,N_11284,N_11285,N_11286,N_11287,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11298,N_11299,N_11300,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11323,N_11324,N_11325,N_11326,N_11327,N_11329,N_11330,N_11333,N_11334,N_11337,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11348,N_11349,N_11350,N_11352,N_11353,N_11354,N_11357,N_11359,N_11361,N_11362,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11373,N_11374,N_11375,N_11376,N_11377,N_11379,N_11381,N_11383,N_11384,N_11389,N_11390,N_11391,N_11393,N_11394,N_11395,N_11396,N_11398,N_11399,N_11400,N_11401,N_11402,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11412,N_11413,N_11414,N_11415,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11443,N_11446,N_11448,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11460,N_11461,N_11463,N_11465,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11491,N_11492,N_11493,N_11494,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11515,N_11516,N_11518,N_11519,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11528,N_11529,N_11530,N_11531,N_11533,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11555,N_11556,N_11557,N_11558,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11584,N_11585,N_11586,N_11587,N_11588,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11602,N_11603,N_11604,N_11605,N_11607,N_11609,N_11610,N_11612,N_11613,N_11615,N_11616,N_11617,N_11619,N_11620,N_11621,N_11622,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11637,N_11640,N_11641,N_11642,N_11644,N_11645,N_11647,N_11648,N_11649,N_11650,N_11651,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11674,N_11675,N_11676,N_11678,N_11679,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11692,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11730,N_11731,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11740,N_11741,N_11742,N_11743,N_11745,N_11746,N_11747,N_11748,N_11749,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11779,N_11780,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11791,N_11792,N_11795,N_11797,N_11798,N_11799,N_11801,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11827,N_11828,N_11829,N_11830,N_11833,N_11834,N_11835,N_11836,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11859,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11884,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11899,N_11900,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11913,N_11914,N_11915,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11928,N_11929,N_11930,N_11931,N_11932,N_11934,N_11935,N_11936,N_11937,N_11939,N_11940,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11949,N_11950,N_11951,N_11953,N_11954,N_11956,N_11957,N_11959,N_11960,N_11961,N_11965,N_11967,N_11968,N_11970,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11989,N_11990,N_11991,N_11994,N_11995,N_11996,N_11997,N_11999,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12009,N_12011,N_12012,N_12013,N_12014,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12023,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12048,N_12049,N_12050,N_12052,N_12055,N_12057,N_12060,N_12061,N_12063,N_12064,N_12065,N_12067,N_12069,N_12070,N_12071,N_12073,N_12074,N_12076,N_12078,N_12079,N_12082,N_12084,N_12085,N_12086,N_12088,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12110,N_12111,N_12112,N_12113,N_12115,N_12116,N_12117,N_12118,N_12120,N_12121,N_12123,N_12125,N_12127,N_12128,N_12129,N_12131,N_12132,N_12133,N_12134,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12155,N_12156,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12186,N_12187,N_12189,N_12191,N_12193,N_12195,N_12196,N_12197,N_12198,N_12199,N_12201,N_12202,N_12203,N_12205,N_12207,N_12208,N_12209,N_12212,N_12213,N_12215,N_12216,N_12217,N_12218,N_12219,N_12221,N_12222,N_12223,N_12224,N_12226,N_12227,N_12228,N_12230,N_12232,N_12234,N_12236,N_12237,N_12238,N_12241,N_12242,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12258,N_12260,N_12261,N_12262,N_12263,N_12264,N_12267,N_12269,N_12270,N_12272,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12281,N_12284,N_12286,N_12287,N_12288,N_12289,N_12291,N_12292,N_12293,N_12295,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12316,N_12317,N_12318,N_12319,N_12320,N_12322,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12331,N_12332,N_12334,N_12335,N_12336,N_12337,N_12339,N_12343,N_12344,N_12345,N_12347,N_12349,N_12351,N_12352,N_12353,N_12354,N_12356,N_12357,N_12358,N_12359,N_12361,N_12362,N_12363,N_12364,N_12365,N_12367,N_12368,N_12369,N_12370,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12396,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12407,N_12408,N_12410,N_12412,N_12413,N_12414,N_12415,N_12416,N_12418,N_12419,N_12420,N_12421,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12431,N_12432,N_12433,N_12434,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12458,N_12459,N_12460,N_12462,N_12463,N_12464,N_12466,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12479,N_12480,N_12481,N_12483,N_12486,N_12487,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12508,N_12509,N_12510,N_12511,N_12512,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12521,N_12522,N_12524,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12560,N_12561,N_12562,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12592,N_12593,N_12594,N_12595,N_12596,N_12598,N_12599,N_12600,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12613,N_12614,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12631,N_12632,N_12633,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12645,N_12647,N_12648,N_12649,N_12651,N_12652,N_12653,N_12654,N_12655,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12666,N_12668,N_12669,N_12670,N_12671,N_12672,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12689,N_12690,N_12691,N_12692,N_12693,N_12695,N_12696,N_12698,N_12699,N_12700,N_12701,N_12703,N_12704,N_12705,N_12707,N_12708,N_12709,N_12710,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12750,N_12753,N_12754,N_12755,N_12756,N_12758,N_12760,N_12761,N_12762,N_12763,N_12765,N_12766,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12790,N_12791,N_12792,N_12795,N_12796,N_12797,N_12798,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12811,N_12812,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12835,N_12836,N_12837,N_12839,N_12840,N_12841,N_12845,N_12846,N_12848,N_12849,N_12851,N_12852,N_12853,N_12854,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12870,N_12871,N_12873,N_12874,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12887,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12898,N_12899,N_12900,N_12902,N_12904,N_12905,N_12907,N_12908,N_12910,N_12911,N_12912,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12965,N_12966,N_12968,N_12969,N_12971,N_12973,N_12974,N_12975,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12984,N_12985,N_12986,N_12987,N_12989,N_12991,N_12992,N_12994,N_12995,N_12996,N_13000,N_13001,N_13002,N_13004,N_13005,N_13006,N_13007,N_13008,N_13010,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13076,N_13077,N_13079,N_13080,N_13081,N_13083,N_13084,N_13086,N_13088,N_13089,N_13090,N_13091,N_13093,N_13094,N_13095,N_13096,N_13097,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13106,N_13108,N_13109,N_13110,N_13112,N_13113,N_13118,N_13119,N_13120,N_13121,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13131,N_13132,N_13133,N_13135,N_13136,N_13137,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13159,N_13161,N_13162,N_13164,N_13165,N_13166,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13176,N_13177,N_13179,N_13180,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13190,N_13192,N_13193,N_13194,N_13195,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13205,N_13206,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13245,N_13247,N_13248,N_13249,N_13250,N_13253,N_13254,N_13255,N_13256,N_13257,N_13260,N_13261,N_13262,N_13264,N_13265,N_13266,N_13267,N_13268,N_13270,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13281,N_13282,N_13283,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13298,N_13299,N_13301,N_13302,N_13304,N_13305,N_13306,N_13307,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13348,N_13350,N_13351,N_13352,N_13354,N_13355,N_13356,N_13357,N_13358,N_13360,N_13361,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13381,N_13382,N_13384,N_13385,N_13386,N_13388,N_13390,N_13391,N_13392,N_13393,N_13394,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13409,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13418,N_13419,N_13420,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13433,N_13434,N_13435,N_13436,N_13437,N_13439,N_13440,N_13441,N_13443,N_13446,N_13447,N_13448,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13459,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13500,N_13501,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13512,N_13514,N_13515,N_13516,N_13517,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13526,N_13529,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13568,N_13569,N_13570,N_13571,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13601,N_13602,N_13603,N_13605,N_13606,N_13607,N_13608,N_13609,N_13611,N_13612,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13625,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13635,N_13636,N_13637,N_13638,N_13639,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13648,N_13649,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13670,N_13671,N_13672,N_13674,N_13675,N_13676,N_13677,N_13682,N_13684,N_13685,N_13686,N_13689,N_13690,N_13691,N_13693,N_13694,N_13695,N_13696,N_13697,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13709,N_13710,N_13711,N_13713,N_13715,N_13716,N_13717,N_13718,N_13719,N_13721,N_13722,N_13723,N_13724,N_13726,N_13727,N_13728,N_13729,N_13730,N_13732,N_13733,N_13734,N_13735,N_13736,N_13738,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13760,N_13761,N_13762,N_13763,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13775,N_13776,N_13777,N_13778,N_13780,N_13781,N_13782,N_13783,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13792,N_13793,N_13794,N_13795,N_13798,N_13799,N_13800,N_13802,N_13803,N_13804,N_13807,N_13808,N_13810,N_13811,N_13813,N_13814,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13824,N_13827,N_13829,N_13830,N_13831,N_13833,N_13835,N_13836,N_13837,N_13839,N_13840,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13917,N_13918,N_13920,N_13921,N_13922,N_13924,N_13926,N_13927,N_13929,N_13930,N_13932,N_13933,N_13935,N_13936,N_13937,N_13938,N_13939,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13974,N_13975,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13986,N_13988,N_13991,N_13992,N_13993,N_13994,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14004,N_14006,N_14008,N_14010,N_14011,N_14012,N_14014,N_14015,N_14016,N_14017,N_14019,N_14020,N_14021,N_14023,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14041,N_14042,N_14044,N_14045,N_14046,N_14047,N_14048,N_14050,N_14051,N_14053,N_14054,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14082,N_14083,N_14084,N_14086,N_14088,N_14091,N_14092,N_14093,N_14094,N_14095,N_14097,N_14098,N_14099,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14160,N_14161,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14181,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14203,N_14205,N_14207,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14244,N_14245,N_14246,N_14248,N_14249,N_14250,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14260,N_14261,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14271,N_14272,N_14273,N_14275,N_14277,N_14278,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14287,N_14288,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14298,N_14299,N_14300,N_14301,N_14303,N_14305,N_14306,N_14307,N_14309,N_14311,N_14312,N_14313,N_14314,N_14315,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14326,N_14328,N_14329,N_14331,N_14334,N_14335,N_14336,N_14337,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14357,N_14358,N_14359,N_14363,N_14364,N_14365,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14402,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14415,N_14417,N_14418,N_14421,N_14422,N_14423,N_14425,N_14426,N_14427,N_14429,N_14430,N_14431,N_14432,N_14434,N_14435,N_14436,N_14437,N_14439,N_14440,N_14441,N_14442,N_14444,N_14445,N_14446,N_14447,N_14448,N_14450,N_14451,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14471,N_14473,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14574,N_14576,N_14578,N_14579,N_14580,N_14581,N_14582,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14620,N_14621,N_14622,N_14623,N_14624,N_14626,N_14627,N_14628,N_14631,N_14632,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14649,N_14650,N_14651,N_14652,N_14654,N_14655,N_14656,N_14657,N_14659,N_14660,N_14662,N_14663,N_14664,N_14665,N_14668,N_14669,N_14670,N_14671,N_14672,N_14674,N_14675,N_14676,N_14677,N_14679,N_14680,N_14681,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14703,N_14704,N_14706,N_14707,N_14709,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14719,N_14721,N_14722,N_14725,N_14726,N_14727,N_14729,N_14731,N_14732,N_14733,N_14734,N_14737,N_14741,N_14742,N_14743,N_14745,N_14746,N_14747,N_14748,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14758,N_14759,N_14760,N_14762,N_14763,N_14766,N_14767,N_14769,N_14771,N_14772,N_14773,N_14774,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14793,N_14794,N_14795,N_14796,N_14797,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14817,N_14818,N_14819,N_14820,N_14821,N_14823,N_14824,N_14825,N_14827,N_14828,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14867,N_14869,N_14870,N_14871,N_14872,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14889,N_14890,N_14891,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14909,N_14910,N_14911,N_14913,N_14914,N_14915,N_14916,N_14917,N_14920,N_14921,N_14922,N_14924,N_14926,N_14927,N_14928,N_14929,N_14930,N_14932,N_14933,N_14934,N_14935,N_14937,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14950,N_14951,N_14952,N_14953,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14972,N_14973,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14997,N_14998;
and U0 (N_0,In_1186,In_1470);
nand U1 (N_1,In_745,In_264);
nor U2 (N_2,In_108,In_534);
nand U3 (N_3,In_1113,In_7);
xnor U4 (N_4,In_933,In_343);
nand U5 (N_5,In_483,In_874);
and U6 (N_6,In_1367,In_1279);
nand U7 (N_7,In_332,In_1436);
or U8 (N_8,In_623,In_928);
and U9 (N_9,In_1346,In_1497);
nor U10 (N_10,In_1339,In_100);
xnor U11 (N_11,In_980,In_1249);
nor U12 (N_12,In_117,In_885);
nand U13 (N_13,In_1387,In_20);
and U14 (N_14,In_67,In_998);
or U15 (N_15,In_76,In_396);
and U16 (N_16,In_1242,In_1163);
nor U17 (N_17,In_95,In_349);
nand U18 (N_18,In_1464,In_345);
nor U19 (N_19,In_378,In_429);
or U20 (N_20,In_704,In_219);
or U21 (N_21,In_42,In_1044);
and U22 (N_22,In_942,In_804);
and U23 (N_23,In_153,In_1384);
and U24 (N_24,In_1465,In_981);
nand U25 (N_25,In_148,In_1471);
nand U26 (N_26,In_247,In_893);
nor U27 (N_27,In_935,In_269);
or U28 (N_28,In_503,In_1385);
xor U29 (N_29,In_927,In_304);
nor U30 (N_30,In_92,In_843);
and U31 (N_31,In_550,In_667);
nand U32 (N_32,In_324,In_1121);
nand U33 (N_33,In_730,In_505);
nor U34 (N_34,In_689,In_810);
nand U35 (N_35,In_682,In_1054);
nand U36 (N_36,In_686,In_1434);
and U37 (N_37,In_169,In_157);
xnor U38 (N_38,In_899,In_1202);
or U39 (N_39,In_685,In_1443);
xnor U40 (N_40,In_1228,In_889);
nor U41 (N_41,In_286,In_109);
nor U42 (N_42,In_1416,In_174);
nand U43 (N_43,In_589,In_641);
xor U44 (N_44,In_1035,In_1167);
nand U45 (N_45,In_1287,In_182);
nand U46 (N_46,In_1134,In_1342);
or U47 (N_47,In_1271,In_526);
and U48 (N_48,In_273,In_989);
nand U49 (N_49,In_767,In_798);
nand U50 (N_50,In_1140,In_13);
nor U51 (N_51,In_578,In_1482);
and U52 (N_52,In_122,In_340);
or U53 (N_53,In_19,In_1042);
xnor U54 (N_54,In_517,In_173);
xnor U55 (N_55,In_339,In_445);
nand U56 (N_56,In_313,In_37);
nor U57 (N_57,In_1127,In_71);
nand U58 (N_58,In_1095,In_1);
or U59 (N_59,In_68,In_650);
nand U60 (N_60,In_175,In_1294);
and U61 (N_61,In_713,In_1239);
and U62 (N_62,In_1336,In_848);
and U63 (N_63,In_61,In_524);
xnor U64 (N_64,In_911,In_1313);
nand U65 (N_65,In_451,In_971);
and U66 (N_66,In_1288,In_1055);
and U67 (N_67,In_1032,In_1439);
and U68 (N_68,In_591,In_338);
nor U69 (N_69,In_797,In_690);
xnor U70 (N_70,In_747,In_777);
and U71 (N_71,In_757,In_739);
nand U72 (N_72,In_1155,In_376);
nand U73 (N_73,In_1096,In_888);
nand U74 (N_74,In_639,In_1029);
and U75 (N_75,In_914,In_211);
or U76 (N_76,In_1437,In_541);
nand U77 (N_77,In_902,In_635);
nand U78 (N_78,In_979,In_1149);
nand U79 (N_79,In_660,In_675);
or U80 (N_80,In_172,In_548);
xnor U81 (N_81,In_612,In_1447);
nand U82 (N_82,In_924,In_358);
or U83 (N_83,In_1438,In_60);
and U84 (N_84,In_401,In_587);
nand U85 (N_85,In_659,In_1115);
nand U86 (N_86,In_152,In_496);
xnor U87 (N_87,In_1479,In_271);
nor U88 (N_88,In_466,In_836);
or U89 (N_89,In_908,In_1089);
xor U90 (N_90,In_1124,In_1411);
nor U91 (N_91,In_937,In_295);
and U92 (N_92,In_1222,In_1252);
and U93 (N_93,In_564,In_918);
and U94 (N_94,In_1307,In_861);
nor U95 (N_95,In_841,In_948);
xor U96 (N_96,In_303,In_1407);
nand U97 (N_97,In_452,In_363);
nand U98 (N_98,In_865,In_543);
nor U99 (N_99,In_178,In_1092);
nor U100 (N_100,In_962,In_905);
xor U101 (N_101,In_1404,In_6);
xnor U102 (N_102,In_1148,In_317);
or U103 (N_103,In_404,In_617);
and U104 (N_104,In_706,In_746);
nor U105 (N_105,In_220,In_1341);
xnor U106 (N_106,In_1024,In_1170);
nor U107 (N_107,In_373,In_70);
or U108 (N_108,In_991,In_693);
xnor U109 (N_109,In_726,In_498);
nand U110 (N_110,In_748,In_977);
xor U111 (N_111,In_856,In_423);
nand U112 (N_112,In_151,In_1211);
or U113 (N_113,In_1273,In_314);
and U114 (N_114,In_129,In_627);
and U115 (N_115,In_1298,In_66);
nand U116 (N_116,In_36,In_1080);
or U117 (N_117,In_1059,In_57);
and U118 (N_118,In_201,In_189);
nand U119 (N_119,In_471,In_293);
and U120 (N_120,In_1281,In_656);
or U121 (N_121,In_593,In_1182);
and U122 (N_122,In_904,In_458);
xor U123 (N_123,In_1119,In_877);
xnor U124 (N_124,In_771,In_728);
or U125 (N_125,In_1023,In_909);
nor U126 (N_126,In_1283,In_1386);
xnor U127 (N_127,In_463,In_862);
nor U128 (N_128,In_1454,In_657);
and U129 (N_129,In_1466,In_28);
and U130 (N_130,In_1215,In_315);
xor U131 (N_131,In_1200,In_691);
and U132 (N_132,In_584,In_1382);
nor U133 (N_133,In_291,In_1176);
or U134 (N_134,In_1133,In_839);
nand U135 (N_135,In_491,In_858);
xor U136 (N_136,In_1378,In_880);
and U137 (N_137,In_828,In_93);
nand U138 (N_138,In_732,In_573);
and U139 (N_139,In_890,In_643);
nand U140 (N_140,In_9,In_1147);
nor U141 (N_141,In_1373,In_692);
xor U142 (N_142,In_1421,In_1338);
nor U143 (N_143,In_38,In_51);
nor U144 (N_144,In_1418,In_1187);
or U145 (N_145,In_280,In_165);
xnor U146 (N_146,In_853,In_711);
and U147 (N_147,In_168,In_360);
nand U148 (N_148,In_258,In_586);
nand U149 (N_149,In_440,In_674);
nand U150 (N_150,In_834,In_259);
xor U151 (N_151,In_167,In_102);
nand U152 (N_152,In_1203,In_1154);
and U153 (N_153,In_951,In_1083);
or U154 (N_154,In_1131,In_735);
nand U155 (N_155,In_16,In_585);
and U156 (N_156,In_1033,In_123);
xnor U157 (N_157,In_1426,In_577);
and U158 (N_158,In_621,In_833);
and U159 (N_159,In_337,In_274);
nand U160 (N_160,In_1364,In_562);
xor U161 (N_161,In_1391,In_14);
nand U162 (N_162,In_910,In_1343);
nor U163 (N_163,In_39,In_956);
and U164 (N_164,In_327,In_857);
xor U165 (N_165,In_619,In_892);
nand U166 (N_166,In_1234,In_23);
and U167 (N_167,In_1104,In_91);
nand U168 (N_168,In_850,In_542);
nand U169 (N_169,In_949,In_1094);
or U170 (N_170,In_1185,In_1039);
nor U171 (N_171,In_1389,In_1414);
or U172 (N_172,In_532,In_1077);
or U173 (N_173,In_1041,In_416);
or U174 (N_174,In_1062,In_139);
and U175 (N_175,In_1358,In_1403);
xnor U176 (N_176,In_243,In_1318);
nand U177 (N_177,In_1011,In_1485);
xnor U178 (N_178,In_1037,In_1312);
nand U179 (N_179,In_945,In_470);
nand U180 (N_180,In_1349,In_855);
or U181 (N_181,In_366,In_1204);
nor U182 (N_182,In_512,In_322);
nor U183 (N_183,In_187,In_257);
xor U184 (N_184,In_137,In_142);
and U185 (N_185,In_871,In_823);
or U186 (N_186,In_465,In_287);
nor U187 (N_187,In_520,In_1276);
xor U188 (N_188,In_903,In_1004);
and U189 (N_189,In_982,In_597);
or U190 (N_190,In_215,In_1016);
nor U191 (N_191,In_1250,In_181);
or U192 (N_192,In_967,In_1157);
or U193 (N_193,In_455,In_1213);
or U194 (N_194,In_1424,In_1458);
xor U195 (N_195,In_188,In_957);
xnor U196 (N_196,In_929,In_1152);
xor U197 (N_197,In_847,In_1245);
and U198 (N_198,In_729,In_1299);
or U199 (N_199,In_74,In_826);
nor U200 (N_200,In_953,In_1028);
and U201 (N_201,In_653,In_377);
xnor U202 (N_202,In_133,In_1067);
nand U203 (N_203,In_164,In_531);
xor U204 (N_204,In_1383,In_1036);
xor U205 (N_205,In_1141,In_1463);
nor U206 (N_206,In_916,In_1164);
xnor U207 (N_207,In_196,In_952);
nand U208 (N_208,In_94,In_321);
xor U209 (N_209,In_556,In_626);
or U210 (N_210,In_759,In_1232);
nor U211 (N_211,In_1345,In_800);
and U212 (N_212,In_947,In_371);
xor U213 (N_213,In_1478,In_563);
or U214 (N_214,In_900,In_387);
and U215 (N_215,In_425,In_1174);
xor U216 (N_216,In_367,In_1160);
or U217 (N_217,In_1189,In_246);
nand U218 (N_218,In_894,In_265);
and U219 (N_219,In_535,In_223);
xnor U220 (N_220,In_365,In_389);
and U221 (N_221,In_1396,In_1330);
nor U222 (N_222,In_966,In_183);
or U223 (N_223,In_642,In_637);
or U224 (N_224,In_940,In_768);
nand U225 (N_225,In_987,In_684);
xnor U226 (N_226,In_1361,In_17);
and U227 (N_227,In_1064,In_783);
xor U228 (N_228,In_1304,In_615);
and U229 (N_229,In_256,In_1293);
xnor U230 (N_230,In_1456,In_624);
nor U231 (N_231,In_791,In_414);
or U232 (N_232,In_1069,In_648);
and U233 (N_233,In_1347,In_676);
nand U234 (N_234,In_1277,In_715);
xor U235 (N_235,In_356,In_551);
nand U236 (N_236,In_1440,In_443);
nor U237 (N_237,In_1199,In_1212);
nor U238 (N_238,In_1168,In_446);
xor U239 (N_239,In_210,In_718);
or U240 (N_240,In_603,In_898);
or U241 (N_241,In_316,In_381);
nand U242 (N_242,In_1297,In_1214);
or U243 (N_243,In_553,In_844);
nand U244 (N_244,In_1181,In_1146);
xor U245 (N_245,In_755,In_453);
xor U246 (N_246,In_85,In_143);
nand U247 (N_247,In_776,In_651);
or U248 (N_248,In_1060,In_427);
nand U249 (N_249,In_868,In_1496);
or U250 (N_250,In_579,In_75);
xnor U251 (N_251,In_695,In_217);
xnor U252 (N_252,In_225,In_1001);
and U253 (N_253,In_753,In_86);
or U254 (N_254,In_230,In_1118);
and U255 (N_255,In_439,In_46);
and U256 (N_256,In_193,In_1244);
and U257 (N_257,In_1315,In_125);
nor U258 (N_258,In_1165,In_906);
nor U259 (N_259,In_1056,In_1260);
and U260 (N_260,In_1498,In_283);
and U261 (N_261,In_409,In_479);
nand U262 (N_262,In_380,In_818);
or U263 (N_263,In_407,In_233);
or U264 (N_264,In_1218,In_368);
xnor U265 (N_265,In_294,In_995);
xor U266 (N_266,In_1449,In_1009);
nor U267 (N_267,In_1153,In_875);
nor U268 (N_268,In_632,In_278);
xnor U269 (N_269,In_803,In_279);
or U270 (N_270,In_1258,In_113);
nand U271 (N_271,In_1284,In_762);
nor U272 (N_272,In_1402,In_752);
nand U273 (N_273,In_618,In_41);
xor U274 (N_274,In_557,In_290);
nand U275 (N_275,In_1427,In_1243);
nor U276 (N_276,In_1494,In_58);
nor U277 (N_277,In_493,In_821);
nand U278 (N_278,In_202,In_395);
nor U279 (N_279,In_1457,In_1455);
or U280 (N_280,In_737,In_406);
nand U281 (N_281,In_282,In_819);
nand U282 (N_282,In_499,In_696);
xor U283 (N_283,In_1005,In_212);
or U284 (N_284,In_239,In_299);
nand U285 (N_285,In_664,In_1107);
nand U286 (N_286,In_214,In_1038);
nor U287 (N_287,In_996,In_1292);
nor U288 (N_288,In_1353,In_592);
nand U289 (N_289,In_318,In_1045);
nor U290 (N_290,In_620,In_1429);
or U291 (N_291,In_529,In_598);
xor U292 (N_292,In_1020,In_866);
nor U293 (N_293,In_1251,In_743);
xor U294 (N_294,In_1130,In_1460);
nand U295 (N_295,In_1159,In_594);
nor U296 (N_296,In_128,In_787);
or U297 (N_297,In_31,In_886);
nor U298 (N_298,In_33,In_922);
and U299 (N_299,In_336,In_519);
nor U300 (N_300,In_540,In_851);
xnor U301 (N_301,In_1231,In_838);
and U302 (N_302,In_1088,In_1324);
and U303 (N_303,In_779,In_528);
and U304 (N_304,In_1070,In_53);
or U305 (N_305,In_758,In_1409);
nand U306 (N_306,In_830,In_870);
nand U307 (N_307,In_1063,In_1310);
xor U308 (N_308,In_1015,In_481);
nor U309 (N_309,In_335,In_530);
nor U310 (N_310,In_357,In_719);
nand U311 (N_311,In_244,In_1380);
xor U312 (N_312,In_634,In_236);
and U313 (N_313,In_802,In_1197);
nand U314 (N_314,In_300,In_1177);
and U315 (N_315,In_1300,In_913);
or U316 (N_316,In_492,In_306);
or U317 (N_317,In_1079,In_724);
and U318 (N_318,In_576,In_677);
nor U319 (N_319,In_687,In_1320);
or U320 (N_320,In_549,In_80);
nand U321 (N_321,In_537,In_527);
xor U322 (N_322,In_932,In_276);
xor U323 (N_323,In_628,In_774);
xnor U324 (N_324,In_958,In_1473);
and U325 (N_325,In_301,In_827);
and U326 (N_326,In_1333,In_794);
and U327 (N_327,In_206,In_1376);
and U328 (N_328,In_504,In_284);
and U329 (N_329,In_272,In_523);
xor U330 (N_330,In_34,In_1366);
xnor U331 (N_331,In_426,In_1481);
xnor U332 (N_332,In_872,In_1040);
xnor U333 (N_333,In_207,In_669);
and U334 (N_334,In_266,In_1493);
and U335 (N_335,In_494,In_896);
nor U336 (N_336,In_1128,In_525);
and U337 (N_337,In_1175,In_792);
xor U338 (N_338,In_78,In_1051);
nand U339 (N_339,In_554,In_428);
nand U340 (N_340,In_984,In_1388);
xnor U341 (N_341,In_934,In_1013);
xor U342 (N_342,In_1375,In_241);
nand U343 (N_343,In_319,In_975);
or U344 (N_344,In_234,In_374);
or U345 (N_345,In_1291,In_296);
nor U346 (N_346,In_369,In_785);
nor U347 (N_347,In_355,In_725);
and U348 (N_348,In_40,In_954);
and U349 (N_349,In_150,In_1467);
nand U350 (N_350,In_1201,In_1049);
nor U351 (N_351,In_569,In_501);
or U352 (N_352,In_775,In_1135);
nor U353 (N_353,In_482,In_285);
nand U354 (N_354,In_221,In_1372);
or U355 (N_355,In_961,In_978);
xnor U356 (N_356,In_490,In_1190);
and U357 (N_357,In_1022,In_372);
and U358 (N_358,In_544,In_1451);
nand U359 (N_359,In_1363,In_789);
or U360 (N_360,In_983,In_976);
nand U361 (N_361,In_8,In_673);
xnor U362 (N_362,In_1359,In_968);
and U363 (N_363,In_24,In_1425);
and U364 (N_364,In_1106,In_795);
or U365 (N_365,In_190,In_62);
nand U366 (N_366,In_438,In_333);
nor U367 (N_367,In_1321,In_629);
nor U368 (N_368,In_55,In_0);
nand U369 (N_369,In_1263,In_1432);
or U370 (N_370,In_418,In_185);
nand U371 (N_371,In_507,In_1205);
or U372 (N_372,In_1445,In_638);
nor U373 (N_373,In_1499,In_235);
nand U374 (N_374,In_30,In_444);
nand U375 (N_375,In_1006,In_1453);
xnor U376 (N_376,In_1109,In_502);
and U377 (N_377,In_744,In_204);
nand U378 (N_378,In_552,In_255);
xnor U379 (N_379,In_1061,In_464);
nor U380 (N_380,In_1129,In_751);
or U381 (N_381,In_156,In_1295);
or U382 (N_382,In_1368,In_1410);
nand U383 (N_383,In_1477,In_1074);
nand U384 (N_384,In_972,In_435);
or U385 (N_385,In_609,In_1166);
nand U386 (N_386,In_588,In_842);
nand U387 (N_387,In_176,In_1351);
xor U388 (N_388,In_506,In_449);
or U389 (N_389,In_678,In_1399);
or U390 (N_390,In_1171,In_1450);
xnor U391 (N_391,In_180,In_897);
or U392 (N_392,In_191,In_82);
or U393 (N_393,In_599,In_668);
nor U394 (N_394,In_1308,In_867);
nor U395 (N_395,In_370,In_415);
and U396 (N_396,In_1272,In_1210);
nor U397 (N_397,In_936,In_1374);
nor U398 (N_398,In_121,In_1145);
and U399 (N_399,In_837,In_1469);
or U400 (N_400,In_388,In_705);
or U401 (N_401,In_649,In_1491);
nor U402 (N_402,In_697,In_662);
nand U403 (N_403,In_993,In_432);
nor U404 (N_404,In_350,In_923);
and U405 (N_405,In_43,In_222);
and U406 (N_406,In_1365,In_965);
or U407 (N_407,In_1401,In_1209);
and U408 (N_408,In_1395,In_116);
or U409 (N_409,In_630,In_1137);
and U410 (N_410,In_666,In_32);
nand U411 (N_411,In_835,In_571);
and U412 (N_412,In_302,In_312);
nand U413 (N_413,In_305,In_1085);
nand U414 (N_414,In_1329,In_197);
and U415 (N_415,In_382,In_1475);
and U416 (N_416,In_846,In_262);
nand U417 (N_417,In_714,In_413);
xnor U418 (N_418,In_700,In_1021);
nor U419 (N_419,In_811,In_763);
and U420 (N_420,In_118,In_1398);
nand U421 (N_421,In_1220,In_1334);
and U422 (N_422,In_484,In_344);
nand U423 (N_423,In_65,In_1068);
or U424 (N_424,In_331,In_655);
and U425 (N_425,In_52,In_805);
xnor U426 (N_426,In_1030,In_394);
nand U427 (N_427,In_773,In_912);
or U428 (N_428,In_722,In_192);
xnor U429 (N_429,In_447,In_1459);
or U430 (N_430,In_570,In_136);
nor U431 (N_431,In_1237,In_539);
xnor U432 (N_432,In_1050,In_1301);
nand U433 (N_433,In_237,In_781);
or U434 (N_434,In_778,In_1224);
nor U435 (N_435,In_334,In_475);
or U436 (N_436,In_1043,In_1267);
and U437 (N_437,In_1240,In_216);
nor U438 (N_438,In_203,In_1125);
and U439 (N_439,In_988,In_1474);
nor U440 (N_440,In_308,In_1317);
nor U441 (N_441,In_390,In_352);
or U442 (N_442,In_309,In_83);
nand U443 (N_443,In_583,In_521);
nand U444 (N_444,In_860,In_734);
nor U445 (N_445,In_27,In_1492);
or U446 (N_446,In_1253,In_699);
xnor U447 (N_447,In_1417,In_1486);
or U448 (N_448,In_249,In_955);
xor U449 (N_449,In_397,In_1423);
nor U450 (N_450,In_383,In_1018);
and U451 (N_451,In_119,In_1256);
xor U452 (N_452,In_298,In_1017);
nand U453 (N_453,In_814,In_1319);
xnor U454 (N_454,In_50,In_1495);
nand U455 (N_455,In_1198,In_680);
and U456 (N_456,In_891,In_104);
and U457 (N_457,In_1322,In_1226);
nand U458 (N_458,In_829,In_1196);
nand U459 (N_459,In_1191,In_963);
or U460 (N_460,In_56,In_433);
xor U461 (N_461,In_96,In_177);
or U462 (N_462,In_1344,In_226);
xor U463 (N_463,In_1241,In_323);
and U464 (N_464,In_654,In_582);
nand U465 (N_465,In_1489,In_1142);
nand U466 (N_466,In_10,In_941);
nand U467 (N_467,In_1078,In_915);
and U468 (N_468,In_252,In_89);
nor U469 (N_469,In_399,In_420);
nor U470 (N_470,In_636,In_1007);
or U471 (N_471,In_1348,In_469);
nand U472 (N_472,In_723,In_1161);
xnor U473 (N_473,In_4,In_901);
or U474 (N_474,In_895,In_717);
xor U475 (N_475,In_111,In_1099);
or U476 (N_476,In_665,In_35);
and U477 (N_477,In_22,In_644);
and U478 (N_478,In_681,In_1326);
xnor U479 (N_479,In_311,In_1394);
or U480 (N_480,In_1173,In_926);
xnor U481 (N_481,In_1025,In_566);
nand U482 (N_482,In_292,In_633);
xnor U483 (N_483,In_1100,In_709);
nand U484 (N_484,In_1370,In_1433);
or U485 (N_485,In_1012,In_248);
nand U486 (N_486,In_267,In_1337);
or U487 (N_487,In_87,In_126);
and U488 (N_488,In_513,In_2);
and U489 (N_489,In_253,In_683);
and U490 (N_490,In_105,In_1105);
nor U491 (N_491,In_1325,In_756);
nor U492 (N_492,In_921,In_883);
nand U493 (N_493,In_1097,In_112);
and U494 (N_494,In_393,In_417);
nand U495 (N_495,In_462,In_876);
nand U496 (N_496,In_386,In_1444);
xor U497 (N_497,In_1031,In_1208);
xnor U498 (N_498,In_1468,In_1430);
xnor U499 (N_499,In_270,In_459);
nand U500 (N_500,In_47,In_1397);
nand U501 (N_501,In_1110,In_646);
or U502 (N_502,In_610,In_1247);
nor U503 (N_503,In_992,In_1255);
xor U504 (N_504,In_581,In_920);
and U505 (N_505,In_760,In_1354);
or U506 (N_506,In_575,In_232);
nor U507 (N_507,In_640,In_974);
and U508 (N_508,In_596,In_478);
xor U509 (N_509,In_144,In_799);
xor U510 (N_510,In_1158,In_1314);
and U511 (N_511,In_1184,In_1227);
nor U512 (N_512,In_845,In_472);
nor U513 (N_513,In_1278,In_392);
or U514 (N_514,In_198,In_454);
or U515 (N_515,In_985,In_146);
xor U516 (N_516,In_1225,In_606);
nor U517 (N_517,In_950,In_1195);
xor U518 (N_518,In_869,In_509);
and U519 (N_519,In_1090,In_1014);
xor U520 (N_520,In_480,In_852);
or U521 (N_521,In_1183,In_547);
and U522 (N_522,In_1233,In_375);
and U523 (N_523,In_1441,In_254);
or U524 (N_524,In_1352,In_1246);
xor U525 (N_525,In_405,In_64);
nor U526 (N_526,In_132,In_1420);
or U527 (N_527,In_275,In_574);
xnor U528 (N_528,In_946,In_661);
nand U529 (N_529,In_1259,In_103);
nor U530 (N_530,In_1270,In_1144);
nor U531 (N_531,In_1066,In_679);
or U532 (N_532,In_515,In_1143);
or U533 (N_533,In_782,In_297);
nand U534 (N_534,In_749,In_1151);
or U535 (N_535,In_120,In_1476);
nand U536 (N_536,In_1328,In_518);
nand U537 (N_537,In_477,In_806);
xnor U538 (N_538,In_809,In_1274);
and U539 (N_539,In_419,In_194);
nand U540 (N_540,In_1126,In_84);
or U541 (N_541,In_184,In_1230);
xnor U542 (N_542,In_1415,In_468);
and U543 (N_543,In_969,In_1408);
xor U544 (N_544,In_326,In_604);
nor U545 (N_545,In_1072,In_663);
nand U546 (N_546,In_1266,In_670);
or U547 (N_547,In_1235,In_793);
nand U548 (N_548,In_268,In_741);
xor U549 (N_549,In_277,In_213);
and U550 (N_550,In_997,In_467);
or U551 (N_551,In_750,In_970);
and U552 (N_552,In_12,In_81);
or U553 (N_553,In_88,In_115);
nand U554 (N_554,In_568,In_702);
or U555 (N_555,In_141,In_1400);
xnor U556 (N_556,In_708,In_769);
or U557 (N_557,In_330,In_720);
or U558 (N_558,In_488,In_224);
nor U559 (N_559,In_1369,In_1091);
or U560 (N_560,In_907,In_884);
and U561 (N_561,In_1223,In_353);
and U562 (N_562,In_1472,In_422);
nand U563 (N_563,In_130,In_1254);
nand U564 (N_564,In_1290,In_261);
and U565 (N_565,In_77,In_79);
nand U566 (N_566,In_69,In_1419);
xor U567 (N_567,In_1162,In_831);
nand U568 (N_568,In_424,In_489);
or U569 (N_569,In_1306,In_1057);
nand U570 (N_570,In_1356,In_1261);
xnor U571 (N_571,In_1178,In_72);
and U572 (N_572,In_508,In_385);
and U573 (N_573,In_195,In_919);
or U574 (N_574,In_325,In_560);
nor U575 (N_575,In_1081,In_18);
nand U576 (N_576,In_825,In_727);
and U577 (N_577,In_461,In_1219);
xor U578 (N_578,In_73,In_1047);
nand U579 (N_579,In_329,In_1108);
xnor U580 (N_580,In_1065,In_179);
xnor U581 (N_581,In_1269,In_1217);
xnor U582 (N_582,In_209,In_770);
and U583 (N_583,In_973,In_960);
xor U584 (N_584,In_595,In_1116);
nor U585 (N_585,In_707,In_567);
and U586 (N_586,In_402,In_1422);
nand U587 (N_587,In_1488,In_944);
nand U588 (N_588,In_1221,In_110);
or U589 (N_589,In_1327,In_1392);
nand U590 (N_590,In_1268,In_1172);
nand U591 (N_591,In_1332,In_959);
nor U592 (N_592,In_815,In_231);
or U593 (N_593,In_90,In_1412);
xnor U594 (N_594,In_672,In_780);
nor U595 (N_595,In_1390,In_124);
or U596 (N_596,In_448,In_1075);
nor U597 (N_597,In_605,In_1265);
xor U598 (N_598,In_1117,In_411);
xnor U599 (N_599,In_1150,In_487);
or U600 (N_600,In_1052,In_613);
or U601 (N_601,In_145,In_764);
nor U602 (N_602,In_1216,In_1393);
nand U603 (N_603,In_1027,In_1275);
or U604 (N_604,In_410,In_474);
nor U605 (N_605,In_1262,In_698);
nand U606 (N_606,In_1305,In_362);
or U607 (N_607,In_688,In_658);
nand U608 (N_608,In_21,In_205);
xnor U609 (N_609,In_625,In_712);
nand U610 (N_610,In_328,In_622);
nor U611 (N_611,In_559,In_647);
xor U612 (N_612,In_1123,In_154);
or U613 (N_613,In_1073,In_98);
nand U614 (N_614,In_1192,In_131);
nor U615 (N_615,In_456,In_160);
or U616 (N_616,In_813,In_45);
nand U617 (N_617,In_1082,In_347);
xor U618 (N_618,In_1193,In_1257);
nor U619 (N_619,In_1010,In_772);
nor U620 (N_620,In_391,In_864);
nand U621 (N_621,In_879,In_421);
xor U622 (N_622,In_1236,In_1406);
and U623 (N_623,In_1136,In_1381);
xor U624 (N_624,In_460,In_1490);
nor U625 (N_625,In_1355,In_652);
or U626 (N_626,In_784,In_457);
nor U627 (N_627,In_607,In_614);
and U628 (N_628,In_590,In_473);
xnor U629 (N_629,In_398,In_788);
nor U630 (N_630,In_384,In_740);
and U631 (N_631,In_878,In_1238);
and U632 (N_632,In_796,In_1452);
and U633 (N_633,In_263,In_1282);
nand U634 (N_634,In_44,In_228);
or U635 (N_635,In_1207,In_1076);
and U636 (N_636,In_859,In_155);
and U637 (N_637,In_930,In_48);
nand U638 (N_638,In_208,In_854);
nand U639 (N_639,In_408,In_1487);
xor U640 (N_640,In_1008,In_495);
and U641 (N_641,In_1138,In_820);
xor U642 (N_642,In_558,In_887);
xnor U643 (N_643,In_436,In_1379);
nand U644 (N_644,In_931,In_516);
and U645 (N_645,In_166,In_754);
or U646 (N_646,In_281,In_1087);
nand U647 (N_647,In_127,In_99);
or U648 (N_648,In_199,In_1002);
nand U649 (N_649,In_943,In_1071);
or U650 (N_650,In_1058,In_533);
nor U651 (N_651,In_538,In_616);
nand U652 (N_652,In_1413,In_1084);
nand U653 (N_653,In_227,In_3);
and U654 (N_654,In_242,In_631);
nor U655 (N_655,In_171,In_1046);
nand U656 (N_656,In_710,In_149);
and U657 (N_657,In_218,In_476);
and U658 (N_658,In_1180,In_1169);
xnor U659 (N_659,In_147,In_97);
nand U660 (N_660,In_1371,In_1360);
nand U661 (N_661,In_1435,In_824);
or U662 (N_662,In_1132,In_546);
nand U663 (N_663,In_1120,In_790);
and U664 (N_664,In_536,In_1405);
nand U665 (N_665,In_882,In_1296);
xnor U666 (N_666,In_1000,In_816);
or U667 (N_667,In_289,In_1048);
or U668 (N_668,In_580,In_437);
nand U669 (N_669,In_694,In_1188);
xor U670 (N_670,In_106,In_1093);
xor U671 (N_671,In_671,In_49);
nor U672 (N_672,In_1302,In_1179);
nand U673 (N_673,In_703,In_54);
nor U674 (N_674,In_1309,In_341);
nand U675 (N_675,In_359,In_348);
or U676 (N_676,In_511,In_817);
nor U677 (N_677,In_135,In_994);
or U678 (N_678,In_822,In_307);
nor U679 (N_679,In_354,In_986);
nor U680 (N_680,In_999,In_807);
nor U681 (N_681,In_1111,In_808);
nor U682 (N_682,In_400,In_1431);
nand U683 (N_683,In_250,In_608);
and U684 (N_684,In_450,In_1229);
xnor U685 (N_685,In_765,In_342);
and U686 (N_686,In_555,In_1316);
nor U687 (N_687,In_361,In_25);
nand U688 (N_688,In_1484,In_1303);
xnor U689 (N_689,In_1331,In_1086);
and U690 (N_690,In_1340,In_600);
and U691 (N_691,In_163,In_736);
xnor U692 (N_692,In_738,In_1289);
nand U693 (N_693,In_364,In_170);
xnor U694 (N_694,In_786,In_1311);
or U695 (N_695,In_733,In_288);
xor U696 (N_696,In_1362,In_500);
and U697 (N_697,In_1461,In_925);
nor U698 (N_698,In_939,In_310);
nor U699 (N_699,In_572,In_260);
nand U700 (N_700,In_1101,In_881);
xor U701 (N_701,In_251,In_1053);
and U702 (N_702,In_510,In_522);
xor U703 (N_703,In_158,In_761);
nand U704 (N_704,In_412,In_545);
and U705 (N_705,In_1446,In_801);
nand U706 (N_706,In_1285,In_716);
nor U707 (N_707,In_863,In_1448);
or U708 (N_708,In_514,In_29);
nor U709 (N_709,In_1122,In_1156);
xnor U710 (N_710,In_1428,In_1248);
and U711 (N_711,In_1003,In_602);
and U712 (N_712,In_107,In_229);
nand U713 (N_713,In_403,In_161);
xnor U714 (N_714,In_441,In_721);
or U715 (N_715,In_486,In_5);
nor U716 (N_716,In_873,In_1206);
nand U717 (N_717,In_497,In_1194);
or U718 (N_718,In_812,In_832);
nor U719 (N_719,In_1442,In_990);
xor U720 (N_720,In_1357,In_742);
or U721 (N_721,In_766,In_731);
and U722 (N_722,In_938,In_59);
xor U723 (N_723,In_1480,In_442);
or U724 (N_724,In_240,In_162);
nand U725 (N_725,In_917,In_101);
and U726 (N_726,In_15,In_1286);
xor U727 (N_727,In_1280,In_561);
and U728 (N_728,In_134,In_964);
nand U729 (N_729,In_1098,In_611);
nand U730 (N_730,In_1335,In_1462);
or U731 (N_731,In_114,In_840);
or U732 (N_732,In_320,In_26);
nand U733 (N_733,In_645,In_63);
or U734 (N_734,In_1350,In_346);
nand U735 (N_735,In_1264,In_1026);
nor U736 (N_736,In_245,In_140);
xnor U737 (N_737,In_485,In_601);
nor U738 (N_738,In_1114,In_186);
nor U739 (N_739,In_434,In_1483);
or U740 (N_740,In_430,In_238);
xnor U741 (N_741,In_849,In_565);
xor U742 (N_742,In_11,In_351);
nor U743 (N_743,In_1377,In_200);
and U744 (N_744,In_1103,In_1323);
or U745 (N_745,In_138,In_1139);
and U746 (N_746,In_701,In_159);
or U747 (N_747,In_1112,In_379);
or U748 (N_748,In_1034,In_431);
and U749 (N_749,In_1019,In_1102);
nor U750 (N_750,In_776,In_1010);
and U751 (N_751,In_543,In_846);
and U752 (N_752,In_259,In_883);
or U753 (N_753,In_1337,In_1158);
and U754 (N_754,In_1044,In_837);
nand U755 (N_755,In_1166,In_1383);
and U756 (N_756,In_1084,In_1294);
xnor U757 (N_757,In_567,In_752);
nor U758 (N_758,In_243,In_1135);
nor U759 (N_759,In_61,In_661);
nor U760 (N_760,In_1330,In_942);
or U761 (N_761,In_790,In_646);
and U762 (N_762,In_908,In_1047);
nand U763 (N_763,In_406,In_11);
nor U764 (N_764,In_1377,In_1464);
nand U765 (N_765,In_57,In_5);
nand U766 (N_766,In_755,In_623);
and U767 (N_767,In_669,In_1292);
nand U768 (N_768,In_401,In_44);
nand U769 (N_769,In_796,In_189);
nand U770 (N_770,In_941,In_585);
nand U771 (N_771,In_45,In_895);
xnor U772 (N_772,In_1044,In_1012);
nor U773 (N_773,In_496,In_1076);
nand U774 (N_774,In_164,In_250);
and U775 (N_775,In_208,In_1483);
xnor U776 (N_776,In_403,In_699);
and U777 (N_777,In_655,In_1276);
or U778 (N_778,In_1097,In_1366);
xor U779 (N_779,In_887,In_1277);
nor U780 (N_780,In_1150,In_807);
or U781 (N_781,In_424,In_1445);
xor U782 (N_782,In_575,In_51);
and U783 (N_783,In_715,In_832);
or U784 (N_784,In_806,In_355);
or U785 (N_785,In_570,In_1230);
nand U786 (N_786,In_1331,In_330);
nand U787 (N_787,In_1405,In_94);
nor U788 (N_788,In_372,In_1269);
nand U789 (N_789,In_430,In_1090);
nor U790 (N_790,In_794,In_852);
nor U791 (N_791,In_396,In_231);
and U792 (N_792,In_128,In_579);
and U793 (N_793,In_832,In_189);
nor U794 (N_794,In_1139,In_520);
xor U795 (N_795,In_336,In_475);
nor U796 (N_796,In_604,In_268);
nor U797 (N_797,In_231,In_1219);
and U798 (N_798,In_413,In_737);
xor U799 (N_799,In_1230,In_265);
nor U800 (N_800,In_1039,In_589);
and U801 (N_801,In_1004,In_1144);
nand U802 (N_802,In_1428,In_522);
nand U803 (N_803,In_653,In_106);
and U804 (N_804,In_580,In_635);
nor U805 (N_805,In_1029,In_316);
and U806 (N_806,In_1374,In_34);
and U807 (N_807,In_732,In_625);
nand U808 (N_808,In_558,In_1045);
nand U809 (N_809,In_1486,In_1239);
or U810 (N_810,In_723,In_862);
or U811 (N_811,In_440,In_1214);
nor U812 (N_812,In_1381,In_775);
nand U813 (N_813,In_535,In_30);
xor U814 (N_814,In_566,In_1331);
xnor U815 (N_815,In_884,In_1046);
and U816 (N_816,In_719,In_352);
and U817 (N_817,In_755,In_50);
xnor U818 (N_818,In_1350,In_40);
xnor U819 (N_819,In_68,In_496);
xor U820 (N_820,In_1088,In_1285);
nor U821 (N_821,In_303,In_758);
and U822 (N_822,In_361,In_478);
and U823 (N_823,In_651,In_1194);
and U824 (N_824,In_227,In_1122);
xor U825 (N_825,In_488,In_593);
nor U826 (N_826,In_1309,In_1486);
nor U827 (N_827,In_1444,In_1112);
nand U828 (N_828,In_986,In_786);
and U829 (N_829,In_1233,In_652);
and U830 (N_830,In_174,In_469);
and U831 (N_831,In_689,In_966);
nor U832 (N_832,In_1361,In_1137);
xor U833 (N_833,In_874,In_855);
xnor U834 (N_834,In_923,In_179);
or U835 (N_835,In_1015,In_1192);
and U836 (N_836,In_968,In_445);
xor U837 (N_837,In_930,In_142);
xor U838 (N_838,In_684,In_570);
nand U839 (N_839,In_174,In_1391);
nand U840 (N_840,In_619,In_381);
and U841 (N_841,In_738,In_644);
nor U842 (N_842,In_1211,In_981);
xor U843 (N_843,In_845,In_380);
and U844 (N_844,In_907,In_275);
and U845 (N_845,In_729,In_1249);
nor U846 (N_846,In_914,In_841);
and U847 (N_847,In_139,In_753);
and U848 (N_848,In_112,In_620);
nand U849 (N_849,In_468,In_1103);
nor U850 (N_850,In_184,In_1078);
nor U851 (N_851,In_1394,In_1437);
xnor U852 (N_852,In_350,In_755);
and U853 (N_853,In_744,In_127);
nand U854 (N_854,In_915,In_236);
or U855 (N_855,In_235,In_1360);
xnor U856 (N_856,In_984,In_369);
nand U857 (N_857,In_674,In_789);
and U858 (N_858,In_302,In_1014);
nor U859 (N_859,In_948,In_568);
and U860 (N_860,In_170,In_571);
and U861 (N_861,In_1185,In_837);
nor U862 (N_862,In_273,In_838);
nand U863 (N_863,In_712,In_503);
and U864 (N_864,In_220,In_660);
nor U865 (N_865,In_864,In_1323);
nand U866 (N_866,In_234,In_86);
or U867 (N_867,In_1007,In_13);
or U868 (N_868,In_631,In_1130);
nand U869 (N_869,In_493,In_990);
nand U870 (N_870,In_1314,In_865);
and U871 (N_871,In_290,In_204);
and U872 (N_872,In_241,In_609);
nor U873 (N_873,In_303,In_140);
or U874 (N_874,In_98,In_1380);
and U875 (N_875,In_903,In_568);
nor U876 (N_876,In_404,In_1325);
or U877 (N_877,In_58,In_1004);
nand U878 (N_878,In_368,In_1029);
xnor U879 (N_879,In_1473,In_51);
nor U880 (N_880,In_513,In_1265);
and U881 (N_881,In_1191,In_267);
nand U882 (N_882,In_81,In_289);
or U883 (N_883,In_1186,In_1462);
and U884 (N_884,In_914,In_943);
or U885 (N_885,In_439,In_451);
xnor U886 (N_886,In_48,In_154);
nand U887 (N_887,In_1473,In_61);
nor U888 (N_888,In_1494,In_1457);
nand U889 (N_889,In_743,In_1093);
xnor U890 (N_890,In_1407,In_452);
xor U891 (N_891,In_768,In_1156);
and U892 (N_892,In_50,In_325);
and U893 (N_893,In_248,In_585);
nand U894 (N_894,In_227,In_1026);
nand U895 (N_895,In_1134,In_784);
xor U896 (N_896,In_1130,In_907);
or U897 (N_897,In_1223,In_18);
nand U898 (N_898,In_168,In_821);
and U899 (N_899,In_1164,In_85);
nand U900 (N_900,In_372,In_301);
or U901 (N_901,In_346,In_194);
xnor U902 (N_902,In_800,In_1427);
xnor U903 (N_903,In_729,In_367);
xor U904 (N_904,In_1,In_1349);
nand U905 (N_905,In_723,In_1223);
and U906 (N_906,In_1296,In_236);
nor U907 (N_907,In_176,In_880);
nor U908 (N_908,In_835,In_647);
or U909 (N_909,In_661,In_975);
or U910 (N_910,In_1243,In_1474);
or U911 (N_911,In_1353,In_158);
nor U912 (N_912,In_1294,In_1055);
nand U913 (N_913,In_722,In_1267);
and U914 (N_914,In_879,In_1325);
and U915 (N_915,In_1038,In_1464);
nor U916 (N_916,In_303,In_1363);
xnor U917 (N_917,In_940,In_531);
nor U918 (N_918,In_1053,In_569);
xnor U919 (N_919,In_541,In_515);
or U920 (N_920,In_742,In_688);
and U921 (N_921,In_1385,In_875);
nor U922 (N_922,In_10,In_314);
and U923 (N_923,In_770,In_505);
nor U924 (N_924,In_1107,In_33);
or U925 (N_925,In_421,In_18);
xnor U926 (N_926,In_1311,In_85);
and U927 (N_927,In_45,In_953);
and U928 (N_928,In_31,In_54);
xor U929 (N_929,In_1225,In_1470);
and U930 (N_930,In_63,In_1220);
nand U931 (N_931,In_601,In_832);
nand U932 (N_932,In_91,In_198);
nand U933 (N_933,In_188,In_753);
nand U934 (N_934,In_314,In_1114);
nor U935 (N_935,In_1127,In_70);
or U936 (N_936,In_1239,In_1383);
nor U937 (N_937,In_346,In_1431);
nand U938 (N_938,In_896,In_1216);
nor U939 (N_939,In_1188,In_376);
nand U940 (N_940,In_689,In_337);
or U941 (N_941,In_1428,In_845);
xor U942 (N_942,In_480,In_825);
and U943 (N_943,In_969,In_531);
or U944 (N_944,In_1181,In_1090);
xnor U945 (N_945,In_1474,In_435);
or U946 (N_946,In_1434,In_1361);
nor U947 (N_947,In_1073,In_1000);
and U948 (N_948,In_147,In_444);
and U949 (N_949,In_867,In_163);
nand U950 (N_950,In_201,In_95);
and U951 (N_951,In_417,In_500);
nand U952 (N_952,In_123,In_1146);
nor U953 (N_953,In_1301,In_314);
and U954 (N_954,In_1125,In_31);
nor U955 (N_955,In_31,In_717);
or U956 (N_956,In_1053,In_642);
and U957 (N_957,In_1436,In_743);
nor U958 (N_958,In_441,In_509);
or U959 (N_959,In_1003,In_1178);
nor U960 (N_960,In_768,In_1296);
and U961 (N_961,In_997,In_273);
nand U962 (N_962,In_453,In_822);
and U963 (N_963,In_917,In_80);
or U964 (N_964,In_319,In_608);
xnor U965 (N_965,In_699,In_117);
or U966 (N_966,In_1471,In_358);
nand U967 (N_967,In_1291,In_963);
xor U968 (N_968,In_975,In_845);
and U969 (N_969,In_872,In_758);
and U970 (N_970,In_660,In_1271);
and U971 (N_971,In_1268,In_534);
and U972 (N_972,In_826,In_943);
or U973 (N_973,In_132,In_921);
and U974 (N_974,In_1235,In_217);
nand U975 (N_975,In_1490,In_1253);
nand U976 (N_976,In_259,In_579);
or U977 (N_977,In_1202,In_264);
nand U978 (N_978,In_841,In_1032);
or U979 (N_979,In_602,In_1313);
nand U980 (N_980,In_289,In_336);
nor U981 (N_981,In_1033,In_1006);
and U982 (N_982,In_496,In_602);
nor U983 (N_983,In_445,In_1208);
nand U984 (N_984,In_468,In_554);
nor U985 (N_985,In_148,In_536);
nor U986 (N_986,In_721,In_461);
nand U987 (N_987,In_229,In_200);
nor U988 (N_988,In_1411,In_650);
or U989 (N_989,In_1404,In_595);
nor U990 (N_990,In_1152,In_988);
nand U991 (N_991,In_1302,In_541);
and U992 (N_992,In_925,In_309);
nand U993 (N_993,In_1258,In_1035);
nand U994 (N_994,In_1290,In_896);
or U995 (N_995,In_271,In_1191);
xnor U996 (N_996,In_239,In_90);
xor U997 (N_997,In_621,In_971);
or U998 (N_998,In_1380,In_1171);
or U999 (N_999,In_951,In_884);
nor U1000 (N_1000,In_1361,In_681);
nand U1001 (N_1001,In_984,In_1277);
and U1002 (N_1002,In_1065,In_1009);
xor U1003 (N_1003,In_495,In_1448);
xnor U1004 (N_1004,In_338,In_832);
and U1005 (N_1005,In_1063,In_355);
nor U1006 (N_1006,In_211,In_536);
nor U1007 (N_1007,In_502,In_137);
or U1008 (N_1008,In_892,In_398);
nand U1009 (N_1009,In_322,In_383);
and U1010 (N_1010,In_449,In_3);
nand U1011 (N_1011,In_1092,In_1159);
and U1012 (N_1012,In_1457,In_378);
nor U1013 (N_1013,In_1205,In_1057);
nor U1014 (N_1014,In_327,In_283);
or U1015 (N_1015,In_425,In_262);
or U1016 (N_1016,In_1321,In_443);
or U1017 (N_1017,In_1115,In_324);
nand U1018 (N_1018,In_1234,In_688);
nand U1019 (N_1019,In_795,In_1034);
xor U1020 (N_1020,In_1224,In_490);
and U1021 (N_1021,In_1149,In_1214);
xnor U1022 (N_1022,In_485,In_489);
or U1023 (N_1023,In_774,In_1461);
xor U1024 (N_1024,In_693,In_284);
nand U1025 (N_1025,In_970,In_1280);
or U1026 (N_1026,In_419,In_1416);
or U1027 (N_1027,In_307,In_667);
xor U1028 (N_1028,In_1231,In_631);
nand U1029 (N_1029,In_970,In_267);
and U1030 (N_1030,In_337,In_479);
or U1031 (N_1031,In_1409,In_1380);
and U1032 (N_1032,In_549,In_497);
nand U1033 (N_1033,In_261,In_1073);
nand U1034 (N_1034,In_411,In_306);
xnor U1035 (N_1035,In_983,In_194);
and U1036 (N_1036,In_458,In_1371);
nand U1037 (N_1037,In_1181,In_568);
and U1038 (N_1038,In_1041,In_1499);
or U1039 (N_1039,In_532,In_842);
or U1040 (N_1040,In_322,In_42);
nor U1041 (N_1041,In_976,In_1088);
or U1042 (N_1042,In_1201,In_517);
nand U1043 (N_1043,In_152,In_716);
or U1044 (N_1044,In_1089,In_395);
and U1045 (N_1045,In_1372,In_869);
nor U1046 (N_1046,In_1347,In_769);
xor U1047 (N_1047,In_595,In_131);
xnor U1048 (N_1048,In_51,In_201);
nand U1049 (N_1049,In_1194,In_133);
nor U1050 (N_1050,In_10,In_446);
nand U1051 (N_1051,In_1082,In_687);
and U1052 (N_1052,In_659,In_285);
nor U1053 (N_1053,In_467,In_61);
or U1054 (N_1054,In_1226,In_528);
xnor U1055 (N_1055,In_789,In_1421);
and U1056 (N_1056,In_1405,In_1395);
nand U1057 (N_1057,In_1300,In_399);
and U1058 (N_1058,In_1353,In_1067);
or U1059 (N_1059,In_906,In_999);
xor U1060 (N_1060,In_687,In_356);
xnor U1061 (N_1061,In_1256,In_507);
nand U1062 (N_1062,In_1159,In_1469);
and U1063 (N_1063,In_372,In_778);
xnor U1064 (N_1064,In_764,In_611);
nand U1065 (N_1065,In_1351,In_1418);
and U1066 (N_1066,In_855,In_1407);
nor U1067 (N_1067,In_853,In_1021);
nor U1068 (N_1068,In_1172,In_1066);
nor U1069 (N_1069,In_908,In_167);
and U1070 (N_1070,In_892,In_520);
or U1071 (N_1071,In_1297,In_728);
nor U1072 (N_1072,In_807,In_141);
nor U1073 (N_1073,In_1383,In_814);
nor U1074 (N_1074,In_373,In_587);
and U1075 (N_1075,In_566,In_0);
or U1076 (N_1076,In_1049,In_581);
and U1077 (N_1077,In_1051,In_629);
xor U1078 (N_1078,In_580,In_355);
and U1079 (N_1079,In_856,In_85);
nand U1080 (N_1080,In_1150,In_293);
or U1081 (N_1081,In_1268,In_547);
xor U1082 (N_1082,In_594,In_713);
nor U1083 (N_1083,In_779,In_502);
or U1084 (N_1084,In_83,In_230);
or U1085 (N_1085,In_906,In_169);
or U1086 (N_1086,In_242,In_977);
nand U1087 (N_1087,In_414,In_546);
or U1088 (N_1088,In_752,In_690);
nor U1089 (N_1089,In_1407,In_298);
nand U1090 (N_1090,In_285,In_479);
nor U1091 (N_1091,In_57,In_0);
or U1092 (N_1092,In_237,In_649);
nor U1093 (N_1093,In_1179,In_817);
or U1094 (N_1094,In_951,In_840);
nor U1095 (N_1095,In_983,In_88);
xnor U1096 (N_1096,In_1369,In_202);
nand U1097 (N_1097,In_1184,In_80);
nor U1098 (N_1098,In_1322,In_1390);
nor U1099 (N_1099,In_143,In_834);
nor U1100 (N_1100,In_859,In_1142);
nor U1101 (N_1101,In_684,In_1131);
or U1102 (N_1102,In_1227,In_5);
and U1103 (N_1103,In_452,In_152);
and U1104 (N_1104,In_1356,In_213);
nand U1105 (N_1105,In_181,In_1310);
and U1106 (N_1106,In_52,In_292);
nand U1107 (N_1107,In_15,In_1006);
xnor U1108 (N_1108,In_1320,In_443);
and U1109 (N_1109,In_1377,In_929);
or U1110 (N_1110,In_1295,In_992);
nor U1111 (N_1111,In_583,In_1093);
nor U1112 (N_1112,In_554,In_342);
nor U1113 (N_1113,In_88,In_426);
and U1114 (N_1114,In_1443,In_159);
nand U1115 (N_1115,In_1269,In_202);
nand U1116 (N_1116,In_408,In_409);
xnor U1117 (N_1117,In_511,In_1003);
xnor U1118 (N_1118,In_731,In_1368);
xnor U1119 (N_1119,In_106,In_382);
nand U1120 (N_1120,In_410,In_1393);
or U1121 (N_1121,In_674,In_1062);
nor U1122 (N_1122,In_544,In_824);
or U1123 (N_1123,In_1307,In_148);
nand U1124 (N_1124,In_837,In_1354);
nand U1125 (N_1125,In_1190,In_1308);
or U1126 (N_1126,In_198,In_949);
nand U1127 (N_1127,In_1482,In_1178);
and U1128 (N_1128,In_816,In_944);
nand U1129 (N_1129,In_32,In_1429);
or U1130 (N_1130,In_189,In_1212);
xor U1131 (N_1131,In_289,In_833);
xor U1132 (N_1132,In_1448,In_797);
and U1133 (N_1133,In_1244,In_75);
and U1134 (N_1134,In_1170,In_1202);
nor U1135 (N_1135,In_430,In_1342);
and U1136 (N_1136,In_849,In_97);
or U1137 (N_1137,In_1274,In_546);
nand U1138 (N_1138,In_1038,In_1177);
or U1139 (N_1139,In_828,In_157);
and U1140 (N_1140,In_476,In_573);
or U1141 (N_1141,In_830,In_308);
xor U1142 (N_1142,In_966,In_1268);
xor U1143 (N_1143,In_14,In_922);
xor U1144 (N_1144,In_308,In_343);
and U1145 (N_1145,In_1375,In_653);
and U1146 (N_1146,In_750,In_804);
nand U1147 (N_1147,In_278,In_118);
nand U1148 (N_1148,In_136,In_546);
xor U1149 (N_1149,In_518,In_693);
and U1150 (N_1150,In_1272,In_1302);
or U1151 (N_1151,In_326,In_191);
nor U1152 (N_1152,In_1301,In_564);
nand U1153 (N_1153,In_979,In_448);
nand U1154 (N_1154,In_268,In_1494);
xnor U1155 (N_1155,In_782,In_61);
and U1156 (N_1156,In_562,In_1005);
and U1157 (N_1157,In_116,In_1406);
and U1158 (N_1158,In_211,In_32);
and U1159 (N_1159,In_49,In_175);
xnor U1160 (N_1160,In_925,In_1262);
nor U1161 (N_1161,In_1073,In_947);
or U1162 (N_1162,In_537,In_600);
nand U1163 (N_1163,In_634,In_738);
xnor U1164 (N_1164,In_984,In_683);
nand U1165 (N_1165,In_695,In_273);
and U1166 (N_1166,In_693,In_1370);
xnor U1167 (N_1167,In_87,In_1454);
nor U1168 (N_1168,In_814,In_312);
nand U1169 (N_1169,In_1180,In_445);
xor U1170 (N_1170,In_1361,In_882);
nand U1171 (N_1171,In_353,In_1144);
and U1172 (N_1172,In_391,In_606);
xnor U1173 (N_1173,In_355,In_249);
nor U1174 (N_1174,In_885,In_685);
nor U1175 (N_1175,In_813,In_1439);
xor U1176 (N_1176,In_1235,In_1287);
and U1177 (N_1177,In_11,In_593);
or U1178 (N_1178,In_970,In_1016);
nor U1179 (N_1179,In_867,In_1003);
nand U1180 (N_1180,In_1239,In_1447);
and U1181 (N_1181,In_550,In_1197);
or U1182 (N_1182,In_1144,In_885);
xor U1183 (N_1183,In_539,In_629);
or U1184 (N_1184,In_276,In_320);
nor U1185 (N_1185,In_360,In_919);
and U1186 (N_1186,In_58,In_1402);
xnor U1187 (N_1187,In_972,In_966);
xnor U1188 (N_1188,In_51,In_1218);
nor U1189 (N_1189,In_1292,In_67);
nand U1190 (N_1190,In_1470,In_957);
and U1191 (N_1191,In_341,In_1221);
nand U1192 (N_1192,In_454,In_1038);
nand U1193 (N_1193,In_778,In_1194);
and U1194 (N_1194,In_686,In_1277);
xnor U1195 (N_1195,In_463,In_966);
nand U1196 (N_1196,In_288,In_694);
nor U1197 (N_1197,In_154,In_149);
xnor U1198 (N_1198,In_975,In_770);
xor U1199 (N_1199,In_151,In_460);
xor U1200 (N_1200,In_434,In_680);
xnor U1201 (N_1201,In_6,In_1042);
or U1202 (N_1202,In_1155,In_40);
nand U1203 (N_1203,In_1236,In_6);
nor U1204 (N_1204,In_954,In_1048);
nor U1205 (N_1205,In_1339,In_1126);
nor U1206 (N_1206,In_119,In_275);
nand U1207 (N_1207,In_1353,In_738);
or U1208 (N_1208,In_709,In_1121);
nand U1209 (N_1209,In_1304,In_185);
nor U1210 (N_1210,In_1114,In_1087);
xnor U1211 (N_1211,In_549,In_189);
xor U1212 (N_1212,In_82,In_869);
and U1213 (N_1213,In_1408,In_114);
xnor U1214 (N_1214,In_420,In_752);
xnor U1215 (N_1215,In_431,In_1207);
nand U1216 (N_1216,In_1206,In_1019);
nor U1217 (N_1217,In_452,In_1488);
and U1218 (N_1218,In_1115,In_289);
nand U1219 (N_1219,In_831,In_733);
or U1220 (N_1220,In_1118,In_183);
and U1221 (N_1221,In_1264,In_379);
and U1222 (N_1222,In_1423,In_829);
nor U1223 (N_1223,In_1389,In_529);
nand U1224 (N_1224,In_860,In_882);
xnor U1225 (N_1225,In_605,In_523);
xor U1226 (N_1226,In_41,In_628);
and U1227 (N_1227,In_1351,In_1347);
nand U1228 (N_1228,In_730,In_160);
xnor U1229 (N_1229,In_621,In_710);
xnor U1230 (N_1230,In_580,In_1132);
and U1231 (N_1231,In_1430,In_894);
nand U1232 (N_1232,In_1164,In_502);
and U1233 (N_1233,In_256,In_186);
nor U1234 (N_1234,In_544,In_153);
nand U1235 (N_1235,In_503,In_1120);
nand U1236 (N_1236,In_523,In_479);
nor U1237 (N_1237,In_648,In_1332);
and U1238 (N_1238,In_665,In_327);
nand U1239 (N_1239,In_1398,In_1390);
or U1240 (N_1240,In_1148,In_177);
nand U1241 (N_1241,In_433,In_711);
nor U1242 (N_1242,In_947,In_605);
and U1243 (N_1243,In_882,In_474);
nor U1244 (N_1244,In_526,In_1443);
and U1245 (N_1245,In_464,In_456);
nand U1246 (N_1246,In_329,In_449);
nand U1247 (N_1247,In_1466,In_405);
nor U1248 (N_1248,In_273,In_3);
xor U1249 (N_1249,In_979,In_1191);
nor U1250 (N_1250,In_365,In_1286);
nand U1251 (N_1251,In_781,In_432);
nand U1252 (N_1252,In_244,In_1488);
nand U1253 (N_1253,In_845,In_1435);
or U1254 (N_1254,In_364,In_373);
and U1255 (N_1255,In_8,In_487);
or U1256 (N_1256,In_686,In_1269);
xor U1257 (N_1257,In_456,In_237);
nor U1258 (N_1258,In_1440,In_204);
or U1259 (N_1259,In_1430,In_644);
xnor U1260 (N_1260,In_248,In_113);
nand U1261 (N_1261,In_1088,In_1499);
and U1262 (N_1262,In_920,In_705);
and U1263 (N_1263,In_680,In_307);
and U1264 (N_1264,In_268,In_54);
or U1265 (N_1265,In_1480,In_1254);
nor U1266 (N_1266,In_99,In_1400);
nor U1267 (N_1267,In_1095,In_712);
nand U1268 (N_1268,In_1424,In_291);
xnor U1269 (N_1269,In_185,In_147);
nand U1270 (N_1270,In_1221,In_1039);
nand U1271 (N_1271,In_362,In_958);
nor U1272 (N_1272,In_1084,In_86);
nor U1273 (N_1273,In_98,In_368);
nand U1274 (N_1274,In_118,In_371);
and U1275 (N_1275,In_1180,In_807);
nor U1276 (N_1276,In_616,In_73);
and U1277 (N_1277,In_201,In_1407);
and U1278 (N_1278,In_451,In_1215);
nor U1279 (N_1279,In_1034,In_705);
xnor U1280 (N_1280,In_609,In_948);
and U1281 (N_1281,In_672,In_956);
nand U1282 (N_1282,In_1119,In_440);
xnor U1283 (N_1283,In_682,In_1438);
and U1284 (N_1284,In_78,In_1455);
xor U1285 (N_1285,In_859,In_16);
xor U1286 (N_1286,In_1488,In_1377);
and U1287 (N_1287,In_1342,In_427);
or U1288 (N_1288,In_970,In_1322);
nor U1289 (N_1289,In_214,In_18);
or U1290 (N_1290,In_973,In_1386);
or U1291 (N_1291,In_1237,In_144);
nand U1292 (N_1292,In_1459,In_111);
nor U1293 (N_1293,In_957,In_1428);
or U1294 (N_1294,In_184,In_153);
or U1295 (N_1295,In_186,In_938);
or U1296 (N_1296,In_157,In_1466);
nand U1297 (N_1297,In_960,In_67);
xnor U1298 (N_1298,In_856,In_466);
xnor U1299 (N_1299,In_246,In_425);
xor U1300 (N_1300,In_1452,In_169);
or U1301 (N_1301,In_1214,In_1093);
nor U1302 (N_1302,In_1079,In_121);
or U1303 (N_1303,In_166,In_900);
nand U1304 (N_1304,In_1079,In_900);
nand U1305 (N_1305,In_1180,In_307);
xnor U1306 (N_1306,In_1461,In_238);
nand U1307 (N_1307,In_1418,In_252);
xor U1308 (N_1308,In_1482,In_1269);
xor U1309 (N_1309,In_1242,In_232);
xor U1310 (N_1310,In_553,In_1056);
xor U1311 (N_1311,In_370,In_1455);
nand U1312 (N_1312,In_471,In_1093);
nor U1313 (N_1313,In_279,In_671);
nand U1314 (N_1314,In_1046,In_128);
nor U1315 (N_1315,In_246,In_743);
and U1316 (N_1316,In_1188,In_897);
and U1317 (N_1317,In_646,In_629);
and U1318 (N_1318,In_492,In_126);
nor U1319 (N_1319,In_495,In_277);
nor U1320 (N_1320,In_482,In_118);
nor U1321 (N_1321,In_968,In_1396);
nand U1322 (N_1322,In_1103,In_1316);
xor U1323 (N_1323,In_458,In_644);
xnor U1324 (N_1324,In_896,In_208);
nor U1325 (N_1325,In_1161,In_1437);
or U1326 (N_1326,In_855,In_480);
nor U1327 (N_1327,In_1366,In_1218);
or U1328 (N_1328,In_54,In_155);
and U1329 (N_1329,In_834,In_1287);
xnor U1330 (N_1330,In_502,In_1359);
and U1331 (N_1331,In_52,In_591);
nor U1332 (N_1332,In_394,In_248);
nor U1333 (N_1333,In_543,In_1113);
xor U1334 (N_1334,In_569,In_605);
xnor U1335 (N_1335,In_1189,In_1114);
and U1336 (N_1336,In_846,In_1285);
nor U1337 (N_1337,In_360,In_808);
nand U1338 (N_1338,In_1261,In_558);
and U1339 (N_1339,In_1456,In_1304);
or U1340 (N_1340,In_1268,In_1376);
or U1341 (N_1341,In_517,In_399);
nand U1342 (N_1342,In_1074,In_897);
xor U1343 (N_1343,In_1080,In_82);
nand U1344 (N_1344,In_26,In_51);
or U1345 (N_1345,In_1284,In_663);
nand U1346 (N_1346,In_77,In_546);
and U1347 (N_1347,In_1408,In_921);
nand U1348 (N_1348,In_635,In_226);
and U1349 (N_1349,In_803,In_1455);
and U1350 (N_1350,In_216,In_250);
xnor U1351 (N_1351,In_880,In_366);
nand U1352 (N_1352,In_515,In_142);
nand U1353 (N_1353,In_1211,In_563);
nand U1354 (N_1354,In_1100,In_601);
nor U1355 (N_1355,In_57,In_1093);
nand U1356 (N_1356,In_13,In_422);
nand U1357 (N_1357,In_321,In_120);
and U1358 (N_1358,In_248,In_1302);
xor U1359 (N_1359,In_226,In_461);
xor U1360 (N_1360,In_461,In_1070);
and U1361 (N_1361,In_475,In_67);
nand U1362 (N_1362,In_127,In_7);
and U1363 (N_1363,In_771,In_408);
nor U1364 (N_1364,In_1353,In_530);
xor U1365 (N_1365,In_1041,In_22);
xnor U1366 (N_1366,In_789,In_1014);
nor U1367 (N_1367,In_589,In_821);
nor U1368 (N_1368,In_510,In_365);
nand U1369 (N_1369,In_608,In_143);
and U1370 (N_1370,In_880,In_1483);
xor U1371 (N_1371,In_884,In_432);
nor U1372 (N_1372,In_1394,In_145);
nand U1373 (N_1373,In_772,In_1476);
nor U1374 (N_1374,In_1135,In_376);
xor U1375 (N_1375,In_81,In_412);
nor U1376 (N_1376,In_959,In_1115);
nand U1377 (N_1377,In_661,In_316);
or U1378 (N_1378,In_1241,In_416);
nand U1379 (N_1379,In_126,In_610);
or U1380 (N_1380,In_1463,In_872);
or U1381 (N_1381,In_1060,In_1464);
or U1382 (N_1382,In_1353,In_1313);
nor U1383 (N_1383,In_613,In_652);
or U1384 (N_1384,In_568,In_631);
nand U1385 (N_1385,In_635,In_114);
or U1386 (N_1386,In_1116,In_305);
and U1387 (N_1387,In_1296,In_301);
or U1388 (N_1388,In_406,In_223);
and U1389 (N_1389,In_181,In_349);
or U1390 (N_1390,In_685,In_1157);
or U1391 (N_1391,In_413,In_1047);
nand U1392 (N_1392,In_1433,In_286);
nor U1393 (N_1393,In_597,In_684);
nand U1394 (N_1394,In_1378,In_899);
and U1395 (N_1395,In_473,In_437);
xnor U1396 (N_1396,In_67,In_1064);
and U1397 (N_1397,In_281,In_90);
nor U1398 (N_1398,In_902,In_906);
or U1399 (N_1399,In_778,In_1141);
or U1400 (N_1400,In_1281,In_1102);
xnor U1401 (N_1401,In_851,In_729);
or U1402 (N_1402,In_1081,In_160);
xor U1403 (N_1403,In_609,In_622);
and U1404 (N_1404,In_1443,In_150);
nor U1405 (N_1405,In_1407,In_944);
or U1406 (N_1406,In_171,In_138);
nor U1407 (N_1407,In_131,In_924);
nand U1408 (N_1408,In_227,In_601);
nand U1409 (N_1409,In_597,In_483);
and U1410 (N_1410,In_839,In_566);
and U1411 (N_1411,In_921,In_1257);
or U1412 (N_1412,In_143,In_1391);
and U1413 (N_1413,In_482,In_543);
nand U1414 (N_1414,In_1100,In_1437);
xor U1415 (N_1415,In_239,In_974);
xor U1416 (N_1416,In_328,In_1253);
or U1417 (N_1417,In_240,In_1313);
xor U1418 (N_1418,In_1156,In_466);
nor U1419 (N_1419,In_824,In_69);
nand U1420 (N_1420,In_1425,In_1071);
or U1421 (N_1421,In_1209,In_893);
xnor U1422 (N_1422,In_521,In_1123);
or U1423 (N_1423,In_1442,In_1117);
nand U1424 (N_1424,In_114,In_557);
nand U1425 (N_1425,In_1327,In_457);
nand U1426 (N_1426,In_419,In_965);
or U1427 (N_1427,In_629,In_322);
or U1428 (N_1428,In_426,In_436);
xnor U1429 (N_1429,In_1227,In_1343);
nor U1430 (N_1430,In_1416,In_1474);
and U1431 (N_1431,In_709,In_955);
nand U1432 (N_1432,In_1254,In_1285);
and U1433 (N_1433,In_1388,In_815);
and U1434 (N_1434,In_1233,In_647);
nand U1435 (N_1435,In_335,In_56);
nor U1436 (N_1436,In_243,In_457);
or U1437 (N_1437,In_980,In_468);
nor U1438 (N_1438,In_1455,In_984);
and U1439 (N_1439,In_198,In_103);
or U1440 (N_1440,In_685,In_974);
nand U1441 (N_1441,In_631,In_24);
or U1442 (N_1442,In_5,In_490);
nor U1443 (N_1443,In_50,In_1489);
xnor U1444 (N_1444,In_903,In_752);
or U1445 (N_1445,In_1185,In_68);
xor U1446 (N_1446,In_1440,In_891);
or U1447 (N_1447,In_859,In_594);
nand U1448 (N_1448,In_815,In_623);
nor U1449 (N_1449,In_1240,In_1066);
and U1450 (N_1450,In_10,In_1346);
or U1451 (N_1451,In_1004,In_615);
and U1452 (N_1452,In_946,In_203);
nand U1453 (N_1453,In_1329,In_816);
nand U1454 (N_1454,In_663,In_1274);
and U1455 (N_1455,In_33,In_610);
xnor U1456 (N_1456,In_413,In_1468);
nor U1457 (N_1457,In_148,In_61);
or U1458 (N_1458,In_916,In_1490);
xnor U1459 (N_1459,In_842,In_1056);
or U1460 (N_1460,In_215,In_325);
nor U1461 (N_1461,In_746,In_667);
nand U1462 (N_1462,In_1473,In_776);
nor U1463 (N_1463,In_1393,In_1295);
nand U1464 (N_1464,In_96,In_940);
xnor U1465 (N_1465,In_44,In_1412);
nor U1466 (N_1466,In_1121,In_831);
nand U1467 (N_1467,In_1194,In_904);
or U1468 (N_1468,In_1237,In_1435);
and U1469 (N_1469,In_258,In_590);
nand U1470 (N_1470,In_252,In_1147);
or U1471 (N_1471,In_1096,In_1124);
and U1472 (N_1472,In_542,In_1454);
nand U1473 (N_1473,In_1377,In_498);
nand U1474 (N_1474,In_740,In_472);
nor U1475 (N_1475,In_189,In_345);
nor U1476 (N_1476,In_1244,In_209);
nand U1477 (N_1477,In_525,In_1368);
and U1478 (N_1478,In_916,In_605);
or U1479 (N_1479,In_138,In_92);
xnor U1480 (N_1480,In_166,In_1392);
or U1481 (N_1481,In_642,In_526);
xnor U1482 (N_1482,In_412,In_561);
and U1483 (N_1483,In_1101,In_462);
nor U1484 (N_1484,In_1230,In_834);
nor U1485 (N_1485,In_980,In_1344);
and U1486 (N_1486,In_1123,In_1385);
and U1487 (N_1487,In_1093,In_1300);
and U1488 (N_1488,In_279,In_64);
or U1489 (N_1489,In_549,In_119);
or U1490 (N_1490,In_1319,In_1239);
nand U1491 (N_1491,In_833,In_425);
or U1492 (N_1492,In_123,In_886);
nand U1493 (N_1493,In_184,In_170);
or U1494 (N_1494,In_1373,In_306);
nor U1495 (N_1495,In_1442,In_505);
or U1496 (N_1496,In_793,In_371);
xor U1497 (N_1497,In_982,In_712);
nor U1498 (N_1498,In_660,In_92);
or U1499 (N_1499,In_907,In_359);
nor U1500 (N_1500,In_841,In_879);
or U1501 (N_1501,In_1243,In_254);
or U1502 (N_1502,In_724,In_1237);
or U1503 (N_1503,In_1477,In_1367);
nor U1504 (N_1504,In_1376,In_917);
or U1505 (N_1505,In_1062,In_612);
nor U1506 (N_1506,In_170,In_349);
nand U1507 (N_1507,In_296,In_255);
nor U1508 (N_1508,In_222,In_835);
nand U1509 (N_1509,In_1454,In_1126);
nor U1510 (N_1510,In_133,In_635);
nor U1511 (N_1511,In_927,In_158);
xor U1512 (N_1512,In_445,In_1327);
xnor U1513 (N_1513,In_483,In_970);
nor U1514 (N_1514,In_1476,In_668);
nand U1515 (N_1515,In_292,In_1318);
and U1516 (N_1516,In_1046,In_271);
nand U1517 (N_1517,In_15,In_577);
xor U1518 (N_1518,In_82,In_370);
nor U1519 (N_1519,In_202,In_466);
xor U1520 (N_1520,In_649,In_383);
xnor U1521 (N_1521,In_1146,In_440);
nor U1522 (N_1522,In_152,In_1047);
xnor U1523 (N_1523,In_552,In_529);
xor U1524 (N_1524,In_76,In_1086);
nand U1525 (N_1525,In_936,In_1034);
or U1526 (N_1526,In_1392,In_807);
or U1527 (N_1527,In_418,In_1308);
xor U1528 (N_1528,In_47,In_195);
nand U1529 (N_1529,In_1219,In_1470);
nor U1530 (N_1530,In_63,In_395);
and U1531 (N_1531,In_282,In_39);
or U1532 (N_1532,In_476,In_1272);
or U1533 (N_1533,In_865,In_432);
and U1534 (N_1534,In_334,In_198);
or U1535 (N_1535,In_95,In_619);
and U1536 (N_1536,In_1490,In_548);
xor U1537 (N_1537,In_41,In_673);
and U1538 (N_1538,In_565,In_1019);
or U1539 (N_1539,In_739,In_854);
or U1540 (N_1540,In_1034,In_787);
xnor U1541 (N_1541,In_431,In_825);
xor U1542 (N_1542,In_207,In_1454);
nand U1543 (N_1543,In_214,In_715);
or U1544 (N_1544,In_1149,In_78);
and U1545 (N_1545,In_718,In_763);
xor U1546 (N_1546,In_174,In_517);
nor U1547 (N_1547,In_1354,In_100);
xor U1548 (N_1548,In_1113,In_36);
or U1549 (N_1549,In_791,In_593);
nor U1550 (N_1550,In_304,In_107);
nor U1551 (N_1551,In_1152,In_486);
nor U1552 (N_1552,In_247,In_914);
xnor U1553 (N_1553,In_998,In_1467);
or U1554 (N_1554,In_1460,In_1297);
or U1555 (N_1555,In_360,In_372);
nor U1556 (N_1556,In_564,In_382);
or U1557 (N_1557,In_810,In_55);
and U1558 (N_1558,In_1077,In_79);
nor U1559 (N_1559,In_77,In_1029);
xnor U1560 (N_1560,In_519,In_111);
nor U1561 (N_1561,In_1350,In_389);
xnor U1562 (N_1562,In_902,In_1054);
and U1563 (N_1563,In_266,In_685);
nand U1564 (N_1564,In_938,In_496);
and U1565 (N_1565,In_1401,In_333);
and U1566 (N_1566,In_14,In_589);
xnor U1567 (N_1567,In_272,In_271);
and U1568 (N_1568,In_874,In_48);
nor U1569 (N_1569,In_1028,In_558);
or U1570 (N_1570,In_1272,In_456);
and U1571 (N_1571,In_1206,In_370);
nor U1572 (N_1572,In_359,In_636);
or U1573 (N_1573,In_1305,In_307);
nand U1574 (N_1574,In_501,In_463);
xor U1575 (N_1575,In_1206,In_1379);
or U1576 (N_1576,In_469,In_1077);
nand U1577 (N_1577,In_329,In_820);
and U1578 (N_1578,In_857,In_619);
and U1579 (N_1579,In_1279,In_482);
nand U1580 (N_1580,In_89,In_278);
xnor U1581 (N_1581,In_975,In_542);
or U1582 (N_1582,In_939,In_1175);
nand U1583 (N_1583,In_352,In_1132);
nand U1584 (N_1584,In_1110,In_980);
nor U1585 (N_1585,In_185,In_1489);
nand U1586 (N_1586,In_1385,In_426);
nand U1587 (N_1587,In_435,In_1422);
and U1588 (N_1588,In_202,In_855);
or U1589 (N_1589,In_1387,In_1413);
and U1590 (N_1590,In_1080,In_277);
xnor U1591 (N_1591,In_714,In_1442);
xor U1592 (N_1592,In_1274,In_501);
nand U1593 (N_1593,In_734,In_578);
or U1594 (N_1594,In_1406,In_383);
xor U1595 (N_1595,In_130,In_1219);
xor U1596 (N_1596,In_499,In_1172);
nand U1597 (N_1597,In_463,In_1410);
or U1598 (N_1598,In_404,In_1039);
xor U1599 (N_1599,In_1403,In_297);
or U1600 (N_1600,In_993,In_386);
nor U1601 (N_1601,In_518,In_43);
xnor U1602 (N_1602,In_780,In_665);
or U1603 (N_1603,In_706,In_1458);
xor U1604 (N_1604,In_1488,In_877);
and U1605 (N_1605,In_405,In_447);
and U1606 (N_1606,In_1368,In_1123);
and U1607 (N_1607,In_1245,In_1014);
or U1608 (N_1608,In_1208,In_703);
xnor U1609 (N_1609,In_1486,In_117);
xnor U1610 (N_1610,In_527,In_160);
nor U1611 (N_1611,In_1045,In_792);
nand U1612 (N_1612,In_1316,In_1391);
nor U1613 (N_1613,In_695,In_334);
xor U1614 (N_1614,In_354,In_493);
and U1615 (N_1615,In_876,In_1331);
nand U1616 (N_1616,In_473,In_1353);
nand U1617 (N_1617,In_87,In_1171);
nand U1618 (N_1618,In_167,In_151);
and U1619 (N_1619,In_1333,In_93);
nor U1620 (N_1620,In_1225,In_573);
xnor U1621 (N_1621,In_272,In_885);
or U1622 (N_1622,In_517,In_477);
xor U1623 (N_1623,In_945,In_641);
xor U1624 (N_1624,In_1265,In_1022);
and U1625 (N_1625,In_800,In_931);
nand U1626 (N_1626,In_530,In_132);
nand U1627 (N_1627,In_993,In_240);
nor U1628 (N_1628,In_1288,In_455);
nor U1629 (N_1629,In_109,In_896);
xor U1630 (N_1630,In_1040,In_295);
nand U1631 (N_1631,In_1192,In_1148);
or U1632 (N_1632,In_500,In_128);
or U1633 (N_1633,In_413,In_1399);
nor U1634 (N_1634,In_1363,In_285);
xor U1635 (N_1635,In_1287,In_743);
xnor U1636 (N_1636,In_1209,In_1080);
nor U1637 (N_1637,In_201,In_7);
nand U1638 (N_1638,In_1220,In_4);
and U1639 (N_1639,In_661,In_784);
or U1640 (N_1640,In_981,In_946);
and U1641 (N_1641,In_1340,In_52);
xnor U1642 (N_1642,In_1170,In_1326);
nor U1643 (N_1643,In_565,In_747);
nor U1644 (N_1644,In_841,In_570);
xor U1645 (N_1645,In_1119,In_956);
nor U1646 (N_1646,In_1077,In_839);
nor U1647 (N_1647,In_807,In_245);
or U1648 (N_1648,In_230,In_150);
and U1649 (N_1649,In_1183,In_980);
and U1650 (N_1650,In_872,In_818);
or U1651 (N_1651,In_301,In_1078);
nand U1652 (N_1652,In_831,In_250);
nand U1653 (N_1653,In_1492,In_37);
nor U1654 (N_1654,In_1241,In_728);
nand U1655 (N_1655,In_797,In_112);
nor U1656 (N_1656,In_359,In_822);
xor U1657 (N_1657,In_12,In_272);
nand U1658 (N_1658,In_139,In_1126);
or U1659 (N_1659,In_1057,In_1318);
or U1660 (N_1660,In_1123,In_103);
or U1661 (N_1661,In_765,In_778);
nor U1662 (N_1662,In_981,In_1293);
nor U1663 (N_1663,In_1034,In_1085);
xor U1664 (N_1664,In_1051,In_1409);
nand U1665 (N_1665,In_425,In_582);
nor U1666 (N_1666,In_55,In_1297);
nor U1667 (N_1667,In_44,In_1046);
and U1668 (N_1668,In_1306,In_1408);
nand U1669 (N_1669,In_1038,In_102);
and U1670 (N_1670,In_1079,In_1476);
and U1671 (N_1671,In_463,In_999);
or U1672 (N_1672,In_1385,In_259);
and U1673 (N_1673,In_1318,In_472);
nor U1674 (N_1674,In_60,In_927);
nor U1675 (N_1675,In_326,In_874);
and U1676 (N_1676,In_1054,In_79);
or U1677 (N_1677,In_359,In_52);
or U1678 (N_1678,In_600,In_1082);
nand U1679 (N_1679,In_720,In_550);
nand U1680 (N_1680,In_508,In_100);
and U1681 (N_1681,In_608,In_304);
nor U1682 (N_1682,In_1112,In_336);
nor U1683 (N_1683,In_745,In_1309);
or U1684 (N_1684,In_563,In_173);
xnor U1685 (N_1685,In_130,In_545);
xnor U1686 (N_1686,In_861,In_1049);
nand U1687 (N_1687,In_943,In_360);
and U1688 (N_1688,In_1057,In_892);
xor U1689 (N_1689,In_950,In_1079);
and U1690 (N_1690,In_1112,In_1344);
or U1691 (N_1691,In_133,In_203);
xnor U1692 (N_1692,In_1348,In_586);
nor U1693 (N_1693,In_190,In_936);
nor U1694 (N_1694,In_341,In_809);
nand U1695 (N_1695,In_1489,In_604);
nor U1696 (N_1696,In_361,In_320);
or U1697 (N_1697,In_552,In_558);
and U1698 (N_1698,In_177,In_273);
xnor U1699 (N_1699,In_606,In_1150);
nand U1700 (N_1700,In_821,In_1189);
or U1701 (N_1701,In_602,In_120);
nand U1702 (N_1702,In_1408,In_372);
and U1703 (N_1703,In_671,In_983);
and U1704 (N_1704,In_722,In_6);
or U1705 (N_1705,In_794,In_950);
nand U1706 (N_1706,In_1038,In_242);
and U1707 (N_1707,In_667,In_936);
nor U1708 (N_1708,In_627,In_767);
or U1709 (N_1709,In_1427,In_916);
and U1710 (N_1710,In_4,In_717);
xor U1711 (N_1711,In_770,In_124);
or U1712 (N_1712,In_1400,In_1329);
or U1713 (N_1713,In_1088,In_188);
xnor U1714 (N_1714,In_853,In_394);
nand U1715 (N_1715,In_1049,In_259);
nor U1716 (N_1716,In_1054,In_692);
and U1717 (N_1717,In_1127,In_153);
and U1718 (N_1718,In_1429,In_594);
and U1719 (N_1719,In_148,In_839);
xor U1720 (N_1720,In_507,In_1456);
nand U1721 (N_1721,In_293,In_870);
and U1722 (N_1722,In_303,In_309);
nor U1723 (N_1723,In_291,In_876);
or U1724 (N_1724,In_83,In_327);
and U1725 (N_1725,In_482,In_283);
nor U1726 (N_1726,In_294,In_1);
and U1727 (N_1727,In_1004,In_241);
nand U1728 (N_1728,In_1158,In_579);
nand U1729 (N_1729,In_733,In_215);
and U1730 (N_1730,In_250,In_856);
nand U1731 (N_1731,In_938,In_1402);
or U1732 (N_1732,In_1497,In_1249);
xor U1733 (N_1733,In_535,In_432);
nor U1734 (N_1734,In_527,In_1120);
nand U1735 (N_1735,In_590,In_527);
nand U1736 (N_1736,In_739,In_483);
xor U1737 (N_1737,In_1167,In_1199);
or U1738 (N_1738,In_1162,In_381);
or U1739 (N_1739,In_190,In_1381);
nand U1740 (N_1740,In_152,In_1408);
nand U1741 (N_1741,In_1048,In_758);
and U1742 (N_1742,In_1154,In_572);
or U1743 (N_1743,In_268,In_67);
and U1744 (N_1744,In_880,In_622);
nand U1745 (N_1745,In_649,In_479);
xor U1746 (N_1746,In_236,In_1262);
or U1747 (N_1747,In_495,In_80);
or U1748 (N_1748,In_165,In_1192);
xor U1749 (N_1749,In_1229,In_1143);
nor U1750 (N_1750,In_1456,In_391);
nand U1751 (N_1751,In_236,In_683);
nand U1752 (N_1752,In_1136,In_599);
or U1753 (N_1753,In_619,In_593);
and U1754 (N_1754,In_1415,In_1441);
and U1755 (N_1755,In_240,In_1454);
or U1756 (N_1756,In_1112,In_1292);
nor U1757 (N_1757,In_943,In_1350);
xnor U1758 (N_1758,In_1338,In_277);
or U1759 (N_1759,In_1212,In_1065);
xnor U1760 (N_1760,In_860,In_733);
or U1761 (N_1761,In_1356,In_179);
nand U1762 (N_1762,In_216,In_1208);
nor U1763 (N_1763,In_280,In_55);
and U1764 (N_1764,In_344,In_612);
or U1765 (N_1765,In_577,In_1269);
nor U1766 (N_1766,In_1385,In_929);
xnor U1767 (N_1767,In_617,In_1498);
and U1768 (N_1768,In_438,In_287);
and U1769 (N_1769,In_742,In_860);
and U1770 (N_1770,In_1413,In_729);
nor U1771 (N_1771,In_686,In_358);
or U1772 (N_1772,In_1053,In_613);
xnor U1773 (N_1773,In_1026,In_586);
nor U1774 (N_1774,In_1458,In_1361);
xor U1775 (N_1775,In_888,In_616);
or U1776 (N_1776,In_1108,In_716);
or U1777 (N_1777,In_495,In_142);
and U1778 (N_1778,In_442,In_1411);
xnor U1779 (N_1779,In_272,In_22);
nor U1780 (N_1780,In_324,In_1399);
nand U1781 (N_1781,In_399,In_1063);
xor U1782 (N_1782,In_101,In_782);
or U1783 (N_1783,In_262,In_127);
and U1784 (N_1784,In_1057,In_476);
nor U1785 (N_1785,In_68,In_146);
nand U1786 (N_1786,In_482,In_1072);
or U1787 (N_1787,In_1227,In_24);
nand U1788 (N_1788,In_341,In_118);
nand U1789 (N_1789,In_1369,In_717);
xor U1790 (N_1790,In_1114,In_579);
nand U1791 (N_1791,In_698,In_124);
or U1792 (N_1792,In_1415,In_217);
nor U1793 (N_1793,In_1290,In_645);
nand U1794 (N_1794,In_1398,In_993);
or U1795 (N_1795,In_598,In_231);
or U1796 (N_1796,In_1318,In_898);
nand U1797 (N_1797,In_399,In_936);
or U1798 (N_1798,In_180,In_59);
xor U1799 (N_1799,In_1129,In_98);
nand U1800 (N_1800,In_860,In_448);
or U1801 (N_1801,In_674,In_1468);
nor U1802 (N_1802,In_1021,In_779);
or U1803 (N_1803,In_1494,In_1340);
nor U1804 (N_1804,In_363,In_658);
or U1805 (N_1805,In_237,In_1183);
and U1806 (N_1806,In_1027,In_171);
nand U1807 (N_1807,In_1236,In_294);
and U1808 (N_1808,In_337,In_970);
or U1809 (N_1809,In_429,In_616);
nand U1810 (N_1810,In_63,In_519);
nor U1811 (N_1811,In_422,In_895);
and U1812 (N_1812,In_1390,In_340);
nand U1813 (N_1813,In_50,In_130);
or U1814 (N_1814,In_1422,In_61);
xor U1815 (N_1815,In_1247,In_1168);
xnor U1816 (N_1816,In_1181,In_423);
nand U1817 (N_1817,In_1260,In_374);
nor U1818 (N_1818,In_565,In_947);
nor U1819 (N_1819,In_1372,In_81);
and U1820 (N_1820,In_543,In_571);
or U1821 (N_1821,In_884,In_1480);
xnor U1822 (N_1822,In_612,In_1393);
and U1823 (N_1823,In_125,In_85);
xor U1824 (N_1824,In_1461,In_762);
xor U1825 (N_1825,In_941,In_688);
and U1826 (N_1826,In_1067,In_344);
nor U1827 (N_1827,In_391,In_1216);
xnor U1828 (N_1828,In_266,In_1134);
nor U1829 (N_1829,In_987,In_790);
nand U1830 (N_1830,In_923,In_833);
xnor U1831 (N_1831,In_1238,In_973);
nand U1832 (N_1832,In_90,In_1197);
nor U1833 (N_1833,In_118,In_1371);
or U1834 (N_1834,In_868,In_1171);
xor U1835 (N_1835,In_1207,In_1395);
and U1836 (N_1836,In_518,In_1057);
xnor U1837 (N_1837,In_995,In_344);
and U1838 (N_1838,In_804,In_1063);
nor U1839 (N_1839,In_573,In_176);
nand U1840 (N_1840,In_1483,In_878);
xor U1841 (N_1841,In_681,In_230);
nor U1842 (N_1842,In_798,In_1327);
nand U1843 (N_1843,In_243,In_1228);
and U1844 (N_1844,In_578,In_812);
xor U1845 (N_1845,In_1009,In_1429);
or U1846 (N_1846,In_329,In_952);
nor U1847 (N_1847,In_260,In_238);
nand U1848 (N_1848,In_1155,In_744);
nand U1849 (N_1849,In_533,In_585);
nor U1850 (N_1850,In_436,In_1038);
or U1851 (N_1851,In_1421,In_959);
or U1852 (N_1852,In_222,In_970);
and U1853 (N_1853,In_468,In_1467);
or U1854 (N_1854,In_1463,In_1473);
nand U1855 (N_1855,In_424,In_283);
nand U1856 (N_1856,In_174,In_408);
xnor U1857 (N_1857,In_510,In_1090);
and U1858 (N_1858,In_436,In_973);
nand U1859 (N_1859,In_1481,In_490);
xor U1860 (N_1860,In_533,In_343);
and U1861 (N_1861,In_1134,In_155);
nand U1862 (N_1862,In_1261,In_313);
nand U1863 (N_1863,In_935,In_1250);
and U1864 (N_1864,In_288,In_1453);
nor U1865 (N_1865,In_1074,In_1331);
or U1866 (N_1866,In_1417,In_823);
nand U1867 (N_1867,In_23,In_903);
nand U1868 (N_1868,In_1468,In_243);
nor U1869 (N_1869,In_1108,In_363);
or U1870 (N_1870,In_1301,In_381);
nor U1871 (N_1871,In_909,In_1303);
xnor U1872 (N_1872,In_892,In_982);
xnor U1873 (N_1873,In_871,In_465);
nand U1874 (N_1874,In_729,In_1372);
nand U1875 (N_1875,In_733,In_1070);
and U1876 (N_1876,In_849,In_216);
nand U1877 (N_1877,In_565,In_1163);
and U1878 (N_1878,In_618,In_268);
nor U1879 (N_1879,In_816,In_131);
xor U1880 (N_1880,In_205,In_1240);
and U1881 (N_1881,In_37,In_784);
nor U1882 (N_1882,In_666,In_400);
xnor U1883 (N_1883,In_182,In_939);
xnor U1884 (N_1884,In_1093,In_792);
nand U1885 (N_1885,In_994,In_1079);
nand U1886 (N_1886,In_857,In_1411);
nor U1887 (N_1887,In_968,In_141);
nand U1888 (N_1888,In_1021,In_422);
or U1889 (N_1889,In_767,In_1480);
nand U1890 (N_1890,In_1283,In_911);
or U1891 (N_1891,In_544,In_380);
xnor U1892 (N_1892,In_325,In_1157);
xor U1893 (N_1893,In_313,In_28);
nand U1894 (N_1894,In_1066,In_480);
xnor U1895 (N_1895,In_634,In_34);
or U1896 (N_1896,In_256,In_1300);
or U1897 (N_1897,In_1383,In_750);
or U1898 (N_1898,In_801,In_1463);
xor U1899 (N_1899,In_282,In_787);
nor U1900 (N_1900,In_1472,In_1194);
and U1901 (N_1901,In_692,In_1254);
nor U1902 (N_1902,In_889,In_762);
or U1903 (N_1903,In_780,In_886);
or U1904 (N_1904,In_945,In_772);
nor U1905 (N_1905,In_1275,In_476);
xnor U1906 (N_1906,In_476,In_550);
xor U1907 (N_1907,In_322,In_268);
xnor U1908 (N_1908,In_1206,In_1390);
xnor U1909 (N_1909,In_1253,In_719);
nand U1910 (N_1910,In_359,In_1364);
xnor U1911 (N_1911,In_445,In_832);
nand U1912 (N_1912,In_646,In_639);
nand U1913 (N_1913,In_699,In_929);
nand U1914 (N_1914,In_219,In_1048);
nand U1915 (N_1915,In_776,In_1413);
nor U1916 (N_1916,In_1301,In_839);
and U1917 (N_1917,In_1267,In_1424);
xor U1918 (N_1918,In_615,In_472);
nand U1919 (N_1919,In_459,In_1273);
xnor U1920 (N_1920,In_560,In_705);
nor U1921 (N_1921,In_784,In_388);
and U1922 (N_1922,In_1065,In_1488);
nand U1923 (N_1923,In_298,In_275);
and U1924 (N_1924,In_1224,In_133);
nand U1925 (N_1925,In_1314,In_907);
and U1926 (N_1926,In_225,In_613);
xnor U1927 (N_1927,In_649,In_722);
and U1928 (N_1928,In_1047,In_664);
xnor U1929 (N_1929,In_1494,In_1464);
nor U1930 (N_1930,In_1027,In_521);
nand U1931 (N_1931,In_812,In_72);
xor U1932 (N_1932,In_1186,In_529);
nand U1933 (N_1933,In_728,In_626);
or U1934 (N_1934,In_86,In_142);
and U1935 (N_1935,In_1195,In_1230);
nand U1936 (N_1936,In_384,In_1020);
nor U1937 (N_1937,In_1403,In_160);
nor U1938 (N_1938,In_1052,In_1141);
and U1939 (N_1939,In_382,In_243);
and U1940 (N_1940,In_868,In_1143);
and U1941 (N_1941,In_29,In_705);
and U1942 (N_1942,In_147,In_1479);
nand U1943 (N_1943,In_450,In_563);
or U1944 (N_1944,In_213,In_390);
or U1945 (N_1945,In_1172,In_216);
or U1946 (N_1946,In_1280,In_1071);
nor U1947 (N_1947,In_1105,In_839);
xnor U1948 (N_1948,In_746,In_749);
nor U1949 (N_1949,In_1066,In_1139);
xnor U1950 (N_1950,In_332,In_1159);
or U1951 (N_1951,In_584,In_1106);
xnor U1952 (N_1952,In_604,In_334);
and U1953 (N_1953,In_172,In_986);
or U1954 (N_1954,In_1382,In_1150);
xor U1955 (N_1955,In_1444,In_764);
xor U1956 (N_1956,In_331,In_796);
nor U1957 (N_1957,In_1080,In_1148);
nand U1958 (N_1958,In_1242,In_327);
and U1959 (N_1959,In_1203,In_1297);
and U1960 (N_1960,In_812,In_1034);
and U1961 (N_1961,In_301,In_585);
and U1962 (N_1962,In_1434,In_1290);
xnor U1963 (N_1963,In_467,In_601);
and U1964 (N_1964,In_166,In_291);
and U1965 (N_1965,In_317,In_372);
nand U1966 (N_1966,In_955,In_701);
nand U1967 (N_1967,In_1390,In_609);
nor U1968 (N_1968,In_882,In_1274);
or U1969 (N_1969,In_682,In_439);
or U1970 (N_1970,In_1,In_932);
nor U1971 (N_1971,In_968,In_245);
xnor U1972 (N_1972,In_766,In_1341);
and U1973 (N_1973,In_562,In_459);
nor U1974 (N_1974,In_1212,In_985);
nor U1975 (N_1975,In_272,In_1039);
or U1976 (N_1976,In_971,In_818);
and U1977 (N_1977,In_1102,In_122);
nand U1978 (N_1978,In_369,In_1026);
nor U1979 (N_1979,In_249,In_166);
nor U1980 (N_1980,In_398,In_1384);
xor U1981 (N_1981,In_1148,In_1291);
and U1982 (N_1982,In_1289,In_356);
and U1983 (N_1983,In_1419,In_1152);
nand U1984 (N_1984,In_526,In_603);
or U1985 (N_1985,In_659,In_378);
or U1986 (N_1986,In_1270,In_1254);
nand U1987 (N_1987,In_615,In_200);
or U1988 (N_1988,In_411,In_248);
and U1989 (N_1989,In_1467,In_420);
nor U1990 (N_1990,In_265,In_1289);
and U1991 (N_1991,In_13,In_548);
or U1992 (N_1992,In_733,In_1065);
nand U1993 (N_1993,In_874,In_122);
or U1994 (N_1994,In_110,In_1029);
nor U1995 (N_1995,In_100,In_58);
and U1996 (N_1996,In_853,In_652);
and U1997 (N_1997,In_515,In_1201);
or U1998 (N_1998,In_1036,In_1457);
nand U1999 (N_1999,In_4,In_1265);
nor U2000 (N_2000,In_749,In_653);
and U2001 (N_2001,In_790,In_543);
nand U2002 (N_2002,In_535,In_1066);
xnor U2003 (N_2003,In_874,In_24);
nand U2004 (N_2004,In_1003,In_1169);
nand U2005 (N_2005,In_531,In_175);
nor U2006 (N_2006,In_1488,In_528);
xor U2007 (N_2007,In_1036,In_865);
nand U2008 (N_2008,In_956,In_32);
nor U2009 (N_2009,In_917,In_930);
and U2010 (N_2010,In_1138,In_469);
xor U2011 (N_2011,In_257,In_19);
xor U2012 (N_2012,In_794,In_253);
and U2013 (N_2013,In_520,In_875);
and U2014 (N_2014,In_392,In_719);
nand U2015 (N_2015,In_637,In_686);
xnor U2016 (N_2016,In_1320,In_86);
xor U2017 (N_2017,In_636,In_792);
or U2018 (N_2018,In_497,In_211);
xor U2019 (N_2019,In_993,In_1097);
and U2020 (N_2020,In_836,In_390);
and U2021 (N_2021,In_123,In_439);
nand U2022 (N_2022,In_921,In_1224);
nor U2023 (N_2023,In_313,In_964);
nor U2024 (N_2024,In_1170,In_223);
nor U2025 (N_2025,In_815,In_70);
and U2026 (N_2026,In_1437,In_1360);
and U2027 (N_2027,In_1414,In_1186);
xnor U2028 (N_2028,In_780,In_205);
nand U2029 (N_2029,In_571,In_251);
nor U2030 (N_2030,In_1371,In_91);
xor U2031 (N_2031,In_976,In_1475);
nand U2032 (N_2032,In_895,In_827);
nand U2033 (N_2033,In_364,In_743);
or U2034 (N_2034,In_681,In_435);
and U2035 (N_2035,In_1291,In_260);
nand U2036 (N_2036,In_790,In_336);
nand U2037 (N_2037,In_1123,In_1431);
nand U2038 (N_2038,In_761,In_581);
and U2039 (N_2039,In_1335,In_1289);
or U2040 (N_2040,In_560,In_348);
and U2041 (N_2041,In_337,In_1401);
or U2042 (N_2042,In_1078,In_8);
or U2043 (N_2043,In_638,In_739);
and U2044 (N_2044,In_1073,In_1191);
xnor U2045 (N_2045,In_508,In_96);
and U2046 (N_2046,In_798,In_346);
nand U2047 (N_2047,In_1377,In_515);
nor U2048 (N_2048,In_1473,In_1394);
and U2049 (N_2049,In_490,In_1041);
xor U2050 (N_2050,In_617,In_702);
or U2051 (N_2051,In_598,In_567);
nor U2052 (N_2052,In_1281,In_771);
xor U2053 (N_2053,In_866,In_738);
nand U2054 (N_2054,In_283,In_558);
xnor U2055 (N_2055,In_510,In_133);
nor U2056 (N_2056,In_377,In_1471);
and U2057 (N_2057,In_815,In_996);
and U2058 (N_2058,In_1094,In_295);
xnor U2059 (N_2059,In_562,In_54);
xor U2060 (N_2060,In_958,In_1180);
nor U2061 (N_2061,In_28,In_1268);
or U2062 (N_2062,In_31,In_23);
or U2063 (N_2063,In_1232,In_1489);
nor U2064 (N_2064,In_99,In_1215);
xnor U2065 (N_2065,In_341,In_71);
nand U2066 (N_2066,In_1022,In_845);
nand U2067 (N_2067,In_1209,In_974);
or U2068 (N_2068,In_755,In_323);
xor U2069 (N_2069,In_536,In_845);
nor U2070 (N_2070,In_198,In_1467);
and U2071 (N_2071,In_969,In_80);
xnor U2072 (N_2072,In_280,In_74);
nor U2073 (N_2073,In_636,In_776);
nor U2074 (N_2074,In_1415,In_1318);
nand U2075 (N_2075,In_779,In_1444);
or U2076 (N_2076,In_667,In_1020);
or U2077 (N_2077,In_30,In_508);
nor U2078 (N_2078,In_1032,In_255);
nand U2079 (N_2079,In_1463,In_1279);
nor U2080 (N_2080,In_1315,In_1395);
or U2081 (N_2081,In_5,In_889);
nor U2082 (N_2082,In_766,In_638);
and U2083 (N_2083,In_222,In_1365);
or U2084 (N_2084,In_787,In_731);
xor U2085 (N_2085,In_163,In_1118);
or U2086 (N_2086,In_186,In_1038);
and U2087 (N_2087,In_526,In_721);
xnor U2088 (N_2088,In_1207,In_142);
nand U2089 (N_2089,In_821,In_1443);
xnor U2090 (N_2090,In_200,In_973);
nand U2091 (N_2091,In_1243,In_134);
xnor U2092 (N_2092,In_1498,In_201);
xor U2093 (N_2093,In_876,In_634);
or U2094 (N_2094,In_1405,In_1435);
xor U2095 (N_2095,In_570,In_115);
xor U2096 (N_2096,In_87,In_1227);
nand U2097 (N_2097,In_921,In_204);
nor U2098 (N_2098,In_284,In_1196);
xnor U2099 (N_2099,In_1159,In_159);
and U2100 (N_2100,In_1494,In_9);
nor U2101 (N_2101,In_45,In_1287);
nand U2102 (N_2102,In_1480,In_1312);
xnor U2103 (N_2103,In_1089,In_1088);
nand U2104 (N_2104,In_1315,In_27);
or U2105 (N_2105,In_519,In_205);
xor U2106 (N_2106,In_322,In_196);
xnor U2107 (N_2107,In_1172,In_688);
xnor U2108 (N_2108,In_414,In_841);
nand U2109 (N_2109,In_1219,In_244);
nand U2110 (N_2110,In_921,In_892);
nor U2111 (N_2111,In_204,In_293);
nand U2112 (N_2112,In_581,In_194);
and U2113 (N_2113,In_368,In_261);
or U2114 (N_2114,In_83,In_879);
or U2115 (N_2115,In_1135,In_267);
or U2116 (N_2116,In_936,In_1150);
nor U2117 (N_2117,In_334,In_230);
and U2118 (N_2118,In_201,In_629);
xnor U2119 (N_2119,In_1330,In_470);
xnor U2120 (N_2120,In_363,In_955);
nand U2121 (N_2121,In_942,In_953);
and U2122 (N_2122,In_727,In_1487);
nor U2123 (N_2123,In_1115,In_1418);
and U2124 (N_2124,In_1071,In_671);
and U2125 (N_2125,In_206,In_878);
or U2126 (N_2126,In_1492,In_920);
nor U2127 (N_2127,In_218,In_426);
and U2128 (N_2128,In_1103,In_447);
or U2129 (N_2129,In_1071,In_1486);
and U2130 (N_2130,In_1479,In_1262);
or U2131 (N_2131,In_400,In_1280);
xor U2132 (N_2132,In_621,In_1193);
xor U2133 (N_2133,In_261,In_1305);
nor U2134 (N_2134,In_904,In_387);
nand U2135 (N_2135,In_798,In_86);
nor U2136 (N_2136,In_133,In_926);
and U2137 (N_2137,In_1004,In_282);
xnor U2138 (N_2138,In_774,In_1373);
and U2139 (N_2139,In_742,In_213);
nor U2140 (N_2140,In_98,In_577);
or U2141 (N_2141,In_130,In_842);
and U2142 (N_2142,In_1122,In_1256);
or U2143 (N_2143,In_359,In_1017);
nor U2144 (N_2144,In_1355,In_1345);
nor U2145 (N_2145,In_417,In_1041);
or U2146 (N_2146,In_1009,In_774);
nand U2147 (N_2147,In_861,In_440);
nand U2148 (N_2148,In_261,In_309);
and U2149 (N_2149,In_355,In_1230);
and U2150 (N_2150,In_533,In_995);
nor U2151 (N_2151,In_385,In_1283);
xor U2152 (N_2152,In_743,In_43);
nor U2153 (N_2153,In_463,In_919);
nand U2154 (N_2154,In_1035,In_1342);
or U2155 (N_2155,In_155,In_1198);
nand U2156 (N_2156,In_639,In_1191);
nand U2157 (N_2157,In_233,In_1360);
nand U2158 (N_2158,In_545,In_264);
or U2159 (N_2159,In_1061,In_1341);
nor U2160 (N_2160,In_1399,In_8);
nor U2161 (N_2161,In_1400,In_1017);
or U2162 (N_2162,In_1406,In_237);
nand U2163 (N_2163,In_902,In_992);
and U2164 (N_2164,In_859,In_1049);
xor U2165 (N_2165,In_1320,In_1258);
and U2166 (N_2166,In_640,In_1240);
nand U2167 (N_2167,In_109,In_694);
and U2168 (N_2168,In_658,In_440);
xnor U2169 (N_2169,In_1438,In_1349);
nor U2170 (N_2170,In_1361,In_684);
nor U2171 (N_2171,In_1452,In_345);
or U2172 (N_2172,In_1401,In_501);
nand U2173 (N_2173,In_453,In_1193);
or U2174 (N_2174,In_1492,In_117);
nand U2175 (N_2175,In_840,In_202);
nor U2176 (N_2176,In_1150,In_1360);
and U2177 (N_2177,In_175,In_729);
and U2178 (N_2178,In_182,In_81);
nor U2179 (N_2179,In_303,In_1215);
nand U2180 (N_2180,In_193,In_1200);
and U2181 (N_2181,In_1050,In_928);
or U2182 (N_2182,In_1152,In_875);
nor U2183 (N_2183,In_1239,In_999);
nand U2184 (N_2184,In_1077,In_1421);
and U2185 (N_2185,In_1101,In_1454);
or U2186 (N_2186,In_1219,In_711);
or U2187 (N_2187,In_315,In_914);
or U2188 (N_2188,In_749,In_1123);
xor U2189 (N_2189,In_264,In_1142);
nor U2190 (N_2190,In_1422,In_568);
xnor U2191 (N_2191,In_1020,In_997);
nand U2192 (N_2192,In_1317,In_876);
nor U2193 (N_2193,In_6,In_725);
or U2194 (N_2194,In_590,In_107);
nor U2195 (N_2195,In_498,In_781);
and U2196 (N_2196,In_644,In_984);
and U2197 (N_2197,In_141,In_889);
nand U2198 (N_2198,In_625,In_724);
and U2199 (N_2199,In_1212,In_1446);
or U2200 (N_2200,In_1180,In_1253);
or U2201 (N_2201,In_873,In_851);
xnor U2202 (N_2202,In_859,In_1125);
xor U2203 (N_2203,In_1314,In_1355);
and U2204 (N_2204,In_1014,In_578);
or U2205 (N_2205,In_1389,In_811);
xor U2206 (N_2206,In_904,In_100);
nor U2207 (N_2207,In_459,In_735);
or U2208 (N_2208,In_1349,In_1312);
nand U2209 (N_2209,In_1001,In_898);
nand U2210 (N_2210,In_1468,In_892);
xnor U2211 (N_2211,In_779,In_122);
or U2212 (N_2212,In_117,In_1102);
and U2213 (N_2213,In_337,In_1318);
nor U2214 (N_2214,In_1278,In_910);
xnor U2215 (N_2215,In_592,In_446);
and U2216 (N_2216,In_779,In_868);
and U2217 (N_2217,In_535,In_531);
or U2218 (N_2218,In_728,In_51);
nand U2219 (N_2219,In_576,In_423);
and U2220 (N_2220,In_987,In_714);
and U2221 (N_2221,In_1249,In_336);
or U2222 (N_2222,In_513,In_209);
xnor U2223 (N_2223,In_145,In_460);
xnor U2224 (N_2224,In_1499,In_830);
xor U2225 (N_2225,In_964,In_1061);
nor U2226 (N_2226,In_1386,In_725);
xor U2227 (N_2227,In_546,In_371);
nor U2228 (N_2228,In_1332,In_1165);
nand U2229 (N_2229,In_605,In_1177);
and U2230 (N_2230,In_200,In_492);
nor U2231 (N_2231,In_905,In_95);
nand U2232 (N_2232,In_1459,In_1180);
or U2233 (N_2233,In_1171,In_807);
nor U2234 (N_2234,In_507,In_720);
xor U2235 (N_2235,In_968,In_1177);
nor U2236 (N_2236,In_981,In_1122);
and U2237 (N_2237,In_1427,In_929);
xor U2238 (N_2238,In_555,In_185);
nor U2239 (N_2239,In_659,In_878);
or U2240 (N_2240,In_1464,In_1420);
nand U2241 (N_2241,In_164,In_731);
or U2242 (N_2242,In_590,In_20);
and U2243 (N_2243,In_1350,In_1186);
xor U2244 (N_2244,In_1240,In_1440);
and U2245 (N_2245,In_22,In_301);
or U2246 (N_2246,In_80,In_222);
or U2247 (N_2247,In_867,In_529);
nor U2248 (N_2248,In_55,In_717);
or U2249 (N_2249,In_852,In_1425);
nor U2250 (N_2250,In_1306,In_113);
nand U2251 (N_2251,In_462,In_854);
nor U2252 (N_2252,In_835,In_632);
or U2253 (N_2253,In_1425,In_363);
or U2254 (N_2254,In_308,In_95);
nand U2255 (N_2255,In_827,In_794);
and U2256 (N_2256,In_1263,In_1361);
and U2257 (N_2257,In_296,In_262);
xnor U2258 (N_2258,In_203,In_436);
or U2259 (N_2259,In_1030,In_37);
and U2260 (N_2260,In_1064,In_864);
xnor U2261 (N_2261,In_1121,In_814);
nand U2262 (N_2262,In_562,In_217);
xnor U2263 (N_2263,In_429,In_382);
nand U2264 (N_2264,In_214,In_50);
nand U2265 (N_2265,In_912,In_918);
and U2266 (N_2266,In_955,In_101);
xnor U2267 (N_2267,In_1417,In_1009);
and U2268 (N_2268,In_1070,In_279);
or U2269 (N_2269,In_881,In_638);
nand U2270 (N_2270,In_1024,In_594);
and U2271 (N_2271,In_325,In_567);
nor U2272 (N_2272,In_2,In_294);
nand U2273 (N_2273,In_814,In_792);
and U2274 (N_2274,In_29,In_551);
nor U2275 (N_2275,In_1429,In_1327);
and U2276 (N_2276,In_23,In_1140);
nand U2277 (N_2277,In_763,In_1146);
or U2278 (N_2278,In_825,In_332);
and U2279 (N_2279,In_625,In_992);
nor U2280 (N_2280,In_559,In_1162);
or U2281 (N_2281,In_1452,In_798);
and U2282 (N_2282,In_807,In_1240);
xor U2283 (N_2283,In_1048,In_1108);
and U2284 (N_2284,In_332,In_336);
xnor U2285 (N_2285,In_974,In_37);
xnor U2286 (N_2286,In_1452,In_1195);
xnor U2287 (N_2287,In_574,In_1387);
and U2288 (N_2288,In_1022,In_337);
or U2289 (N_2289,In_1322,In_481);
and U2290 (N_2290,In_93,In_596);
nand U2291 (N_2291,In_560,In_1465);
or U2292 (N_2292,In_1154,In_1215);
nand U2293 (N_2293,In_332,In_523);
xor U2294 (N_2294,In_121,In_1006);
nor U2295 (N_2295,In_727,In_259);
or U2296 (N_2296,In_262,In_1470);
xor U2297 (N_2297,In_73,In_950);
xor U2298 (N_2298,In_497,In_958);
xnor U2299 (N_2299,In_11,In_572);
or U2300 (N_2300,In_300,In_1302);
or U2301 (N_2301,In_744,In_1494);
and U2302 (N_2302,In_1277,In_1146);
and U2303 (N_2303,In_760,In_168);
or U2304 (N_2304,In_658,In_886);
nor U2305 (N_2305,In_1288,In_770);
or U2306 (N_2306,In_1037,In_132);
nand U2307 (N_2307,In_1271,In_1321);
xnor U2308 (N_2308,In_969,In_53);
or U2309 (N_2309,In_889,In_297);
nor U2310 (N_2310,In_198,In_1090);
xnor U2311 (N_2311,In_1353,In_339);
xnor U2312 (N_2312,In_582,In_445);
or U2313 (N_2313,In_1157,In_946);
xor U2314 (N_2314,In_639,In_835);
or U2315 (N_2315,In_727,In_1085);
xor U2316 (N_2316,In_110,In_50);
nor U2317 (N_2317,In_1169,In_678);
and U2318 (N_2318,In_821,In_449);
nor U2319 (N_2319,In_1131,In_312);
or U2320 (N_2320,In_686,In_58);
xor U2321 (N_2321,In_478,In_968);
nor U2322 (N_2322,In_318,In_965);
or U2323 (N_2323,In_781,In_182);
nand U2324 (N_2324,In_934,In_745);
or U2325 (N_2325,In_284,In_245);
or U2326 (N_2326,In_111,In_1339);
or U2327 (N_2327,In_1410,In_141);
and U2328 (N_2328,In_1157,In_219);
nand U2329 (N_2329,In_1473,In_236);
xnor U2330 (N_2330,In_791,In_950);
xor U2331 (N_2331,In_533,In_878);
and U2332 (N_2332,In_726,In_840);
or U2333 (N_2333,In_150,In_584);
xor U2334 (N_2334,In_328,In_1277);
and U2335 (N_2335,In_156,In_899);
nor U2336 (N_2336,In_217,In_393);
nand U2337 (N_2337,In_1211,In_915);
and U2338 (N_2338,In_555,In_458);
or U2339 (N_2339,In_429,In_1142);
xor U2340 (N_2340,In_867,In_617);
nand U2341 (N_2341,In_661,In_615);
nor U2342 (N_2342,In_477,In_785);
or U2343 (N_2343,In_1263,In_914);
nand U2344 (N_2344,In_698,In_490);
or U2345 (N_2345,In_399,In_1073);
nand U2346 (N_2346,In_715,In_290);
nand U2347 (N_2347,In_1493,In_1037);
and U2348 (N_2348,In_944,In_1493);
or U2349 (N_2349,In_1457,In_1090);
or U2350 (N_2350,In_140,In_1176);
nor U2351 (N_2351,In_564,In_1195);
or U2352 (N_2352,In_543,In_490);
or U2353 (N_2353,In_441,In_464);
xnor U2354 (N_2354,In_163,In_838);
xnor U2355 (N_2355,In_592,In_1463);
and U2356 (N_2356,In_1269,In_874);
or U2357 (N_2357,In_957,In_908);
or U2358 (N_2358,In_254,In_1449);
nand U2359 (N_2359,In_1401,In_249);
nor U2360 (N_2360,In_418,In_1416);
xnor U2361 (N_2361,In_1471,In_304);
or U2362 (N_2362,In_757,In_381);
xnor U2363 (N_2363,In_230,In_1242);
and U2364 (N_2364,In_1476,In_828);
nand U2365 (N_2365,In_1002,In_316);
nor U2366 (N_2366,In_57,In_541);
nand U2367 (N_2367,In_1192,In_764);
and U2368 (N_2368,In_1128,In_325);
nor U2369 (N_2369,In_1370,In_407);
nand U2370 (N_2370,In_1262,In_957);
xor U2371 (N_2371,In_668,In_896);
nand U2372 (N_2372,In_436,In_1463);
and U2373 (N_2373,In_244,In_1005);
and U2374 (N_2374,In_1148,In_1222);
and U2375 (N_2375,In_429,In_479);
nor U2376 (N_2376,In_1435,In_579);
or U2377 (N_2377,In_39,In_658);
xor U2378 (N_2378,In_1471,In_349);
or U2379 (N_2379,In_1186,In_1399);
or U2380 (N_2380,In_246,In_1058);
xor U2381 (N_2381,In_122,In_1269);
and U2382 (N_2382,In_1348,In_1154);
or U2383 (N_2383,In_1048,In_440);
nor U2384 (N_2384,In_285,In_771);
xnor U2385 (N_2385,In_1187,In_97);
nand U2386 (N_2386,In_614,In_115);
nand U2387 (N_2387,In_441,In_573);
nand U2388 (N_2388,In_1305,In_917);
or U2389 (N_2389,In_453,In_1382);
and U2390 (N_2390,In_381,In_984);
nand U2391 (N_2391,In_692,In_148);
nor U2392 (N_2392,In_622,In_519);
or U2393 (N_2393,In_1324,In_1401);
nor U2394 (N_2394,In_1398,In_572);
nor U2395 (N_2395,In_1091,In_505);
xnor U2396 (N_2396,In_41,In_664);
or U2397 (N_2397,In_1231,In_866);
nor U2398 (N_2398,In_423,In_974);
and U2399 (N_2399,In_1136,In_1238);
and U2400 (N_2400,In_634,In_1317);
xnor U2401 (N_2401,In_236,In_312);
or U2402 (N_2402,In_789,In_267);
nand U2403 (N_2403,In_482,In_359);
xor U2404 (N_2404,In_1119,In_1291);
nor U2405 (N_2405,In_805,In_1455);
and U2406 (N_2406,In_1101,In_162);
and U2407 (N_2407,In_1439,In_707);
nor U2408 (N_2408,In_1143,In_769);
and U2409 (N_2409,In_1217,In_1496);
or U2410 (N_2410,In_1098,In_755);
and U2411 (N_2411,In_583,In_182);
or U2412 (N_2412,In_930,In_85);
nor U2413 (N_2413,In_1234,In_396);
and U2414 (N_2414,In_1158,In_1495);
nand U2415 (N_2415,In_1342,In_1071);
nor U2416 (N_2416,In_878,In_1323);
and U2417 (N_2417,In_394,In_865);
nand U2418 (N_2418,In_1361,In_1410);
nand U2419 (N_2419,In_1369,In_1412);
nand U2420 (N_2420,In_997,In_1292);
xnor U2421 (N_2421,In_438,In_1470);
xnor U2422 (N_2422,In_526,In_320);
xor U2423 (N_2423,In_1310,In_1420);
nand U2424 (N_2424,In_939,In_226);
and U2425 (N_2425,In_1217,In_1138);
xnor U2426 (N_2426,In_871,In_121);
xor U2427 (N_2427,In_1338,In_814);
and U2428 (N_2428,In_361,In_953);
and U2429 (N_2429,In_320,In_60);
xnor U2430 (N_2430,In_548,In_971);
nor U2431 (N_2431,In_359,In_1480);
or U2432 (N_2432,In_352,In_310);
nor U2433 (N_2433,In_434,In_1090);
and U2434 (N_2434,In_592,In_633);
nor U2435 (N_2435,In_1376,In_63);
nand U2436 (N_2436,In_767,In_580);
or U2437 (N_2437,In_1280,In_778);
xor U2438 (N_2438,In_46,In_433);
and U2439 (N_2439,In_1144,In_1230);
and U2440 (N_2440,In_1374,In_51);
or U2441 (N_2441,In_137,In_1363);
and U2442 (N_2442,In_1195,In_139);
nor U2443 (N_2443,In_695,In_397);
or U2444 (N_2444,In_628,In_1283);
and U2445 (N_2445,In_1280,In_776);
nor U2446 (N_2446,In_730,In_1301);
nand U2447 (N_2447,In_1025,In_88);
and U2448 (N_2448,In_6,In_374);
or U2449 (N_2449,In_705,In_525);
nand U2450 (N_2450,In_1073,In_267);
xnor U2451 (N_2451,In_580,In_1066);
nor U2452 (N_2452,In_1380,In_137);
nor U2453 (N_2453,In_1102,In_408);
xor U2454 (N_2454,In_1446,In_1493);
xor U2455 (N_2455,In_764,In_1324);
and U2456 (N_2456,In_11,In_85);
xor U2457 (N_2457,In_665,In_1257);
or U2458 (N_2458,In_617,In_621);
nor U2459 (N_2459,In_1293,In_704);
nor U2460 (N_2460,In_1173,In_995);
nor U2461 (N_2461,In_495,In_420);
nand U2462 (N_2462,In_348,In_977);
xor U2463 (N_2463,In_1042,In_606);
xor U2464 (N_2464,In_1289,In_763);
nor U2465 (N_2465,In_787,In_266);
xor U2466 (N_2466,In_1254,In_216);
and U2467 (N_2467,In_984,In_675);
nand U2468 (N_2468,In_1215,In_248);
and U2469 (N_2469,In_1297,In_155);
or U2470 (N_2470,In_588,In_264);
and U2471 (N_2471,In_47,In_78);
nand U2472 (N_2472,In_852,In_350);
or U2473 (N_2473,In_319,In_252);
and U2474 (N_2474,In_651,In_271);
nor U2475 (N_2475,In_1265,In_1372);
xnor U2476 (N_2476,In_510,In_421);
or U2477 (N_2477,In_1220,In_842);
or U2478 (N_2478,In_902,In_736);
or U2479 (N_2479,In_850,In_1081);
or U2480 (N_2480,In_717,In_206);
xnor U2481 (N_2481,In_172,In_899);
nand U2482 (N_2482,In_1195,In_671);
xnor U2483 (N_2483,In_1144,In_828);
nand U2484 (N_2484,In_356,In_919);
and U2485 (N_2485,In_1394,In_413);
nand U2486 (N_2486,In_883,In_1247);
nor U2487 (N_2487,In_635,In_1470);
xor U2488 (N_2488,In_230,In_303);
nor U2489 (N_2489,In_36,In_176);
or U2490 (N_2490,In_1304,In_1298);
nor U2491 (N_2491,In_18,In_546);
or U2492 (N_2492,In_1085,In_890);
nand U2493 (N_2493,In_213,In_395);
and U2494 (N_2494,In_371,In_1012);
nand U2495 (N_2495,In_15,In_1329);
nor U2496 (N_2496,In_1389,In_720);
xnor U2497 (N_2497,In_925,In_114);
xnor U2498 (N_2498,In_773,In_871);
or U2499 (N_2499,In_241,In_1478);
and U2500 (N_2500,In_166,In_1415);
or U2501 (N_2501,In_292,In_1467);
nor U2502 (N_2502,In_42,In_75);
nand U2503 (N_2503,In_637,In_76);
xnor U2504 (N_2504,In_1024,In_1006);
nand U2505 (N_2505,In_596,In_1297);
and U2506 (N_2506,In_900,In_1329);
xnor U2507 (N_2507,In_901,In_776);
nor U2508 (N_2508,In_1315,In_10);
xnor U2509 (N_2509,In_1345,In_860);
nand U2510 (N_2510,In_891,In_258);
and U2511 (N_2511,In_119,In_559);
xor U2512 (N_2512,In_906,In_874);
and U2513 (N_2513,In_793,In_29);
xor U2514 (N_2514,In_1409,In_123);
xnor U2515 (N_2515,In_1401,In_794);
xor U2516 (N_2516,In_138,In_298);
and U2517 (N_2517,In_1272,In_1042);
nor U2518 (N_2518,In_1411,In_237);
or U2519 (N_2519,In_78,In_1146);
and U2520 (N_2520,In_512,In_2);
nor U2521 (N_2521,In_861,In_1410);
xor U2522 (N_2522,In_145,In_334);
nor U2523 (N_2523,In_870,In_714);
or U2524 (N_2524,In_1028,In_9);
nand U2525 (N_2525,In_1442,In_417);
nor U2526 (N_2526,In_654,In_1412);
xor U2527 (N_2527,In_1132,In_463);
xnor U2528 (N_2528,In_1473,In_526);
or U2529 (N_2529,In_295,In_1318);
or U2530 (N_2530,In_243,In_269);
xnor U2531 (N_2531,In_922,In_148);
nand U2532 (N_2532,In_1474,In_1475);
and U2533 (N_2533,In_514,In_197);
or U2534 (N_2534,In_1325,In_1116);
nand U2535 (N_2535,In_208,In_44);
nand U2536 (N_2536,In_569,In_1120);
and U2537 (N_2537,In_10,In_835);
xnor U2538 (N_2538,In_901,In_441);
xnor U2539 (N_2539,In_212,In_516);
and U2540 (N_2540,In_1284,In_832);
xnor U2541 (N_2541,In_787,In_1206);
nor U2542 (N_2542,In_24,In_822);
nor U2543 (N_2543,In_1134,In_488);
nor U2544 (N_2544,In_548,In_178);
and U2545 (N_2545,In_1453,In_523);
xnor U2546 (N_2546,In_483,In_393);
xor U2547 (N_2547,In_445,In_874);
and U2548 (N_2548,In_1351,In_921);
and U2549 (N_2549,In_284,In_866);
nor U2550 (N_2550,In_1198,In_1138);
or U2551 (N_2551,In_802,In_96);
and U2552 (N_2552,In_195,In_1153);
xor U2553 (N_2553,In_849,In_459);
nand U2554 (N_2554,In_23,In_1467);
nand U2555 (N_2555,In_1262,In_207);
and U2556 (N_2556,In_1413,In_253);
and U2557 (N_2557,In_1008,In_663);
and U2558 (N_2558,In_650,In_1211);
xor U2559 (N_2559,In_721,In_905);
or U2560 (N_2560,In_1427,In_879);
nor U2561 (N_2561,In_314,In_408);
or U2562 (N_2562,In_728,In_1228);
xor U2563 (N_2563,In_847,In_447);
nor U2564 (N_2564,In_255,In_1193);
or U2565 (N_2565,In_792,In_260);
nor U2566 (N_2566,In_1327,In_262);
nor U2567 (N_2567,In_1217,In_1012);
and U2568 (N_2568,In_1064,In_731);
xor U2569 (N_2569,In_74,In_1090);
nand U2570 (N_2570,In_1125,In_1147);
and U2571 (N_2571,In_1415,In_441);
and U2572 (N_2572,In_863,In_283);
and U2573 (N_2573,In_1232,In_1371);
or U2574 (N_2574,In_479,In_924);
or U2575 (N_2575,In_79,In_136);
nand U2576 (N_2576,In_1481,In_953);
xnor U2577 (N_2577,In_1088,In_815);
or U2578 (N_2578,In_132,In_688);
nor U2579 (N_2579,In_486,In_15);
nand U2580 (N_2580,In_8,In_746);
nand U2581 (N_2581,In_779,In_332);
nand U2582 (N_2582,In_545,In_823);
xnor U2583 (N_2583,In_412,In_390);
nor U2584 (N_2584,In_601,In_1309);
and U2585 (N_2585,In_504,In_1362);
nor U2586 (N_2586,In_484,In_32);
and U2587 (N_2587,In_750,In_41);
nor U2588 (N_2588,In_1094,In_1062);
xor U2589 (N_2589,In_271,In_338);
or U2590 (N_2590,In_1174,In_68);
or U2591 (N_2591,In_427,In_1472);
and U2592 (N_2592,In_1166,In_1240);
or U2593 (N_2593,In_320,In_192);
xor U2594 (N_2594,In_1472,In_171);
or U2595 (N_2595,In_1215,In_626);
or U2596 (N_2596,In_1145,In_6);
nand U2597 (N_2597,In_309,In_748);
and U2598 (N_2598,In_1300,In_1097);
nor U2599 (N_2599,In_353,In_92);
and U2600 (N_2600,In_482,In_600);
nor U2601 (N_2601,In_794,In_1301);
xnor U2602 (N_2602,In_202,In_1147);
or U2603 (N_2603,In_715,In_1269);
nand U2604 (N_2604,In_27,In_264);
nor U2605 (N_2605,In_455,In_679);
and U2606 (N_2606,In_1483,In_1007);
nand U2607 (N_2607,In_1226,In_873);
xnor U2608 (N_2608,In_624,In_701);
and U2609 (N_2609,In_82,In_668);
nor U2610 (N_2610,In_967,In_1247);
nand U2611 (N_2611,In_712,In_1319);
xor U2612 (N_2612,In_736,In_576);
nand U2613 (N_2613,In_738,In_836);
or U2614 (N_2614,In_166,In_1423);
xnor U2615 (N_2615,In_580,In_1114);
and U2616 (N_2616,In_751,In_710);
or U2617 (N_2617,In_511,In_1233);
or U2618 (N_2618,In_921,In_1220);
nand U2619 (N_2619,In_425,In_1150);
and U2620 (N_2620,In_1174,In_1303);
or U2621 (N_2621,In_1407,In_1236);
nand U2622 (N_2622,In_1139,In_660);
and U2623 (N_2623,In_1070,In_302);
nor U2624 (N_2624,In_1448,In_1491);
or U2625 (N_2625,In_1332,In_1029);
or U2626 (N_2626,In_756,In_1173);
nand U2627 (N_2627,In_1152,In_620);
or U2628 (N_2628,In_1101,In_493);
xor U2629 (N_2629,In_333,In_31);
and U2630 (N_2630,In_340,In_314);
and U2631 (N_2631,In_806,In_122);
nor U2632 (N_2632,In_839,In_751);
nand U2633 (N_2633,In_1282,In_1212);
xnor U2634 (N_2634,In_460,In_566);
nand U2635 (N_2635,In_69,In_540);
or U2636 (N_2636,In_202,In_962);
and U2637 (N_2637,In_137,In_1393);
nor U2638 (N_2638,In_952,In_832);
and U2639 (N_2639,In_597,In_1211);
nor U2640 (N_2640,In_1263,In_758);
xor U2641 (N_2641,In_914,In_267);
nand U2642 (N_2642,In_1247,In_1266);
nor U2643 (N_2643,In_92,In_312);
nand U2644 (N_2644,In_73,In_460);
xnor U2645 (N_2645,In_321,In_35);
and U2646 (N_2646,In_1162,In_1018);
xnor U2647 (N_2647,In_376,In_868);
xor U2648 (N_2648,In_319,In_1168);
nand U2649 (N_2649,In_1201,In_726);
nand U2650 (N_2650,In_13,In_82);
and U2651 (N_2651,In_1462,In_1348);
nand U2652 (N_2652,In_621,In_550);
and U2653 (N_2653,In_341,In_193);
or U2654 (N_2654,In_585,In_430);
nor U2655 (N_2655,In_307,In_15);
or U2656 (N_2656,In_220,In_906);
xor U2657 (N_2657,In_1063,In_944);
or U2658 (N_2658,In_1145,In_1108);
and U2659 (N_2659,In_1114,In_1429);
xnor U2660 (N_2660,In_1362,In_952);
nor U2661 (N_2661,In_426,In_226);
nand U2662 (N_2662,In_682,In_1250);
or U2663 (N_2663,In_771,In_898);
and U2664 (N_2664,In_819,In_1246);
nand U2665 (N_2665,In_141,In_540);
nor U2666 (N_2666,In_1315,In_1443);
nand U2667 (N_2667,In_52,In_1126);
xnor U2668 (N_2668,In_997,In_1386);
nand U2669 (N_2669,In_1309,In_1005);
and U2670 (N_2670,In_587,In_884);
xor U2671 (N_2671,In_1036,In_409);
nand U2672 (N_2672,In_393,In_166);
or U2673 (N_2673,In_827,In_545);
nor U2674 (N_2674,In_1064,In_781);
and U2675 (N_2675,In_414,In_1239);
xor U2676 (N_2676,In_833,In_274);
or U2677 (N_2677,In_1295,In_14);
xnor U2678 (N_2678,In_146,In_1233);
or U2679 (N_2679,In_1405,In_385);
and U2680 (N_2680,In_889,In_950);
xor U2681 (N_2681,In_400,In_1348);
nand U2682 (N_2682,In_873,In_664);
nor U2683 (N_2683,In_67,In_598);
nand U2684 (N_2684,In_31,In_514);
nor U2685 (N_2685,In_389,In_117);
and U2686 (N_2686,In_906,In_1032);
xor U2687 (N_2687,In_407,In_1288);
and U2688 (N_2688,In_828,In_1213);
or U2689 (N_2689,In_261,In_1176);
nand U2690 (N_2690,In_946,In_1167);
nor U2691 (N_2691,In_327,In_279);
nand U2692 (N_2692,In_1450,In_1463);
nor U2693 (N_2693,In_180,In_1088);
or U2694 (N_2694,In_92,In_403);
nor U2695 (N_2695,In_1350,In_1389);
and U2696 (N_2696,In_786,In_1344);
xor U2697 (N_2697,In_1380,In_1304);
or U2698 (N_2698,In_1365,In_877);
xnor U2699 (N_2699,In_23,In_404);
nand U2700 (N_2700,In_582,In_1112);
nor U2701 (N_2701,In_847,In_413);
nand U2702 (N_2702,In_324,In_857);
nor U2703 (N_2703,In_332,In_1434);
or U2704 (N_2704,In_586,In_1392);
or U2705 (N_2705,In_291,In_762);
and U2706 (N_2706,In_17,In_675);
and U2707 (N_2707,In_421,In_509);
nor U2708 (N_2708,In_800,In_284);
or U2709 (N_2709,In_211,In_472);
or U2710 (N_2710,In_273,In_1165);
and U2711 (N_2711,In_24,In_1437);
or U2712 (N_2712,In_1281,In_1470);
and U2713 (N_2713,In_13,In_1233);
nor U2714 (N_2714,In_292,In_494);
nor U2715 (N_2715,In_1218,In_573);
and U2716 (N_2716,In_1340,In_10);
or U2717 (N_2717,In_777,In_448);
or U2718 (N_2718,In_1030,In_366);
nor U2719 (N_2719,In_1038,In_826);
nand U2720 (N_2720,In_845,In_528);
and U2721 (N_2721,In_1402,In_937);
or U2722 (N_2722,In_217,In_45);
or U2723 (N_2723,In_1151,In_1273);
and U2724 (N_2724,In_1079,In_1305);
nand U2725 (N_2725,In_4,In_1480);
xor U2726 (N_2726,In_1487,In_91);
nor U2727 (N_2727,In_112,In_582);
nand U2728 (N_2728,In_1024,In_48);
xor U2729 (N_2729,In_702,In_1102);
or U2730 (N_2730,In_1393,In_1088);
xor U2731 (N_2731,In_1423,In_129);
nor U2732 (N_2732,In_38,In_410);
and U2733 (N_2733,In_1149,In_544);
or U2734 (N_2734,In_1473,In_655);
or U2735 (N_2735,In_1267,In_1206);
xor U2736 (N_2736,In_1080,In_352);
nand U2737 (N_2737,In_229,In_1210);
nor U2738 (N_2738,In_1088,In_1220);
nor U2739 (N_2739,In_1299,In_764);
nand U2740 (N_2740,In_1121,In_345);
xor U2741 (N_2741,In_1147,In_569);
and U2742 (N_2742,In_1476,In_598);
and U2743 (N_2743,In_991,In_1435);
nand U2744 (N_2744,In_41,In_1403);
xnor U2745 (N_2745,In_41,In_364);
or U2746 (N_2746,In_840,In_598);
nand U2747 (N_2747,In_193,In_92);
nand U2748 (N_2748,In_367,In_97);
nor U2749 (N_2749,In_1307,In_51);
or U2750 (N_2750,In_747,In_770);
or U2751 (N_2751,In_1482,In_84);
or U2752 (N_2752,In_500,In_1222);
or U2753 (N_2753,In_567,In_360);
nor U2754 (N_2754,In_1359,In_798);
xor U2755 (N_2755,In_291,In_1403);
and U2756 (N_2756,In_548,In_1331);
or U2757 (N_2757,In_723,In_702);
and U2758 (N_2758,In_995,In_712);
xor U2759 (N_2759,In_1400,In_440);
xnor U2760 (N_2760,In_155,In_586);
xnor U2761 (N_2761,In_319,In_509);
xor U2762 (N_2762,In_338,In_928);
nor U2763 (N_2763,In_702,In_211);
nor U2764 (N_2764,In_804,In_484);
or U2765 (N_2765,In_802,In_690);
and U2766 (N_2766,In_1173,In_1287);
or U2767 (N_2767,In_165,In_1419);
nor U2768 (N_2768,In_872,In_457);
nand U2769 (N_2769,In_735,In_929);
and U2770 (N_2770,In_159,In_1267);
xnor U2771 (N_2771,In_453,In_804);
or U2772 (N_2772,In_1282,In_1429);
xnor U2773 (N_2773,In_431,In_226);
or U2774 (N_2774,In_140,In_971);
or U2775 (N_2775,In_284,In_158);
xnor U2776 (N_2776,In_1038,In_481);
nand U2777 (N_2777,In_1314,In_370);
nor U2778 (N_2778,In_89,In_1086);
nand U2779 (N_2779,In_91,In_164);
nand U2780 (N_2780,In_946,In_494);
and U2781 (N_2781,In_1433,In_460);
or U2782 (N_2782,In_793,In_251);
or U2783 (N_2783,In_194,In_789);
and U2784 (N_2784,In_716,In_1234);
or U2785 (N_2785,In_718,In_347);
nor U2786 (N_2786,In_1146,In_386);
nor U2787 (N_2787,In_1433,In_208);
xor U2788 (N_2788,In_1424,In_43);
or U2789 (N_2789,In_1324,In_178);
xor U2790 (N_2790,In_1062,In_1028);
and U2791 (N_2791,In_1247,In_1354);
nand U2792 (N_2792,In_99,In_956);
or U2793 (N_2793,In_990,In_1254);
or U2794 (N_2794,In_1458,In_382);
nor U2795 (N_2795,In_1166,In_902);
and U2796 (N_2796,In_628,In_239);
and U2797 (N_2797,In_620,In_704);
nand U2798 (N_2798,In_257,In_799);
or U2799 (N_2799,In_907,In_1293);
nand U2800 (N_2800,In_500,In_1475);
and U2801 (N_2801,In_196,In_709);
nand U2802 (N_2802,In_242,In_819);
and U2803 (N_2803,In_1162,In_385);
or U2804 (N_2804,In_939,In_1259);
nor U2805 (N_2805,In_345,In_1398);
nor U2806 (N_2806,In_828,In_5);
and U2807 (N_2807,In_782,In_49);
nand U2808 (N_2808,In_362,In_881);
xnor U2809 (N_2809,In_1118,In_851);
and U2810 (N_2810,In_691,In_27);
or U2811 (N_2811,In_955,In_799);
nand U2812 (N_2812,In_134,In_1307);
xnor U2813 (N_2813,In_650,In_780);
or U2814 (N_2814,In_262,In_623);
nor U2815 (N_2815,In_1463,In_35);
nand U2816 (N_2816,In_1142,In_1002);
and U2817 (N_2817,In_1484,In_4);
nand U2818 (N_2818,In_1385,In_371);
nand U2819 (N_2819,In_1273,In_41);
nand U2820 (N_2820,In_701,In_1306);
and U2821 (N_2821,In_1366,In_601);
nand U2822 (N_2822,In_308,In_1464);
or U2823 (N_2823,In_814,In_248);
and U2824 (N_2824,In_1420,In_1026);
nor U2825 (N_2825,In_228,In_847);
xor U2826 (N_2826,In_124,In_1121);
or U2827 (N_2827,In_101,In_89);
xnor U2828 (N_2828,In_940,In_311);
xor U2829 (N_2829,In_741,In_1334);
xor U2830 (N_2830,In_1205,In_447);
or U2831 (N_2831,In_170,In_126);
nor U2832 (N_2832,In_561,In_1284);
or U2833 (N_2833,In_50,In_950);
nor U2834 (N_2834,In_801,In_1100);
nand U2835 (N_2835,In_588,In_1060);
nor U2836 (N_2836,In_730,In_1314);
and U2837 (N_2837,In_934,In_505);
nand U2838 (N_2838,In_1347,In_888);
nor U2839 (N_2839,In_1418,In_1400);
xnor U2840 (N_2840,In_308,In_261);
nand U2841 (N_2841,In_945,In_799);
xnor U2842 (N_2842,In_389,In_1178);
and U2843 (N_2843,In_531,In_634);
xnor U2844 (N_2844,In_572,In_556);
or U2845 (N_2845,In_377,In_1274);
xnor U2846 (N_2846,In_335,In_1181);
or U2847 (N_2847,In_361,In_998);
and U2848 (N_2848,In_245,In_671);
nor U2849 (N_2849,In_903,In_234);
nor U2850 (N_2850,In_1117,In_748);
nor U2851 (N_2851,In_109,In_1014);
nand U2852 (N_2852,In_110,In_1332);
nor U2853 (N_2853,In_544,In_285);
nor U2854 (N_2854,In_717,In_1163);
nor U2855 (N_2855,In_391,In_600);
and U2856 (N_2856,In_931,In_1395);
xnor U2857 (N_2857,In_692,In_824);
nand U2858 (N_2858,In_823,In_103);
or U2859 (N_2859,In_215,In_452);
nand U2860 (N_2860,In_895,In_662);
nand U2861 (N_2861,In_1038,In_1332);
nand U2862 (N_2862,In_1100,In_1327);
or U2863 (N_2863,In_262,In_18);
xor U2864 (N_2864,In_95,In_978);
xnor U2865 (N_2865,In_501,In_1427);
xor U2866 (N_2866,In_277,In_1170);
nor U2867 (N_2867,In_116,In_520);
or U2868 (N_2868,In_469,In_494);
nor U2869 (N_2869,In_1445,In_879);
nand U2870 (N_2870,In_557,In_555);
nor U2871 (N_2871,In_1095,In_561);
and U2872 (N_2872,In_887,In_1267);
xor U2873 (N_2873,In_1093,In_282);
nor U2874 (N_2874,In_264,In_1313);
and U2875 (N_2875,In_325,In_1243);
and U2876 (N_2876,In_39,In_678);
xor U2877 (N_2877,In_263,In_1202);
xnor U2878 (N_2878,In_722,In_1446);
and U2879 (N_2879,In_397,In_242);
and U2880 (N_2880,In_764,In_547);
nor U2881 (N_2881,In_858,In_567);
or U2882 (N_2882,In_1217,In_527);
nand U2883 (N_2883,In_26,In_435);
xor U2884 (N_2884,In_577,In_1174);
and U2885 (N_2885,In_271,In_180);
or U2886 (N_2886,In_449,In_1044);
nand U2887 (N_2887,In_979,In_830);
xor U2888 (N_2888,In_1493,In_1379);
or U2889 (N_2889,In_1465,In_1327);
or U2890 (N_2890,In_1218,In_768);
xor U2891 (N_2891,In_395,In_1000);
xor U2892 (N_2892,In_1081,In_1398);
nor U2893 (N_2893,In_1438,In_1125);
nand U2894 (N_2894,In_663,In_590);
nor U2895 (N_2895,In_1076,In_389);
xor U2896 (N_2896,In_286,In_553);
xnor U2897 (N_2897,In_239,In_475);
xor U2898 (N_2898,In_784,In_435);
nand U2899 (N_2899,In_530,In_742);
xnor U2900 (N_2900,In_1471,In_706);
nand U2901 (N_2901,In_93,In_1257);
or U2902 (N_2902,In_304,In_216);
nor U2903 (N_2903,In_717,In_252);
or U2904 (N_2904,In_530,In_1126);
xnor U2905 (N_2905,In_1209,In_749);
nor U2906 (N_2906,In_189,In_696);
nand U2907 (N_2907,In_1314,In_1249);
and U2908 (N_2908,In_1211,In_228);
nor U2909 (N_2909,In_10,In_1045);
nand U2910 (N_2910,In_660,In_1096);
and U2911 (N_2911,In_195,In_1022);
and U2912 (N_2912,In_1202,In_12);
nor U2913 (N_2913,In_1448,In_414);
and U2914 (N_2914,In_1301,In_445);
or U2915 (N_2915,In_1190,In_791);
nand U2916 (N_2916,In_765,In_1399);
nor U2917 (N_2917,In_1169,In_974);
nor U2918 (N_2918,In_350,In_895);
or U2919 (N_2919,In_1092,In_791);
and U2920 (N_2920,In_767,In_1414);
nor U2921 (N_2921,In_1497,In_431);
nand U2922 (N_2922,In_404,In_321);
and U2923 (N_2923,In_1338,In_872);
nand U2924 (N_2924,In_175,In_668);
and U2925 (N_2925,In_958,In_273);
and U2926 (N_2926,In_1450,In_902);
xnor U2927 (N_2927,In_471,In_1035);
nand U2928 (N_2928,In_982,In_502);
and U2929 (N_2929,In_997,In_117);
nand U2930 (N_2930,In_276,In_1339);
nor U2931 (N_2931,In_1123,In_733);
and U2932 (N_2932,In_1163,In_967);
xor U2933 (N_2933,In_1454,In_471);
xor U2934 (N_2934,In_45,In_966);
nand U2935 (N_2935,In_181,In_414);
and U2936 (N_2936,In_231,In_1431);
or U2937 (N_2937,In_1312,In_405);
nor U2938 (N_2938,In_1133,In_1017);
xor U2939 (N_2939,In_723,In_1002);
nand U2940 (N_2940,In_1242,In_755);
and U2941 (N_2941,In_701,In_184);
nor U2942 (N_2942,In_730,In_532);
nand U2943 (N_2943,In_1405,In_392);
and U2944 (N_2944,In_542,In_715);
and U2945 (N_2945,In_1027,In_563);
and U2946 (N_2946,In_1148,In_686);
nand U2947 (N_2947,In_77,In_287);
nor U2948 (N_2948,In_19,In_606);
nor U2949 (N_2949,In_962,In_686);
nand U2950 (N_2950,In_488,In_524);
and U2951 (N_2951,In_1072,In_262);
and U2952 (N_2952,In_1231,In_521);
nor U2953 (N_2953,In_1228,In_1084);
or U2954 (N_2954,In_249,In_368);
xor U2955 (N_2955,In_1407,In_993);
nand U2956 (N_2956,In_1213,In_816);
nor U2957 (N_2957,In_200,In_1234);
and U2958 (N_2958,In_139,In_633);
nor U2959 (N_2959,In_1148,In_667);
nor U2960 (N_2960,In_660,In_457);
xnor U2961 (N_2961,In_72,In_299);
xnor U2962 (N_2962,In_22,In_1194);
or U2963 (N_2963,In_1441,In_800);
and U2964 (N_2964,In_1459,In_94);
and U2965 (N_2965,In_259,In_71);
or U2966 (N_2966,In_1410,In_961);
nor U2967 (N_2967,In_1346,In_1255);
and U2968 (N_2968,In_820,In_668);
nor U2969 (N_2969,In_602,In_1265);
xor U2970 (N_2970,In_841,In_1429);
or U2971 (N_2971,In_1036,In_175);
nand U2972 (N_2972,In_840,In_769);
xor U2973 (N_2973,In_562,In_621);
nor U2974 (N_2974,In_1343,In_1423);
or U2975 (N_2975,In_313,In_1332);
or U2976 (N_2976,In_300,In_326);
nand U2977 (N_2977,In_1053,In_1234);
nand U2978 (N_2978,In_1349,In_535);
nor U2979 (N_2979,In_1019,In_300);
nor U2980 (N_2980,In_826,In_68);
nor U2981 (N_2981,In_767,In_818);
or U2982 (N_2982,In_513,In_1256);
nand U2983 (N_2983,In_206,In_535);
or U2984 (N_2984,In_462,In_843);
and U2985 (N_2985,In_162,In_1489);
xor U2986 (N_2986,In_694,In_1235);
nor U2987 (N_2987,In_1359,In_965);
nand U2988 (N_2988,In_120,In_165);
xnor U2989 (N_2989,In_897,In_950);
or U2990 (N_2990,In_566,In_699);
and U2991 (N_2991,In_836,In_1492);
xor U2992 (N_2992,In_638,In_600);
xor U2993 (N_2993,In_366,In_689);
xor U2994 (N_2994,In_1071,In_247);
xor U2995 (N_2995,In_349,In_253);
nand U2996 (N_2996,In_424,In_508);
xnor U2997 (N_2997,In_908,In_835);
or U2998 (N_2998,In_1385,In_882);
nand U2999 (N_2999,In_912,In_1380);
xor U3000 (N_3000,In_854,In_1320);
xor U3001 (N_3001,In_1309,In_1051);
nand U3002 (N_3002,In_1405,In_346);
nor U3003 (N_3003,In_318,In_1446);
and U3004 (N_3004,In_127,In_1284);
nor U3005 (N_3005,In_1115,In_1125);
or U3006 (N_3006,In_1078,In_101);
and U3007 (N_3007,In_1290,In_421);
xor U3008 (N_3008,In_373,In_258);
xnor U3009 (N_3009,In_1264,In_1109);
nor U3010 (N_3010,In_167,In_1177);
nor U3011 (N_3011,In_71,In_715);
nor U3012 (N_3012,In_764,In_1134);
and U3013 (N_3013,In_1497,In_996);
nor U3014 (N_3014,In_1402,In_949);
and U3015 (N_3015,In_60,In_655);
nand U3016 (N_3016,In_1140,In_377);
or U3017 (N_3017,In_1152,In_731);
nand U3018 (N_3018,In_535,In_87);
and U3019 (N_3019,In_1398,In_1214);
nor U3020 (N_3020,In_700,In_493);
and U3021 (N_3021,In_685,In_1259);
nor U3022 (N_3022,In_1370,In_1249);
xor U3023 (N_3023,In_15,In_630);
nor U3024 (N_3024,In_366,In_241);
nand U3025 (N_3025,In_979,In_350);
nor U3026 (N_3026,In_1229,In_889);
nand U3027 (N_3027,In_969,In_15);
and U3028 (N_3028,In_644,In_388);
and U3029 (N_3029,In_1319,In_522);
nor U3030 (N_3030,In_728,In_299);
nor U3031 (N_3031,In_537,In_699);
xor U3032 (N_3032,In_406,In_814);
xnor U3033 (N_3033,In_1368,In_446);
nor U3034 (N_3034,In_1470,In_1326);
and U3035 (N_3035,In_562,In_1054);
xor U3036 (N_3036,In_482,In_414);
and U3037 (N_3037,In_1247,In_1239);
or U3038 (N_3038,In_863,In_288);
nand U3039 (N_3039,In_1387,In_1001);
nor U3040 (N_3040,In_1305,In_562);
nand U3041 (N_3041,In_379,In_1037);
or U3042 (N_3042,In_1218,In_685);
and U3043 (N_3043,In_753,In_319);
and U3044 (N_3044,In_304,In_503);
nand U3045 (N_3045,In_166,In_1087);
and U3046 (N_3046,In_430,In_894);
xor U3047 (N_3047,In_1473,In_1114);
nand U3048 (N_3048,In_664,In_1137);
nor U3049 (N_3049,In_1139,In_473);
and U3050 (N_3050,In_1115,In_745);
nor U3051 (N_3051,In_223,In_1039);
nand U3052 (N_3052,In_463,In_99);
nor U3053 (N_3053,In_396,In_605);
xor U3054 (N_3054,In_1214,In_122);
or U3055 (N_3055,In_1203,In_375);
and U3056 (N_3056,In_361,In_462);
nor U3057 (N_3057,In_519,In_525);
nor U3058 (N_3058,In_1398,In_755);
xor U3059 (N_3059,In_624,In_1328);
xor U3060 (N_3060,In_1415,In_466);
or U3061 (N_3061,In_1490,In_84);
nor U3062 (N_3062,In_1315,In_1095);
or U3063 (N_3063,In_118,In_896);
xor U3064 (N_3064,In_382,In_865);
xor U3065 (N_3065,In_902,In_1254);
xnor U3066 (N_3066,In_1183,In_560);
or U3067 (N_3067,In_1455,In_906);
xor U3068 (N_3068,In_476,In_360);
nor U3069 (N_3069,In_825,In_476);
nor U3070 (N_3070,In_1299,In_342);
or U3071 (N_3071,In_651,In_299);
or U3072 (N_3072,In_1249,In_1143);
nand U3073 (N_3073,In_647,In_761);
and U3074 (N_3074,In_1200,In_651);
or U3075 (N_3075,In_1134,In_249);
nor U3076 (N_3076,In_48,In_806);
nor U3077 (N_3077,In_375,In_1462);
nand U3078 (N_3078,In_434,In_1041);
nand U3079 (N_3079,In_813,In_1369);
or U3080 (N_3080,In_671,In_308);
and U3081 (N_3081,In_9,In_1136);
or U3082 (N_3082,In_65,In_546);
nand U3083 (N_3083,In_1236,In_439);
nor U3084 (N_3084,In_1407,In_1171);
or U3085 (N_3085,In_851,In_1427);
and U3086 (N_3086,In_1112,In_1200);
nor U3087 (N_3087,In_675,In_403);
nor U3088 (N_3088,In_208,In_1248);
nand U3089 (N_3089,In_1330,In_514);
and U3090 (N_3090,In_51,In_1359);
xnor U3091 (N_3091,In_38,In_1280);
nand U3092 (N_3092,In_259,In_449);
or U3093 (N_3093,In_1483,In_1345);
xor U3094 (N_3094,In_573,In_1452);
nor U3095 (N_3095,In_1146,In_533);
or U3096 (N_3096,In_1214,In_670);
or U3097 (N_3097,In_1149,In_49);
nor U3098 (N_3098,In_229,In_428);
nand U3099 (N_3099,In_1022,In_354);
nand U3100 (N_3100,In_342,In_710);
nand U3101 (N_3101,In_1375,In_411);
nor U3102 (N_3102,In_206,In_621);
nor U3103 (N_3103,In_1135,In_1179);
xnor U3104 (N_3104,In_9,In_226);
nor U3105 (N_3105,In_465,In_305);
or U3106 (N_3106,In_319,In_1431);
nor U3107 (N_3107,In_414,In_677);
and U3108 (N_3108,In_510,In_228);
nor U3109 (N_3109,In_405,In_603);
and U3110 (N_3110,In_1324,In_30);
xnor U3111 (N_3111,In_510,In_550);
or U3112 (N_3112,In_770,In_1372);
nand U3113 (N_3113,In_443,In_1372);
xnor U3114 (N_3114,In_149,In_323);
or U3115 (N_3115,In_175,In_1281);
nand U3116 (N_3116,In_1134,In_97);
and U3117 (N_3117,In_741,In_501);
xor U3118 (N_3118,In_333,In_1198);
xnor U3119 (N_3119,In_293,In_1390);
nor U3120 (N_3120,In_946,In_1093);
nor U3121 (N_3121,In_856,In_17);
xor U3122 (N_3122,In_302,In_840);
or U3123 (N_3123,In_178,In_286);
xnor U3124 (N_3124,In_236,In_1244);
nor U3125 (N_3125,In_482,In_40);
or U3126 (N_3126,In_202,In_1495);
and U3127 (N_3127,In_615,In_1102);
nand U3128 (N_3128,In_786,In_464);
or U3129 (N_3129,In_616,In_1385);
xnor U3130 (N_3130,In_600,In_516);
and U3131 (N_3131,In_1460,In_784);
or U3132 (N_3132,In_803,In_1121);
nand U3133 (N_3133,In_1144,In_1494);
nand U3134 (N_3134,In_780,In_1469);
xnor U3135 (N_3135,In_368,In_1143);
nor U3136 (N_3136,In_610,In_1084);
nor U3137 (N_3137,In_951,In_404);
nor U3138 (N_3138,In_13,In_758);
or U3139 (N_3139,In_1344,In_1309);
nand U3140 (N_3140,In_801,In_713);
and U3141 (N_3141,In_1205,In_641);
xor U3142 (N_3142,In_938,In_74);
or U3143 (N_3143,In_687,In_374);
xor U3144 (N_3144,In_1033,In_1063);
nand U3145 (N_3145,In_1357,In_206);
nor U3146 (N_3146,In_14,In_125);
and U3147 (N_3147,In_990,In_645);
xor U3148 (N_3148,In_409,In_1268);
nor U3149 (N_3149,In_88,In_978);
and U3150 (N_3150,In_56,In_453);
nor U3151 (N_3151,In_515,In_1020);
xor U3152 (N_3152,In_1060,In_147);
and U3153 (N_3153,In_1116,In_309);
and U3154 (N_3154,In_706,In_365);
or U3155 (N_3155,In_807,In_74);
xnor U3156 (N_3156,In_1080,In_1216);
xor U3157 (N_3157,In_1166,In_60);
or U3158 (N_3158,In_1444,In_255);
xnor U3159 (N_3159,In_1172,In_505);
nand U3160 (N_3160,In_701,In_107);
nand U3161 (N_3161,In_1022,In_679);
or U3162 (N_3162,In_1315,In_1092);
nand U3163 (N_3163,In_330,In_22);
nor U3164 (N_3164,In_1443,In_836);
or U3165 (N_3165,In_208,In_406);
nor U3166 (N_3166,In_1013,In_1201);
xor U3167 (N_3167,In_1182,In_261);
and U3168 (N_3168,In_1207,In_645);
or U3169 (N_3169,In_161,In_485);
xnor U3170 (N_3170,In_1441,In_1201);
xor U3171 (N_3171,In_407,In_899);
xnor U3172 (N_3172,In_609,In_895);
and U3173 (N_3173,In_949,In_429);
nor U3174 (N_3174,In_240,In_172);
xnor U3175 (N_3175,In_484,In_435);
nand U3176 (N_3176,In_1456,In_960);
nand U3177 (N_3177,In_657,In_212);
or U3178 (N_3178,In_903,In_1495);
nand U3179 (N_3179,In_1141,In_603);
and U3180 (N_3180,In_1201,In_290);
nand U3181 (N_3181,In_879,In_1394);
or U3182 (N_3182,In_1182,In_461);
nor U3183 (N_3183,In_870,In_60);
and U3184 (N_3184,In_282,In_904);
or U3185 (N_3185,In_571,In_190);
nor U3186 (N_3186,In_1202,In_996);
nand U3187 (N_3187,In_888,In_944);
nor U3188 (N_3188,In_88,In_700);
or U3189 (N_3189,In_691,In_1218);
or U3190 (N_3190,In_1063,In_983);
nor U3191 (N_3191,In_1080,In_847);
and U3192 (N_3192,In_343,In_1497);
xnor U3193 (N_3193,In_782,In_622);
xor U3194 (N_3194,In_314,In_688);
nand U3195 (N_3195,In_636,In_337);
or U3196 (N_3196,In_42,In_380);
or U3197 (N_3197,In_721,In_32);
or U3198 (N_3198,In_339,In_21);
nand U3199 (N_3199,In_519,In_256);
or U3200 (N_3200,In_1247,In_142);
xor U3201 (N_3201,In_405,In_356);
nand U3202 (N_3202,In_257,In_1019);
and U3203 (N_3203,In_975,In_392);
xnor U3204 (N_3204,In_1428,In_521);
nor U3205 (N_3205,In_1012,In_1070);
and U3206 (N_3206,In_1252,In_1223);
nor U3207 (N_3207,In_54,In_676);
nor U3208 (N_3208,In_473,In_1110);
and U3209 (N_3209,In_331,In_876);
and U3210 (N_3210,In_426,In_1474);
nand U3211 (N_3211,In_438,In_1103);
nand U3212 (N_3212,In_990,In_828);
and U3213 (N_3213,In_1483,In_719);
xnor U3214 (N_3214,In_858,In_358);
nand U3215 (N_3215,In_965,In_329);
nor U3216 (N_3216,In_280,In_335);
or U3217 (N_3217,In_1086,In_663);
and U3218 (N_3218,In_1341,In_400);
nand U3219 (N_3219,In_429,In_598);
and U3220 (N_3220,In_879,In_1087);
and U3221 (N_3221,In_932,In_131);
and U3222 (N_3222,In_224,In_617);
nor U3223 (N_3223,In_67,In_810);
nor U3224 (N_3224,In_9,In_1151);
and U3225 (N_3225,In_918,In_593);
nand U3226 (N_3226,In_648,In_1248);
nand U3227 (N_3227,In_254,In_912);
or U3228 (N_3228,In_34,In_1303);
nor U3229 (N_3229,In_19,In_400);
xor U3230 (N_3230,In_280,In_261);
nand U3231 (N_3231,In_805,In_30);
and U3232 (N_3232,In_625,In_623);
or U3233 (N_3233,In_847,In_663);
or U3234 (N_3234,In_132,In_1235);
nor U3235 (N_3235,In_1395,In_501);
nor U3236 (N_3236,In_479,In_683);
and U3237 (N_3237,In_792,In_739);
nand U3238 (N_3238,In_287,In_458);
xor U3239 (N_3239,In_1060,In_1369);
and U3240 (N_3240,In_301,In_1262);
and U3241 (N_3241,In_1350,In_187);
and U3242 (N_3242,In_1156,In_969);
nor U3243 (N_3243,In_935,In_1094);
nor U3244 (N_3244,In_1460,In_180);
nor U3245 (N_3245,In_1114,In_849);
xor U3246 (N_3246,In_1434,In_61);
or U3247 (N_3247,In_1403,In_209);
and U3248 (N_3248,In_360,In_287);
or U3249 (N_3249,In_647,In_231);
nor U3250 (N_3250,In_963,In_537);
and U3251 (N_3251,In_84,In_1097);
or U3252 (N_3252,In_675,In_1373);
nand U3253 (N_3253,In_1118,In_682);
nand U3254 (N_3254,In_364,In_129);
nor U3255 (N_3255,In_125,In_366);
xor U3256 (N_3256,In_222,In_759);
nor U3257 (N_3257,In_433,In_132);
nor U3258 (N_3258,In_514,In_466);
xnor U3259 (N_3259,In_189,In_718);
or U3260 (N_3260,In_485,In_1237);
nor U3261 (N_3261,In_451,In_639);
nor U3262 (N_3262,In_594,In_499);
xnor U3263 (N_3263,In_1418,In_1258);
nand U3264 (N_3264,In_537,In_1073);
or U3265 (N_3265,In_1331,In_1431);
nor U3266 (N_3266,In_1059,In_795);
xor U3267 (N_3267,In_445,In_923);
xnor U3268 (N_3268,In_707,In_582);
or U3269 (N_3269,In_1203,In_1365);
or U3270 (N_3270,In_708,In_262);
xnor U3271 (N_3271,In_1046,In_16);
nand U3272 (N_3272,In_914,In_1260);
nand U3273 (N_3273,In_847,In_893);
nor U3274 (N_3274,In_1032,In_257);
nor U3275 (N_3275,In_974,In_818);
or U3276 (N_3276,In_876,In_1309);
and U3277 (N_3277,In_910,In_1391);
and U3278 (N_3278,In_773,In_1461);
xnor U3279 (N_3279,In_751,In_1113);
xor U3280 (N_3280,In_366,In_1106);
nor U3281 (N_3281,In_457,In_56);
and U3282 (N_3282,In_915,In_269);
xnor U3283 (N_3283,In_342,In_619);
and U3284 (N_3284,In_270,In_1380);
or U3285 (N_3285,In_542,In_308);
nand U3286 (N_3286,In_195,In_512);
nor U3287 (N_3287,In_396,In_1058);
or U3288 (N_3288,In_988,In_474);
nand U3289 (N_3289,In_1155,In_137);
and U3290 (N_3290,In_1465,In_22);
nor U3291 (N_3291,In_1445,In_919);
xnor U3292 (N_3292,In_76,In_856);
and U3293 (N_3293,In_1388,In_102);
and U3294 (N_3294,In_1000,In_1476);
nor U3295 (N_3295,In_471,In_1455);
xnor U3296 (N_3296,In_1106,In_671);
nand U3297 (N_3297,In_1388,In_1278);
and U3298 (N_3298,In_1091,In_1351);
or U3299 (N_3299,In_764,In_1163);
and U3300 (N_3300,In_1250,In_527);
or U3301 (N_3301,In_1287,In_945);
nor U3302 (N_3302,In_822,In_1247);
nor U3303 (N_3303,In_247,In_1018);
or U3304 (N_3304,In_347,In_1074);
and U3305 (N_3305,In_267,In_347);
and U3306 (N_3306,In_1042,In_122);
nor U3307 (N_3307,In_801,In_978);
xor U3308 (N_3308,In_976,In_1287);
nor U3309 (N_3309,In_695,In_1235);
and U3310 (N_3310,In_1111,In_927);
and U3311 (N_3311,In_756,In_169);
or U3312 (N_3312,In_854,In_1147);
xor U3313 (N_3313,In_890,In_1333);
xnor U3314 (N_3314,In_28,In_577);
and U3315 (N_3315,In_723,In_1270);
nand U3316 (N_3316,In_1365,In_837);
and U3317 (N_3317,In_230,In_1354);
nand U3318 (N_3318,In_916,In_1196);
or U3319 (N_3319,In_1179,In_122);
and U3320 (N_3320,In_504,In_1314);
nand U3321 (N_3321,In_448,In_1399);
nand U3322 (N_3322,In_632,In_593);
and U3323 (N_3323,In_471,In_707);
and U3324 (N_3324,In_525,In_1389);
xnor U3325 (N_3325,In_546,In_804);
and U3326 (N_3326,In_461,In_598);
or U3327 (N_3327,In_1249,In_813);
and U3328 (N_3328,In_1478,In_400);
nand U3329 (N_3329,In_1359,In_60);
nor U3330 (N_3330,In_284,In_482);
xnor U3331 (N_3331,In_277,In_53);
or U3332 (N_3332,In_3,In_163);
and U3333 (N_3333,In_1300,In_429);
xor U3334 (N_3334,In_686,In_1158);
and U3335 (N_3335,In_259,In_666);
nand U3336 (N_3336,In_361,In_322);
xnor U3337 (N_3337,In_829,In_1064);
nor U3338 (N_3338,In_473,In_674);
xnor U3339 (N_3339,In_1421,In_1099);
and U3340 (N_3340,In_1255,In_186);
xor U3341 (N_3341,In_139,In_724);
xor U3342 (N_3342,In_717,In_620);
xnor U3343 (N_3343,In_7,In_537);
nand U3344 (N_3344,In_811,In_1322);
and U3345 (N_3345,In_1118,In_182);
xnor U3346 (N_3346,In_1449,In_1394);
nor U3347 (N_3347,In_166,In_1282);
and U3348 (N_3348,In_1021,In_996);
nor U3349 (N_3349,In_1281,In_1357);
and U3350 (N_3350,In_544,In_1306);
and U3351 (N_3351,In_795,In_77);
nand U3352 (N_3352,In_1227,In_680);
and U3353 (N_3353,In_396,In_599);
or U3354 (N_3354,In_24,In_1463);
nor U3355 (N_3355,In_1378,In_1063);
nand U3356 (N_3356,In_184,In_204);
and U3357 (N_3357,In_321,In_995);
nor U3358 (N_3358,In_1035,In_425);
nand U3359 (N_3359,In_1,In_745);
xnor U3360 (N_3360,In_326,In_1083);
xor U3361 (N_3361,In_990,In_664);
or U3362 (N_3362,In_46,In_854);
and U3363 (N_3363,In_1365,In_226);
xnor U3364 (N_3364,In_862,In_1338);
and U3365 (N_3365,In_911,In_1380);
and U3366 (N_3366,In_693,In_1166);
and U3367 (N_3367,In_64,In_391);
xnor U3368 (N_3368,In_1360,In_177);
and U3369 (N_3369,In_1263,In_618);
or U3370 (N_3370,In_594,In_237);
xnor U3371 (N_3371,In_766,In_1395);
and U3372 (N_3372,In_767,In_1368);
or U3373 (N_3373,In_1077,In_978);
xor U3374 (N_3374,In_442,In_837);
nand U3375 (N_3375,In_861,In_49);
nor U3376 (N_3376,In_1071,In_1325);
and U3377 (N_3377,In_478,In_15);
nand U3378 (N_3378,In_1171,In_124);
nor U3379 (N_3379,In_1175,In_26);
and U3380 (N_3380,In_1033,In_497);
nand U3381 (N_3381,In_1364,In_570);
nor U3382 (N_3382,In_708,In_501);
nand U3383 (N_3383,In_984,In_499);
nand U3384 (N_3384,In_1484,In_106);
nor U3385 (N_3385,In_886,In_470);
nor U3386 (N_3386,In_1215,In_441);
nand U3387 (N_3387,In_623,In_610);
nand U3388 (N_3388,In_549,In_876);
and U3389 (N_3389,In_835,In_3);
or U3390 (N_3390,In_678,In_355);
or U3391 (N_3391,In_1216,In_953);
or U3392 (N_3392,In_743,In_1222);
nand U3393 (N_3393,In_175,In_1319);
nor U3394 (N_3394,In_1236,In_1043);
xor U3395 (N_3395,In_1402,In_1113);
nor U3396 (N_3396,In_893,In_491);
nor U3397 (N_3397,In_1113,In_834);
nor U3398 (N_3398,In_238,In_211);
xnor U3399 (N_3399,In_1256,In_1208);
nor U3400 (N_3400,In_634,In_792);
and U3401 (N_3401,In_232,In_167);
and U3402 (N_3402,In_225,In_1435);
nor U3403 (N_3403,In_356,In_512);
nor U3404 (N_3404,In_1040,In_1343);
and U3405 (N_3405,In_322,In_1411);
and U3406 (N_3406,In_467,In_1444);
and U3407 (N_3407,In_1442,In_1299);
or U3408 (N_3408,In_1483,In_198);
and U3409 (N_3409,In_1098,In_747);
nand U3410 (N_3410,In_331,In_216);
or U3411 (N_3411,In_769,In_1186);
and U3412 (N_3412,In_58,In_966);
and U3413 (N_3413,In_537,In_1224);
and U3414 (N_3414,In_991,In_1449);
or U3415 (N_3415,In_818,In_32);
nor U3416 (N_3416,In_1271,In_948);
nand U3417 (N_3417,In_1264,In_67);
and U3418 (N_3418,In_1107,In_952);
nor U3419 (N_3419,In_1376,In_1465);
or U3420 (N_3420,In_234,In_355);
or U3421 (N_3421,In_999,In_1293);
nor U3422 (N_3422,In_728,In_325);
nand U3423 (N_3423,In_906,In_452);
xor U3424 (N_3424,In_1314,In_520);
nand U3425 (N_3425,In_1235,In_680);
nor U3426 (N_3426,In_119,In_501);
nand U3427 (N_3427,In_1329,In_28);
xor U3428 (N_3428,In_560,In_429);
or U3429 (N_3429,In_502,In_1330);
nor U3430 (N_3430,In_811,In_1454);
and U3431 (N_3431,In_821,In_780);
nor U3432 (N_3432,In_1004,In_1094);
or U3433 (N_3433,In_238,In_716);
or U3434 (N_3434,In_1418,In_223);
nand U3435 (N_3435,In_772,In_211);
xnor U3436 (N_3436,In_20,In_1141);
and U3437 (N_3437,In_734,In_546);
xnor U3438 (N_3438,In_302,In_375);
xnor U3439 (N_3439,In_1156,In_814);
nand U3440 (N_3440,In_1490,In_953);
or U3441 (N_3441,In_722,In_92);
nand U3442 (N_3442,In_67,In_895);
nor U3443 (N_3443,In_1265,In_761);
xor U3444 (N_3444,In_479,In_1335);
nand U3445 (N_3445,In_442,In_540);
nand U3446 (N_3446,In_1218,In_240);
or U3447 (N_3447,In_628,In_948);
xor U3448 (N_3448,In_1092,In_829);
nor U3449 (N_3449,In_1342,In_792);
or U3450 (N_3450,In_519,In_740);
xor U3451 (N_3451,In_333,In_270);
nand U3452 (N_3452,In_981,In_1044);
or U3453 (N_3453,In_1499,In_753);
nor U3454 (N_3454,In_1234,In_1061);
nor U3455 (N_3455,In_1252,In_1081);
or U3456 (N_3456,In_983,In_1101);
xor U3457 (N_3457,In_566,In_1254);
xor U3458 (N_3458,In_8,In_1110);
or U3459 (N_3459,In_745,In_505);
or U3460 (N_3460,In_1133,In_1117);
and U3461 (N_3461,In_1457,In_752);
nand U3462 (N_3462,In_256,In_900);
xnor U3463 (N_3463,In_1278,In_780);
or U3464 (N_3464,In_498,In_32);
or U3465 (N_3465,In_26,In_878);
nor U3466 (N_3466,In_1484,In_1077);
nor U3467 (N_3467,In_635,In_232);
nand U3468 (N_3468,In_392,In_646);
xnor U3469 (N_3469,In_279,In_145);
nand U3470 (N_3470,In_1259,In_843);
or U3471 (N_3471,In_1332,In_1010);
and U3472 (N_3472,In_1115,In_1473);
and U3473 (N_3473,In_1407,In_885);
nor U3474 (N_3474,In_1074,In_272);
xor U3475 (N_3475,In_1111,In_364);
nor U3476 (N_3476,In_1378,In_845);
and U3477 (N_3477,In_578,In_1324);
xor U3478 (N_3478,In_620,In_742);
and U3479 (N_3479,In_324,In_572);
xor U3480 (N_3480,In_986,In_195);
nor U3481 (N_3481,In_1150,In_1021);
or U3482 (N_3482,In_1326,In_205);
nand U3483 (N_3483,In_632,In_563);
nor U3484 (N_3484,In_503,In_1376);
nor U3485 (N_3485,In_876,In_313);
or U3486 (N_3486,In_946,In_1274);
nand U3487 (N_3487,In_728,In_1123);
nor U3488 (N_3488,In_644,In_771);
and U3489 (N_3489,In_1049,In_1396);
nor U3490 (N_3490,In_1312,In_237);
and U3491 (N_3491,In_1047,In_564);
or U3492 (N_3492,In_1218,In_709);
and U3493 (N_3493,In_381,In_71);
and U3494 (N_3494,In_1481,In_1165);
nand U3495 (N_3495,In_47,In_421);
and U3496 (N_3496,In_1081,In_610);
and U3497 (N_3497,In_698,In_267);
xor U3498 (N_3498,In_1058,In_291);
and U3499 (N_3499,In_425,In_802);
nor U3500 (N_3500,In_875,In_414);
or U3501 (N_3501,In_226,In_1206);
nor U3502 (N_3502,In_1398,In_1466);
and U3503 (N_3503,In_863,In_949);
nand U3504 (N_3504,In_135,In_875);
nor U3505 (N_3505,In_194,In_106);
xnor U3506 (N_3506,In_947,In_573);
xnor U3507 (N_3507,In_123,In_538);
nor U3508 (N_3508,In_833,In_1182);
and U3509 (N_3509,In_119,In_1423);
and U3510 (N_3510,In_691,In_840);
and U3511 (N_3511,In_516,In_1482);
or U3512 (N_3512,In_477,In_843);
xnor U3513 (N_3513,In_442,In_1454);
or U3514 (N_3514,In_1283,In_252);
and U3515 (N_3515,In_1203,In_1354);
nor U3516 (N_3516,In_878,In_364);
nor U3517 (N_3517,In_1452,In_928);
or U3518 (N_3518,In_860,In_587);
and U3519 (N_3519,In_625,In_1134);
and U3520 (N_3520,In_980,In_368);
xnor U3521 (N_3521,In_811,In_134);
and U3522 (N_3522,In_303,In_638);
xor U3523 (N_3523,In_336,In_924);
nor U3524 (N_3524,In_455,In_402);
xor U3525 (N_3525,In_89,In_679);
nor U3526 (N_3526,In_336,In_194);
or U3527 (N_3527,In_331,In_390);
and U3528 (N_3528,In_399,In_183);
nor U3529 (N_3529,In_46,In_341);
and U3530 (N_3530,In_630,In_779);
and U3531 (N_3531,In_163,In_322);
and U3532 (N_3532,In_781,In_375);
nor U3533 (N_3533,In_145,In_182);
and U3534 (N_3534,In_77,In_59);
or U3535 (N_3535,In_891,In_147);
and U3536 (N_3536,In_1379,In_1143);
xor U3537 (N_3537,In_773,In_1196);
and U3538 (N_3538,In_853,In_682);
and U3539 (N_3539,In_885,In_581);
or U3540 (N_3540,In_452,In_912);
nand U3541 (N_3541,In_654,In_21);
or U3542 (N_3542,In_256,In_620);
nand U3543 (N_3543,In_560,In_754);
or U3544 (N_3544,In_199,In_1272);
nand U3545 (N_3545,In_634,In_315);
nand U3546 (N_3546,In_773,In_27);
and U3547 (N_3547,In_856,In_1129);
or U3548 (N_3548,In_568,In_1136);
and U3549 (N_3549,In_1049,In_1453);
xnor U3550 (N_3550,In_847,In_291);
nor U3551 (N_3551,In_470,In_588);
and U3552 (N_3552,In_1192,In_478);
nand U3553 (N_3553,In_1349,In_1279);
and U3554 (N_3554,In_431,In_7);
nor U3555 (N_3555,In_1444,In_187);
nor U3556 (N_3556,In_1325,In_1460);
xor U3557 (N_3557,In_335,In_832);
and U3558 (N_3558,In_1271,In_841);
nand U3559 (N_3559,In_398,In_708);
nor U3560 (N_3560,In_1224,In_1491);
and U3561 (N_3561,In_212,In_1055);
nor U3562 (N_3562,In_759,In_987);
xnor U3563 (N_3563,In_1051,In_59);
nor U3564 (N_3564,In_371,In_532);
or U3565 (N_3565,In_1068,In_1131);
or U3566 (N_3566,In_1396,In_523);
xor U3567 (N_3567,In_1026,In_457);
nand U3568 (N_3568,In_464,In_82);
xor U3569 (N_3569,In_23,In_602);
nor U3570 (N_3570,In_210,In_1237);
or U3571 (N_3571,In_244,In_1362);
nor U3572 (N_3572,In_1178,In_1001);
or U3573 (N_3573,In_1040,In_684);
and U3574 (N_3574,In_1486,In_228);
and U3575 (N_3575,In_49,In_328);
nor U3576 (N_3576,In_1348,In_125);
xor U3577 (N_3577,In_603,In_142);
nand U3578 (N_3578,In_546,In_1036);
or U3579 (N_3579,In_36,In_1017);
nor U3580 (N_3580,In_521,In_11);
nor U3581 (N_3581,In_1423,In_141);
or U3582 (N_3582,In_1247,In_440);
nor U3583 (N_3583,In_98,In_1095);
nand U3584 (N_3584,In_480,In_424);
and U3585 (N_3585,In_501,In_1429);
nand U3586 (N_3586,In_791,In_1014);
nor U3587 (N_3587,In_515,In_1332);
and U3588 (N_3588,In_1379,In_403);
nor U3589 (N_3589,In_858,In_836);
xnor U3590 (N_3590,In_807,In_1223);
or U3591 (N_3591,In_594,In_1207);
and U3592 (N_3592,In_564,In_204);
nand U3593 (N_3593,In_1168,In_1155);
nor U3594 (N_3594,In_1013,In_537);
nand U3595 (N_3595,In_1174,In_177);
and U3596 (N_3596,In_297,In_499);
and U3597 (N_3597,In_1004,In_318);
nor U3598 (N_3598,In_1383,In_497);
and U3599 (N_3599,In_1263,In_857);
nor U3600 (N_3600,In_274,In_467);
xnor U3601 (N_3601,In_900,In_715);
nor U3602 (N_3602,In_340,In_178);
xnor U3603 (N_3603,In_1093,In_1012);
xor U3604 (N_3604,In_525,In_675);
and U3605 (N_3605,In_281,In_414);
or U3606 (N_3606,In_921,In_1124);
and U3607 (N_3607,In_156,In_280);
xor U3608 (N_3608,In_223,In_541);
xnor U3609 (N_3609,In_1457,In_581);
xnor U3610 (N_3610,In_582,In_1155);
or U3611 (N_3611,In_302,In_1479);
and U3612 (N_3612,In_1051,In_1195);
nor U3613 (N_3613,In_1061,In_746);
xor U3614 (N_3614,In_964,In_209);
nand U3615 (N_3615,In_1126,In_444);
or U3616 (N_3616,In_1148,In_1437);
nor U3617 (N_3617,In_469,In_1017);
xor U3618 (N_3618,In_326,In_973);
xor U3619 (N_3619,In_1185,In_1213);
xor U3620 (N_3620,In_1206,In_496);
nand U3621 (N_3621,In_126,In_917);
xor U3622 (N_3622,In_285,In_639);
nor U3623 (N_3623,In_772,In_607);
xor U3624 (N_3624,In_759,In_1374);
nor U3625 (N_3625,In_666,In_30);
xnor U3626 (N_3626,In_41,In_494);
nand U3627 (N_3627,In_1007,In_1129);
or U3628 (N_3628,In_736,In_652);
and U3629 (N_3629,In_1253,In_459);
nand U3630 (N_3630,In_390,In_562);
xnor U3631 (N_3631,In_579,In_528);
nor U3632 (N_3632,In_372,In_1132);
or U3633 (N_3633,In_1425,In_816);
and U3634 (N_3634,In_1486,In_13);
or U3635 (N_3635,In_705,In_1164);
nand U3636 (N_3636,In_1074,In_1124);
or U3637 (N_3637,In_513,In_1129);
or U3638 (N_3638,In_1346,In_297);
or U3639 (N_3639,In_98,In_856);
nor U3640 (N_3640,In_938,In_206);
xor U3641 (N_3641,In_1255,In_985);
xnor U3642 (N_3642,In_355,In_980);
and U3643 (N_3643,In_220,In_701);
or U3644 (N_3644,In_857,In_628);
xor U3645 (N_3645,In_289,In_982);
or U3646 (N_3646,In_599,In_324);
and U3647 (N_3647,In_1418,In_123);
and U3648 (N_3648,In_455,In_1352);
or U3649 (N_3649,In_1433,In_129);
nand U3650 (N_3650,In_772,In_141);
and U3651 (N_3651,In_661,In_20);
xor U3652 (N_3652,In_1378,In_746);
and U3653 (N_3653,In_604,In_1285);
nand U3654 (N_3654,In_1353,In_630);
or U3655 (N_3655,In_265,In_884);
nand U3656 (N_3656,In_166,In_1080);
or U3657 (N_3657,In_1167,In_768);
xor U3658 (N_3658,In_588,In_58);
and U3659 (N_3659,In_23,In_277);
or U3660 (N_3660,In_568,In_870);
nor U3661 (N_3661,In_1209,In_813);
xnor U3662 (N_3662,In_1143,In_1360);
nand U3663 (N_3663,In_1003,In_933);
xnor U3664 (N_3664,In_540,In_201);
xnor U3665 (N_3665,In_1318,In_25);
xnor U3666 (N_3666,In_790,In_770);
xor U3667 (N_3667,In_1446,In_1272);
nor U3668 (N_3668,In_300,In_46);
xor U3669 (N_3669,In_1350,In_1169);
and U3670 (N_3670,In_52,In_133);
xor U3671 (N_3671,In_698,In_1448);
nand U3672 (N_3672,In_1109,In_1025);
and U3673 (N_3673,In_281,In_255);
or U3674 (N_3674,In_884,In_1076);
and U3675 (N_3675,In_1097,In_1016);
nor U3676 (N_3676,In_817,In_670);
or U3677 (N_3677,In_831,In_281);
nor U3678 (N_3678,In_764,In_1347);
and U3679 (N_3679,In_1298,In_1329);
nor U3680 (N_3680,In_394,In_257);
or U3681 (N_3681,In_462,In_1051);
or U3682 (N_3682,In_1168,In_923);
xnor U3683 (N_3683,In_880,In_665);
and U3684 (N_3684,In_264,In_436);
or U3685 (N_3685,In_802,In_589);
xor U3686 (N_3686,In_31,In_1000);
nor U3687 (N_3687,In_36,In_517);
nor U3688 (N_3688,In_1110,In_242);
and U3689 (N_3689,In_771,In_1044);
xor U3690 (N_3690,In_265,In_268);
and U3691 (N_3691,In_34,In_561);
nor U3692 (N_3692,In_832,In_1474);
nor U3693 (N_3693,In_966,In_1185);
nand U3694 (N_3694,In_59,In_474);
and U3695 (N_3695,In_1351,In_645);
nor U3696 (N_3696,In_1474,In_830);
xnor U3697 (N_3697,In_493,In_964);
xnor U3698 (N_3698,In_287,In_50);
nand U3699 (N_3699,In_584,In_1307);
nand U3700 (N_3700,In_565,In_334);
nand U3701 (N_3701,In_920,In_191);
xnor U3702 (N_3702,In_465,In_1478);
and U3703 (N_3703,In_564,In_125);
nand U3704 (N_3704,In_140,In_1393);
nand U3705 (N_3705,In_280,In_528);
xor U3706 (N_3706,In_308,In_767);
and U3707 (N_3707,In_1204,In_1487);
nand U3708 (N_3708,In_1221,In_1321);
nand U3709 (N_3709,In_836,In_0);
xnor U3710 (N_3710,In_918,In_459);
or U3711 (N_3711,In_1266,In_1318);
and U3712 (N_3712,In_791,In_1143);
xnor U3713 (N_3713,In_1366,In_359);
nor U3714 (N_3714,In_331,In_1162);
nand U3715 (N_3715,In_183,In_1442);
and U3716 (N_3716,In_1045,In_348);
or U3717 (N_3717,In_42,In_820);
or U3718 (N_3718,In_950,In_494);
or U3719 (N_3719,In_1477,In_652);
and U3720 (N_3720,In_198,In_1);
nor U3721 (N_3721,In_704,In_1448);
nor U3722 (N_3722,In_780,In_500);
or U3723 (N_3723,In_760,In_388);
or U3724 (N_3724,In_238,In_1103);
nand U3725 (N_3725,In_224,In_87);
nand U3726 (N_3726,In_393,In_926);
or U3727 (N_3727,In_665,In_685);
nor U3728 (N_3728,In_486,In_1193);
and U3729 (N_3729,In_944,In_685);
nand U3730 (N_3730,In_1317,In_1230);
xnor U3731 (N_3731,In_292,In_923);
nand U3732 (N_3732,In_482,In_1005);
nand U3733 (N_3733,In_1229,In_366);
nor U3734 (N_3734,In_615,In_666);
nand U3735 (N_3735,In_94,In_151);
nand U3736 (N_3736,In_164,In_1270);
or U3737 (N_3737,In_29,In_1061);
nor U3738 (N_3738,In_399,In_1026);
nand U3739 (N_3739,In_1399,In_1364);
or U3740 (N_3740,In_894,In_837);
or U3741 (N_3741,In_362,In_601);
nand U3742 (N_3742,In_1343,In_879);
xor U3743 (N_3743,In_965,In_1056);
nor U3744 (N_3744,In_876,In_379);
nor U3745 (N_3745,In_696,In_759);
or U3746 (N_3746,In_1143,In_239);
or U3747 (N_3747,In_1430,In_1001);
or U3748 (N_3748,In_471,In_1133);
and U3749 (N_3749,In_566,In_445);
and U3750 (N_3750,In_766,In_796);
xnor U3751 (N_3751,In_827,In_920);
xnor U3752 (N_3752,In_1096,In_1107);
nor U3753 (N_3753,In_301,In_173);
and U3754 (N_3754,In_689,In_473);
nand U3755 (N_3755,In_577,In_1241);
nor U3756 (N_3756,In_547,In_123);
nand U3757 (N_3757,In_1006,In_793);
nor U3758 (N_3758,In_13,In_1448);
or U3759 (N_3759,In_641,In_1039);
and U3760 (N_3760,In_921,In_231);
nor U3761 (N_3761,In_394,In_1127);
nand U3762 (N_3762,In_529,In_606);
or U3763 (N_3763,In_1068,In_1224);
or U3764 (N_3764,In_820,In_348);
xor U3765 (N_3765,In_168,In_975);
and U3766 (N_3766,In_625,In_962);
nand U3767 (N_3767,In_891,In_236);
xnor U3768 (N_3768,In_411,In_294);
nand U3769 (N_3769,In_396,In_977);
or U3770 (N_3770,In_435,In_717);
and U3771 (N_3771,In_150,In_1383);
nand U3772 (N_3772,In_251,In_911);
or U3773 (N_3773,In_1141,In_751);
or U3774 (N_3774,In_369,In_395);
nand U3775 (N_3775,In_733,In_1263);
or U3776 (N_3776,In_624,In_1015);
xnor U3777 (N_3777,In_381,In_166);
nand U3778 (N_3778,In_280,In_589);
or U3779 (N_3779,In_786,In_1372);
and U3780 (N_3780,In_766,In_53);
and U3781 (N_3781,In_687,In_1138);
or U3782 (N_3782,In_165,In_240);
and U3783 (N_3783,In_169,In_1490);
or U3784 (N_3784,In_142,In_434);
or U3785 (N_3785,In_880,In_539);
or U3786 (N_3786,In_647,In_1092);
nand U3787 (N_3787,In_728,In_917);
nand U3788 (N_3788,In_1344,In_577);
nor U3789 (N_3789,In_1299,In_140);
xnor U3790 (N_3790,In_1009,In_245);
nand U3791 (N_3791,In_1284,In_129);
xor U3792 (N_3792,In_114,In_1199);
and U3793 (N_3793,In_214,In_1003);
nand U3794 (N_3794,In_1291,In_1200);
and U3795 (N_3795,In_722,In_474);
and U3796 (N_3796,In_631,In_998);
and U3797 (N_3797,In_984,In_1243);
xor U3798 (N_3798,In_89,In_152);
nor U3799 (N_3799,In_1470,In_675);
nand U3800 (N_3800,In_1339,In_691);
and U3801 (N_3801,In_1389,In_1374);
and U3802 (N_3802,In_301,In_278);
nand U3803 (N_3803,In_1270,In_155);
and U3804 (N_3804,In_403,In_626);
nor U3805 (N_3805,In_1391,In_214);
nand U3806 (N_3806,In_64,In_1004);
nand U3807 (N_3807,In_265,In_17);
and U3808 (N_3808,In_1421,In_1024);
or U3809 (N_3809,In_941,In_551);
nand U3810 (N_3810,In_353,In_885);
xor U3811 (N_3811,In_41,In_1158);
xnor U3812 (N_3812,In_1191,In_1120);
and U3813 (N_3813,In_1491,In_973);
nand U3814 (N_3814,In_866,In_1126);
and U3815 (N_3815,In_340,In_1384);
nor U3816 (N_3816,In_1379,In_1336);
or U3817 (N_3817,In_1121,In_879);
nor U3818 (N_3818,In_215,In_778);
nor U3819 (N_3819,In_646,In_997);
nor U3820 (N_3820,In_292,In_949);
xnor U3821 (N_3821,In_864,In_804);
and U3822 (N_3822,In_643,In_887);
and U3823 (N_3823,In_153,In_938);
xnor U3824 (N_3824,In_680,In_333);
nor U3825 (N_3825,In_1233,In_805);
or U3826 (N_3826,In_1497,In_667);
xnor U3827 (N_3827,In_677,In_590);
and U3828 (N_3828,In_66,In_52);
nor U3829 (N_3829,In_1468,In_189);
nand U3830 (N_3830,In_1012,In_1262);
or U3831 (N_3831,In_240,In_1235);
and U3832 (N_3832,In_1151,In_544);
xor U3833 (N_3833,In_497,In_1316);
nand U3834 (N_3834,In_380,In_547);
nand U3835 (N_3835,In_162,In_1279);
and U3836 (N_3836,In_558,In_1126);
xor U3837 (N_3837,In_1163,In_1368);
xor U3838 (N_3838,In_1353,In_1193);
and U3839 (N_3839,In_388,In_1352);
or U3840 (N_3840,In_473,In_516);
nand U3841 (N_3841,In_1199,In_476);
or U3842 (N_3842,In_22,In_357);
or U3843 (N_3843,In_1018,In_549);
and U3844 (N_3844,In_212,In_1388);
or U3845 (N_3845,In_1184,In_354);
xnor U3846 (N_3846,In_218,In_87);
nor U3847 (N_3847,In_231,In_610);
nor U3848 (N_3848,In_225,In_1454);
nor U3849 (N_3849,In_933,In_1155);
xor U3850 (N_3850,In_1156,In_824);
nor U3851 (N_3851,In_1462,In_920);
or U3852 (N_3852,In_474,In_1115);
xor U3853 (N_3853,In_40,In_1121);
xnor U3854 (N_3854,In_865,In_1357);
and U3855 (N_3855,In_242,In_483);
nor U3856 (N_3856,In_1268,In_882);
nor U3857 (N_3857,In_1361,In_28);
nor U3858 (N_3858,In_1348,In_298);
xor U3859 (N_3859,In_96,In_141);
xor U3860 (N_3860,In_406,In_571);
and U3861 (N_3861,In_1224,In_813);
nand U3862 (N_3862,In_753,In_326);
nor U3863 (N_3863,In_1370,In_782);
or U3864 (N_3864,In_143,In_690);
xor U3865 (N_3865,In_657,In_1411);
and U3866 (N_3866,In_722,In_1167);
nor U3867 (N_3867,In_520,In_283);
nor U3868 (N_3868,In_1024,In_578);
xor U3869 (N_3869,In_183,In_752);
and U3870 (N_3870,In_445,In_191);
and U3871 (N_3871,In_522,In_1276);
nor U3872 (N_3872,In_643,In_41);
or U3873 (N_3873,In_1312,In_133);
nor U3874 (N_3874,In_970,In_1298);
nand U3875 (N_3875,In_214,In_1129);
nor U3876 (N_3876,In_449,In_717);
nor U3877 (N_3877,In_1407,In_1459);
or U3878 (N_3878,In_908,In_563);
nor U3879 (N_3879,In_140,In_532);
xor U3880 (N_3880,In_398,In_1386);
xor U3881 (N_3881,In_56,In_1291);
or U3882 (N_3882,In_142,In_1191);
nand U3883 (N_3883,In_329,In_231);
nand U3884 (N_3884,In_1288,In_1418);
and U3885 (N_3885,In_1196,In_1228);
and U3886 (N_3886,In_1222,In_714);
or U3887 (N_3887,In_491,In_821);
xor U3888 (N_3888,In_1087,In_1084);
and U3889 (N_3889,In_160,In_763);
xor U3890 (N_3890,In_1207,In_465);
or U3891 (N_3891,In_406,In_197);
nand U3892 (N_3892,In_325,In_472);
nor U3893 (N_3893,In_1198,In_1173);
nand U3894 (N_3894,In_523,In_411);
xor U3895 (N_3895,In_178,In_36);
and U3896 (N_3896,In_69,In_689);
xor U3897 (N_3897,In_1200,In_402);
nor U3898 (N_3898,In_1465,In_580);
nand U3899 (N_3899,In_7,In_1407);
xnor U3900 (N_3900,In_1191,In_80);
nand U3901 (N_3901,In_846,In_502);
nor U3902 (N_3902,In_1344,In_1212);
and U3903 (N_3903,In_900,In_41);
or U3904 (N_3904,In_1185,In_147);
or U3905 (N_3905,In_703,In_1441);
or U3906 (N_3906,In_756,In_229);
xor U3907 (N_3907,In_1226,In_878);
nand U3908 (N_3908,In_1178,In_170);
xor U3909 (N_3909,In_359,In_602);
and U3910 (N_3910,In_15,In_82);
xnor U3911 (N_3911,In_1488,In_68);
nand U3912 (N_3912,In_1418,In_824);
xnor U3913 (N_3913,In_911,In_670);
nand U3914 (N_3914,In_1134,In_936);
or U3915 (N_3915,In_562,In_406);
xnor U3916 (N_3916,In_1044,In_170);
and U3917 (N_3917,In_296,In_316);
nand U3918 (N_3918,In_580,In_870);
xor U3919 (N_3919,In_4,In_1492);
or U3920 (N_3920,In_341,In_982);
nor U3921 (N_3921,In_604,In_619);
nor U3922 (N_3922,In_755,In_545);
nor U3923 (N_3923,In_553,In_287);
or U3924 (N_3924,In_913,In_1095);
or U3925 (N_3925,In_1060,In_1238);
nand U3926 (N_3926,In_1362,In_829);
and U3927 (N_3927,In_315,In_57);
or U3928 (N_3928,In_892,In_438);
nor U3929 (N_3929,In_121,In_34);
nand U3930 (N_3930,In_700,In_1188);
and U3931 (N_3931,In_483,In_713);
nand U3932 (N_3932,In_734,In_67);
and U3933 (N_3933,In_188,In_611);
nor U3934 (N_3934,In_237,In_875);
xor U3935 (N_3935,In_972,In_1338);
nand U3936 (N_3936,In_494,In_1285);
nor U3937 (N_3937,In_1150,In_1306);
nor U3938 (N_3938,In_7,In_225);
xor U3939 (N_3939,In_867,In_1035);
nor U3940 (N_3940,In_1312,In_398);
and U3941 (N_3941,In_803,In_289);
nand U3942 (N_3942,In_1084,In_1207);
nand U3943 (N_3943,In_1350,In_1181);
and U3944 (N_3944,In_984,In_172);
nand U3945 (N_3945,In_702,In_522);
nand U3946 (N_3946,In_364,In_1056);
or U3947 (N_3947,In_1477,In_113);
or U3948 (N_3948,In_112,In_784);
nor U3949 (N_3949,In_634,In_166);
and U3950 (N_3950,In_850,In_1355);
and U3951 (N_3951,In_494,In_479);
xor U3952 (N_3952,In_888,In_200);
xnor U3953 (N_3953,In_1460,In_55);
and U3954 (N_3954,In_1121,In_888);
nor U3955 (N_3955,In_1286,In_1472);
and U3956 (N_3956,In_438,In_655);
and U3957 (N_3957,In_71,In_765);
xor U3958 (N_3958,In_1456,In_800);
and U3959 (N_3959,In_425,In_937);
or U3960 (N_3960,In_347,In_368);
nor U3961 (N_3961,In_1064,In_610);
xnor U3962 (N_3962,In_394,In_420);
and U3963 (N_3963,In_727,In_741);
or U3964 (N_3964,In_843,In_558);
xor U3965 (N_3965,In_343,In_361);
xnor U3966 (N_3966,In_870,In_1471);
nor U3967 (N_3967,In_6,In_149);
or U3968 (N_3968,In_370,In_1087);
xnor U3969 (N_3969,In_126,In_921);
xor U3970 (N_3970,In_163,In_856);
xnor U3971 (N_3971,In_1261,In_701);
nor U3972 (N_3972,In_256,In_1121);
nor U3973 (N_3973,In_633,In_42);
nand U3974 (N_3974,In_1267,In_1147);
nand U3975 (N_3975,In_617,In_57);
xor U3976 (N_3976,In_196,In_234);
xor U3977 (N_3977,In_421,In_1277);
and U3978 (N_3978,In_327,In_471);
nor U3979 (N_3979,In_937,In_1245);
or U3980 (N_3980,In_568,In_141);
xor U3981 (N_3981,In_1340,In_933);
or U3982 (N_3982,In_1082,In_814);
xor U3983 (N_3983,In_1328,In_1022);
xnor U3984 (N_3984,In_152,In_507);
nor U3985 (N_3985,In_813,In_692);
and U3986 (N_3986,In_73,In_650);
and U3987 (N_3987,In_538,In_657);
nand U3988 (N_3988,In_1027,In_761);
nand U3989 (N_3989,In_916,In_829);
and U3990 (N_3990,In_717,In_3);
or U3991 (N_3991,In_775,In_948);
nand U3992 (N_3992,In_1433,In_624);
and U3993 (N_3993,In_563,In_429);
nor U3994 (N_3994,In_1279,In_457);
nor U3995 (N_3995,In_1231,In_248);
nand U3996 (N_3996,In_16,In_318);
nor U3997 (N_3997,In_1475,In_401);
and U3998 (N_3998,In_323,In_1169);
nand U3999 (N_3999,In_1464,In_865);
nand U4000 (N_4000,In_649,In_457);
xnor U4001 (N_4001,In_739,In_421);
or U4002 (N_4002,In_810,In_1296);
xnor U4003 (N_4003,In_1264,In_324);
nand U4004 (N_4004,In_1431,In_1280);
and U4005 (N_4005,In_1170,In_1477);
xnor U4006 (N_4006,In_1248,In_861);
and U4007 (N_4007,In_611,In_1394);
xnor U4008 (N_4008,In_1189,In_1374);
nand U4009 (N_4009,In_18,In_638);
xor U4010 (N_4010,In_1299,In_739);
and U4011 (N_4011,In_845,In_803);
nor U4012 (N_4012,In_1349,In_170);
or U4013 (N_4013,In_102,In_218);
xor U4014 (N_4014,In_650,In_1252);
or U4015 (N_4015,In_152,In_199);
xor U4016 (N_4016,In_1159,In_1283);
or U4017 (N_4017,In_460,In_421);
nor U4018 (N_4018,In_680,In_667);
xnor U4019 (N_4019,In_342,In_84);
nor U4020 (N_4020,In_1185,In_98);
or U4021 (N_4021,In_1435,In_1145);
xnor U4022 (N_4022,In_260,In_1311);
or U4023 (N_4023,In_1028,In_1363);
nor U4024 (N_4024,In_1490,In_553);
nand U4025 (N_4025,In_1029,In_853);
xor U4026 (N_4026,In_1463,In_1240);
nor U4027 (N_4027,In_564,In_210);
nor U4028 (N_4028,In_1218,In_1276);
and U4029 (N_4029,In_682,In_1322);
nand U4030 (N_4030,In_96,In_1319);
or U4031 (N_4031,In_767,In_1176);
and U4032 (N_4032,In_1179,In_374);
xor U4033 (N_4033,In_8,In_1229);
nor U4034 (N_4034,In_508,In_71);
xor U4035 (N_4035,In_1275,In_522);
and U4036 (N_4036,In_1252,In_263);
nand U4037 (N_4037,In_845,In_408);
nor U4038 (N_4038,In_828,In_122);
xor U4039 (N_4039,In_1247,In_993);
xnor U4040 (N_4040,In_722,In_103);
or U4041 (N_4041,In_1254,In_1164);
nand U4042 (N_4042,In_1292,In_1493);
nand U4043 (N_4043,In_533,In_1246);
xor U4044 (N_4044,In_551,In_1414);
xnor U4045 (N_4045,In_1494,In_936);
nor U4046 (N_4046,In_38,In_505);
and U4047 (N_4047,In_1298,In_673);
xnor U4048 (N_4048,In_1133,In_1385);
xor U4049 (N_4049,In_412,In_358);
and U4050 (N_4050,In_1364,In_542);
xor U4051 (N_4051,In_1394,In_617);
xor U4052 (N_4052,In_295,In_625);
and U4053 (N_4053,In_1470,In_982);
or U4054 (N_4054,In_438,In_1116);
nor U4055 (N_4055,In_861,In_1419);
nor U4056 (N_4056,In_185,In_950);
and U4057 (N_4057,In_990,In_50);
xor U4058 (N_4058,In_96,In_7);
nor U4059 (N_4059,In_1382,In_450);
nand U4060 (N_4060,In_1197,In_1429);
or U4061 (N_4061,In_1169,In_284);
nor U4062 (N_4062,In_761,In_1071);
or U4063 (N_4063,In_1087,In_1332);
nand U4064 (N_4064,In_419,In_1306);
nand U4065 (N_4065,In_1398,In_887);
nor U4066 (N_4066,In_485,In_910);
and U4067 (N_4067,In_1000,In_390);
xnor U4068 (N_4068,In_375,In_999);
or U4069 (N_4069,In_1229,In_194);
nand U4070 (N_4070,In_365,In_308);
or U4071 (N_4071,In_1028,In_839);
and U4072 (N_4072,In_295,In_736);
and U4073 (N_4073,In_1242,In_1122);
nor U4074 (N_4074,In_1099,In_940);
or U4075 (N_4075,In_339,In_734);
nor U4076 (N_4076,In_1179,In_972);
and U4077 (N_4077,In_1468,In_517);
or U4078 (N_4078,In_462,In_1078);
and U4079 (N_4079,In_611,In_772);
nand U4080 (N_4080,In_780,In_756);
and U4081 (N_4081,In_1053,In_243);
and U4082 (N_4082,In_1029,In_615);
or U4083 (N_4083,In_703,In_236);
and U4084 (N_4084,In_1209,In_1420);
xnor U4085 (N_4085,In_292,In_183);
nor U4086 (N_4086,In_1048,In_272);
xor U4087 (N_4087,In_1056,In_1488);
nor U4088 (N_4088,In_881,In_1371);
or U4089 (N_4089,In_24,In_496);
nand U4090 (N_4090,In_452,In_303);
nand U4091 (N_4091,In_559,In_457);
or U4092 (N_4092,In_182,In_1013);
nor U4093 (N_4093,In_763,In_1153);
xor U4094 (N_4094,In_334,In_922);
nor U4095 (N_4095,In_1181,In_61);
nor U4096 (N_4096,In_555,In_1318);
or U4097 (N_4097,In_633,In_1428);
nor U4098 (N_4098,In_1325,In_624);
and U4099 (N_4099,In_802,In_1468);
xnor U4100 (N_4100,In_82,In_903);
or U4101 (N_4101,In_1332,In_1033);
and U4102 (N_4102,In_75,In_972);
nand U4103 (N_4103,In_554,In_989);
or U4104 (N_4104,In_710,In_760);
nand U4105 (N_4105,In_1207,In_577);
nor U4106 (N_4106,In_453,In_53);
or U4107 (N_4107,In_336,In_693);
nor U4108 (N_4108,In_1004,In_98);
xor U4109 (N_4109,In_1331,In_1255);
xnor U4110 (N_4110,In_711,In_444);
nor U4111 (N_4111,In_481,In_535);
nor U4112 (N_4112,In_1423,In_575);
nand U4113 (N_4113,In_1084,In_243);
nor U4114 (N_4114,In_1149,In_1479);
and U4115 (N_4115,In_1102,In_299);
nand U4116 (N_4116,In_1436,In_256);
nor U4117 (N_4117,In_54,In_735);
nand U4118 (N_4118,In_742,In_980);
nor U4119 (N_4119,In_28,In_851);
and U4120 (N_4120,In_1479,In_860);
nor U4121 (N_4121,In_13,In_957);
nor U4122 (N_4122,In_188,In_1472);
xor U4123 (N_4123,In_767,In_415);
nor U4124 (N_4124,In_1225,In_1088);
xor U4125 (N_4125,In_301,In_1352);
or U4126 (N_4126,In_385,In_844);
or U4127 (N_4127,In_907,In_1205);
nand U4128 (N_4128,In_228,In_1259);
nand U4129 (N_4129,In_811,In_646);
nand U4130 (N_4130,In_480,In_1245);
and U4131 (N_4131,In_1323,In_533);
and U4132 (N_4132,In_400,In_562);
xor U4133 (N_4133,In_107,In_799);
nand U4134 (N_4134,In_1213,In_1463);
xnor U4135 (N_4135,In_104,In_449);
nor U4136 (N_4136,In_958,In_546);
or U4137 (N_4137,In_137,In_351);
and U4138 (N_4138,In_349,In_1218);
nand U4139 (N_4139,In_1161,In_1373);
or U4140 (N_4140,In_363,In_1386);
nand U4141 (N_4141,In_1147,In_911);
nand U4142 (N_4142,In_963,In_586);
or U4143 (N_4143,In_720,In_853);
nand U4144 (N_4144,In_1375,In_232);
nand U4145 (N_4145,In_782,In_986);
xor U4146 (N_4146,In_1320,In_1247);
nand U4147 (N_4147,In_394,In_70);
and U4148 (N_4148,In_898,In_1315);
nand U4149 (N_4149,In_267,In_922);
and U4150 (N_4150,In_726,In_354);
or U4151 (N_4151,In_523,In_715);
nor U4152 (N_4152,In_41,In_132);
and U4153 (N_4153,In_1289,In_166);
xnor U4154 (N_4154,In_298,In_419);
xor U4155 (N_4155,In_563,In_555);
or U4156 (N_4156,In_1258,In_399);
and U4157 (N_4157,In_628,In_913);
nand U4158 (N_4158,In_303,In_237);
nor U4159 (N_4159,In_177,In_1490);
nor U4160 (N_4160,In_41,In_1373);
or U4161 (N_4161,In_1310,In_1323);
nor U4162 (N_4162,In_100,In_880);
or U4163 (N_4163,In_241,In_722);
xnor U4164 (N_4164,In_1452,In_386);
nor U4165 (N_4165,In_341,In_575);
nand U4166 (N_4166,In_444,In_1283);
nor U4167 (N_4167,In_173,In_1132);
xnor U4168 (N_4168,In_1491,In_540);
nand U4169 (N_4169,In_1158,In_62);
and U4170 (N_4170,In_895,In_1263);
xnor U4171 (N_4171,In_1361,In_1310);
or U4172 (N_4172,In_902,In_1039);
nor U4173 (N_4173,In_1260,In_32);
or U4174 (N_4174,In_170,In_1358);
nand U4175 (N_4175,In_100,In_787);
nor U4176 (N_4176,In_496,In_614);
xnor U4177 (N_4177,In_1265,In_150);
or U4178 (N_4178,In_985,In_547);
nand U4179 (N_4179,In_123,In_35);
and U4180 (N_4180,In_872,In_166);
nand U4181 (N_4181,In_1068,In_1354);
or U4182 (N_4182,In_911,In_659);
or U4183 (N_4183,In_918,In_813);
nor U4184 (N_4184,In_944,In_805);
or U4185 (N_4185,In_1121,In_302);
nand U4186 (N_4186,In_9,In_139);
nor U4187 (N_4187,In_488,In_462);
and U4188 (N_4188,In_797,In_724);
and U4189 (N_4189,In_1040,In_402);
xnor U4190 (N_4190,In_1446,In_940);
or U4191 (N_4191,In_282,In_1402);
xor U4192 (N_4192,In_1484,In_1029);
nor U4193 (N_4193,In_1414,In_801);
nand U4194 (N_4194,In_660,In_382);
nor U4195 (N_4195,In_868,In_613);
nor U4196 (N_4196,In_289,In_1003);
and U4197 (N_4197,In_110,In_1111);
nand U4198 (N_4198,In_1277,In_619);
xnor U4199 (N_4199,In_1099,In_1153);
nand U4200 (N_4200,In_743,In_990);
nand U4201 (N_4201,In_707,In_114);
nand U4202 (N_4202,In_199,In_1053);
nand U4203 (N_4203,In_1425,In_659);
nor U4204 (N_4204,In_133,In_1208);
nor U4205 (N_4205,In_1129,In_819);
and U4206 (N_4206,In_1386,In_20);
nand U4207 (N_4207,In_1460,In_818);
xnor U4208 (N_4208,In_536,In_712);
or U4209 (N_4209,In_67,In_1144);
nor U4210 (N_4210,In_646,In_546);
xnor U4211 (N_4211,In_402,In_1413);
and U4212 (N_4212,In_905,In_957);
or U4213 (N_4213,In_172,In_865);
nor U4214 (N_4214,In_477,In_618);
nand U4215 (N_4215,In_983,In_1469);
nor U4216 (N_4216,In_81,In_1178);
nand U4217 (N_4217,In_676,In_91);
nor U4218 (N_4218,In_514,In_673);
nor U4219 (N_4219,In_1339,In_1315);
or U4220 (N_4220,In_439,In_977);
nor U4221 (N_4221,In_993,In_1062);
or U4222 (N_4222,In_1023,In_692);
nand U4223 (N_4223,In_221,In_215);
nand U4224 (N_4224,In_1447,In_1342);
or U4225 (N_4225,In_391,In_379);
or U4226 (N_4226,In_1407,In_735);
xor U4227 (N_4227,In_522,In_98);
xnor U4228 (N_4228,In_696,In_879);
nor U4229 (N_4229,In_996,In_807);
xnor U4230 (N_4230,In_1446,In_41);
or U4231 (N_4231,In_268,In_181);
or U4232 (N_4232,In_1,In_472);
nor U4233 (N_4233,In_1493,In_597);
nand U4234 (N_4234,In_1434,In_1297);
or U4235 (N_4235,In_498,In_1245);
nand U4236 (N_4236,In_651,In_663);
and U4237 (N_4237,In_1386,In_245);
nor U4238 (N_4238,In_1176,In_49);
or U4239 (N_4239,In_459,In_585);
nor U4240 (N_4240,In_116,In_640);
nand U4241 (N_4241,In_923,In_1033);
or U4242 (N_4242,In_1441,In_338);
nand U4243 (N_4243,In_318,In_342);
nand U4244 (N_4244,In_1492,In_968);
nor U4245 (N_4245,In_1495,In_453);
and U4246 (N_4246,In_1004,In_1303);
xor U4247 (N_4247,In_654,In_1177);
xor U4248 (N_4248,In_315,In_972);
nand U4249 (N_4249,In_8,In_1070);
nor U4250 (N_4250,In_1307,In_615);
and U4251 (N_4251,In_856,In_793);
xor U4252 (N_4252,In_972,In_1377);
nor U4253 (N_4253,In_554,In_355);
and U4254 (N_4254,In_1270,In_745);
and U4255 (N_4255,In_365,In_446);
nor U4256 (N_4256,In_1355,In_451);
nand U4257 (N_4257,In_1153,In_317);
nor U4258 (N_4258,In_1333,In_1205);
nand U4259 (N_4259,In_144,In_705);
nor U4260 (N_4260,In_1203,In_328);
nor U4261 (N_4261,In_653,In_621);
nor U4262 (N_4262,In_154,In_991);
xnor U4263 (N_4263,In_1276,In_1341);
or U4264 (N_4264,In_1085,In_594);
and U4265 (N_4265,In_23,In_767);
nor U4266 (N_4266,In_1454,In_1070);
nor U4267 (N_4267,In_519,In_185);
nand U4268 (N_4268,In_709,In_1327);
nor U4269 (N_4269,In_200,In_1452);
xnor U4270 (N_4270,In_503,In_661);
nand U4271 (N_4271,In_993,In_422);
and U4272 (N_4272,In_807,In_417);
nand U4273 (N_4273,In_989,In_973);
nand U4274 (N_4274,In_435,In_571);
and U4275 (N_4275,In_708,In_1064);
xor U4276 (N_4276,In_830,In_426);
nand U4277 (N_4277,In_1342,In_276);
and U4278 (N_4278,In_972,In_321);
or U4279 (N_4279,In_582,In_529);
and U4280 (N_4280,In_850,In_333);
nor U4281 (N_4281,In_554,In_526);
and U4282 (N_4282,In_447,In_1011);
or U4283 (N_4283,In_247,In_920);
xor U4284 (N_4284,In_888,In_897);
nand U4285 (N_4285,In_423,In_255);
and U4286 (N_4286,In_427,In_1300);
nand U4287 (N_4287,In_26,In_1468);
or U4288 (N_4288,In_25,In_279);
and U4289 (N_4289,In_930,In_1264);
and U4290 (N_4290,In_841,In_279);
xor U4291 (N_4291,In_769,In_889);
or U4292 (N_4292,In_84,In_469);
nand U4293 (N_4293,In_332,In_1189);
nand U4294 (N_4294,In_140,In_801);
or U4295 (N_4295,In_1339,In_486);
or U4296 (N_4296,In_1080,In_939);
nand U4297 (N_4297,In_940,In_989);
or U4298 (N_4298,In_71,In_353);
nand U4299 (N_4299,In_1419,In_276);
or U4300 (N_4300,In_1197,In_1302);
nor U4301 (N_4301,In_318,In_426);
or U4302 (N_4302,In_1230,In_370);
nand U4303 (N_4303,In_552,In_882);
xnor U4304 (N_4304,In_558,In_889);
nand U4305 (N_4305,In_1469,In_536);
and U4306 (N_4306,In_877,In_644);
or U4307 (N_4307,In_353,In_657);
xnor U4308 (N_4308,In_902,In_836);
or U4309 (N_4309,In_340,In_880);
or U4310 (N_4310,In_143,In_584);
nand U4311 (N_4311,In_231,In_1051);
or U4312 (N_4312,In_244,In_1048);
xor U4313 (N_4313,In_401,In_1066);
and U4314 (N_4314,In_570,In_434);
nor U4315 (N_4315,In_263,In_910);
and U4316 (N_4316,In_481,In_1205);
xor U4317 (N_4317,In_611,In_1405);
nor U4318 (N_4318,In_904,In_107);
and U4319 (N_4319,In_850,In_1269);
nand U4320 (N_4320,In_630,In_376);
nor U4321 (N_4321,In_635,In_981);
or U4322 (N_4322,In_649,In_1135);
xnor U4323 (N_4323,In_952,In_728);
or U4324 (N_4324,In_553,In_1278);
or U4325 (N_4325,In_810,In_545);
nor U4326 (N_4326,In_1000,In_535);
or U4327 (N_4327,In_1453,In_1260);
xor U4328 (N_4328,In_277,In_219);
nand U4329 (N_4329,In_1026,In_698);
nor U4330 (N_4330,In_409,In_844);
nor U4331 (N_4331,In_1016,In_877);
nor U4332 (N_4332,In_982,In_1101);
nor U4333 (N_4333,In_136,In_1333);
and U4334 (N_4334,In_1155,In_539);
or U4335 (N_4335,In_1027,In_284);
nor U4336 (N_4336,In_617,In_51);
nand U4337 (N_4337,In_336,In_1299);
and U4338 (N_4338,In_1393,In_1366);
xnor U4339 (N_4339,In_214,In_357);
nor U4340 (N_4340,In_385,In_1456);
xnor U4341 (N_4341,In_1365,In_239);
nor U4342 (N_4342,In_1401,In_644);
nor U4343 (N_4343,In_1052,In_657);
nand U4344 (N_4344,In_1328,In_1165);
and U4345 (N_4345,In_952,In_1428);
and U4346 (N_4346,In_982,In_868);
xor U4347 (N_4347,In_798,In_606);
nor U4348 (N_4348,In_1361,In_771);
or U4349 (N_4349,In_1188,In_943);
xor U4350 (N_4350,In_78,In_771);
or U4351 (N_4351,In_548,In_409);
xnor U4352 (N_4352,In_494,In_1169);
or U4353 (N_4353,In_699,In_101);
nand U4354 (N_4354,In_947,In_787);
and U4355 (N_4355,In_1380,In_1308);
and U4356 (N_4356,In_983,In_931);
nor U4357 (N_4357,In_777,In_757);
xnor U4358 (N_4358,In_479,In_1210);
nand U4359 (N_4359,In_272,In_598);
nor U4360 (N_4360,In_1300,In_1443);
and U4361 (N_4361,In_1379,In_1008);
nor U4362 (N_4362,In_741,In_954);
xor U4363 (N_4363,In_1223,In_469);
nand U4364 (N_4364,In_538,In_59);
and U4365 (N_4365,In_1144,In_862);
nor U4366 (N_4366,In_994,In_623);
and U4367 (N_4367,In_1454,In_536);
xnor U4368 (N_4368,In_460,In_1463);
or U4369 (N_4369,In_404,In_894);
and U4370 (N_4370,In_609,In_1401);
xor U4371 (N_4371,In_379,In_1143);
nor U4372 (N_4372,In_1175,In_772);
nor U4373 (N_4373,In_150,In_976);
nor U4374 (N_4374,In_839,In_1455);
nand U4375 (N_4375,In_1304,In_882);
xor U4376 (N_4376,In_1048,In_1347);
or U4377 (N_4377,In_1051,In_903);
nor U4378 (N_4378,In_1107,In_67);
and U4379 (N_4379,In_1206,In_930);
nor U4380 (N_4380,In_221,In_295);
or U4381 (N_4381,In_842,In_345);
nor U4382 (N_4382,In_141,In_1038);
nor U4383 (N_4383,In_1463,In_1144);
nand U4384 (N_4384,In_152,In_1115);
and U4385 (N_4385,In_324,In_391);
xnor U4386 (N_4386,In_1112,In_1012);
xnor U4387 (N_4387,In_815,In_452);
or U4388 (N_4388,In_692,In_1466);
and U4389 (N_4389,In_182,In_586);
nand U4390 (N_4390,In_1024,In_753);
xnor U4391 (N_4391,In_1388,In_1341);
xor U4392 (N_4392,In_515,In_514);
nor U4393 (N_4393,In_909,In_1457);
nand U4394 (N_4394,In_929,In_1062);
xnor U4395 (N_4395,In_799,In_239);
nand U4396 (N_4396,In_1024,In_186);
and U4397 (N_4397,In_73,In_927);
xnor U4398 (N_4398,In_410,In_1231);
and U4399 (N_4399,In_1258,In_721);
and U4400 (N_4400,In_1436,In_1387);
xor U4401 (N_4401,In_1090,In_907);
or U4402 (N_4402,In_1199,In_1455);
nor U4403 (N_4403,In_693,In_1437);
xor U4404 (N_4404,In_1351,In_1049);
or U4405 (N_4405,In_1288,In_818);
nor U4406 (N_4406,In_990,In_138);
and U4407 (N_4407,In_626,In_711);
nor U4408 (N_4408,In_318,In_1058);
or U4409 (N_4409,In_1205,In_981);
nand U4410 (N_4410,In_1402,In_729);
nand U4411 (N_4411,In_910,In_249);
nand U4412 (N_4412,In_886,In_904);
or U4413 (N_4413,In_1451,In_896);
and U4414 (N_4414,In_170,In_377);
and U4415 (N_4415,In_151,In_1391);
xnor U4416 (N_4416,In_1434,In_552);
xor U4417 (N_4417,In_933,In_60);
nand U4418 (N_4418,In_645,In_541);
nor U4419 (N_4419,In_1473,In_703);
or U4420 (N_4420,In_285,In_229);
nor U4421 (N_4421,In_402,In_63);
nor U4422 (N_4422,In_1275,In_1273);
nor U4423 (N_4423,In_413,In_962);
xor U4424 (N_4424,In_586,In_841);
and U4425 (N_4425,In_1467,In_466);
or U4426 (N_4426,In_498,In_56);
xnor U4427 (N_4427,In_990,In_1149);
nor U4428 (N_4428,In_897,In_1474);
nand U4429 (N_4429,In_998,In_1234);
nand U4430 (N_4430,In_1007,In_947);
or U4431 (N_4431,In_749,In_134);
or U4432 (N_4432,In_745,In_952);
nand U4433 (N_4433,In_1118,In_1112);
xnor U4434 (N_4434,In_329,In_1064);
and U4435 (N_4435,In_1459,In_830);
nor U4436 (N_4436,In_312,In_9);
nor U4437 (N_4437,In_495,In_389);
and U4438 (N_4438,In_263,In_653);
or U4439 (N_4439,In_1186,In_182);
nor U4440 (N_4440,In_1076,In_610);
nor U4441 (N_4441,In_928,In_1134);
and U4442 (N_4442,In_1395,In_1015);
xnor U4443 (N_4443,In_211,In_387);
xor U4444 (N_4444,In_343,In_179);
nor U4445 (N_4445,In_1443,In_1202);
or U4446 (N_4446,In_756,In_171);
and U4447 (N_4447,In_900,In_80);
xnor U4448 (N_4448,In_1157,In_665);
or U4449 (N_4449,In_925,In_837);
or U4450 (N_4450,In_1109,In_22);
nand U4451 (N_4451,In_197,In_95);
and U4452 (N_4452,In_684,In_715);
and U4453 (N_4453,In_1458,In_195);
or U4454 (N_4454,In_481,In_929);
nand U4455 (N_4455,In_1055,In_431);
nor U4456 (N_4456,In_927,In_1480);
or U4457 (N_4457,In_711,In_1196);
nand U4458 (N_4458,In_512,In_723);
or U4459 (N_4459,In_201,In_960);
xor U4460 (N_4460,In_742,In_474);
xor U4461 (N_4461,In_807,In_126);
nor U4462 (N_4462,In_582,In_931);
nand U4463 (N_4463,In_1488,In_642);
nand U4464 (N_4464,In_1352,In_1058);
nor U4465 (N_4465,In_218,In_235);
nand U4466 (N_4466,In_78,In_1162);
nor U4467 (N_4467,In_80,In_735);
nand U4468 (N_4468,In_944,In_650);
and U4469 (N_4469,In_301,In_101);
xnor U4470 (N_4470,In_1301,In_422);
nor U4471 (N_4471,In_973,In_202);
nand U4472 (N_4472,In_79,In_1185);
or U4473 (N_4473,In_472,In_627);
nand U4474 (N_4474,In_124,In_131);
and U4475 (N_4475,In_236,In_839);
or U4476 (N_4476,In_1382,In_1348);
xnor U4477 (N_4477,In_1301,In_1438);
or U4478 (N_4478,In_872,In_116);
nor U4479 (N_4479,In_317,In_504);
nand U4480 (N_4480,In_1129,In_552);
nand U4481 (N_4481,In_990,In_1143);
xnor U4482 (N_4482,In_1023,In_423);
nor U4483 (N_4483,In_503,In_619);
xnor U4484 (N_4484,In_1027,In_260);
xor U4485 (N_4485,In_690,In_190);
nand U4486 (N_4486,In_495,In_1125);
and U4487 (N_4487,In_1322,In_1476);
nor U4488 (N_4488,In_177,In_227);
nor U4489 (N_4489,In_341,In_236);
nor U4490 (N_4490,In_344,In_387);
xor U4491 (N_4491,In_508,In_826);
or U4492 (N_4492,In_981,In_986);
or U4493 (N_4493,In_528,In_1060);
xnor U4494 (N_4494,In_77,In_539);
and U4495 (N_4495,In_1211,In_688);
nand U4496 (N_4496,In_215,In_234);
and U4497 (N_4497,In_903,In_90);
xor U4498 (N_4498,In_1406,In_208);
nand U4499 (N_4499,In_103,In_283);
nor U4500 (N_4500,In_1412,In_1135);
xor U4501 (N_4501,In_1302,In_1281);
xnor U4502 (N_4502,In_687,In_1114);
or U4503 (N_4503,In_1108,In_887);
and U4504 (N_4504,In_280,In_7);
nand U4505 (N_4505,In_1194,In_871);
and U4506 (N_4506,In_1217,In_326);
nand U4507 (N_4507,In_71,In_1120);
nand U4508 (N_4508,In_1299,In_218);
nor U4509 (N_4509,In_601,In_981);
nand U4510 (N_4510,In_336,In_533);
nand U4511 (N_4511,In_64,In_559);
xor U4512 (N_4512,In_1362,In_1221);
and U4513 (N_4513,In_176,In_859);
nand U4514 (N_4514,In_1031,In_662);
or U4515 (N_4515,In_586,In_448);
and U4516 (N_4516,In_465,In_647);
xnor U4517 (N_4517,In_1431,In_61);
nand U4518 (N_4518,In_1308,In_19);
nor U4519 (N_4519,In_419,In_410);
nand U4520 (N_4520,In_142,In_810);
or U4521 (N_4521,In_291,In_267);
nor U4522 (N_4522,In_729,In_894);
and U4523 (N_4523,In_235,In_333);
and U4524 (N_4524,In_1372,In_928);
and U4525 (N_4525,In_999,In_376);
xnor U4526 (N_4526,In_1464,In_397);
xnor U4527 (N_4527,In_236,In_124);
nand U4528 (N_4528,In_410,In_607);
xnor U4529 (N_4529,In_649,In_495);
xor U4530 (N_4530,In_1050,In_264);
nor U4531 (N_4531,In_397,In_730);
nor U4532 (N_4532,In_453,In_1115);
or U4533 (N_4533,In_1256,In_475);
nand U4534 (N_4534,In_151,In_1022);
or U4535 (N_4535,In_1032,In_736);
and U4536 (N_4536,In_917,In_366);
and U4537 (N_4537,In_188,In_421);
or U4538 (N_4538,In_500,In_286);
nand U4539 (N_4539,In_228,In_1326);
and U4540 (N_4540,In_87,In_834);
xnor U4541 (N_4541,In_373,In_1055);
nor U4542 (N_4542,In_993,In_328);
nand U4543 (N_4543,In_1106,In_1100);
and U4544 (N_4544,In_1386,In_1389);
nor U4545 (N_4545,In_1439,In_231);
and U4546 (N_4546,In_1045,In_1125);
and U4547 (N_4547,In_132,In_270);
xor U4548 (N_4548,In_1493,In_802);
and U4549 (N_4549,In_1264,In_97);
or U4550 (N_4550,In_724,In_1302);
or U4551 (N_4551,In_115,In_835);
nor U4552 (N_4552,In_1281,In_820);
xnor U4553 (N_4553,In_215,In_714);
or U4554 (N_4554,In_1453,In_964);
and U4555 (N_4555,In_1095,In_274);
and U4556 (N_4556,In_751,In_915);
nand U4557 (N_4557,In_608,In_693);
or U4558 (N_4558,In_411,In_768);
and U4559 (N_4559,In_1305,In_1300);
nand U4560 (N_4560,In_995,In_690);
nor U4561 (N_4561,In_134,In_268);
and U4562 (N_4562,In_645,In_1484);
or U4563 (N_4563,In_1058,In_528);
xnor U4564 (N_4564,In_691,In_1349);
nor U4565 (N_4565,In_790,In_1053);
or U4566 (N_4566,In_1115,In_760);
and U4567 (N_4567,In_47,In_1320);
xnor U4568 (N_4568,In_1073,In_1197);
xor U4569 (N_4569,In_391,In_1064);
nand U4570 (N_4570,In_383,In_1015);
xor U4571 (N_4571,In_1476,In_1290);
xor U4572 (N_4572,In_1068,In_623);
or U4573 (N_4573,In_1016,In_968);
xnor U4574 (N_4574,In_637,In_215);
xnor U4575 (N_4575,In_1290,In_573);
xnor U4576 (N_4576,In_1129,In_428);
and U4577 (N_4577,In_1272,In_1096);
nor U4578 (N_4578,In_362,In_482);
xor U4579 (N_4579,In_1264,In_1154);
and U4580 (N_4580,In_1090,In_1077);
nor U4581 (N_4581,In_415,In_1376);
or U4582 (N_4582,In_389,In_853);
or U4583 (N_4583,In_177,In_454);
or U4584 (N_4584,In_1449,In_307);
nand U4585 (N_4585,In_1190,In_1231);
and U4586 (N_4586,In_652,In_30);
nor U4587 (N_4587,In_604,In_11);
or U4588 (N_4588,In_1434,In_1335);
nor U4589 (N_4589,In_757,In_74);
or U4590 (N_4590,In_974,In_797);
xnor U4591 (N_4591,In_238,In_1101);
nor U4592 (N_4592,In_747,In_482);
nor U4593 (N_4593,In_868,In_1062);
nor U4594 (N_4594,In_1145,In_279);
nand U4595 (N_4595,In_333,In_120);
nand U4596 (N_4596,In_793,In_654);
nor U4597 (N_4597,In_1263,In_1492);
nand U4598 (N_4598,In_873,In_268);
nor U4599 (N_4599,In_481,In_519);
nand U4600 (N_4600,In_1081,In_1201);
and U4601 (N_4601,In_861,In_1019);
nand U4602 (N_4602,In_622,In_500);
and U4603 (N_4603,In_134,In_768);
nor U4604 (N_4604,In_1082,In_1217);
nor U4605 (N_4605,In_1395,In_428);
and U4606 (N_4606,In_223,In_187);
nand U4607 (N_4607,In_1150,In_1422);
and U4608 (N_4608,In_1225,In_404);
or U4609 (N_4609,In_173,In_1046);
nor U4610 (N_4610,In_439,In_1185);
xnor U4611 (N_4611,In_529,In_834);
or U4612 (N_4612,In_895,In_867);
and U4613 (N_4613,In_1132,In_1374);
or U4614 (N_4614,In_321,In_1499);
nor U4615 (N_4615,In_1045,In_964);
nor U4616 (N_4616,In_1133,In_872);
or U4617 (N_4617,In_1130,In_89);
nor U4618 (N_4618,In_1248,In_701);
nand U4619 (N_4619,In_723,In_146);
or U4620 (N_4620,In_345,In_1302);
and U4621 (N_4621,In_465,In_1055);
xnor U4622 (N_4622,In_462,In_672);
and U4623 (N_4623,In_1308,In_276);
and U4624 (N_4624,In_846,In_338);
and U4625 (N_4625,In_692,In_178);
or U4626 (N_4626,In_694,In_1321);
nand U4627 (N_4627,In_454,In_1246);
and U4628 (N_4628,In_48,In_819);
or U4629 (N_4629,In_1006,In_437);
and U4630 (N_4630,In_1377,In_828);
and U4631 (N_4631,In_132,In_1074);
xnor U4632 (N_4632,In_1171,In_603);
nor U4633 (N_4633,In_684,In_38);
nand U4634 (N_4634,In_503,In_1419);
xor U4635 (N_4635,In_378,In_808);
or U4636 (N_4636,In_247,In_1353);
nor U4637 (N_4637,In_232,In_1095);
or U4638 (N_4638,In_1227,In_226);
xor U4639 (N_4639,In_292,In_1217);
nand U4640 (N_4640,In_0,In_1361);
or U4641 (N_4641,In_747,In_844);
and U4642 (N_4642,In_33,In_664);
nor U4643 (N_4643,In_1474,In_1483);
nand U4644 (N_4644,In_321,In_447);
and U4645 (N_4645,In_396,In_809);
xnor U4646 (N_4646,In_1355,In_271);
and U4647 (N_4647,In_971,In_833);
nand U4648 (N_4648,In_174,In_1338);
and U4649 (N_4649,In_1088,In_145);
and U4650 (N_4650,In_578,In_694);
and U4651 (N_4651,In_449,In_1398);
xnor U4652 (N_4652,In_175,In_344);
and U4653 (N_4653,In_1099,In_7);
or U4654 (N_4654,In_1288,In_55);
xor U4655 (N_4655,In_1175,In_947);
nor U4656 (N_4656,In_479,In_1232);
xor U4657 (N_4657,In_1107,In_736);
nor U4658 (N_4658,In_719,In_1472);
xnor U4659 (N_4659,In_308,In_960);
nor U4660 (N_4660,In_406,In_118);
nor U4661 (N_4661,In_449,In_371);
or U4662 (N_4662,In_1195,In_886);
nor U4663 (N_4663,In_358,In_1279);
nor U4664 (N_4664,In_375,In_648);
nand U4665 (N_4665,In_658,In_731);
xor U4666 (N_4666,In_505,In_1312);
xor U4667 (N_4667,In_1166,In_840);
and U4668 (N_4668,In_856,In_530);
nand U4669 (N_4669,In_52,In_99);
nor U4670 (N_4670,In_792,In_1180);
and U4671 (N_4671,In_762,In_1485);
or U4672 (N_4672,In_1071,In_1184);
nor U4673 (N_4673,In_1356,In_550);
xnor U4674 (N_4674,In_253,In_4);
xnor U4675 (N_4675,In_1242,In_148);
nor U4676 (N_4676,In_467,In_1485);
nand U4677 (N_4677,In_622,In_985);
nor U4678 (N_4678,In_153,In_30);
or U4679 (N_4679,In_651,In_241);
or U4680 (N_4680,In_144,In_569);
or U4681 (N_4681,In_159,In_900);
or U4682 (N_4682,In_860,In_1196);
or U4683 (N_4683,In_332,In_106);
and U4684 (N_4684,In_307,In_630);
nor U4685 (N_4685,In_527,In_390);
or U4686 (N_4686,In_554,In_606);
and U4687 (N_4687,In_1497,In_799);
xor U4688 (N_4688,In_1432,In_1143);
nor U4689 (N_4689,In_130,In_518);
and U4690 (N_4690,In_1145,In_207);
and U4691 (N_4691,In_1195,In_35);
or U4692 (N_4692,In_197,In_771);
or U4693 (N_4693,In_587,In_596);
nand U4694 (N_4694,In_1010,In_1435);
and U4695 (N_4695,In_219,In_450);
and U4696 (N_4696,In_40,In_781);
xnor U4697 (N_4697,In_1464,In_436);
nand U4698 (N_4698,In_198,In_249);
nand U4699 (N_4699,In_1170,In_1125);
xor U4700 (N_4700,In_1221,In_622);
nand U4701 (N_4701,In_1321,In_1378);
or U4702 (N_4702,In_1315,In_355);
or U4703 (N_4703,In_483,In_1179);
nand U4704 (N_4704,In_1085,In_425);
xor U4705 (N_4705,In_224,In_181);
nand U4706 (N_4706,In_20,In_855);
and U4707 (N_4707,In_1058,In_496);
or U4708 (N_4708,In_639,In_132);
or U4709 (N_4709,In_790,In_1095);
or U4710 (N_4710,In_796,In_1483);
and U4711 (N_4711,In_1081,In_336);
nor U4712 (N_4712,In_1017,In_1281);
nor U4713 (N_4713,In_1353,In_593);
xor U4714 (N_4714,In_858,In_1219);
nand U4715 (N_4715,In_977,In_319);
xnor U4716 (N_4716,In_652,In_1304);
nand U4717 (N_4717,In_928,In_954);
or U4718 (N_4718,In_738,In_489);
and U4719 (N_4719,In_1292,In_792);
or U4720 (N_4720,In_1360,In_520);
nand U4721 (N_4721,In_1306,In_666);
nand U4722 (N_4722,In_131,In_198);
or U4723 (N_4723,In_1244,In_970);
nand U4724 (N_4724,In_663,In_1041);
or U4725 (N_4725,In_164,In_163);
xnor U4726 (N_4726,In_1127,In_1413);
nand U4727 (N_4727,In_385,In_1073);
or U4728 (N_4728,In_1387,In_1148);
and U4729 (N_4729,In_44,In_114);
nand U4730 (N_4730,In_829,In_1492);
or U4731 (N_4731,In_886,In_874);
nand U4732 (N_4732,In_562,In_939);
xor U4733 (N_4733,In_1003,In_732);
nand U4734 (N_4734,In_1369,In_79);
xor U4735 (N_4735,In_393,In_1029);
nand U4736 (N_4736,In_518,In_812);
or U4737 (N_4737,In_221,In_287);
or U4738 (N_4738,In_367,In_612);
or U4739 (N_4739,In_231,In_59);
or U4740 (N_4740,In_743,In_992);
nand U4741 (N_4741,In_543,In_67);
nand U4742 (N_4742,In_582,In_1212);
nor U4743 (N_4743,In_770,In_1056);
nand U4744 (N_4744,In_124,In_1438);
nand U4745 (N_4745,In_746,In_160);
xnor U4746 (N_4746,In_538,In_917);
xnor U4747 (N_4747,In_8,In_1369);
and U4748 (N_4748,In_779,In_573);
nor U4749 (N_4749,In_960,In_305);
nand U4750 (N_4750,In_1257,In_1349);
nand U4751 (N_4751,In_642,In_234);
xnor U4752 (N_4752,In_440,In_895);
nor U4753 (N_4753,In_1080,In_486);
nor U4754 (N_4754,In_1212,In_9);
or U4755 (N_4755,In_987,In_1054);
xor U4756 (N_4756,In_934,In_548);
and U4757 (N_4757,In_330,In_155);
nand U4758 (N_4758,In_859,In_1366);
xnor U4759 (N_4759,In_330,In_635);
xnor U4760 (N_4760,In_1090,In_1249);
xor U4761 (N_4761,In_303,In_1143);
nor U4762 (N_4762,In_46,In_16);
nor U4763 (N_4763,In_552,In_202);
and U4764 (N_4764,In_163,In_1367);
xnor U4765 (N_4765,In_1048,In_1157);
nand U4766 (N_4766,In_255,In_196);
nor U4767 (N_4767,In_138,In_1235);
nor U4768 (N_4768,In_55,In_1206);
or U4769 (N_4769,In_1303,In_1011);
or U4770 (N_4770,In_657,In_552);
nor U4771 (N_4771,In_457,In_878);
xnor U4772 (N_4772,In_1018,In_705);
nor U4773 (N_4773,In_936,In_617);
xor U4774 (N_4774,In_1495,In_175);
nor U4775 (N_4775,In_545,In_1029);
nand U4776 (N_4776,In_65,In_586);
or U4777 (N_4777,In_1309,In_550);
xor U4778 (N_4778,In_787,In_1256);
nand U4779 (N_4779,In_602,In_1413);
nand U4780 (N_4780,In_857,In_21);
and U4781 (N_4781,In_1395,In_101);
or U4782 (N_4782,In_885,In_1265);
and U4783 (N_4783,In_25,In_1344);
nor U4784 (N_4784,In_366,In_377);
nor U4785 (N_4785,In_503,In_949);
nand U4786 (N_4786,In_489,In_1426);
nand U4787 (N_4787,In_936,In_471);
or U4788 (N_4788,In_909,In_367);
xor U4789 (N_4789,In_651,In_105);
nand U4790 (N_4790,In_1021,In_1123);
and U4791 (N_4791,In_512,In_645);
xnor U4792 (N_4792,In_555,In_1489);
xor U4793 (N_4793,In_1404,In_1149);
xor U4794 (N_4794,In_1021,In_801);
nand U4795 (N_4795,In_633,In_527);
nor U4796 (N_4796,In_709,In_1451);
nand U4797 (N_4797,In_1329,In_356);
or U4798 (N_4798,In_713,In_195);
xnor U4799 (N_4799,In_840,In_1498);
xor U4800 (N_4800,In_946,In_91);
or U4801 (N_4801,In_122,In_759);
and U4802 (N_4802,In_548,In_958);
or U4803 (N_4803,In_1433,In_783);
nand U4804 (N_4804,In_85,In_1059);
nand U4805 (N_4805,In_795,In_231);
or U4806 (N_4806,In_710,In_993);
xor U4807 (N_4807,In_1185,In_864);
nor U4808 (N_4808,In_1154,In_818);
and U4809 (N_4809,In_1329,In_1161);
nor U4810 (N_4810,In_928,In_1298);
nor U4811 (N_4811,In_658,In_232);
or U4812 (N_4812,In_303,In_232);
and U4813 (N_4813,In_867,In_551);
nor U4814 (N_4814,In_991,In_602);
and U4815 (N_4815,In_1339,In_277);
xor U4816 (N_4816,In_1264,In_901);
xnor U4817 (N_4817,In_152,In_1068);
nor U4818 (N_4818,In_332,In_1276);
nor U4819 (N_4819,In_1204,In_1450);
xor U4820 (N_4820,In_695,In_47);
nor U4821 (N_4821,In_1465,In_421);
or U4822 (N_4822,In_692,In_782);
or U4823 (N_4823,In_382,In_350);
and U4824 (N_4824,In_768,In_264);
xor U4825 (N_4825,In_173,In_1238);
nor U4826 (N_4826,In_613,In_639);
and U4827 (N_4827,In_996,In_804);
or U4828 (N_4828,In_896,In_742);
nand U4829 (N_4829,In_1406,In_1043);
nand U4830 (N_4830,In_969,In_1114);
nand U4831 (N_4831,In_82,In_1077);
nor U4832 (N_4832,In_716,In_930);
xnor U4833 (N_4833,In_1343,In_162);
or U4834 (N_4834,In_293,In_24);
nand U4835 (N_4835,In_604,In_1264);
or U4836 (N_4836,In_1382,In_1036);
or U4837 (N_4837,In_285,In_657);
and U4838 (N_4838,In_449,In_44);
and U4839 (N_4839,In_395,In_272);
or U4840 (N_4840,In_370,In_172);
nand U4841 (N_4841,In_1101,In_1278);
xor U4842 (N_4842,In_454,In_1030);
nand U4843 (N_4843,In_875,In_405);
and U4844 (N_4844,In_171,In_1416);
and U4845 (N_4845,In_1373,In_540);
xnor U4846 (N_4846,In_1067,In_291);
nor U4847 (N_4847,In_410,In_1472);
nand U4848 (N_4848,In_942,In_1358);
and U4849 (N_4849,In_96,In_1279);
and U4850 (N_4850,In_1410,In_1420);
nor U4851 (N_4851,In_1060,In_1244);
nand U4852 (N_4852,In_1453,In_1315);
nand U4853 (N_4853,In_342,In_1166);
nand U4854 (N_4854,In_1011,In_850);
nand U4855 (N_4855,In_22,In_1352);
or U4856 (N_4856,In_20,In_921);
xnor U4857 (N_4857,In_92,In_1172);
nor U4858 (N_4858,In_889,In_296);
nor U4859 (N_4859,In_615,In_258);
nand U4860 (N_4860,In_502,In_1423);
nor U4861 (N_4861,In_1319,In_145);
or U4862 (N_4862,In_552,In_48);
nand U4863 (N_4863,In_204,In_114);
xnor U4864 (N_4864,In_1326,In_255);
nor U4865 (N_4865,In_769,In_692);
nand U4866 (N_4866,In_579,In_512);
xor U4867 (N_4867,In_1030,In_45);
xnor U4868 (N_4868,In_1124,In_548);
nor U4869 (N_4869,In_99,In_710);
nor U4870 (N_4870,In_105,In_849);
xor U4871 (N_4871,In_769,In_1169);
xor U4872 (N_4872,In_173,In_1005);
or U4873 (N_4873,In_423,In_1454);
xnor U4874 (N_4874,In_201,In_916);
nor U4875 (N_4875,In_1172,In_181);
xnor U4876 (N_4876,In_1084,In_1270);
and U4877 (N_4877,In_1066,In_6);
and U4878 (N_4878,In_168,In_303);
and U4879 (N_4879,In_908,In_242);
nor U4880 (N_4880,In_669,In_1186);
xor U4881 (N_4881,In_675,In_1103);
or U4882 (N_4882,In_112,In_990);
nand U4883 (N_4883,In_722,In_1279);
and U4884 (N_4884,In_1414,In_194);
xor U4885 (N_4885,In_512,In_1106);
nor U4886 (N_4886,In_1274,In_820);
nand U4887 (N_4887,In_951,In_579);
or U4888 (N_4888,In_223,In_1169);
xnor U4889 (N_4889,In_1481,In_726);
xor U4890 (N_4890,In_1300,In_45);
or U4891 (N_4891,In_1332,In_298);
or U4892 (N_4892,In_998,In_403);
nor U4893 (N_4893,In_172,In_421);
and U4894 (N_4894,In_345,In_318);
nand U4895 (N_4895,In_739,In_335);
nand U4896 (N_4896,In_1287,In_765);
and U4897 (N_4897,In_224,In_1117);
nand U4898 (N_4898,In_1378,In_586);
or U4899 (N_4899,In_1194,In_111);
or U4900 (N_4900,In_455,In_737);
xor U4901 (N_4901,In_254,In_790);
and U4902 (N_4902,In_1172,In_197);
xnor U4903 (N_4903,In_1276,In_560);
or U4904 (N_4904,In_1061,In_259);
nor U4905 (N_4905,In_115,In_1355);
and U4906 (N_4906,In_1066,In_894);
nand U4907 (N_4907,In_252,In_1106);
and U4908 (N_4908,In_608,In_334);
xor U4909 (N_4909,In_1400,In_241);
nor U4910 (N_4910,In_121,In_1179);
or U4911 (N_4911,In_1410,In_437);
nor U4912 (N_4912,In_759,In_1125);
nor U4913 (N_4913,In_1239,In_1204);
or U4914 (N_4914,In_559,In_452);
xnor U4915 (N_4915,In_562,In_1446);
nand U4916 (N_4916,In_198,In_1131);
or U4917 (N_4917,In_1233,In_1219);
or U4918 (N_4918,In_955,In_663);
nand U4919 (N_4919,In_566,In_784);
nor U4920 (N_4920,In_489,In_1375);
or U4921 (N_4921,In_105,In_232);
xnor U4922 (N_4922,In_374,In_220);
or U4923 (N_4923,In_1187,In_696);
nand U4924 (N_4924,In_315,In_1403);
nor U4925 (N_4925,In_960,In_873);
nor U4926 (N_4926,In_867,In_118);
or U4927 (N_4927,In_826,In_428);
xor U4928 (N_4928,In_1127,In_953);
nor U4929 (N_4929,In_1384,In_741);
nand U4930 (N_4930,In_1206,In_13);
nand U4931 (N_4931,In_501,In_904);
or U4932 (N_4932,In_889,In_632);
and U4933 (N_4933,In_1303,In_1383);
and U4934 (N_4934,In_680,In_249);
nor U4935 (N_4935,In_276,In_1288);
xor U4936 (N_4936,In_837,In_726);
xnor U4937 (N_4937,In_501,In_1026);
or U4938 (N_4938,In_83,In_454);
or U4939 (N_4939,In_796,In_1415);
and U4940 (N_4940,In_403,In_976);
or U4941 (N_4941,In_1155,In_591);
or U4942 (N_4942,In_634,In_894);
xnor U4943 (N_4943,In_1359,In_222);
or U4944 (N_4944,In_1161,In_126);
xor U4945 (N_4945,In_920,In_482);
or U4946 (N_4946,In_1299,In_876);
nand U4947 (N_4947,In_989,In_1216);
and U4948 (N_4948,In_425,In_763);
and U4949 (N_4949,In_583,In_1215);
xnor U4950 (N_4950,In_750,In_1224);
and U4951 (N_4951,In_1277,In_1236);
or U4952 (N_4952,In_531,In_1435);
or U4953 (N_4953,In_849,In_464);
xnor U4954 (N_4954,In_968,In_481);
xor U4955 (N_4955,In_114,In_597);
nor U4956 (N_4956,In_1451,In_512);
nand U4957 (N_4957,In_1324,In_1069);
nor U4958 (N_4958,In_824,In_968);
xnor U4959 (N_4959,In_931,In_77);
or U4960 (N_4960,In_874,In_137);
and U4961 (N_4961,In_5,In_216);
xnor U4962 (N_4962,In_938,In_83);
nor U4963 (N_4963,In_1065,In_575);
xor U4964 (N_4964,In_367,In_835);
or U4965 (N_4965,In_4,In_848);
and U4966 (N_4966,In_500,In_826);
and U4967 (N_4967,In_612,In_1019);
or U4968 (N_4968,In_550,In_1071);
nor U4969 (N_4969,In_1308,In_1413);
nand U4970 (N_4970,In_1408,In_218);
and U4971 (N_4971,In_724,In_952);
xnor U4972 (N_4972,In_851,In_1440);
or U4973 (N_4973,In_802,In_558);
and U4974 (N_4974,In_1075,In_648);
nand U4975 (N_4975,In_904,In_761);
nand U4976 (N_4976,In_776,In_1441);
nor U4977 (N_4977,In_1262,In_1398);
xnor U4978 (N_4978,In_872,In_1102);
xnor U4979 (N_4979,In_1329,In_807);
nand U4980 (N_4980,In_1151,In_337);
or U4981 (N_4981,In_1381,In_1128);
or U4982 (N_4982,In_309,In_862);
nand U4983 (N_4983,In_688,In_516);
nand U4984 (N_4984,In_9,In_1114);
or U4985 (N_4985,In_114,In_99);
nand U4986 (N_4986,In_67,In_1026);
xnor U4987 (N_4987,In_1300,In_1059);
nand U4988 (N_4988,In_418,In_1211);
nand U4989 (N_4989,In_404,In_994);
or U4990 (N_4990,In_952,In_229);
nand U4991 (N_4991,In_146,In_1366);
nand U4992 (N_4992,In_577,In_1243);
or U4993 (N_4993,In_938,In_975);
xnor U4994 (N_4994,In_1098,In_281);
or U4995 (N_4995,In_1140,In_1247);
and U4996 (N_4996,In_746,In_633);
nor U4997 (N_4997,In_71,In_1240);
xor U4998 (N_4998,In_492,In_473);
nand U4999 (N_4999,In_514,In_250);
or U5000 (N_5000,N_2076,N_3350);
nor U5001 (N_5001,N_3755,N_3261);
xor U5002 (N_5002,N_3733,N_275);
nor U5003 (N_5003,N_1250,N_553);
or U5004 (N_5004,N_3782,N_4683);
nor U5005 (N_5005,N_4788,N_3775);
and U5006 (N_5006,N_4860,N_1592);
and U5007 (N_5007,N_1413,N_3814);
nand U5008 (N_5008,N_3723,N_4569);
xnor U5009 (N_5009,N_4337,N_649);
nor U5010 (N_5010,N_1173,N_4892);
nor U5011 (N_5011,N_2171,N_4499);
xnor U5012 (N_5012,N_4707,N_406);
nand U5013 (N_5013,N_4110,N_3749);
nor U5014 (N_5014,N_185,N_4100);
and U5015 (N_5015,N_4019,N_2640);
xor U5016 (N_5016,N_1615,N_2251);
nand U5017 (N_5017,N_1837,N_601);
nand U5018 (N_5018,N_4671,N_549);
xor U5019 (N_5019,N_3793,N_2086);
or U5020 (N_5020,N_1417,N_3416);
nor U5021 (N_5021,N_2091,N_2921);
nand U5022 (N_5022,N_731,N_814);
xnor U5023 (N_5023,N_4547,N_2328);
and U5024 (N_5024,N_2914,N_2273);
nand U5025 (N_5025,N_4712,N_4343);
or U5026 (N_5026,N_3007,N_3560);
or U5027 (N_5027,N_3461,N_458);
or U5028 (N_5028,N_984,N_4317);
and U5029 (N_5029,N_3288,N_3199);
or U5030 (N_5030,N_1727,N_2505);
or U5031 (N_5031,N_1560,N_328);
nand U5032 (N_5032,N_4801,N_4239);
nor U5033 (N_5033,N_811,N_1405);
or U5034 (N_5034,N_3044,N_2429);
nor U5035 (N_5035,N_292,N_3791);
nand U5036 (N_5036,N_3349,N_1677);
xor U5037 (N_5037,N_1061,N_1717);
and U5038 (N_5038,N_3215,N_4280);
or U5039 (N_5039,N_1194,N_3283);
xor U5040 (N_5040,N_3668,N_1799);
xor U5041 (N_5041,N_212,N_4886);
or U5042 (N_5042,N_2025,N_283);
or U5043 (N_5043,N_2306,N_4898);
and U5044 (N_5044,N_3996,N_3903);
nand U5045 (N_5045,N_2634,N_2063);
nand U5046 (N_5046,N_2973,N_4717);
nor U5047 (N_5047,N_4615,N_96);
nor U5048 (N_5048,N_1334,N_1768);
nand U5049 (N_5049,N_914,N_815);
nand U5050 (N_5050,N_3824,N_2827);
xnor U5051 (N_5051,N_3522,N_4639);
xor U5052 (N_5052,N_4956,N_4245);
or U5053 (N_5053,N_3969,N_390);
nor U5054 (N_5054,N_1458,N_1190);
and U5055 (N_5055,N_2998,N_4274);
and U5056 (N_5056,N_1374,N_4688);
or U5057 (N_5057,N_4799,N_2960);
nor U5058 (N_5058,N_4390,N_2682);
nor U5059 (N_5059,N_104,N_1776);
nor U5060 (N_5060,N_2678,N_371);
nor U5061 (N_5061,N_2800,N_1761);
nand U5062 (N_5062,N_1435,N_1611);
xor U5063 (N_5063,N_4939,N_3123);
or U5064 (N_5064,N_3615,N_3130);
xnor U5065 (N_5065,N_3605,N_4980);
xnor U5066 (N_5066,N_1702,N_643);
nor U5067 (N_5067,N_1311,N_1527);
nor U5068 (N_5068,N_4722,N_1397);
or U5069 (N_5069,N_3997,N_1986);
nor U5070 (N_5070,N_1286,N_732);
nor U5071 (N_5071,N_950,N_2695);
nand U5072 (N_5072,N_173,N_4310);
or U5073 (N_5073,N_1925,N_1453);
nand U5074 (N_5074,N_4412,N_2624);
and U5075 (N_5075,N_2233,N_3492);
or U5076 (N_5076,N_4052,N_3392);
and U5077 (N_5077,N_2408,N_40);
or U5078 (N_5078,N_1132,N_2984);
and U5079 (N_5079,N_4861,N_1525);
nand U5080 (N_5080,N_2106,N_2254);
and U5081 (N_5081,N_4125,N_317);
or U5082 (N_5082,N_2206,N_4432);
nand U5083 (N_5083,N_2940,N_502);
nand U5084 (N_5084,N_2475,N_531);
nor U5085 (N_5085,N_3906,N_452);
or U5086 (N_5086,N_1310,N_2279);
xnor U5087 (N_5087,N_1995,N_4562);
and U5088 (N_5088,N_2765,N_3558);
xnor U5089 (N_5089,N_4525,N_2889);
nand U5090 (N_5090,N_4720,N_1695);
and U5091 (N_5091,N_2882,N_1756);
nand U5092 (N_5092,N_3256,N_1680);
nand U5093 (N_5093,N_1967,N_740);
or U5094 (N_5094,N_2437,N_4395);
and U5095 (N_5095,N_3355,N_1539);
or U5096 (N_5096,N_78,N_1123);
and U5097 (N_5097,N_1635,N_1801);
nor U5098 (N_5098,N_3002,N_4992);
nand U5099 (N_5099,N_2215,N_3189);
nand U5100 (N_5100,N_3157,N_1876);
and U5101 (N_5101,N_1710,N_791);
xor U5102 (N_5102,N_3999,N_1326);
and U5103 (N_5103,N_841,N_1213);
nor U5104 (N_5104,N_4355,N_385);
xnor U5105 (N_5105,N_230,N_2824);
nor U5106 (N_5106,N_1728,N_600);
nor U5107 (N_5107,N_4117,N_478);
nand U5108 (N_5108,N_4560,N_4794);
nor U5109 (N_5109,N_403,N_4542);
nor U5110 (N_5110,N_3340,N_4650);
or U5111 (N_5111,N_3036,N_4571);
nor U5112 (N_5112,N_4001,N_2690);
or U5113 (N_5113,N_3704,N_3736);
and U5114 (N_5114,N_623,N_3436);
nor U5115 (N_5115,N_113,N_4630);
nor U5116 (N_5116,N_2459,N_3014);
nand U5117 (N_5117,N_2418,N_3665);
nor U5118 (N_5118,N_1751,N_1038);
nand U5119 (N_5119,N_3098,N_3404);
nand U5120 (N_5120,N_312,N_3487);
nor U5121 (N_5121,N_439,N_1234);
or U5122 (N_5122,N_1515,N_1016);
or U5123 (N_5123,N_621,N_1044);
nor U5124 (N_5124,N_2795,N_2278);
nor U5125 (N_5125,N_1272,N_3391);
or U5126 (N_5126,N_3105,N_2718);
nor U5127 (N_5127,N_4619,N_509);
nand U5128 (N_5128,N_1519,N_960);
nor U5129 (N_5129,N_1419,N_1073);
or U5130 (N_5130,N_2806,N_3710);
or U5131 (N_5131,N_4006,N_1386);
or U5132 (N_5132,N_1284,N_1468);
nand U5133 (N_5133,N_3735,N_4585);
nor U5134 (N_5134,N_2517,N_1307);
xnor U5135 (N_5135,N_3221,N_2180);
and U5136 (N_5136,N_4523,N_1464);
nor U5137 (N_5137,N_1873,N_3718);
nand U5138 (N_5138,N_443,N_4561);
xor U5139 (N_5139,N_3318,N_622);
nor U5140 (N_5140,N_4544,N_2837);
and U5141 (N_5141,N_842,N_2691);
nor U5142 (N_5142,N_4051,N_1993);
xnor U5143 (N_5143,N_4495,N_4709);
nor U5144 (N_5144,N_2699,N_758);
and U5145 (N_5145,N_466,N_614);
nand U5146 (N_5146,N_3981,N_4577);
and U5147 (N_5147,N_2404,N_4424);
or U5148 (N_5148,N_350,N_1989);
nand U5149 (N_5149,N_4084,N_615);
nor U5150 (N_5150,N_4692,N_1654);
or U5151 (N_5151,N_3308,N_2573);
or U5152 (N_5152,N_1834,N_124);
nor U5153 (N_5153,N_4821,N_65);
nand U5154 (N_5154,N_3109,N_4697);
xor U5155 (N_5155,N_2083,N_3973);
nand U5156 (N_5156,N_874,N_1590);
and U5157 (N_5157,N_2116,N_1809);
and U5158 (N_5158,N_2348,N_4475);
or U5159 (N_5159,N_1984,N_3582);
nand U5160 (N_5160,N_3376,N_2117);
and U5161 (N_5161,N_2567,N_3863);
xnor U5162 (N_5162,N_581,N_3621);
nor U5163 (N_5163,N_2426,N_4737);
and U5164 (N_5164,N_433,N_3167);
xnor U5165 (N_5165,N_3013,N_1257);
and U5166 (N_5166,N_2876,N_2399);
nand U5167 (N_5167,N_3887,N_2257);
or U5168 (N_5168,N_802,N_1109);
and U5169 (N_5169,N_4854,N_4604);
or U5170 (N_5170,N_2022,N_4696);
or U5171 (N_5171,N_4748,N_2637);
xor U5172 (N_5172,N_3222,N_2043);
or U5173 (N_5173,N_3609,N_4220);
and U5174 (N_5174,N_3364,N_1080);
and U5175 (N_5175,N_4864,N_1953);
nand U5176 (N_5176,N_2137,N_2146);
and U5177 (N_5177,N_3656,N_477);
or U5178 (N_5178,N_2230,N_2518);
nand U5179 (N_5179,N_3988,N_1549);
xor U5180 (N_5180,N_2884,N_3190);
xnor U5181 (N_5181,N_1529,N_866);
xor U5182 (N_5182,N_3385,N_778);
xor U5183 (N_5183,N_98,N_1682);
or U5184 (N_5184,N_1960,N_4134);
or U5185 (N_5185,N_1156,N_498);
nand U5186 (N_5186,N_2458,N_4917);
or U5187 (N_5187,N_1671,N_2142);
xnor U5188 (N_5188,N_1785,N_450);
or U5189 (N_5189,N_3020,N_3091);
xor U5190 (N_5190,N_2357,N_1747);
nand U5191 (N_5191,N_2187,N_4570);
or U5192 (N_5192,N_869,N_2340);
or U5193 (N_5193,N_4434,N_481);
nor U5194 (N_5194,N_4775,N_1588);
xnor U5195 (N_5195,N_770,N_1906);
and U5196 (N_5196,N_933,N_789);
and U5197 (N_5197,N_1301,N_4059);
or U5198 (N_5198,N_1455,N_1322);
or U5199 (N_5199,N_3546,N_4279);
xnor U5200 (N_5200,N_1782,N_4676);
or U5201 (N_5201,N_998,N_3849);
nor U5202 (N_5202,N_3462,N_339);
nand U5203 (N_5203,N_2968,N_3207);
nor U5204 (N_5204,N_3942,N_3305);
and U5205 (N_5205,N_2620,N_497);
xnor U5206 (N_5206,N_3620,N_62);
nor U5207 (N_5207,N_4290,N_3345);
and U5208 (N_5208,N_4575,N_4930);
or U5209 (N_5209,N_4330,N_3822);
xnor U5210 (N_5210,N_579,N_1885);
and U5211 (N_5211,N_3081,N_2727);
and U5212 (N_5212,N_3696,N_3317);
or U5213 (N_5213,N_1649,N_2420);
and U5214 (N_5214,N_3511,N_763);
nand U5215 (N_5215,N_3515,N_1442);
or U5216 (N_5216,N_784,N_1806);
and U5217 (N_5217,N_4485,N_4361);
and U5218 (N_5218,N_4158,N_2021);
nand U5219 (N_5219,N_3227,N_47);
xnor U5220 (N_5220,N_3096,N_1443);
nand U5221 (N_5221,N_4987,N_1872);
xnor U5222 (N_5222,N_3417,N_4625);
and U5223 (N_5223,N_2006,N_3631);
nand U5224 (N_5224,N_4477,N_3662);
or U5225 (N_5225,N_4471,N_2170);
and U5226 (N_5226,N_1495,N_3667);
xor U5227 (N_5227,N_3532,N_4715);
nor U5228 (N_5228,N_229,N_3770);
nand U5229 (N_5229,N_4282,N_979);
nor U5230 (N_5230,N_1570,N_1632);
and U5231 (N_5231,N_4098,N_4305);
nand U5232 (N_5232,N_2852,N_2675);
nor U5233 (N_5233,N_3984,N_3917);
nor U5234 (N_5234,N_454,N_3865);
and U5235 (N_5235,N_4512,N_3049);
nand U5236 (N_5236,N_2923,N_4368);
xor U5237 (N_5237,N_1857,N_1875);
xor U5238 (N_5238,N_2160,N_1520);
xnor U5239 (N_5239,N_902,N_4701);
nand U5240 (N_5240,N_4918,N_1970);
nand U5241 (N_5241,N_1990,N_4469);
nand U5242 (N_5242,N_1431,N_3242);
nand U5243 (N_5243,N_1302,N_4408);
nor U5244 (N_5244,N_1790,N_3720);
nand U5245 (N_5245,N_4359,N_4350);
xor U5246 (N_5246,N_1911,N_2445);
xor U5247 (N_5247,N_2834,N_424);
or U5248 (N_5248,N_2297,N_3080);
and U5249 (N_5249,N_3274,N_2093);
xor U5250 (N_5250,N_4587,N_3071);
nand U5251 (N_5251,N_1623,N_8);
nand U5252 (N_5252,N_4165,N_1124);
nor U5253 (N_5253,N_2967,N_3692);
or U5254 (N_5254,N_3832,N_1506);
nand U5255 (N_5255,N_1810,N_3562);
or U5256 (N_5256,N_1805,N_1736);
xnor U5257 (N_5257,N_1867,N_1916);
or U5258 (N_5258,N_2349,N_4186);
and U5259 (N_5259,N_2683,N_3358);
or U5260 (N_5260,N_3373,N_3471);
and U5261 (N_5261,N_2312,N_1434);
nor U5262 (N_5262,N_4196,N_2268);
or U5263 (N_5263,N_1254,N_1847);
or U5264 (N_5264,N_1369,N_2151);
nor U5265 (N_5265,N_1533,N_2771);
xor U5266 (N_5266,N_3874,N_2071);
or U5267 (N_5267,N_2059,N_1343);
xor U5268 (N_5268,N_2961,N_868);
xnor U5269 (N_5269,N_4442,N_4143);
or U5270 (N_5270,N_3410,N_9);
xnor U5271 (N_5271,N_3622,N_4747);
and U5272 (N_5272,N_3729,N_1764);
xor U5273 (N_5273,N_3425,N_728);
or U5274 (N_5274,N_3528,N_2139);
and U5275 (N_5275,N_2177,N_1412);
xor U5276 (N_5276,N_4822,N_1147);
xnor U5277 (N_5277,N_3208,N_852);
and U5278 (N_5278,N_1192,N_4530);
or U5279 (N_5279,N_3559,N_965);
nand U5280 (N_5280,N_4172,N_2596);
xnor U5281 (N_5281,N_4470,N_3165);
and U5282 (N_5282,N_4520,N_701);
nor U5283 (N_5283,N_1071,N_1952);
or U5284 (N_5284,N_1796,N_800);
nor U5285 (N_5285,N_3217,N_2199);
xnor U5286 (N_5286,N_2088,N_4629);
nor U5287 (N_5287,N_1774,N_2702);
and U5288 (N_5288,N_2748,N_4855);
nand U5289 (N_5289,N_1981,N_3498);
nand U5290 (N_5290,N_4986,N_2195);
xnor U5291 (N_5291,N_1472,N_75);
and U5292 (N_5292,N_311,N_3494);
nand U5293 (N_5293,N_2974,N_1196);
and U5294 (N_5294,N_3001,N_4675);
or U5295 (N_5295,N_3534,N_4246);
nand U5296 (N_5296,N_4035,N_1932);
xor U5297 (N_5297,N_990,N_4095);
xor U5298 (N_5298,N_3690,N_447);
or U5299 (N_5299,N_3257,N_2997);
or U5300 (N_5300,N_266,N_2052);
and U5301 (N_5301,N_2149,N_915);
or U5302 (N_5302,N_1200,N_2582);
xor U5303 (N_5303,N_3188,N_1714);
nand U5304 (N_5304,N_4459,N_2466);
nand U5305 (N_5305,N_3581,N_107);
or U5306 (N_5306,N_1400,N_4654);
nand U5307 (N_5307,N_3037,N_118);
or U5308 (N_5308,N_1188,N_4580);
or U5309 (N_5309,N_734,N_3160);
nor U5310 (N_5310,N_2693,N_4056);
or U5311 (N_5311,N_3170,N_2299);
nand U5312 (N_5312,N_1202,N_3435);
xor U5313 (N_5313,N_1441,N_508);
nand U5314 (N_5314,N_810,N_4677);
or U5315 (N_5315,N_4309,N_3264);
nor U5316 (N_5316,N_2965,N_2330);
nand U5317 (N_5317,N_894,N_123);
nor U5318 (N_5318,N_3053,N_1377);
or U5319 (N_5319,N_144,N_1933);
or U5320 (N_5320,N_20,N_2887);
or U5321 (N_5321,N_1956,N_1807);
nor U5322 (N_5322,N_2506,N_3677);
nor U5323 (N_5323,N_560,N_4094);
or U5324 (N_5324,N_1026,N_704);
nor U5325 (N_5325,N_652,N_343);
or U5326 (N_5326,N_1328,N_3252);
nor U5327 (N_5327,N_535,N_840);
nor U5328 (N_5328,N_1891,N_3235);
xnor U5329 (N_5329,N_4136,N_3951);
nand U5330 (N_5330,N_3544,N_4155);
nand U5331 (N_5331,N_1079,N_4262);
xor U5332 (N_5332,N_3919,N_4414);
and U5333 (N_5333,N_891,N_364);
nor U5334 (N_5334,N_3218,N_922);
and U5335 (N_5335,N_2794,N_3888);
xnor U5336 (N_5336,N_1365,N_259);
nand U5337 (N_5337,N_1424,N_72);
xor U5338 (N_5338,N_4809,N_2947);
nand U5339 (N_5339,N_883,N_1329);
or U5340 (N_5340,N_3458,N_3553);
or U5341 (N_5341,N_4071,N_4230);
nand U5342 (N_5342,N_1423,N_611);
or U5343 (N_5343,N_4429,N_2939);
nor U5344 (N_5344,N_2452,N_4351);
nand U5345 (N_5345,N_335,N_4876);
and U5346 (N_5346,N_2026,N_4732);
or U5347 (N_5347,N_220,N_4759);
nand U5348 (N_5348,N_2724,N_214);
nor U5349 (N_5349,N_356,N_2432);
xnor U5350 (N_5350,N_1998,N_1593);
xor U5351 (N_5351,N_3666,N_799);
or U5352 (N_5352,N_3563,N_4405);
or U5353 (N_5353,N_2296,N_3589);
xnor U5354 (N_5354,N_4138,N_4693);
xor U5355 (N_5355,N_2435,N_386);
and U5356 (N_5356,N_1220,N_2148);
nor U5357 (N_5357,N_774,N_2867);
nor U5358 (N_5358,N_4959,N_781);
xor U5359 (N_5359,N_2104,N_2809);
xor U5360 (N_5360,N_825,N_4597);
or U5361 (N_5361,N_2542,N_573);
nand U5362 (N_5362,N_1040,N_1171);
and U5363 (N_5363,N_700,N_3);
xnor U5364 (N_5364,N_854,N_3859);
nor U5365 (N_5365,N_1685,N_2666);
nor U5366 (N_5366,N_3805,N_867);
or U5367 (N_5367,N_566,N_1069);
xor U5368 (N_5368,N_876,N_4229);
nor U5369 (N_5369,N_2274,N_3073);
nand U5370 (N_5370,N_968,N_2775);
nor U5371 (N_5371,N_4631,N_2654);
and U5372 (N_5372,N_3867,N_4257);
or U5373 (N_5373,N_2388,N_3518);
xor U5374 (N_5374,N_2796,N_2167);
or U5375 (N_5375,N_2628,N_4616);
or U5376 (N_5376,N_3357,N_1313);
and U5377 (N_5377,N_4106,N_175);
and U5378 (N_5378,N_4289,N_2912);
or U5379 (N_5379,N_1603,N_1186);
xnor U5380 (N_5380,N_1606,N_4481);
or U5381 (N_5381,N_1036,N_2526);
nor U5382 (N_5382,N_2182,N_4632);
and U5383 (N_5383,N_2287,N_598);
nand U5384 (N_5384,N_1544,N_1007);
xor U5385 (N_5385,N_1056,N_2038);
nor U5386 (N_5386,N_1612,N_3974);
and U5387 (N_5387,N_1499,N_3638);
xnor U5388 (N_5388,N_4425,N_4595);
xnor U5389 (N_5389,N_3482,N_1237);
xor U5390 (N_5390,N_3716,N_161);
nand U5391 (N_5391,N_2598,N_315);
or U5392 (N_5392,N_3882,N_4658);
nor U5393 (N_5393,N_2770,N_3079);
and U5394 (N_5394,N_596,N_1251);
nand U5395 (N_5395,N_861,N_1347);
or U5396 (N_5396,N_583,N_771);
or U5397 (N_5397,N_1162,N_1881);
nand U5398 (N_5398,N_4154,N_4912);
nand U5399 (N_5399,N_2872,N_483);
nand U5400 (N_5400,N_3672,N_3398);
nand U5401 (N_5401,N_4124,N_524);
or U5402 (N_5402,N_2041,N_402);
or U5403 (N_5403,N_3426,N_1022);
or U5404 (N_5404,N_1771,N_3178);
nand U5405 (N_5405,N_1822,N_325);
and U5406 (N_5406,N_2720,N_1909);
nor U5407 (N_5407,N_1296,N_4506);
nor U5408 (N_5408,N_479,N_3139);
or U5409 (N_5409,N_4275,N_1391);
xor U5410 (N_5410,N_1898,N_994);
nor U5411 (N_5411,N_4652,N_4844);
or U5412 (N_5412,N_1426,N_3322);
or U5413 (N_5413,N_2845,N_1346);
nand U5414 (N_5414,N_102,N_297);
nand U5415 (N_5415,N_4311,N_2134);
or U5416 (N_5416,N_3005,N_2808);
and U5417 (N_5417,N_140,N_4335);
nand U5418 (N_5418,N_4925,N_4823);
nor U5419 (N_5419,N_4741,N_1081);
or U5420 (N_5420,N_3852,N_1380);
xnor U5421 (N_5421,N_862,N_61);
and U5422 (N_5422,N_4492,N_2407);
nand U5423 (N_5423,N_2838,N_827);
nand U5424 (N_5424,N_1877,N_3493);
nand U5425 (N_5425,N_4769,N_2092);
nor U5426 (N_5426,N_900,N_1824);
nor U5427 (N_5427,N_3034,N_4030);
nor U5428 (N_5428,N_1724,N_2712);
xnor U5429 (N_5429,N_81,N_2613);
xnor U5430 (N_5430,N_4270,N_73);
and U5431 (N_5431,N_1140,N_4315);
or U5432 (N_5432,N_1339,N_4932);
nor U5433 (N_5433,N_4089,N_2860);
nand U5434 (N_5434,N_3259,N_1367);
nand U5435 (N_5435,N_1798,N_2111);
nor U5436 (N_5436,N_3590,N_831);
or U5437 (N_5437,N_2057,N_3653);
xor U5438 (N_5438,N_1735,N_1829);
and U5439 (N_5439,N_280,N_1314);
nand U5440 (N_5440,N_2866,N_2721);
xnor U5441 (N_5441,N_3226,N_690);
nor U5442 (N_5442,N_2497,N_3442);
nor U5443 (N_5443,N_2970,N_1031);
and U5444 (N_5444,N_219,N_3172);
and U5445 (N_5445,N_3606,N_1144);
nand U5446 (N_5446,N_2164,N_194);
and U5447 (N_5447,N_2283,N_1559);
xnor U5448 (N_5448,N_193,N_673);
nor U5449 (N_5449,N_2050,N_4008);
or U5450 (N_5450,N_797,N_1248);
or U5451 (N_5451,N_1550,N_459);
xnor U5452 (N_5452,N_3192,N_4914);
xnor U5453 (N_5453,N_4736,N_4074);
nand U5454 (N_5454,N_3925,N_2723);
or U5455 (N_5455,N_1586,N_4944);
and U5456 (N_5456,N_3248,N_4713);
nor U5457 (N_5457,N_4226,N_3597);
xor U5458 (N_5458,N_1762,N_4097);
nand U5459 (N_5459,N_4785,N_204);
nand U5460 (N_5460,N_2861,N_23);
nor U5461 (N_5461,N_1573,N_4116);
nand U5462 (N_5462,N_3086,N_4611);
nand U5463 (N_5463,N_2925,N_3128);
nand U5464 (N_5464,N_3296,N_3163);
xnor U5465 (N_5465,N_4958,N_3871);
and U5466 (N_5466,N_4271,N_3712);
or U5467 (N_5467,N_4762,N_4133);
nand U5468 (N_5468,N_1502,N_1224);
and U5469 (N_5469,N_482,N_3564);
and U5470 (N_5470,N_966,N_441);
or U5471 (N_5471,N_2439,N_3754);
xnor U5472 (N_5472,N_3801,N_3649);
and U5473 (N_5473,N_1214,N_235);
nand U5474 (N_5474,N_2292,N_1097);
xor U5475 (N_5475,N_4160,N_2286);
nand U5476 (N_5476,N_3354,N_4563);
or U5477 (N_5477,N_4935,N_2096);
and U5478 (N_5478,N_2764,N_249);
and U5479 (N_5479,N_3070,N_4897);
nand U5480 (N_5480,N_2152,N_2653);
and U5481 (N_5481,N_2243,N_2544);
xnor U5482 (N_5482,N_2554,N_4387);
nor U5483 (N_5483,N_4127,N_1759);
nor U5484 (N_5484,N_3224,N_1731);
and U5485 (N_5485,N_3778,N_2519);
nand U5486 (N_5486,N_4260,N_3780);
or U5487 (N_5487,N_119,N_3279);
and U5488 (N_5488,N_822,N_1134);
or U5489 (N_5489,N_2803,N_1045);
and U5490 (N_5490,N_1425,N_2431);
or U5491 (N_5491,N_3454,N_4248);
and U5492 (N_5492,N_2419,N_561);
nor U5493 (N_5493,N_331,N_1161);
or U5494 (N_5494,N_2652,N_3989);
and U5495 (N_5495,N_1792,N_3790);
nand U5496 (N_5496,N_4787,N_1690);
xor U5497 (N_5497,N_263,N_1420);
and U5498 (N_5498,N_4567,N_3877);
or U5499 (N_5499,N_2983,N_4233);
nand U5500 (N_5500,N_4907,N_2358);
nand U5501 (N_5501,N_225,N_326);
xnor U5502 (N_5502,N_425,N_4754);
xnor U5503 (N_5503,N_1631,N_4483);
nand U5504 (N_5504,N_4755,N_730);
nand U5505 (N_5505,N_3823,N_957);
and U5506 (N_5506,N_3727,N_1866);
nand U5507 (N_5507,N_2515,N_1725);
or U5508 (N_5508,N_949,N_4719);
nand U5509 (N_5509,N_1922,N_2389);
or U5510 (N_5510,N_1291,N_3861);
nand U5511 (N_5511,N_1940,N_1467);
and U5512 (N_5512,N_1901,N_4291);
nand U5513 (N_5513,N_3807,N_2423);
and U5514 (N_5514,N_1107,N_4963);
nor U5515 (N_5515,N_1878,N_3505);
and U5516 (N_5516,N_1800,N_1924);
nor U5517 (N_5517,N_3846,N_4394);
or U5518 (N_5518,N_3552,N_4076);
nand U5519 (N_5519,N_2898,N_2009);
nor U5520 (N_5520,N_3403,N_3043);
nor U5521 (N_5521,N_1083,N_3635);
or U5522 (N_5522,N_4764,N_1067);
nand U5523 (N_5523,N_2001,N_4557);
nand U5524 (N_5524,N_27,N_2324);
nor U5525 (N_5525,N_3228,N_1804);
nor U5526 (N_5526,N_4072,N_1803);
nor U5527 (N_5527,N_455,N_2669);
and U5528 (N_5528,N_4321,N_830);
or U5529 (N_5529,N_1490,N_3250);
and U5530 (N_5530,N_3858,N_4657);
xor U5531 (N_5531,N_1641,N_2015);
and U5532 (N_5532,N_3113,N_1235);
nand U5533 (N_5533,N_377,N_2670);
xnor U5534 (N_5534,N_309,N_2759);
and U5535 (N_5535,N_2725,N_2455);
or U5536 (N_5536,N_2290,N_1914);
nand U5537 (N_5537,N_1966,N_1258);
nor U5538 (N_5538,N_837,N_2143);
xnor U5539 (N_5539,N_4295,N_3521);
nand U5540 (N_5540,N_3839,N_794);
nand U5541 (N_5541,N_158,N_3757);
and U5542 (N_5542,N_3689,N_378);
xnor U5543 (N_5543,N_637,N_4392);
and U5544 (N_5544,N_3437,N_2562);
nor U5545 (N_5545,N_4507,N_3298);
nor U5546 (N_5546,N_4264,N_1227);
and U5547 (N_5547,N_1910,N_1851);
nor U5548 (N_5548,N_1253,N_4009);
nor U5549 (N_5549,N_2788,N_924);
and U5550 (N_5550,N_4659,N_340);
xnor U5551 (N_5551,N_3448,N_4955);
or U5552 (N_5552,N_1651,N_2603);
and U5553 (N_5553,N_3598,N_4645);
nand U5554 (N_5554,N_3360,N_3844);
nor U5555 (N_5555,N_1485,N_4763);
or U5556 (N_5556,N_790,N_170);
xnor U5557 (N_5557,N_2208,N_4204);
xnor U5558 (N_5558,N_4064,N_57);
or U5559 (N_5559,N_824,N_1575);
nand U5560 (N_5560,N_2097,N_3162);
or U5561 (N_5561,N_67,N_3066);
or U5562 (N_5562,N_3876,N_702);
xor U5563 (N_5563,N_1630,N_3230);
xor U5564 (N_5564,N_4043,N_591);
nor U5565 (N_5565,N_3985,N_1949);
nor U5566 (N_5566,N_426,N_2988);
or U5567 (N_5567,N_4760,N_1935);
or U5568 (N_5568,N_1681,N_4792);
nand U5569 (N_5569,N_1514,N_1563);
xor U5570 (N_5570,N_4894,N_255);
and U5571 (N_5571,N_2556,N_4366);
xor U5572 (N_5572,N_1927,N_2642);
nand U5573 (N_5573,N_1243,N_4943);
or U5574 (N_5574,N_242,N_4213);
xnor U5575 (N_5575,N_2696,N_1408);
and U5576 (N_5576,N_4396,N_4433);
nand U5577 (N_5577,N_1662,N_1551);
nor U5578 (N_5578,N_3960,N_4480);
nand U5579 (N_5579,N_1154,N_1555);
xnor U5580 (N_5580,N_2830,N_2661);
and U5581 (N_5581,N_3928,N_3082);
and U5582 (N_5582,N_3205,N_4589);
and U5583 (N_5583,N_3023,N_247);
or U5584 (N_5584,N_4786,N_4024);
nor U5585 (N_5585,N_86,N_1151);
and U5586 (N_5586,N_1241,N_1013);
nor U5587 (N_5587,N_608,N_2665);
nor U5588 (N_5588,N_3978,N_1047);
and U5589 (N_5589,N_3701,N_3746);
and U5590 (N_5590,N_2561,N_3278);
or U5591 (N_5591,N_327,N_4417);
xor U5592 (N_5592,N_1627,N_4803);
nand U5593 (N_5593,N_200,N_3625);
xnor U5594 (N_5594,N_3545,N_3862);
or U5595 (N_5595,N_3549,N_3926);
and U5596 (N_5596,N_4926,N_4496);
nand U5597 (N_5597,N_2090,N_4551);
and U5598 (N_5598,N_2917,N_2710);
xnor U5599 (N_5599,N_3099,N_4256);
xnor U5600 (N_5600,N_2060,N_4105);
and U5601 (N_5601,N_3307,N_1183);
and U5602 (N_5602,N_400,N_3135);
and U5603 (N_5603,N_4746,N_1091);
and U5604 (N_5604,N_709,N_3835);
nor U5605 (N_5605,N_1687,N_1064);
or U5606 (N_5606,N_2793,N_4142);
xnor U5607 (N_5607,N_1958,N_783);
nand U5608 (N_5608,N_1709,N_3808);
nor U5609 (N_5609,N_4814,N_3963);
nor U5610 (N_5610,N_780,N_3837);
and U5611 (N_5611,N_1480,N_3470);
and U5612 (N_5612,N_337,N_4126);
xor U5613 (N_5613,N_3580,N_2522);
and U5614 (N_5614,N_1526,N_4320);
or U5615 (N_5615,N_4118,N_3131);
nor U5616 (N_5616,N_3281,N_2786);
or U5617 (N_5617,N_4872,N_1325);
or U5618 (N_5618,N_1043,N_4448);
nor U5619 (N_5619,N_2531,N_2401);
nand U5620 (N_5620,N_3468,N_1167);
nor U5621 (N_5621,N_1655,N_1860);
nand U5622 (N_5622,N_2713,N_1379);
nand U5623 (N_5623,N_4430,N_708);
and U5624 (N_5624,N_1861,N_176);
xor U5625 (N_5625,N_3406,N_559);
nor U5626 (N_5626,N_2591,N_2843);
and U5627 (N_5627,N_3753,N_1133);
or U5628 (N_5628,N_884,N_2863);
xor U5629 (N_5629,N_4695,N_3347);
xnor U5630 (N_5630,N_1948,N_4357);
or U5631 (N_5631,N_391,N_4789);
and U5632 (N_5632,N_4422,N_3830);
xor U5633 (N_5633,N_1492,N_4191);
xnor U5634 (N_5634,N_2463,N_2572);
or U5635 (N_5635,N_3295,N_2311);
or U5636 (N_5636,N_2301,N_4928);
nor U5637 (N_5637,N_2959,N_1583);
or U5638 (N_5638,N_2886,N_1078);
or U5639 (N_5639,N_460,N_992);
or U5640 (N_5640,N_2446,N_4656);
or U5641 (N_5641,N_3460,N_2535);
nand U5642 (N_5642,N_2881,N_4088);
or U5643 (N_5643,N_1475,N_4038);
nor U5644 (N_5644,N_417,N_826);
xnor U5645 (N_5645,N_892,N_4140);
nand U5646 (N_5646,N_3247,N_2018);
xor U5647 (N_5647,N_3077,N_953);
xnor U5648 (N_5648,N_1991,N_419);
nor U5649 (N_5649,N_4624,N_2173);
and U5650 (N_5650,N_1208,N_3596);
or U5651 (N_5651,N_2468,N_2717);
nand U5652 (N_5652,N_2651,N_605);
xnor U5653 (N_5653,N_370,N_375);
and U5654 (N_5654,N_2361,N_1090);
and U5655 (N_5655,N_4850,N_4203);
xor U5656 (N_5656,N_4841,N_3399);
nand U5657 (N_5657,N_3161,N_4808);
nand U5658 (N_5658,N_1268,N_4610);
or U5659 (N_5659,N_1629,N_3765);
nor U5660 (N_5660,N_159,N_2757);
nor U5661 (N_5661,N_3149,N_1247);
nand U5662 (N_5662,N_1516,N_3380);
nor U5663 (N_5663,N_3845,N_4960);
nor U5664 (N_5664,N_1230,N_2857);
and U5665 (N_5665,N_786,N_1609);
nand U5666 (N_5666,N_132,N_1359);
nand U5667 (N_5667,N_1784,N_752);
and U5668 (N_5668,N_4251,N_773);
nor U5669 (N_5669,N_2481,N_4488);
xnor U5670 (N_5670,N_4498,N_4674);
xnor U5671 (N_5671,N_1633,N_0);
xnor U5672 (N_5672,N_2600,N_1169);
or U5673 (N_5673,N_4528,N_3719);
or U5674 (N_5674,N_1141,N_648);
and U5675 (N_5675,N_299,N_4016);
or U5676 (N_5676,N_2135,N_3838);
nor U5677 (N_5677,N_4050,N_2714);
or U5678 (N_5678,N_112,N_4132);
or U5679 (N_5679,N_3616,N_1111);
and U5680 (N_5680,N_4445,N_4119);
nand U5681 (N_5681,N_3320,N_2291);
or U5682 (N_5682,N_1832,N_3272);
and U5683 (N_5683,N_307,N_4416);
nand U5684 (N_5684,N_1179,N_3503);
nor U5685 (N_5685,N_3232,N_681);
xor U5686 (N_5686,N_3731,N_4607);
nand U5687 (N_5687,N_712,N_1017);
and U5688 (N_5688,N_4129,N_2000);
xor U5689 (N_5689,N_1817,N_4847);
nand U5690 (N_5690,N_2275,N_3991);
or U5691 (N_5691,N_93,N_2858);
or U5692 (N_5692,N_4021,N_4168);
and U5693 (N_5693,N_4478,N_506);
and U5694 (N_5694,N_484,N_2364);
and U5695 (N_5695,N_429,N_738);
nand U5696 (N_5696,N_1205,N_1309);
and U5697 (N_5697,N_4997,N_3554);
and U5698 (N_5698,N_1285,N_1460);
and U5699 (N_5699,N_1136,N_3277);
xnor U5700 (N_5700,N_4238,N_231);
nor U5701 (N_5701,N_1034,N_3419);
nand U5702 (N_5702,N_1269,N_1149);
xor U5703 (N_5703,N_3567,N_2456);
or U5704 (N_5704,N_527,N_788);
and U5705 (N_5705,N_507,N_2996);
nand U5706 (N_5706,N_1401,N_4862);
and U5707 (N_5707,N_2847,N_3112);
nor U5708 (N_5708,N_4767,N_612);
xnor U5709 (N_5709,N_3591,N_1010);
xnor U5710 (N_5710,N_618,N_2003);
and U5711 (N_5711,N_4161,N_3367);
and U5712 (N_5712,N_3977,N_3697);
nand U5713 (N_5713,N_2797,N_4596);
or U5714 (N_5714,N_362,N_2581);
nand U5715 (N_5715,N_4364,N_2490);
xnor U5716 (N_5716,N_4871,N_1907);
and U5717 (N_5717,N_3268,N_1504);
and U5718 (N_5718,N_2460,N_2469);
xnor U5719 (N_5719,N_2918,N_3467);
and U5720 (N_5720,N_3745,N_555);
xor U5721 (N_5721,N_389,N_541);
or U5722 (N_5722,N_691,N_2049);
xor U5723 (N_5723,N_2472,N_3240);
nor U5724 (N_5724,N_547,N_904);
nor U5725 (N_5725,N_746,N_3378);
or U5726 (N_5726,N_351,N_3525);
nand U5727 (N_5727,N_3641,N_3156);
or U5728 (N_5728,N_1596,N_670);
nand U5729 (N_5729,N_1862,N_1518);
xor U5730 (N_5730,N_847,N_2667);
and U5731 (N_5731,N_766,N_3869);
and U5732 (N_5732,N_3936,N_4893);
or U5733 (N_5733,N_4919,N_3475);
xor U5734 (N_5734,N_576,N_3931);
or U5735 (N_5735,N_1820,N_3106);
xnor U5736 (N_5736,N_4781,N_655);
xnor U5737 (N_5737,N_3107,N_2948);
or U5738 (N_5738,N_4180,N_3853);
xnor U5739 (N_5739,N_2447,N_4995);
nor U5740 (N_5740,N_2780,N_3602);
and U5741 (N_5741,N_4586,N_2074);
or U5742 (N_5742,N_2343,N_4621);
nor U5743 (N_5743,N_4399,N_451);
xnor U5744 (N_5744,N_4831,N_306);
nor U5745 (N_5745,N_2825,N_4866);
nor U5746 (N_5746,N_1896,N_846);
nand U5747 (N_5747,N_110,N_4592);
nor U5748 (N_5748,N_4176,N_3968);
or U5749 (N_5749,N_3108,N_982);
nand U5750 (N_5750,N_476,N_4984);
or U5751 (N_5751,N_4163,N_521);
nand U5752 (N_5752,N_1137,N_3927);
nand U5753 (N_5753,N_2248,N_988);
and U5754 (N_5754,N_4128,N_358);
xnor U5755 (N_5755,N_2256,N_30);
or U5756 (N_5756,N_3371,N_1075);
or U5757 (N_5757,N_2442,N_3121);
nor U5758 (N_5758,N_4345,N_839);
nor U5759 (N_5759,N_3556,N_1338);
nor U5760 (N_5760,N_3490,N_2660);
and U5761 (N_5761,N_4950,N_3114);
and U5762 (N_5762,N_2123,N_523);
nand U5763 (N_5763,N_3206,N_3390);
and U5764 (N_5764,N_910,N_775);
or U5765 (N_5765,N_1738,N_3759);
xor U5766 (N_5766,N_1100,N_2779);
xor U5767 (N_5767,N_2110,N_3085);
or U5768 (N_5768,N_2915,N_1025);
nand U5769 (N_5769,N_2227,N_1395);
or U5770 (N_5770,N_4063,N_2743);
or U5771 (N_5771,N_4806,N_4559);
or U5772 (N_5772,N_4423,N_3975);
nor U5773 (N_5773,N_3185,N_2084);
or U5774 (N_5774,N_392,N_3747);
xnor U5775 (N_5775,N_3302,N_4644);
nand U5776 (N_5776,N_4020,N_4490);
nor U5777 (N_5777,N_1657,N_4464);
nor U5778 (N_5778,N_1092,N_4348);
and U5779 (N_5779,N_3335,N_3587);
and U5780 (N_5780,N_3312,N_644);
or U5781 (N_5781,N_3875,N_1348);
nor U5782 (N_5782,N_4007,N_2729);
nand U5783 (N_5783,N_1432,N_2975);
nor U5784 (N_5784,N_4946,N_2849);
nor U5785 (N_5785,N_4463,N_4385);
nor U5786 (N_5786,N_3348,N_3422);
or U5787 (N_5787,N_638,N_1840);
nand U5788 (N_5788,N_1604,N_4468);
nand U5789 (N_5789,N_2196,N_1070);
or U5790 (N_5790,N_3326,N_4484);
or U5791 (N_5791,N_772,N_872);
and U5792 (N_5792,N_3455,N_3812);
nor U5793 (N_5793,N_1944,N_4774);
nor U5794 (N_5794,N_2424,N_265);
nor U5795 (N_5795,N_1418,N_2396);
and U5796 (N_5796,N_4576,N_4772);
or U5797 (N_5797,N_993,N_3741);
nor U5798 (N_5798,N_809,N_3709);
nand U5799 (N_5799,N_835,N_80);
or U5800 (N_5800,N_2470,N_1084);
nand U5801 (N_5801,N_4948,N_3713);
nand U5802 (N_5802,N_1062,N_1233);
xor U5803 (N_5803,N_2258,N_4455);
xor U5804 (N_5804,N_2266,N_2557);
xor U5805 (N_5805,N_684,N_1941);
and U5806 (N_5806,N_787,N_324);
xnor U5807 (N_5807,N_4193,N_3794);
xor U5808 (N_5808,N_3495,N_911);
nor U5809 (N_5809,N_3714,N_1163);
nand U5810 (N_5810,N_959,N_376);
or U5811 (N_5811,N_551,N_4389);
and U5812 (N_5812,N_4819,N_3145);
nand U5813 (N_5813,N_2119,N_1488);
and U5814 (N_5814,N_4673,N_2741);
xor U5815 (N_5815,N_1244,N_689);
nor U5816 (N_5816,N_887,N_2169);
nor U5817 (N_5817,N_1351,N_238);
xnor U5818 (N_5818,N_2840,N_2909);
or U5819 (N_5819,N_3413,N_4979);
nor U5820 (N_5820,N_2244,N_4323);
xnor U5821 (N_5821,N_2673,N_4916);
nor U5822 (N_5822,N_1145,N_2118);
and U5823 (N_5823,N_2676,N_248);
and U5824 (N_5824,N_2597,N_849);
nor U5825 (N_5825,N_4421,N_3900);
or U5826 (N_5826,N_1858,N_4510);
nand U5827 (N_5827,N_3138,N_4045);
nand U5828 (N_5828,N_3191,N_947);
and U5829 (N_5829,N_632,N_3284);
nand U5830 (N_5830,N_723,N_4500);
nand U5831 (N_5831,N_1757,N_332);
nand U5832 (N_5832,N_1267,N_4933);
xor U5833 (N_5833,N_937,N_4970);
and U5834 (N_5834,N_2680,N_733);
and U5835 (N_5835,N_1945,N_1886);
nor U5836 (N_5836,N_4055,N_92);
or U5837 (N_5837,N_223,N_4891);
nand U5838 (N_5838,N_4843,N_1579);
and U5839 (N_5839,N_2412,N_2502);
and U5840 (N_5840,N_1713,N_1854);
nand U5841 (N_5841,N_3024,N_2482);
nor U5842 (N_5842,N_2768,N_1482);
xnor U5843 (N_5843,N_1053,N_142);
nand U5844 (N_5844,N_149,N_3244);
xnor U5845 (N_5845,N_951,N_2478);
nand U5846 (N_5846,N_3918,N_1496);
and U5847 (N_5847,N_4750,N_2955);
nor U5848 (N_5848,N_4150,N_4730);
nand U5849 (N_5849,N_703,N_1745);
or U5850 (N_5850,N_1174,N_3703);
nor U5851 (N_5851,N_1009,N_4174);
or U5852 (N_5852,N_4023,N_889);
xor U5853 (N_5853,N_1410,N_4091);
xnor U5854 (N_5854,N_1779,N_2089);
nand U5855 (N_5855,N_168,N_888);
and U5856 (N_5856,N_3950,N_4931);
and U5857 (N_5857,N_658,N_3397);
and U5858 (N_5858,N_1848,N_4346);
xor U5859 (N_5859,N_890,N_4870);
and U5860 (N_5860,N_2144,N_3764);
or U5861 (N_5861,N_4600,N_3449);
xnor U5862 (N_5862,N_4096,N_2744);
and U5863 (N_5863,N_188,N_545);
or U5864 (N_5864,N_1584,N_4664);
xor U5865 (N_5865,N_3233,N_1060);
and U5866 (N_5866,N_3286,N_1992);
xnor U5867 (N_5867,N_4046,N_3388);
and U5868 (N_5868,N_1571,N_2159);
nor U5869 (N_5869,N_586,N_1678);
and U5870 (N_5870,N_713,N_4103);
nand U5871 (N_5871,N_4286,N_3512);
and U5872 (N_5872,N_4824,N_3947);
nor U5873 (N_5873,N_1259,N_3198);
nor U5874 (N_5874,N_3898,N_2817);
and U5875 (N_5875,N_1780,N_3118);
nor U5876 (N_5876,N_4784,N_2560);
nand U5877 (N_5877,N_593,N_4937);
xnor U5878 (N_5878,N_3592,N_599);
nand U5879 (N_5879,N_3241,N_3694);
xor U5880 (N_5880,N_1148,N_3010);
and U5881 (N_5881,N_2457,N_1684);
nand U5882 (N_5882,N_500,N_3756);
or U5883 (N_5883,N_3894,N_55);
nand U5884 (N_5884,N_2212,N_3211);
or U5885 (N_5885,N_3630,N_2109);
nand U5886 (N_5886,N_1542,N_1650);
nand U5887 (N_5887,N_4685,N_4151);
xor U5888 (N_5888,N_1105,N_267);
nor U5889 (N_5889,N_329,N_4519);
nand U5890 (N_5890,N_2236,N_1098);
nand U5891 (N_5891,N_3026,N_226);
nand U5892 (N_5892,N_2635,N_1277);
xor U5893 (N_5893,N_3964,N_2246);
nand U5894 (N_5894,N_352,N_2668);
nor U5895 (N_5895,N_2643,N_3076);
xnor U5896 (N_5896,N_1416,N_4418);
nor U5897 (N_5897,N_4393,N_1330);
and U5898 (N_5898,N_806,N_4579);
and U5899 (N_5899,N_2625,N_2594);
nand U5900 (N_5900,N_2332,N_206);
nor U5901 (N_5901,N_3032,N_1928);
and U5902 (N_5902,N_2663,N_626);
nor U5903 (N_5903,N_1773,N_4031);
nor U5904 (N_5904,N_1324,N_3087);
and U5905 (N_5905,N_1749,N_422);
nand U5906 (N_5906,N_1308,N_4243);
nor U5907 (N_5907,N_4214,N_2674);
or U5908 (N_5908,N_2777,N_4002);
nand U5909 (N_5909,N_4635,N_3088);
nor U5910 (N_5910,N_71,N_4376);
nor U5911 (N_5911,N_1598,N_669);
or U5912 (N_5912,N_490,N_177);
or U5913 (N_5913,N_2484,N_489);
xnor U5914 (N_5914,N_291,N_1696);
nand U5915 (N_5915,N_679,N_2226);
xor U5916 (N_5916,N_3565,N_4797);
xor U5917 (N_5917,N_68,N_428);
and U5918 (N_5918,N_4524,N_1947);
and U5919 (N_5919,N_264,N_4815);
and U5920 (N_5920,N_2391,N_3446);
or U5921 (N_5921,N_3195,N_3332);
or U5922 (N_5922,N_1113,N_1605);
or U5923 (N_5923,N_3873,N_2913);
nor U5924 (N_5924,N_1880,N_4027);
nand U5925 (N_5925,N_368,N_711);
or U5926 (N_5926,N_1312,N_795);
and U5927 (N_5927,N_2066,N_899);
nor U5928 (N_5928,N_294,N_2990);
nor U5929 (N_5929,N_384,N_4556);
xnor U5930 (N_5930,N_26,N_533);
nor U5931 (N_5931,N_4816,N_3201);
or U5932 (N_5932,N_4093,N_1980);
nor U5933 (N_5933,N_2697,N_3478);
nor U5934 (N_5934,N_2395,N_14);
and U5935 (N_5935,N_261,N_2732);
nor U5936 (N_5936,N_4192,N_1368);
xnor U5937 (N_5937,N_1997,N_2008);
nor U5938 (N_5938,N_3618,N_434);
or U5939 (N_5939,N_2738,N_657);
nor U5940 (N_5940,N_2934,N_519);
xor U5941 (N_5941,N_2130,N_4472);
or U5942 (N_5942,N_685,N_2558);
xor U5943 (N_5943,N_2028,N_1128);
xor U5944 (N_5944,N_4678,N_2755);
and U5945 (N_5945,N_4662,N_197);
and U5946 (N_5946,N_1406,N_4164);
nand U5947 (N_5947,N_1054,N_1811);
nor U5948 (N_5948,N_2747,N_1117);
and U5949 (N_5949,N_3140,N_4758);
or U5950 (N_5950,N_582,N_3760);
and U5951 (N_5951,N_4840,N_4241);
nor U5952 (N_5952,N_3896,N_3995);
xor U5953 (N_5953,N_4451,N_2007);
nor U5954 (N_5954,N_2687,N_1883);
nand U5955 (N_5955,N_1512,N_3429);
nand U5956 (N_5956,N_2605,N_3040);
nand U5957 (N_5957,N_1238,N_1294);
nand U5958 (N_5958,N_4489,N_4909);
and U5959 (N_5959,N_4725,N_3450);
or U5960 (N_5960,N_3647,N_3949);
nor U5961 (N_5961,N_3944,N_3219);
or U5962 (N_5962,N_1321,N_3501);
nand U5963 (N_5963,N_1152,N_1894);
xnor U5964 (N_5964,N_2020,N_1963);
and U5965 (N_5965,N_1793,N_3127);
nor U5966 (N_5966,N_1912,N_757);
and U5967 (N_5967,N_4386,N_4953);
xnor U5968 (N_5968,N_619,N_4162);
nand U5969 (N_5969,N_2877,N_2308);
and U5970 (N_5970,N_4306,N_3932);
and U5971 (N_5971,N_4011,N_4648);
nor U5972 (N_5972,N_4646,N_796);
and U5973 (N_5973,N_755,N_864);
nor U5974 (N_5974,N_514,N_3430);
xor U5975 (N_5975,N_3225,N_1120);
nand U5976 (N_5976,N_4318,N_2263);
or U5977 (N_5977,N_4791,N_1086);
nor U5978 (N_5978,N_4179,N_160);
nor U5979 (N_5979,N_413,N_2017);
nor U5980 (N_5980,N_1279,N_3411);
or U5981 (N_5981,N_360,N_2155);
nor U5982 (N_5982,N_1964,N_2282);
and U5983 (N_5983,N_2039,N_1288);
nand U5984 (N_5984,N_1094,N_804);
or U5985 (N_5985,N_692,N_1703);
or U5986 (N_5986,N_520,N_3389);
and U5987 (N_5987,N_3769,N_3686);
and U5988 (N_5988,N_3657,N_2054);
nand U5989 (N_5989,N_1437,N_1833);
nand U5990 (N_5990,N_2441,N_4706);
xor U5991 (N_5991,N_1870,N_2341);
xor U5992 (N_5992,N_2971,N_3517);
nand U5993 (N_5993,N_1168,N_3474);
nor U5994 (N_5994,N_985,N_1146);
xor U5995 (N_5995,N_2417,N_2671);
or U5996 (N_5996,N_3825,N_1270);
and U5997 (N_5997,N_4591,N_1445);
nor U5998 (N_5998,N_3779,N_405);
xnor U5999 (N_5999,N_3074,N_2168);
nand U6000 (N_6000,N_2956,N_919);
nor U6001 (N_6001,N_2815,N_4833);
or U6002 (N_6002,N_89,N_2811);
or U6003 (N_6003,N_2126,N_536);
xor U6004 (N_6004,N_1902,N_4210);
nand U6005 (N_6005,N_4623,N_1943);
xnor U6006 (N_6006,N_1305,N_2073);
or U6007 (N_6007,N_3829,N_41);
xnor U6008 (N_6008,N_4427,N_1846);
and U6009 (N_6009,N_1965,N_4798);
nand U6010 (N_6010,N_4040,N_2985);
nor U6011 (N_6011,N_1219,N_1189);
and U6012 (N_6012,N_2739,N_1987);
or U6013 (N_6013,N_4349,N_4339);
and U6014 (N_6014,N_2632,N_4852);
nand U6015 (N_6015,N_4531,N_3619);
xnor U6016 (N_6016,N_693,N_4829);
or U6017 (N_6017,N_1436,N_2530);
and U6018 (N_6018,N_1166,N_1620);
nand U6019 (N_6019,N_1077,N_971);
or U6020 (N_6020,N_4473,N_2329);
nor U6021 (N_6021,N_1315,N_3484);
or U6022 (N_6022,N_3282,N_2352);
and U6023 (N_6023,N_906,N_2397);
or U6024 (N_6024,N_2211,N_2477);
nor U6025 (N_6025,N_2751,N_1349);
or U6026 (N_6026,N_1704,N_1177);
nand U6027 (N_6027,N_4508,N_4965);
xnor U6028 (N_6028,N_1530,N_4521);
xnor U6029 (N_6029,N_1414,N_1125);
xor U6030 (N_6030,N_3008,N_5);
nand U6031 (N_6031,N_1831,N_2314);
and U6032 (N_6032,N_1498,N_1469);
or U6033 (N_6033,N_3826,N_3881);
or U6034 (N_6034,N_882,N_1587);
nand U6035 (N_6035,N_2951,N_2772);
nand U6036 (N_6036,N_3129,N_3508);
nor U6037 (N_6037,N_257,N_245);
nor U6038 (N_6038,N_597,N_3006);
or U6039 (N_6039,N_4294,N_2464);
nand U6040 (N_6040,N_4649,N_1931);
xor U6041 (N_6041,N_2791,N_2494);
nor U6042 (N_6042,N_162,N_3970);
nand U6043 (N_6043,N_396,N_4982);
nand U6044 (N_6044,N_2434,N_415);
or U6045 (N_6045,N_3489,N_296);
or U6046 (N_6046,N_672,N_2416);
or U6047 (N_6047,N_2260,N_4853);
or U6048 (N_6048,N_4742,N_293);
xor U6049 (N_6049,N_671,N_4839);
xor U6050 (N_6050,N_3526,N_3650);
or U6051 (N_6051,N_2604,N_3773);
nand U6052 (N_6052,N_845,N_3083);
nand U6053 (N_6053,N_3547,N_1548);
nand U6054 (N_6054,N_3507,N_2862);
xor U6055 (N_6055,N_2835,N_66);
nand U6056 (N_6056,N_4543,N_1844);
nand U6057 (N_6057,N_2085,N_4242);
nor U6058 (N_6058,N_1005,N_4450);
nor U6059 (N_6059,N_4702,N_172);
nor U6060 (N_6060,N_1789,N_2069);
nand U6061 (N_6061,N_4329,N_767);
nand U6062 (N_6062,N_829,N_3270);
nor U6063 (N_6063,N_4565,N_3972);
nand U6064 (N_6064,N_1645,N_4590);
xor U6065 (N_6065,N_3346,N_1249);
nor U6066 (N_6066,N_3033,N_2608);
or U6067 (N_6067,N_4197,N_2031);
xor U6068 (N_6068,N_2105,N_2931);
nor U6069 (N_6069,N_2374,N_35);
or U6070 (N_6070,N_3120,N_724);
nor U6071 (N_6071,N_631,N_3634);
nand U6072 (N_6072,N_1589,N_1197);
or U6073 (N_6073,N_4526,N_3101);
xnor U6074 (N_6074,N_496,N_2242);
nand U6075 (N_6075,N_3424,N_1879);
nand U6076 (N_6076,N_1528,N_1261);
xor U6077 (N_6077,N_2510,N_853);
nand U6078 (N_6078,N_1394,N_2612);
and U6079 (N_6079,N_2754,N_3229);
and U6080 (N_6080,N_2509,N_2381);
and U6081 (N_6081,N_881,N_77);
and U6082 (N_6082,N_1676,N_1116);
or U6083 (N_6083,N_1783,N_871);
xor U6084 (N_6084,N_3016,N_4426);
and U6085 (N_6085,N_4884,N_143);
xnor U6086 (N_6086,N_4601,N_666);
xor U6087 (N_6087,N_2377,N_2075);
xor U6088 (N_6088,N_1576,N_363);
xor U6089 (N_6089,N_4102,N_1795);
or U6090 (N_6090,N_727,N_1666);
nor U6091 (N_6091,N_166,N_1734);
or U6092 (N_6092,N_2543,N_3420);
nor U6093 (N_6093,N_1404,N_3089);
nor U6094 (N_6094,N_4818,N_3679);
nor U6095 (N_6095,N_4413,N_4691);
xor U6096 (N_6096,N_1547,N_744);
and U6097 (N_6097,N_4217,N_4328);
nor U6098 (N_6098,N_817,N_1946);
nand U6099 (N_6099,N_2529,N_409);
or U6100 (N_6100,N_4205,N_3194);
nor U6101 (N_6101,N_3693,N_1222);
and U6102 (N_6102,N_2491,N_3246);
and U6103 (N_6103,N_4684,N_208);
nor U6104 (N_6104,N_17,N_4278);
nand U6105 (N_6105,N_3786,N_3935);
xor U6106 (N_6106,N_1127,N_4487);
and U6107 (N_6107,N_3571,N_3943);
nand U6108 (N_6108,N_4896,N_316);
or U6109 (N_6109,N_3323,N_246);
and U6110 (N_6110,N_1729,N_1808);
nor U6111 (N_6111,N_4111,N_2430);
or U6112 (N_6112,N_2492,N_1849);
xor U6113 (N_6113,N_1299,N_3394);
xnor U6114 (N_6114,N_3164,N_217);
and U6115 (N_6115,N_3414,N_1553);
or U6116 (N_6116,N_1890,N_676);
nand U6117 (N_6117,N_1263,N_1827);
or U6118 (N_6118,N_617,N_1639);
or U6119 (N_6119,N_3891,N_171);
xor U6120 (N_6120,N_518,N_3251);
nand U6121 (N_6121,N_2790,N_1342);
nand U6122 (N_6122,N_764,N_2905);
or U6123 (N_6123,N_2883,N_474);
nand U6124 (N_6124,N_1850,N_1888);
nor U6125 (N_6125,N_2945,N_1660);
nand U6126 (N_6126,N_3637,N_1919);
or U6127 (N_6127,N_4149,N_1552);
xnor U6128 (N_6128,N_3183,N_1694);
or U6129 (N_6129,N_4269,N_1362);
nor U6130 (N_6130,N_3204,N_577);
xnor U6131 (N_6131,N_2157,N_1289);
nor U6132 (N_6132,N_133,N_2024);
nor U6133 (N_6133,N_2136,N_3137);
or U6134 (N_6134,N_2823,N_2873);
nand U6135 (N_6135,N_1741,N_592);
xor U6136 (N_6136,N_3459,N_572);
and U6137 (N_6137,N_2415,N_737);
nand U6138 (N_6138,N_3529,N_580);
nor U6139 (N_6139,N_3263,N_1523);
nand U6140 (N_6140,N_4672,N_397);
or U6141 (N_6141,N_3181,N_3758);
and U6142 (N_6142,N_1884,N_2120);
xor U6143 (N_6143,N_3147,N_1753);
xnor U6144 (N_6144,N_819,N_4332);
or U6145 (N_6145,N_3652,N_2108);
and U6146 (N_6146,N_747,N_2574);
nor U6147 (N_6147,N_4913,N_3344);
xnor U6148 (N_6148,N_4790,N_3646);
and U6149 (N_6149,N_1843,N_4114);
nand U6150 (N_6150,N_1142,N_3831);
xor U6151 (N_6151,N_463,N_2949);
nor U6152 (N_6152,N_3734,N_2201);
and U6153 (N_6153,N_290,N_4325);
and U6154 (N_6154,N_879,N_716);
or U6155 (N_6155,N_1046,N_920);
or U6156 (N_6156,N_3514,N_921);
nor U6157 (N_6157,N_3003,N_1797);
or U6158 (N_6158,N_3994,N_427);
nand U6159 (N_6159,N_4380,N_1921);
nand U6160 (N_6160,N_2776,N_1225);
and U6161 (N_6161,N_2129,N_3945);
nand U6162 (N_6162,N_762,N_2709);
and U6163 (N_6163,N_2615,N_2659);
nor U6164 (N_6164,N_1712,N_1900);
nor U6165 (N_6165,N_4402,N_3642);
xnor U6166 (N_6166,N_4206,N_1613);
nand U6167 (N_6167,N_4216,N_4049);
nor U6168 (N_6168,N_1865,N_1895);
nor U6169 (N_6169,N_3509,N_2223);
xnor U6170 (N_6170,N_1276,N_2735);
nor U6171 (N_6171,N_1191,N_1438);
nand U6172 (N_6172,N_2102,N_2593);
nor U6173 (N_6173,N_3767,N_499);
xnor U6174 (N_6174,N_1706,N_472);
and U6175 (N_6175,N_1638,N_4075);
nor U6176 (N_6176,N_504,N_1255);
or U6177 (N_6177,N_4888,N_4934);
and U6178 (N_6178,N_4353,N_4352);
or U6179 (N_6179,N_4297,N_941);
and U6180 (N_6180,N_3557,N_2692);
and U6181 (N_6181,N_4068,N_2927);
and U6182 (N_6182,N_2536,N_1769);
xor U6183 (N_6183,N_2864,N_218);
and U6184 (N_6184,N_4626,N_1698);
nor U6185 (N_6185,N_4228,N_179);
nand U6186 (N_6186,N_3352,N_163);
nor U6187 (N_6187,N_10,N_95);
xnor U6188 (N_6188,N_2288,N_3060);
nor U6189 (N_6189,N_4085,N_2400);
and U6190 (N_6190,N_250,N_4457);
nand U6191 (N_6191,N_2954,N_2952);
xnor U6192 (N_6192,N_278,N_4887);
and U6193 (N_6193,N_2132,N_22);
nand U6194 (N_6194,N_2234,N_1918);
or U6195 (N_6195,N_557,N_1524);
and U6196 (N_6196,N_1050,N_2977);
nand U6197 (N_6197,N_659,N_3055);
or U6198 (N_6198,N_3965,N_2174);
xnor U6199 (N_6199,N_1354,N_2933);
or U6200 (N_6200,N_2205,N_4334);
xnor U6201 (N_6201,N_2495,N_3271);
and U6202 (N_6202,N_750,N_1663);
nor U6203 (N_6203,N_3441,N_4170);
nand U6204 (N_6204,N_3699,N_4740);
or U6205 (N_6205,N_721,N_3732);
xnor U6206 (N_6206,N_192,N_4698);
or U6207 (N_6207,N_1178,N_2926);
or U6208 (N_6208,N_776,N_2068);
and U6209 (N_6209,N_1181,N_1199);
nand U6210 (N_6210,N_1697,N_2322);
xnor U6211 (N_6211,N_2540,N_945);
nand U6212 (N_6212,N_2488,N_1767);
nor U6213 (N_6213,N_510,N_3570);
nand U6214 (N_6214,N_4240,N_4090);
xor U6215 (N_6215,N_3586,N_1449);
or U6216 (N_6216,N_2095,N_857);
or U6217 (N_6217,N_2125,N_4223);
and U6218 (N_6218,N_4012,N_1532);
nor U6219 (N_6219,N_4073,N_3499);
nand U6220 (N_6220,N_1905,N_3214);
or U6221 (N_6221,N_97,N_1510);
or U6222 (N_6222,N_91,N_4647);
nand U6223 (N_6223,N_2336,N_3116);
nor U6224 (N_6224,N_1701,N_3496);
nor U6225 (N_6225,N_2999,N_2023);
nand U6226 (N_6226,N_2762,N_2101);
or U6227 (N_6227,N_3285,N_3636);
and U6228 (N_6228,N_4018,N_1859);
nor U6229 (N_6229,N_457,N_4453);
nor U6230 (N_6230,N_1157,N_1370);
xor U6231 (N_6231,N_227,N_2222);
xnor U6232 (N_6232,N_3457,N_2220);
nor U6233 (N_6233,N_955,N_4388);
nand U6234 (N_6234,N_3800,N_435);
xor U6235 (N_6235,N_2737,N_63);
xor U6236 (N_6236,N_1387,N_3628);
nand U6237 (N_6237,N_4194,N_2081);
nand U6238 (N_6238,N_4222,N_1008);
nor U6239 (N_6239,N_3851,N_2261);
and U6240 (N_6240,N_1340,N_207);
nor U6241 (N_6241,N_3648,N_607);
nand U6242 (N_6242,N_3377,N_525);
and U6243 (N_6243,N_201,N_4004);
and U6244 (N_6244,N_4175,N_334);
and U6245 (N_6245,N_4437,N_438);
nor U6246 (N_6246,N_3431,N_3890);
or U6247 (N_6247,N_2708,N_4391);
and U6248 (N_6248,N_1962,N_3762);
nor U6249 (N_6249,N_2590,N_109);
nand U6250 (N_6250,N_1821,N_1534);
xnor U6251 (N_6251,N_241,N_1304);
nor U6252 (N_6252,N_901,N_4267);
nand U6253 (N_6253,N_2742,N_116);
nand U6254 (N_6254,N_2225,N_4370);
or U6255 (N_6255,N_4541,N_4780);
nand U6256 (N_6256,N_1027,N_3303);
xnor U6257 (N_6257,N_4232,N_1719);
nor U6258 (N_6258,N_49,N_4536);
nor U6259 (N_6259,N_4666,N_3711);
xor U6260 (N_6260,N_3134,N_366);
or U6261 (N_6261,N_83,N_2380);
nand U6262 (N_6262,N_1223,N_2454);
and U6263 (N_6263,N_4985,N_517);
xnor U6264 (N_6264,N_1231,N_4183);
or U6265 (N_6265,N_3669,N_3069);
xnor U6266 (N_6266,N_725,N_3828);
nand U6267 (N_6267,N_1275,N_228);
xnor U6268 (N_6268,N_656,N_2056);
nor U6269 (N_6269,N_349,N_3309);
xor U6270 (N_6270,N_1093,N_1129);
and U6271 (N_6271,N_4494,N_863);
nor U6272 (N_6272,N_2147,N_1647);
nor U6273 (N_6273,N_4112,N_3907);
xnor U6274 (N_6274,N_4436,N_3387);
and U6275 (N_6275,N_4895,N_3169);
xnor U6276 (N_6276,N_1937,N_3019);
nor U6277 (N_6277,N_3184,N_3269);
and U6278 (N_6278,N_2972,N_276);
and U6279 (N_6279,N_2217,N_2513);
nand U6280 (N_6280,N_1390,N_2524);
or U6281 (N_6281,N_1450,N_1558);
xnor U6282 (N_6282,N_3691,N_1355);
nand U6283 (N_6283,N_537,N_4966);
nand U6284 (N_6284,N_1838,N_2338);
nand U6285 (N_6285,N_3421,N_3361);
and U6286 (N_6286,N_3056,N_668);
or U6287 (N_6287,N_2740,N_180);
nand U6288 (N_6288,N_630,N_1384);
or U6289 (N_6289,N_3028,N_2325);
or U6290 (N_6290,N_11,N_678);
or U6291 (N_6291,N_33,N_99);
nor U6292 (N_6292,N_1874,N_2115);
nor U6293 (N_6293,N_1076,N_3439);
and U6294 (N_6294,N_3768,N_4535);
xor U6295 (N_6295,N_1337,N_2922);
nor U6296 (N_6296,N_1538,N_2592);
xor U6297 (N_6297,N_3601,N_995);
nand U6298 (N_6298,N_1617,N_2385);
xor U6299 (N_6299,N_2467,N_2479);
xor U6300 (N_6300,N_4377,N_253);
nor U6301 (N_6301,N_2326,N_1176);
xor U6302 (N_6302,N_2521,N_2080);
or U6303 (N_6303,N_395,N_1746);
and U6304 (N_6304,N_1033,N_146);
or U6305 (N_6305,N_4991,N_1982);
nand U6306 (N_6306,N_4744,N_2294);
nand U6307 (N_6307,N_1561,N_3456);
nor U6308 (N_6308,N_3031,N_2036);
or U6309 (N_6309,N_2916,N_4397);
and U6310 (N_6310,N_485,N_3415);
and U6311 (N_6311,N_4680,N_2619);
and U6312 (N_6312,N_2082,N_3383);
xor U6313 (N_6313,N_4299,N_2941);
nor U6314 (N_6314,N_1444,N_2162);
nor U6315 (N_6315,N_660,N_2367);
xor U6316 (N_6316,N_720,N_4873);
or U6317 (N_6317,N_401,N_2525);
xnor U6318 (N_6318,N_4779,N_640);
and U6319 (N_6319,N_3119,N_1508);
and U6320 (N_6320,N_926,N_873);
or U6321 (N_6321,N_300,N_2087);
nand U6322 (N_6322,N_387,N_4148);
nand U6323 (N_6323,N_4041,N_3428);
xnor U6324 (N_6324,N_1642,N_165);
xnor U6325 (N_6325,N_2281,N_1201);
nor U6326 (N_6326,N_2853,N_4554);
xor U6327 (N_6327,N_3186,N_4796);
nor U6328 (N_6328,N_589,N_4805);
or U6329 (N_6329,N_1236,N_4144);
and U6330 (N_6330,N_4838,N_2566);
or U6331 (N_6331,N_1118,N_2269);
or U6332 (N_6332,N_1024,N_1904);
nor U6333 (N_6333,N_3097,N_4177);
nand U6334 (N_6334,N_3046,N_4447);
nand U6335 (N_6335,N_3820,N_1814);
nor U6336 (N_6336,N_4407,N_4344);
or U6337 (N_6337,N_2356,N_3583);
nand U6338 (N_6338,N_2438,N_3897);
and U6339 (N_6339,N_4518,N_628);
xor U6340 (N_6340,N_436,N_1618);
nor U6341 (N_6341,N_1646,N_233);
or U6342 (N_6342,N_1957,N_3798);
nand U6343 (N_6343,N_2911,N_3982);
and U6344 (N_6344,N_3154,N_4545);
xnor U6345 (N_6345,N_1491,N_1852);
xor U6346 (N_6346,N_461,N_4293);
or U6347 (N_6347,N_2360,N_714);
or U6348 (N_6348,N_749,N_1936);
or U6349 (N_6349,N_1102,N_211);
nand U6350 (N_6350,N_742,N_4527);
nor U6351 (N_6351,N_319,N_3551);
and U6352 (N_6352,N_967,N_1954);
xnor U6353 (N_6353,N_106,N_2607);
or U6354 (N_6354,N_1018,N_473);
and U6355 (N_6355,N_4921,N_1206);
xor U6356 (N_6356,N_4440,N_3576);
nor U6357 (N_6357,N_3817,N_4904);
and U6358 (N_6358,N_2474,N_935);
xnor U6359 (N_6359,N_538,N_1439);
and U6360 (N_6360,N_962,N_2070);
nor U6361 (N_6361,N_1066,N_4358);
or U6362 (N_6362,N_1021,N_2450);
nand U6363 (N_6363,N_505,N_4842);
xor U6364 (N_6364,N_554,N_929);
nor U6365 (N_6365,N_4283,N_431);
xnor U6366 (N_6366,N_3797,N_961);
nand U6367 (N_6367,N_2821,N_782);
or U6368 (N_6368,N_3045,N_3427);
or U6369 (N_6369,N_3239,N_1121);
nor U6370 (N_6370,N_2679,N_515);
xnor U6371 (N_6371,N_928,N_4066);
and U6372 (N_6372,N_568,N_190);
and U6373 (N_6373,N_4687,N_2285);
nor U6374 (N_6374,N_4514,N_4327);
xor U6375 (N_6375,N_3688,N_423);
xor U6376 (N_6376,N_2133,N_2122);
xnor U6377 (N_6377,N_661,N_2346);
xnor U6378 (N_6378,N_4265,N_4022);
and U6379 (N_6379,N_1373,N_2920);
nor U6380 (N_6380,N_4849,N_2178);
nand U6381 (N_6381,N_2190,N_4968);
and U6382 (N_6382,N_1483,N_1476);
xor U6383 (N_6383,N_3267,N_347);
nor U6384 (N_6384,N_2662,N_54);
nor U6385 (N_6385,N_4501,N_1126);
or U6386 (N_6386,N_2354,N_3568);
and U6387 (N_6387,N_1540,N_3940);
and U6388 (N_6388,N_2270,N_3372);
and U6389 (N_6389,N_4877,N_4259);
nor U6390 (N_6390,N_3575,N_2942);
nor U6391 (N_6391,N_2403,N_4857);
and U6392 (N_6392,N_3039,N_2067);
and U6393 (N_6393,N_182,N_4800);
nor U6394 (N_6394,N_3933,N_4537);
xor U6395 (N_6395,N_381,N_3200);
or U6396 (N_6396,N_1122,N_2773);
xnor U6397 (N_6397,N_7,N_2785);
xor U6398 (N_6398,N_2953,N_2677);
and U6399 (N_6399,N_4178,N_2820);
or U6400 (N_6400,N_1170,N_548);
xor U6401 (N_6401,N_4832,N_4660);
xor U6402 (N_6402,N_1457,N_1572);
or U6403 (N_6403,N_4371,N_3090);
and U6404 (N_6404,N_2181,N_446);
and U6405 (N_6405,N_1969,N_3168);
xnor U6406 (N_6406,N_3730,N_2855);
nand U6407 (N_6407,N_2189,N_2962);
and U6408 (N_6408,N_2871,N_4638);
nor U6409 (N_6409,N_270,N_3535);
nand U6410 (N_6410,N_3293,N_1788);
xor U6411 (N_6411,N_1509,N_1739);
or U6412 (N_6412,N_3986,N_304);
and U6413 (N_6413,N_2584,N_2138);
nor U6414 (N_6414,N_4285,N_3015);
or U6415 (N_6415,N_2019,N_2032);
xnor U6416 (N_6416,N_4065,N_556);
or U6417 (N_6417,N_4304,N_1020);
xor U6418 (N_6418,N_793,N_1887);
and U6419 (N_6419,N_4634,N_4593);
nor U6420 (N_6420,N_131,N_4699);
xnor U6421 (N_6421,N_128,N_3393);
nor U6422 (N_6422,N_1961,N_1459);
nor U6423 (N_6423,N_1802,N_4187);
and U6424 (N_6424,N_2339,N_1693);
nand U6425 (N_6425,N_2850,N_4978);
nor U6426 (N_6426,N_1556,N_2539);
or U6427 (N_6427,N_2386,N_3761);
and U6428 (N_6428,N_768,N_2298);
xor U6429 (N_6429,N_1072,N_2810);
and U6430 (N_6430,N_354,N_3533);
nor U6431 (N_6431,N_2004,N_210);
or U6432 (N_6432,N_4081,N_3892);
nor U6433 (N_6433,N_1055,N_4147);
or U6434 (N_6434,N_3645,N_4181);
xor U6435 (N_6435,N_2749,N_1644);
xnor U6436 (N_6436,N_838,N_1217);
xor U6437 (N_6437,N_3510,N_305);
and U6438 (N_6438,N_503,N_4301);
xor U6439 (N_6439,N_4770,N_4039);
and U6440 (N_6440,N_2551,N_2303);
and U6441 (N_6441,N_3400,N_550);
nor U6442 (N_6442,N_513,N_1740);
nor U6443 (N_6443,N_3708,N_372);
nor U6444 (N_6444,N_4974,N_1626);
or U6445 (N_6445,N_893,N_2228);
and U6446 (N_6446,N_2444,N_3141);
or U6447 (N_6447,N_2207,N_3771);
and U6448 (N_6448,N_1758,N_4903);
xor U6449 (N_6449,N_3453,N_3153);
nor U6450 (N_6450,N_634,N_585);
nor U6451 (N_6451,N_2473,N_2656);
or U6452 (N_6452,N_3351,N_3479);
nor U6453 (N_6453,N_3275,N_3914);
or U6454 (N_6454,N_4190,N_3785);
xnor U6455 (N_6455,N_3276,N_4858);
nand U6456 (N_6456,N_2595,N_629);
and U6457 (N_6457,N_1845,N_1930);
nor U6458 (N_6458,N_2276,N_2305);
and U6459 (N_6459,N_1983,N_2859);
nand U6460 (N_6460,N_4171,N_4539);
nor U6461 (N_6461,N_606,N_4263);
xnor U6462 (N_6462,N_3611,N_2553);
nor U6463 (N_6463,N_2127,N_4765);
and U6464 (N_6464,N_2943,N_3472);
and U6465 (N_6465,N_1164,N_2633);
nand U6466 (N_6466,N_1569,N_821);
nor U6467 (N_6467,N_1085,N_2649);
xnor U6468 (N_6468,N_3833,N_4628);
and U6469 (N_6469,N_3573,N_3683);
or U6470 (N_6470,N_2156,N_4123);
and U6471 (N_6471,N_3705,N_2792);
xor U6472 (N_6472,N_832,N_3663);
and U6473 (N_6473,N_4195,N_2705);
and U6474 (N_6474,N_2896,N_3197);
or U6475 (N_6475,N_313,N_602);
nand U6476 (N_6476,N_2323,N_4509);
or U6477 (N_6477,N_3294,N_2440);
nor U6478 (N_6478,N_2499,N_2746);
xnor U6479 (N_6479,N_651,N_696);
and U6480 (N_6480,N_342,N_1830);
xor U6481 (N_6481,N_2150,N_2398);
nor U6482 (N_6482,N_380,N_3763);
nor U6483 (N_6483,N_3774,N_3976);
nand U6484 (N_6484,N_3816,N_2504);
nor U6485 (N_6485,N_3030,N_2874);
nand U6486 (N_6486,N_1229,N_4374);
or U6487 (N_6487,N_798,N_516);
and U6488 (N_6488,N_4885,N_3803);
or U6489 (N_6489,N_365,N_2982);
or U6490 (N_6490,N_748,N_2267);
nand U6491 (N_6491,N_1096,N_174);
nor U6492 (N_6492,N_4710,N_1052);
or U6493 (N_6493,N_1868,N_70);
xnor U6494 (N_6494,N_3993,N_3555);
or U6495 (N_6495,N_3885,N_1923);
or U6496 (N_6496,N_4572,N_221);
nand U6497 (N_6497,N_462,N_4723);
nand U6498 (N_6498,N_3260,N_2839);
nand U6499 (N_6499,N_534,N_2252);
or U6500 (N_6500,N_491,N_338);
xnor U6501 (N_6501,N_1521,N_286);
or U6502 (N_6502,N_284,N_3506);
nor U6503 (N_6503,N_3610,N_2798);
and U6504 (N_6504,N_4731,N_855);
nor U6505 (N_6505,N_58,N_2436);
nand U6506 (N_6506,N_2571,N_972);
nand U6507 (N_6507,N_2078,N_1290);
nand U6508 (N_6508,N_646,N_4078);
or U6509 (N_6509,N_974,N_1913);
nor U6510 (N_6510,N_624,N_1185);
and U6511 (N_6511,N_3676,N_3196);
xnor U6512 (N_6512,N_3864,N_4341);
or U6513 (N_6513,N_843,N_3297);
nand U6514 (N_6514,N_4599,N_917);
nand U6515 (N_6515,N_2694,N_3174);
and U6516 (N_6516,N_3804,N_3477);
or U6517 (N_6517,N_2383,N_699);
nand U6518 (N_6518,N_449,N_683);
and U6519 (N_6519,N_4996,N_3480);
xor U6520 (N_6520,N_4015,N_3599);
nand U6521 (N_6521,N_3633,N_4883);
nor U6522 (N_6522,N_1608,N_2903);
nor U6523 (N_6523,N_2631,N_688);
and U6524 (N_6524,N_4443,N_2570);
or U6525 (N_6525,N_2875,N_818);
or U6526 (N_6526,N_1065,N_1392);
xnor U6527 (N_6527,N_2235,N_2421);
nand U6528 (N_6528,N_2655,N_2061);
xnor U6529 (N_6529,N_987,N_4189);
nor U6530 (N_6530,N_4714,N_726);
nand U6531 (N_6531,N_1511,N_4836);
nand U6532 (N_6532,N_1487,N_3962);
or U6533 (N_6533,N_754,N_2011);
and U6534 (N_6534,N_2901,N_4947);
xor U6535 (N_6535,N_4047,N_4428);
and U6536 (N_6536,N_1082,N_3905);
nand U6537 (N_6537,N_2413,N_3075);
xnor U6538 (N_6538,N_1908,N_2158);
or U6539 (N_6539,N_4578,N_2363);
nor U6540 (N_6540,N_2904,N_1634);
and U6541 (N_6541,N_1341,N_4048);
nor U6542 (N_6542,N_1135,N_1319);
nand U6543 (N_6543,N_923,N_3889);
nand U6544 (N_6544,N_3236,N_2878);
and U6545 (N_6545,N_2546,N_3886);
nand U6546 (N_6546,N_2221,N_4466);
or U6547 (N_6547,N_2994,N_1281);
nor U6548 (N_6548,N_4135,N_4080);
nor U6549 (N_6549,N_3744,N_3929);
nor U6550 (N_6550,N_2658,N_3262);
nor U6551 (N_6551,N_4503,N_2734);
nor U6552 (N_6552,N_215,N_3203);
or U6553 (N_6553,N_3177,N_90);
xor U6554 (N_6554,N_2523,N_4938);
nor U6555 (N_6555,N_642,N_4082);
and U6556 (N_6556,N_2555,N_4070);
nor U6557 (N_6557,N_571,N_4867);
nor U6558 (N_6558,N_934,N_4404);
nand U6559 (N_6559,N_4258,N_3359);
and U6560 (N_6560,N_1172,N_4060);
nand U6561 (N_6561,N_4467,N_2114);
or U6562 (N_6562,N_4620,N_321);
and U6563 (N_6563,N_2179,N_3093);
nor U6564 (N_6564,N_151,N_2715);
xnor U6565 (N_6565,N_878,N_1486);
xor U6566 (N_6566,N_2219,N_2698);
and U6567 (N_6567,N_539,N_3238);
nand U6568 (N_6568,N_1744,N_2533);
or U6569 (N_6569,N_3444,N_4905);
and U6570 (N_6570,N_3909,N_3368);
or U6571 (N_6571,N_3148,N_3715);
and U6572 (N_6572,N_2833,N_2568);
nor U6573 (N_6573,N_4681,N_1835);
or U6574 (N_6574,N_4548,N_1461);
xor U6575 (N_6575,N_4296,N_1673);
nor U6576 (N_6576,N_2277,N_464);
or U6577 (N_6577,N_4753,N_4033);
and U6578 (N_6578,N_1674,N_2932);
xor U6579 (N_6579,N_4782,N_875);
and U6580 (N_6580,N_3052,N_2516);
or U6581 (N_6581,N_4502,N_1332);
or U6582 (N_6582,N_918,N_2906);
nor U6583 (N_6583,N_4653,N_4749);
nand U6584 (N_6584,N_3539,N_1577);
xnor U6585 (N_6585,N_289,N_2194);
or U6586 (N_6586,N_885,N_4773);
and U6587 (N_6587,N_3674,N_3231);
xor U6588 (N_6588,N_1282,N_2646);
xor U6589 (N_6589,N_964,N_3253);
or U6590 (N_6590,N_154,N_4314);
nand U6591 (N_6591,N_1451,N_2801);
nand U6592 (N_6592,N_4617,N_970);
nand U6593 (N_6593,N_3901,N_1750);
or U6594 (N_6594,N_2103,N_856);
or U6595 (N_6595,N_1535,N_4594);
nand U6596 (N_6596,N_3466,N_3481);
and U6597 (N_6597,N_2370,N_4287);
nand U6598 (N_6598,N_1155,N_2548);
nand U6599 (N_6599,N_3678,N_2366);
xnor U6600 (N_6600,N_2844,N_3524);
nand U6601 (N_6601,N_2371,N_4255);
nand U6602 (N_6602,N_1240,N_3902);
xnor U6603 (N_6603,N_2485,N_710);
or U6604 (N_6604,N_1035,N_3572);
nand U6605 (N_6605,N_2250,N_4553);
and U6606 (N_6606,N_4522,N_3607);
nand U6607 (N_6607,N_205,N_2641);
nor U6608 (N_6608,N_3912,N_4881);
nor U6609 (N_6609,N_1565,N_2828);
and U6610 (N_6610,N_3144,N_2935);
nand U6611 (N_6611,N_4642,N_978);
nand U6612 (N_6612,N_4993,N_2293);
xnor U6613 (N_6613,N_759,N_665);
nor U6614 (N_6614,N_3941,N_4532);
and U6615 (N_6615,N_2758,N_2736);
and U6616 (N_6616,N_3125,N_4101);
xor U6617 (N_6617,N_13,N_4037);
xor U6618 (N_6618,N_136,N_3497);
nand U6619 (N_6619,N_2335,N_2029);
and U6620 (N_6620,N_330,N_475);
or U6621 (N_6621,N_3396,N_1763);
nand U6622 (N_6622,N_675,N_187);
or U6623 (N_6623,N_2213,N_2958);
or U6624 (N_6624,N_4184,N_2320);
nor U6625 (N_6625,N_3038,N_4827);
nor U6626 (N_6626,N_1130,N_3374);
nor U6627 (N_6627,N_3857,N_4726);
nand U6628 (N_6628,N_4409,N_1361);
nor U6629 (N_6629,N_1711,N_1889);
and U6630 (N_6630,N_3465,N_3325);
xnor U6631 (N_6631,N_4964,N_139);
nand U6632 (N_6632,N_2184,N_4612);
nor U6633 (N_6633,N_25,N_85);
xor U6634 (N_6634,N_269,N_1371);
xnor U6635 (N_6635,N_3574,N_741);
nand U6636 (N_6636,N_3815,N_1182);
and U6637 (N_6637,N_1968,N_394);
nand U6638 (N_6638,N_3721,N_1580);
xnor U6639 (N_6639,N_4868,N_3210);
and U6640 (N_6640,N_50,N_3395);
nand U6641 (N_6641,N_936,N_4952);
xnor U6642 (N_6642,N_4633,N_2304);
nor U6643 (N_6643,N_996,N_650);
nand U6644 (N_6644,N_2393,N_1971);
and U6645 (N_6645,N_735,N_353);
nand U6646 (N_6646,N_3110,N_488);
nand U6647 (N_6647,N_3409,N_1473);
nand U6648 (N_6648,N_1622,N_2778);
or U6649 (N_6649,N_4751,N_4807);
xnor U6650 (N_6650,N_1754,N_4410);
nor U6651 (N_6651,N_126,N_3655);
nor U6652 (N_6652,N_4446,N_760);
nor U6653 (N_6653,N_3213,N_4444);
nor U6654 (N_6654,N_4640,N_1988);
nor U6655 (N_6655,N_117,N_1344);
or U6656 (N_6656,N_1546,N_4244);
or U6657 (N_6657,N_3362,N_2767);
xnor U6658 (N_6658,N_2265,N_4319);
nand U6659 (N_6659,N_4605,N_3054);
nor U6660 (N_6660,N_2198,N_4811);
nand U6661 (N_6661,N_345,N_4173);
and U6662 (N_6662,N_4250,N_1659);
nor U6663 (N_6663,N_1562,N_1280);
and U6664 (N_6664,N_2508,N_4284);
and U6665 (N_6665,N_382,N_411);
xor U6666 (N_6666,N_850,N_1942);
or U6667 (N_6667,N_1226,N_1293);
and U6668 (N_6668,N_3819,N_1585);
nand U6669 (N_6669,N_1689,N_195);
nor U6670 (N_6670,N_1692,N_178);
nand U6671 (N_6671,N_1658,N_1737);
and U6672 (N_6672,N_4716,N_410);
nor U6673 (N_6673,N_2703,N_2814);
or U6674 (N_6674,N_2688,N_4911);
or U6675 (N_6675,N_3516,N_4462);
or U6676 (N_6676,N_1839,N_717);
nor U6677 (N_6677,N_4990,N_4752);
xor U6678 (N_6678,N_3540,N_2010);
nand U6679 (N_6679,N_4908,N_3860);
nor U6680 (N_6680,N_3333,N_232);
nand U6681 (N_6681,N_2585,N_108);
xnor U6682 (N_6682,N_336,N_4812);
xnor U6683 (N_6683,N_298,N_4655);
and U6684 (N_6684,N_3856,N_4273);
xnor U6685 (N_6685,N_2579,N_1316);
xnor U6686 (N_6686,N_101,N_2527);
nor U6687 (N_6687,N_1616,N_3934);
and U6688 (N_6688,N_4036,N_2989);
nor U6689 (N_6689,N_138,N_805);
and U6690 (N_6690,N_4369,N_986);
and U6691 (N_6691,N_2589,N_147);
or U6692 (N_6692,N_2756,N_3685);
nor U6693 (N_6693,N_3438,N_1393);
and U6694 (N_6694,N_1101,N_3700);
nor U6695 (N_6695,N_543,N_1039);
nand U6696 (N_6696,N_4546,N_12);
xnor U6697 (N_6697,N_2728,N_907);
and U6698 (N_6698,N_1378,N_2331);
nor U6699 (N_6699,N_1977,N_2610);
and U6700 (N_6700,N_2245,N_198);
and U6701 (N_6701,N_1825,N_4734);
nor U6702 (N_6702,N_3220,N_801);
xnor U6703 (N_6703,N_155,N_983);
or U6704 (N_6704,N_4254,N_4231);
nand U6705 (N_6705,N_4449,N_469);
and U6706 (N_6706,N_3051,N_3366);
nor U6707 (N_6707,N_2231,N_314);
or U6708 (N_6708,N_2317,N_1218);
and U6709 (N_6709,N_4998,N_3408);
and U6710 (N_6710,N_184,N_1826);
nor U6711 (N_6711,N_1661,N_1601);
xnor U6712 (N_6712,N_2241,N_2752);
xor U6713 (N_6713,N_1686,N_3519);
nor U6714 (N_6714,N_3659,N_2601);
nand U6715 (N_6715,N_3868,N_4665);
nor U6716 (N_6716,N_2722,N_2950);
and U6717 (N_6717,N_2648,N_74);
and U6718 (N_6718,N_48,N_3904);
or U6719 (N_6719,N_1766,N_1656);
nor U6720 (N_6720,N_3675,N_4252);
and U6721 (N_6721,N_2271,N_272);
or U6722 (N_6722,N_4292,N_3319);
nand U6723 (N_6723,N_3365,N_1212);
or U6724 (N_6724,N_3608,N_3847);
or U6725 (N_6725,N_4669,N_120);
nand U6726 (N_6726,N_4044,N_4983);
nand U6727 (N_6727,N_301,N_4874);
nor U6728 (N_6728,N_4810,N_2449);
and U6729 (N_6729,N_3783,N_3992);
nor U6730 (N_6730,N_4431,N_361);
or U6731 (N_6731,N_3058,N_4951);
xor U6732 (N_6732,N_3883,N_2033);
nand U6733 (N_6733,N_3603,N_558);
and U6734 (N_6734,N_111,N_2991);
xor U6735 (N_6735,N_4826,N_3182);
xnor U6736 (N_6736,N_4700,N_3739);
nor U6737 (N_6737,N_37,N_1004);
nor U6738 (N_6738,N_4686,N_1920);
and U6739 (N_6739,N_4875,N_2027);
and U6740 (N_6740,N_2240,N_2726);
nor U6741 (N_6741,N_2802,N_134);
xnor U6742 (N_6742,N_3327,N_707);
and U6743 (N_6743,N_4458,N_1479);
nand U6744 (N_6744,N_3143,N_4003);
xnor U6745 (N_6745,N_3834,N_3948);
and U6746 (N_6746,N_3027,N_4705);
xnor U6747 (N_6747,N_932,N_3370);
nor U6748 (N_6748,N_52,N_4000);
nor U6749 (N_6749,N_2681,N_1503);
and U6750 (N_6750,N_779,N_2894);
nor U6751 (N_6751,N_2145,N_4340);
nand U6752 (N_6752,N_3111,N_2900);
xnor U6753 (N_6753,N_739,N_4641);
xor U6754 (N_6754,N_3243,N_3673);
and U6755 (N_6755,N_4209,N_877);
and U6756 (N_6756,N_1363,N_56);
xnor U6757 (N_6757,N_1287,N_2302);
xnor U6758 (N_6758,N_2042,N_3375);
nor U6759 (N_6759,N_4957,N_1336);
or U6760 (N_6760,N_28,N_2902);
nor U6761 (N_6761,N_4219,N_1517);
nand U6762 (N_6762,N_4756,N_991);
and U6763 (N_6763,N_493,N_209);
and U6764 (N_6764,N_4682,N_1715);
nor U6765 (N_6765,N_1497,N_4869);
and U6766 (N_6766,N_3584,N_2799);
xnor U6767 (N_6767,N_4316,N_2964);
xor U6768 (N_6768,N_2910,N_3401);
xor U6769 (N_6769,N_2121,N_3878);
or U6770 (N_6770,N_2204,N_4967);
xnor U6771 (N_6771,N_1143,N_4347);
nand U6772 (N_6772,N_1643,N_3643);
or U6773 (N_6773,N_2700,N_567);
nand U6774 (N_6774,N_2362,N_1869);
and U6775 (N_6775,N_2616,N_2831);
nand U6776 (N_6776,N_1440,N_4281);
and U6777 (N_6777,N_1748,N_4738);
and U6778 (N_6778,N_3531,N_1415);
or U6779 (N_6779,N_121,N_2203);
xnor U6780 (N_6780,N_4086,N_2183);
xor U6781 (N_6781,N_3566,N_1743);
nand U6782 (N_6782,N_2868,N_2100);
or U6783 (N_6783,N_3381,N_2185);
nor U6784 (N_6784,N_3799,N_3687);
nand U6785 (N_6785,N_367,N_1994);
or U6786 (N_6786,N_4131,N_2565);
and U6787 (N_6787,N_705,N_1447);
xor U6788 (N_6788,N_4533,N_2310);
xnor U6789 (N_6789,N_3724,N_2848);
or U6790 (N_6790,N_2175,N_167);
and U6791 (N_6791,N_1462,N_1760);
xnor U6792 (N_6792,N_2537,N_3369);
and U6793 (N_6793,N_976,N_414);
or U6794 (N_6794,N_2957,N_1203);
nor U6795 (N_6795,N_925,N_1564);
xnor U6796 (N_6796,N_467,N_3788);
and U6797 (N_6797,N_4504,N_2099);
or U6798 (N_6798,N_445,N_1360);
nor U6799 (N_6799,N_3311,N_186);
or U6800 (N_6800,N_948,N_1193);
and U6801 (N_6801,N_2599,N_3922);
or U6802 (N_6802,N_1318,N_2731);
and U6803 (N_6803,N_736,N_913);
and U6804 (N_6804,N_181,N_4961);
and U6805 (N_6805,N_2924,N_4212);
nor U6806 (N_6806,N_2532,N_191);
and U6807 (N_6807,N_886,N_4338);
nor U6808 (N_6808,N_3939,N_1996);
and U6809 (N_6809,N_1011,N_3772);
or U6810 (N_6810,N_3752,N_471);
nand U6811 (N_6811,N_1153,N_3966);
xnor U6812 (N_6812,N_1899,N_1119);
and U6813 (N_6813,N_4026,N_1454);
or U6814 (N_6814,N_1209,N_3173);
nor U6815 (N_6815,N_408,N_302);
nor U6816 (N_6816,N_2321,N_3795);
xor U6817 (N_6817,N_4828,N_1841);
or U6818 (N_6818,N_3151,N_3843);
nand U6819 (N_6819,N_1335,N_1317);
nor U6820 (N_6820,N_2035,N_2392);
xor U6821 (N_6821,N_2880,N_2812);
and U6822 (N_6822,N_2760,N_344);
or U6823 (N_6823,N_4482,N_2587);
or U6824 (N_6824,N_1481,N_4977);
nand U6825 (N_6825,N_2611,N_4029);
or U6826 (N_6826,N_2062,N_4215);
xor U6827 (N_6827,N_3464,N_3725);
and U6828 (N_6828,N_3004,N_2969);
or U6829 (N_6829,N_448,N_2486);
nor U6830 (N_6830,N_4010,N_1679);
or U6831 (N_6831,N_2869,N_310);
nor U6832 (N_6832,N_4936,N_281);
and U6833 (N_6833,N_1882,N_4889);
nand U6834 (N_6834,N_2575,N_4141);
nor U6835 (N_6835,N_4381,N_4529);
xnor U6836 (N_6836,N_2580,N_3115);
nor U6837 (N_6837,N_103,N_4461);
xor U6838 (N_6838,N_833,N_4859);
nor U6839 (N_6839,N_2559,N_1353);
or U6840 (N_6840,N_3245,N_912);
or U6841 (N_6841,N_3443,N_609);
or U6842 (N_6842,N_2368,N_820);
and U6843 (N_6843,N_3310,N_1264);
nand U6844 (N_6844,N_2865,N_4690);
and U6845 (N_6845,N_1216,N_2353);
nand U6846 (N_6846,N_1465,N_4005);
xnor U6847 (N_6847,N_3684,N_2382);
or U6848 (N_6848,N_346,N_3971);
nand U6849 (N_6849,N_4941,N_1448);
nand U6850 (N_6850,N_1610,N_2344);
or U6851 (N_6851,N_3179,N_4360);
and U6852 (N_6852,N_4237,N_398);
or U6853 (N_6853,N_4972,N_2425);
nor U6854 (N_6854,N_4922,N_3336);
xnor U6855 (N_6855,N_243,N_2272);
nor U6856 (N_6856,N_1411,N_4949);
xor U6857 (N_6857,N_610,N_4288);
xnor U6858 (N_6858,N_3612,N_4643);
nor U6859 (N_6859,N_695,N_125);
nand U6860 (N_6860,N_3237,N_3654);
nor U6861 (N_6861,N_3569,N_3150);
or U6862 (N_6862,N_3021,N_3063);
xnor U6863 (N_6863,N_1115,N_4375);
and U6864 (N_6864,N_1331,N_3059);
or U6865 (N_6865,N_1356,N_3536);
nand U6866 (N_6866,N_388,N_3434);
nand U6867 (N_6867,N_1366,N_3463);
or U6868 (N_6868,N_4689,N_15);
and U6869 (N_6869,N_3432,N_4419);
nor U6870 (N_6870,N_2483,N_1675);
and U6871 (N_6871,N_4247,N_4034);
and U6872 (N_6872,N_4479,N_1999);
nand U6873 (N_6873,N_2044,N_3543);
or U6874 (N_6874,N_4153,N_2888);
and U6875 (N_6875,N_2351,N_4906);
nor U6876 (N_6876,N_4308,N_3938);
nor U6877 (N_6877,N_199,N_4169);
and U6878 (N_6878,N_3476,N_1975);
nand U6879 (N_6879,N_4566,N_4971);
nand U6880 (N_6880,N_4718,N_4486);
nor U6881 (N_6881,N_4837,N_3047);
nand U6882 (N_6882,N_1582,N_2012);
or U6883 (N_6883,N_1051,N_4159);
xnor U6884 (N_6884,N_3537,N_4618);
xnor U6885 (N_6885,N_2789,N_4139);
xnor U6886 (N_6886,N_244,N_3806);
or U6887 (N_6887,N_2707,N_2034);
or U6888 (N_6888,N_2197,N_2140);
nand U6889 (N_6889,N_3743,N_88);
nand U6890 (N_6890,N_1099,N_2390);
nand U6891 (N_6891,N_1030,N_2701);
nand U6892 (N_6892,N_4804,N_3117);
nand U6893 (N_6893,N_1705,N_2210);
nand U6894 (N_6894,N_2541,N_3331);
and U6895 (N_6895,N_153,N_3158);
and U6896 (N_6896,N_2048,N_3538);
nand U6897 (N_6897,N_82,N_105);
or U6898 (N_6898,N_3386,N_4899);
nand U6899 (N_6899,N_3122,N_3742);
and U6900 (N_6900,N_2805,N_2787);
nor U6901 (N_6901,N_4583,N_4609);
xnor U6902 (N_6902,N_4555,N_938);
xnor U6903 (N_6903,N_4793,N_4200);
or U6904 (N_6904,N_2512,N_2511);
and U6905 (N_6905,N_677,N_2987);
or U6906 (N_6906,N_3483,N_29);
nand U6907 (N_6907,N_745,N_1463);
and U6908 (N_6908,N_4277,N_858);
xnor U6909 (N_6909,N_942,N_4079);
or U6910 (N_6910,N_1320,N_647);
nor U6911 (N_6911,N_3848,N_64);
xor U6912 (N_6912,N_1531,N_963);
nor U6913 (N_6913,N_3595,N_1812);
xor U6914 (N_6914,N_807,N_4661);
nor U6915 (N_6915,N_4973,N_202);
and U6916 (N_6916,N_1298,N_3491);
nor U6917 (N_6917,N_3884,N_1187);
and U6918 (N_6918,N_4711,N_130);
or U6919 (N_6919,N_4668,N_1926);
and U6920 (N_6920,N_2928,N_2626);
xor U6921 (N_6921,N_2856,N_3212);
xnor U6922 (N_6922,N_1892,N_2829);
or U6923 (N_6923,N_1306,N_1578);
or U6924 (N_6924,N_1716,N_2569);
and U6925 (N_6925,N_4379,N_295);
nand U6926 (N_6926,N_3802,N_4516);
nor U6927 (N_6927,N_1721,N_2307);
nor U6928 (N_6928,N_2870,N_3680);
and U6929 (N_6929,N_4954,N_664);
and U6930 (N_6930,N_1815,N_39);
nand U6931 (N_6931,N_952,N_1292);
or U6932 (N_6932,N_1648,N_1707);
nand U6933 (N_6933,N_1407,N_2576);
nand U6934 (N_6934,N_418,N_4945);
xnor U6935 (N_6935,N_1672,N_3078);
or U6936 (N_6936,N_975,N_2193);
nor U6937 (N_6937,N_1628,N_1787);
nand U6938 (N_6938,N_836,N_1723);
nand U6939 (N_6939,N_3092,N_909);
and U6940 (N_6940,N_4920,N_1429);
or U6941 (N_6941,N_2232,N_2316);
nor U6942 (N_6942,N_333,N_3722);
or U6943 (N_6943,N_3146,N_3639);
xnor U6944 (N_6944,N_1667,N_1358);
nand U6945 (N_6945,N_2264,N_3338);
and U6946 (N_6946,N_3787,N_2577);
and U6947 (N_6947,N_2545,N_2528);
and U6948 (N_6948,N_87,N_2514);
and U6949 (N_6949,N_3670,N_2549);
nand U6950 (N_6950,N_1452,N_813);
xnor U6951 (N_6951,N_4667,N_1614);
and U6952 (N_6952,N_3750,N_2411);
nor U6953 (N_6953,N_1427,N_1256);
xor U6954 (N_6954,N_903,N_1089);
or U6955 (N_6955,N_3166,N_2053);
nand U6956 (N_6956,N_4540,N_1242);
and U6957 (N_6957,N_1057,N_3613);
or U6958 (N_6958,N_1652,N_2763);
and U6959 (N_6959,N_251,N_127);
nor U6960 (N_6960,N_32,N_2583);
nor U6961 (N_6961,N_4825,N_940);
and U6962 (N_6962,N_3737,N_4497);
nor U6963 (N_6963,N_3841,N_2334);
nand U6964 (N_6964,N_4777,N_3299);
nor U6965 (N_6965,N_1691,N_4152);
nand U6966 (N_6966,N_2373,N_3328);
nand U6967 (N_6967,N_2153,N_3924);
xor U6968 (N_6968,N_4929,N_1621);
and U6969 (N_6969,N_4025,N_1074);
and U6970 (N_6970,N_196,N_1972);
xor U6971 (N_6971,N_3342,N_383);
nor U6972 (N_6972,N_4298,N_3341);
or U6973 (N_6973,N_3915,N_2630);
and U6974 (N_6974,N_2617,N_44);
and U6975 (N_6975,N_3042,N_2372);
and U6976 (N_6976,N_4188,N_2394);
nand U6977 (N_6977,N_4976,N_564);
xnor U6978 (N_6978,N_115,N_989);
nor U6979 (N_6979,N_2782,N_4145);
and U6980 (N_6980,N_4198,N_1557);
or U6981 (N_6981,N_282,N_4083);
nor U6982 (N_6982,N_4411,N_1184);
or U6983 (N_6983,N_2064,N_2498);
nor U6984 (N_6984,N_2783,N_430);
and U6985 (N_6985,N_4054,N_2588);
nor U6986 (N_6986,N_2315,N_4491);
nand U6987 (N_6987,N_3062,N_1554);
xor U6988 (N_6988,N_823,N_2946);
or U6989 (N_6989,N_2550,N_3273);
xnor U6990 (N_6990,N_1816,N_2981);
nand U6991 (N_6991,N_2192,N_3094);
and U6992 (N_6992,N_4367,N_1974);
nor U6993 (N_6993,N_997,N_2769);
nor U6994 (N_6994,N_4739,N_4365);
and U6995 (N_6995,N_1,N_542);
and U6996 (N_6996,N_4733,N_3266);
nor U6997 (N_6997,N_274,N_2214);
nor U6998 (N_6998,N_765,N_1049);
nand U6999 (N_6999,N_3009,N_3041);
nor U7000 (N_7000,N_3872,N_3664);
xor U7001 (N_7001,N_254,N_501);
xnor U7002 (N_7002,N_3176,N_4201);
nand U7003 (N_7003,N_1210,N_3363);
xnor U7004 (N_7004,N_4476,N_1104);
and U7005 (N_7005,N_4156,N_36);
nand U7006 (N_7006,N_1006,N_1068);
nand U7007 (N_7007,N_4378,N_3541);
nor U7008 (N_7008,N_1003,N_3265);
nand U7009 (N_7009,N_3682,N_4099);
or U7010 (N_7010,N_240,N_2899);
and U7011 (N_7011,N_440,N_973);
nand U7012 (N_7012,N_1095,N_2014);
xnor U7013 (N_7013,N_1221,N_2191);
and U7014 (N_7014,N_432,N_374);
or U7015 (N_7015,N_3234,N_2480);
xor U7016 (N_7016,N_2224,N_2448);
and U7017 (N_7017,N_3132,N_2065);
or U7018 (N_7018,N_1383,N_4923);
nor U7019 (N_7019,N_3792,N_4454);
or U7020 (N_7020,N_3180,N_3136);
nor U7021 (N_7021,N_1274,N_3961);
nor U7022 (N_7022,N_3124,N_2402);
nor U7023 (N_7023,N_2822,N_1388);
or U7024 (N_7024,N_3061,N_1158);
nor U7025 (N_7025,N_1110,N_3651);
nand U7026 (N_7026,N_4057,N_1246);
nor U7027 (N_7027,N_916,N_31);
or U7028 (N_7028,N_2113,N_719);
and U7029 (N_7029,N_4768,N_4704);
and U7030 (N_7030,N_4092,N_2172);
xor U7031 (N_7031,N_2355,N_236);
nor U7032 (N_7032,N_1389,N_3290);
and U7033 (N_7033,N_1568,N_2013);
xor U7034 (N_7034,N_421,N_4342);
and U7035 (N_7035,N_2963,N_341);
xnor U7036 (N_7036,N_3908,N_1114);
nor U7037 (N_7037,N_625,N_486);
xor U7038 (N_7038,N_1600,N_529);
or U7039 (N_7039,N_3025,N_3315);
nor U7040 (N_7040,N_1688,N_1180);
xor U7041 (N_7041,N_2295,N_18);
or U7042 (N_7042,N_468,N_3600);
xor U7043 (N_7043,N_271,N_653);
nand U7044 (N_7044,N_4743,N_1385);
and U7045 (N_7045,N_1303,N_3578);
or U7046 (N_7046,N_4312,N_1446);
nand U7047 (N_7047,N_2609,N_3530);
and U7048 (N_7048,N_1670,N_2578);
or U7049 (N_7049,N_1938,N_24);
and U7050 (N_7050,N_3445,N_4817);
or U7051 (N_7051,N_816,N_1333);
nor U7052 (N_7052,N_3893,N_355);
nand U7053 (N_7053,N_4940,N_2689);
nand U7054 (N_7054,N_3337,N_412);
or U7055 (N_7055,N_1283,N_1653);
xnor U7056 (N_7056,N_4121,N_4902);
and U7057 (N_7057,N_2209,N_2622);
nand U7058 (N_7058,N_1357,N_3579);
nor U7059 (N_7059,N_1599,N_1636);
or U7060 (N_7060,N_4107,N_2154);
or U7061 (N_7061,N_4372,N_137);
xor U7062 (N_7062,N_1607,N_4331);
nand U7063 (N_7063,N_45,N_1001);
xor U7064 (N_7064,N_1566,N_4728);
xor U7065 (N_7065,N_2686,N_2487);
nor U7066 (N_7066,N_2319,N_2895);
nand U7067 (N_7067,N_3740,N_718);
or U7068 (N_7068,N_3796,N_1708);
or U7069 (N_7069,N_667,N_3469);
xor U7070 (N_7070,N_359,N_4962);
xnor U7071 (N_7071,N_956,N_3956);
nand U7072 (N_7072,N_1791,N_3594);
nor U7073 (N_7073,N_530,N_1014);
nor U7074 (N_7074,N_4574,N_2262);
xor U7075 (N_7075,N_2842,N_148);
nand U7076 (N_7076,N_3254,N_1823);
or U7077 (N_7077,N_3316,N_1421);
and U7078 (N_7078,N_3629,N_3957);
or U7079 (N_7079,N_1856,N_4622);
or U7080 (N_7080,N_3895,N_2247);
nand U7081 (N_7081,N_1402,N_620);
and U7082 (N_7082,N_1765,N_4679);
nand U7083 (N_7083,N_3527,N_3627);
or U7084 (N_7084,N_2409,N_522);
or U7085 (N_7085,N_3661,N_2342);
and U7086 (N_7086,N_2202,N_2500);
xnor U7087 (N_7087,N_4077,N_3624);
nor U7088 (N_7088,N_4028,N_1059);
nor U7089 (N_7089,N_1979,N_1273);
nand U7090 (N_7090,N_53,N_4820);
xnor U7091 (N_7091,N_3330,N_3923);
nor U7092 (N_7092,N_3930,N_4975);
xnor U7093 (N_7093,N_2186,N_4757);
xor U7094 (N_7094,N_3324,N_1260);
xnor U7095 (N_7095,N_1637,N_1500);
nor U7096 (N_7096,N_1195,N_1350);
nand U7097 (N_7097,N_2077,N_323);
xnor U7098 (N_7098,N_1478,N_2476);
nor U7099 (N_7099,N_2976,N_2879);
or U7100 (N_7100,N_4783,N_3811);
and U7101 (N_7101,N_4637,N_1903);
nor U7102 (N_7102,N_687,N_2128);
nor U7103 (N_7103,N_2538,N_277);
nand U7104 (N_7104,N_1139,N_2309);
or U7105 (N_7105,N_4362,N_4878);
nand U7106 (N_7106,N_1732,N_416);
or U7107 (N_7107,N_2493,N_2730);
nor U7108 (N_7108,N_1494,N_2602);
nor U7109 (N_7109,N_859,N_587);
xnor U7110 (N_7110,N_2891,N_1522);
nor U7111 (N_7111,N_3821,N_3287);
nand U7112 (N_7112,N_3623,N_3343);
or U7113 (N_7113,N_1396,N_2237);
nand U7114 (N_7114,N_1245,N_3920);
xnor U7115 (N_7115,N_4266,N_3958);
or U7116 (N_7116,N_633,N_129);
and U7117 (N_7117,N_2614,N_3980);
nand U7118 (N_7118,N_570,N_865);
xnor U7119 (N_7119,N_540,N_761);
and U7120 (N_7120,N_4999,N_1794);
and U7121 (N_7121,N_1048,N_2745);
xnor U7122 (N_7122,N_135,N_4333);
nand U7123 (N_7123,N_546,N_3953);
nand U7124 (N_7124,N_2280,N_1836);
or U7125 (N_7125,N_3695,N_1772);
xor U7126 (N_7126,N_3954,N_21);
or U7127 (N_7127,N_4856,N_4234);
nor U7128 (N_7128,N_2337,N_4272);
or U7129 (N_7129,N_4108,N_2284);
nand U7130 (N_7130,N_3952,N_1786);
nor U7131 (N_7131,N_2650,N_1228);
and U7132 (N_7132,N_2239,N_4225);
and U7133 (N_7133,N_3738,N_3485);
xor U7134 (N_7134,N_2200,N_4994);
and U7135 (N_7135,N_3854,N_4564);
or U7136 (N_7136,N_2040,N_4013);
and U7137 (N_7137,N_1726,N_3102);
xor U7138 (N_7138,N_4606,N_4724);
nor U7139 (N_7139,N_2893,N_1594);
xnor U7140 (N_7140,N_2929,N_2704);
xor U7141 (N_7141,N_4558,N_2979);
or U7142 (N_7142,N_3644,N_3751);
or U7143 (N_7143,N_3447,N_3095);
and U7144 (N_7144,N_3255,N_4435);
and U7145 (N_7145,N_1106,N_526);
xor U7146 (N_7146,N_1733,N_3500);
nand U7147 (N_7147,N_686,N_1382);
or U7148 (N_7148,N_777,N_2627);
nand U7149 (N_7149,N_46,N_512);
nand U7150 (N_7150,N_1505,N_977);
nor U7151 (N_7151,N_4420,N_931);
nor U7152 (N_7152,N_4465,N_60);
or U7153 (N_7153,N_4550,N_84);
nand U7154 (N_7154,N_4130,N_1160);
nand U7155 (N_7155,N_1131,N_2410);
xor U7156 (N_7156,N_2832,N_3451);
nor U7157 (N_7157,N_279,N_1755);
nand U7158 (N_7158,N_258,N_2826);
and U7159 (N_7159,N_4882,N_2107);
nor U7160 (N_7160,N_2892,N_2807);
and U7161 (N_7161,N_2055,N_2318);
or U7162 (N_7162,N_635,N_803);
nand U7163 (N_7163,N_2684,N_1973);
and U7164 (N_7164,N_3959,N_980);
and U7165 (N_7165,N_3910,N_3412);
nor U7166 (N_7166,N_4474,N_322);
xnor U7167 (N_7167,N_3035,N_2621);
and U7168 (N_7168,N_645,N_4942);
or U7169 (N_7169,N_4113,N_1818);
and U7170 (N_7170,N_4534,N_4846);
and U7171 (N_7171,N_4415,N_1770);
xnor U7172 (N_7172,N_2098,N_1537);
and U7173 (N_7173,N_3068,N_2836);
nor U7174 (N_7174,N_3990,N_4515);
nand U7175 (N_7175,N_100,N_2623);
and U7176 (N_7176,N_2471,N_6);
xnor U7177 (N_7177,N_1477,N_114);
nand U7178 (N_7178,N_4383,N_2166);
nand U7179 (N_7179,N_3379,N_2761);
xnor U7180 (N_7180,N_604,N_3301);
and U7181 (N_7181,N_4795,N_3304);
nor U7182 (N_7182,N_2733,N_3152);
and U7183 (N_7183,N_2938,N_2462);
nor U7184 (N_7184,N_1399,N_1019);
and U7185 (N_7185,N_4032,N_851);
or U7186 (N_7186,N_3866,N_697);
xor U7187 (N_7187,N_2496,N_16);
or U7188 (N_7188,N_2037,N_420);
and U7189 (N_7189,N_3550,N_2854);
nand U7190 (N_7190,N_3216,N_1430);
nor U7191 (N_7191,N_627,N_939);
and U7192 (N_7192,N_4776,N_3103);
or U7193 (N_7193,N_3855,N_2259);
or U7194 (N_7194,N_2443,N_1058);
or U7195 (N_7195,N_1352,N_3011);
nand U7196 (N_7196,N_4670,N_4813);
xnor U7197 (N_7197,N_4651,N_3983);
and U7198 (N_7198,N_169,N_3329);
and U7199 (N_7199,N_4441,N_34);
nand U7200 (N_7200,N_1664,N_4452);
or U7201 (N_7201,N_2379,N_1893);
nor U7202 (N_7202,N_3405,N_4663);
xor U7203 (N_7203,N_2422,N_38);
xor U7204 (N_7204,N_4307,N_636);
xnor U7205 (N_7205,N_1300,N_2);
xor U7206 (N_7206,N_4268,N_3850);
xor U7207 (N_7207,N_552,N_3840);
or U7208 (N_7208,N_2333,N_1959);
xor U7209 (N_7209,N_3784,N_4208);
nand U7210 (N_7210,N_150,N_756);
nand U7211 (N_7211,N_1917,N_4224);
or U7212 (N_7212,N_3133,N_2507);
and U7213 (N_7213,N_3334,N_357);
nand U7214 (N_7214,N_3660,N_4890);
nor U7215 (N_7215,N_908,N_2218);
or U7216 (N_7216,N_3050,N_152);
nand U7217 (N_7217,N_584,N_4581);
xnor U7218 (N_7218,N_2253,N_1375);
nand U7219 (N_7219,N_3880,N_682);
xnor U7220 (N_7220,N_4745,N_2978);
nor U7221 (N_7221,N_1063,N_3072);
and U7222 (N_7222,N_1204,N_4552);
xnor U7223 (N_7223,N_2161,N_4927);
and U7224 (N_7224,N_1323,N_1252);
or U7225 (N_7225,N_1198,N_2908);
xor U7226 (N_7226,N_1929,N_3818);
and U7227 (N_7227,N_4249,N_3321);
or U7228 (N_7228,N_4729,N_1265);
or U7229 (N_7229,N_808,N_4401);
and U7230 (N_7230,N_4120,N_1669);
or U7231 (N_7231,N_3223,N_1484);
and U7232 (N_7232,N_4236,N_285);
or U7233 (N_7233,N_1409,N_2503);
and U7234 (N_7234,N_2846,N_2079);
nand U7235 (N_7235,N_1262,N_79);
nand U7236 (N_7236,N_1863,N_3513);
nand U7237 (N_7237,N_2347,N_2813);
and U7238 (N_7238,N_1159,N_3588);
nor U7239 (N_7239,N_3827,N_1777);
or U7240 (N_7240,N_4989,N_3911);
nor U7241 (N_7241,N_674,N_3979);
nor U7242 (N_7242,N_4614,N_4703);
nand U7243 (N_7243,N_2563,N_1088);
nand U7244 (N_7244,N_4613,N_3585);
or U7245 (N_7245,N_1015,N_4403);
and U7246 (N_7246,N_2405,N_1819);
and U7247 (N_7247,N_189,N_51);
and U7248 (N_7248,N_2465,N_2930);
nand U7249 (N_7249,N_4584,N_4185);
nor U7250 (N_7250,N_860,N_1398);
or U7251 (N_7251,N_2051,N_999);
xor U7252 (N_7252,N_1828,N_442);
nor U7253 (N_7253,N_2030,N_4053);
and U7254 (N_7254,N_2406,N_511);
or U7255 (N_7255,N_3836,N_3899);
and U7256 (N_7256,N_4603,N_722);
or U7257 (N_7257,N_2255,N_1108);
xnor U7258 (N_7258,N_812,N_2520);
and U7259 (N_7259,N_844,N_2501);
xnor U7260 (N_7260,N_3313,N_3258);
xnor U7261 (N_7261,N_4438,N_1211);
or U7262 (N_7262,N_1381,N_680);
and U7263 (N_7263,N_3306,N_3766);
and U7264 (N_7264,N_3548,N_2176);
xor U7265 (N_7265,N_1950,N_3433);
and U7266 (N_7266,N_373,N_1103);
nand U7267 (N_7267,N_4211,N_2188);
xnor U7268 (N_7268,N_3810,N_4324);
and U7269 (N_7269,N_2753,N_1032);
or U7270 (N_7270,N_954,N_2427);
and U7271 (N_7271,N_4761,N_1489);
nor U7272 (N_7272,N_654,N_2433);
nor U7273 (N_7273,N_318,N_1700);
nand U7274 (N_7274,N_2378,N_3776);
xor U7275 (N_7275,N_3209,N_1474);
nor U7276 (N_7276,N_3937,N_3452);
nor U7277 (N_7277,N_4253,N_4336);
nor U7278 (N_7278,N_1327,N_4924);
nand U7279 (N_7279,N_1278,N_1042);
and U7280 (N_7280,N_1742,N_487);
and U7281 (N_7281,N_2451,N_958);
or U7282 (N_7282,N_3193,N_897);
nand U7283 (N_7283,N_2534,N_2986);
nor U7284 (N_7284,N_1028,N_1403);
xor U7285 (N_7285,N_43,N_2165);
or U7286 (N_7286,N_2163,N_59);
or U7287 (N_7287,N_2112,N_2638);
and U7288 (N_7288,N_753,N_495);
or U7289 (N_7289,N_4598,N_4834);
and U7290 (N_7290,N_222,N_4879);
nor U7291 (N_7291,N_4235,N_4863);
and U7292 (N_7292,N_4602,N_4227);
xnor U7293 (N_7293,N_2094,N_76);
or U7294 (N_7294,N_3423,N_3614);
xor U7295 (N_7295,N_1507,N_603);
nor U7296 (N_7296,N_3777,N_870);
or U7297 (N_7297,N_1683,N_641);
or U7298 (N_7298,N_1207,N_69);
and U7299 (N_7299,N_2345,N_2216);
and U7300 (N_7300,N_4910,N_4900);
and U7301 (N_7301,N_1470,N_4313);
and U7302 (N_7302,N_1752,N_3155);
nor U7303 (N_7303,N_2369,N_4398);
xor U7304 (N_7304,N_4460,N_4493);
and U7305 (N_7305,N_2818,N_141);
nand U7306 (N_7306,N_662,N_544);
nor U7307 (N_7307,N_3473,N_3407);
and U7308 (N_7308,N_3249,N_2289);
nand U7309 (N_7309,N_3671,N_4582);
and U7310 (N_7310,N_616,N_3402);
nand U7311 (N_7311,N_4778,N_1536);
or U7312 (N_7312,N_3681,N_465);
nand U7313 (N_7313,N_3789,N_4830);
xnor U7314 (N_7314,N_2647,N_927);
nand U7315 (N_7315,N_3314,N_157);
xnor U7316 (N_7316,N_3202,N_2897);
and U7317 (N_7317,N_1150,N_1574);
and U7318 (N_7318,N_213,N_4069);
nand U7319 (N_7319,N_3382,N_1665);
xor U7320 (N_7320,N_848,N_590);
or U7321 (N_7321,N_1012,N_470);
nor U7322 (N_7322,N_4326,N_3640);
xor U7323 (N_7323,N_4721,N_252);
xnor U7324 (N_7324,N_1541,N_480);
xnor U7325 (N_7325,N_1602,N_2944);
or U7326 (N_7326,N_2636,N_1625);
nand U7327 (N_7327,N_3175,N_4517);
nand U7328 (N_7328,N_1002,N_4014);
nor U7329 (N_7329,N_3726,N_4802);
nor U7330 (N_7330,N_3879,N_4261);
nand U7331 (N_7331,N_3542,N_1775);
xor U7332 (N_7332,N_3126,N_595);
nor U7333 (N_7333,N_2300,N_4608);
nand U7334 (N_7334,N_4505,N_308);
nand U7335 (N_7335,N_4062,N_1466);
nor U7336 (N_7336,N_4,N_4166);
and U7337 (N_7337,N_3809,N_528);
and U7338 (N_7338,N_2672,N_4104);
or U7339 (N_7339,N_2327,N_287);
nand U7340 (N_7340,N_2453,N_3084);
and U7341 (N_7341,N_3012,N_1232);
xnor U7342 (N_7342,N_569,N_379);
and U7343 (N_7343,N_3967,N_895);
or U7344 (N_7344,N_3617,N_224);
nor U7345 (N_7345,N_3870,N_4538);
xnor U7346 (N_7346,N_3913,N_3702);
or U7347 (N_7347,N_1855,N_663);
or U7348 (N_7348,N_1985,N_2966);
xor U7349 (N_7349,N_2629,N_4207);
or U7350 (N_7350,N_565,N_2131);
nand U7351 (N_7351,N_3706,N_1239);
xor U7352 (N_7352,N_2657,N_4146);
nor U7353 (N_7353,N_2461,N_2414);
and U7354 (N_7354,N_3504,N_145);
or U7355 (N_7355,N_3781,N_3946);
nand U7356 (N_7356,N_237,N_1543);
xnor U7357 (N_7357,N_532,N_2072);
xnor U7358 (N_7358,N_2716,N_4109);
and U7359 (N_7359,N_2249,N_1000);
nor U7360 (N_7360,N_1297,N_3171);
and U7361 (N_7361,N_3728,N_2002);
xnor U7362 (N_7362,N_2706,N_203);
and U7363 (N_7363,N_4766,N_456);
nand U7364 (N_7364,N_4588,N_19);
xnor U7365 (N_7365,N_4880,N_1175);
nand U7366 (N_7366,N_369,N_164);
nor U7367 (N_7367,N_3998,N_4058);
or U7368 (N_7368,N_1951,N_42);
xnor U7369 (N_7369,N_4901,N_4915);
xor U7370 (N_7370,N_2238,N_4456);
nand U7371 (N_7371,N_1699,N_4157);
and U7372 (N_7372,N_4042,N_3029);
or U7373 (N_7373,N_1619,N_3488);
nor U7374 (N_7374,N_3280,N_2992);
or U7375 (N_7375,N_1471,N_2919);
nor U7376 (N_7376,N_3440,N_4406);
xor U7377 (N_7377,N_2547,N_3065);
nor U7378 (N_7378,N_4182,N_1640);
and U7379 (N_7379,N_2980,N_4988);
nand U7380 (N_7380,N_348,N_1456);
xnor U7381 (N_7381,N_4851,N_4568);
and U7382 (N_7382,N_1864,N_4771);
or U7383 (N_7383,N_1978,N_4835);
nor U7384 (N_7384,N_1730,N_575);
or U7385 (N_7385,N_1939,N_453);
nor U7386 (N_7386,N_743,N_2890);
or U7387 (N_7387,N_2645,N_4513);
and U7388 (N_7388,N_2816,N_2350);
nor U7389 (N_7389,N_3707,N_969);
or U7390 (N_7390,N_1545,N_1720);
nand U7391 (N_7391,N_1624,N_2376);
nor U7392 (N_7392,N_1023,N_2365);
nor U7393 (N_7393,N_4845,N_2046);
xnor U7394 (N_7394,N_2606,N_588);
nand U7395 (N_7395,N_563,N_1513);
nand U7396 (N_7396,N_1976,N_1718);
nand U7397 (N_7397,N_3048,N_2841);
xor U7398 (N_7398,N_2711,N_1581);
nor U7399 (N_7399,N_2016,N_4137);
and U7400 (N_7400,N_3187,N_2995);
nor U7401 (N_7401,N_2005,N_3698);
nor U7402 (N_7402,N_4627,N_2851);
nor U7403 (N_7403,N_828,N_2766);
xnor U7404 (N_7404,N_2750,N_3017);
nor U7405 (N_7405,N_3057,N_1041);
and U7406 (N_7406,N_268,N_715);
or U7407 (N_7407,N_4400,N_1897);
or U7408 (N_7408,N_1037,N_1215);
nand U7409 (N_7409,N_3748,N_2058);
xor U7410 (N_7410,N_2781,N_1955);
and U7411 (N_7411,N_930,N_4373);
and U7412 (N_7412,N_2936,N_3717);
and U7413 (N_7413,N_3289,N_2229);
nand U7414 (N_7414,N_262,N_393);
xor U7415 (N_7415,N_3353,N_494);
nand U7416 (N_7416,N_1871,N_3921);
or U7417 (N_7417,N_834,N_273);
or U7418 (N_7418,N_2141,N_4865);
or U7419 (N_7419,N_3339,N_3561);
nor U7420 (N_7420,N_2489,N_751);
xor U7421 (N_7421,N_2618,N_769);
nand U7422 (N_7422,N_3291,N_2907);
and U7423 (N_7423,N_880,N_3523);
and U7424 (N_7424,N_3632,N_698);
or U7425 (N_7425,N_1813,N_122);
or U7426 (N_7426,N_2885,N_1029);
nand U7427 (N_7427,N_1853,N_2375);
nor U7428 (N_7428,N_4439,N_4276);
xnor U7429 (N_7429,N_3384,N_613);
or U7430 (N_7430,N_3000,N_156);
xor U7431 (N_7431,N_4735,N_2664);
xnor U7432 (N_7432,N_3593,N_2804);
xnor U7433 (N_7433,N_303,N_4115);
and U7434 (N_7434,N_3022,N_2719);
xnor U7435 (N_7435,N_3520,N_1376);
or U7436 (N_7436,N_4356,N_4303);
nor U7437 (N_7437,N_578,N_4017);
nor U7438 (N_7438,N_4302,N_3292);
and U7439 (N_7439,N_3987,N_3159);
or U7440 (N_7440,N_981,N_1364);
or U7441 (N_7441,N_1087,N_1295);
nor U7442 (N_7442,N_3604,N_1493);
and U7443 (N_7443,N_3916,N_2313);
nand U7444 (N_7444,N_239,N_3626);
nor U7445 (N_7445,N_4122,N_4848);
nor U7446 (N_7446,N_256,N_4636);
xnor U7447 (N_7447,N_562,N_2384);
xnor U7448 (N_7448,N_3658,N_4087);
and U7449 (N_7449,N_2993,N_1781);
nand U7450 (N_7450,N_1722,N_4981);
xor U7451 (N_7451,N_492,N_2644);
xnor U7452 (N_7452,N_3418,N_216);
or U7453 (N_7453,N_2937,N_3067);
nand U7454 (N_7454,N_2586,N_1345);
nor U7455 (N_7455,N_1595,N_4511);
or U7456 (N_7456,N_1934,N_574);
nor U7457 (N_7457,N_946,N_1271);
or U7458 (N_7458,N_706,N_2047);
nand U7459 (N_7459,N_944,N_4969);
xor U7460 (N_7460,N_3104,N_943);
or U7461 (N_7461,N_1138,N_2774);
and U7462 (N_7462,N_1165,N_4727);
xor U7463 (N_7463,N_3955,N_2552);
nand U7464 (N_7464,N_4363,N_234);
nor U7465 (N_7465,N_3018,N_4382);
nand U7466 (N_7466,N_639,N_2428);
nand U7467 (N_7467,N_1591,N_694);
nand U7468 (N_7468,N_3842,N_3300);
xor U7469 (N_7469,N_4708,N_407);
nor U7470 (N_7470,N_399,N_4384);
nor U7471 (N_7471,N_260,N_898);
nand U7472 (N_7472,N_3100,N_1372);
and U7473 (N_7473,N_4694,N_444);
nand U7474 (N_7474,N_4549,N_792);
xnor U7475 (N_7475,N_1433,N_3577);
nor U7476 (N_7476,N_2685,N_4067);
xor U7477 (N_7477,N_1567,N_4221);
xor U7478 (N_7478,N_3486,N_3502);
xnor U7479 (N_7479,N_4573,N_4322);
xor U7480 (N_7480,N_1428,N_4167);
nand U7481 (N_7481,N_3356,N_2819);
nor U7482 (N_7482,N_3142,N_1112);
nor U7483 (N_7483,N_4354,N_1842);
or U7484 (N_7484,N_2359,N_437);
and U7485 (N_7485,N_896,N_594);
or U7486 (N_7486,N_2784,N_2639);
and U7487 (N_7487,N_94,N_288);
xor U7488 (N_7488,N_183,N_3813);
xor U7489 (N_7489,N_2564,N_1668);
xnor U7490 (N_7490,N_1778,N_4199);
nor U7491 (N_7491,N_1597,N_4218);
xor U7492 (N_7492,N_404,N_4202);
and U7493 (N_7493,N_2124,N_320);
xnor U7494 (N_7494,N_2387,N_2045);
or U7495 (N_7495,N_1915,N_1266);
nand U7496 (N_7496,N_3064,N_4300);
xor U7497 (N_7497,N_4061,N_785);
nand U7498 (N_7498,N_1422,N_729);
nor U7499 (N_7499,N_905,N_1501);
xor U7500 (N_7500,N_1080,N_247);
or U7501 (N_7501,N_586,N_3316);
or U7502 (N_7502,N_2814,N_380);
nor U7503 (N_7503,N_2992,N_4437);
nand U7504 (N_7504,N_517,N_991);
nor U7505 (N_7505,N_338,N_4107);
or U7506 (N_7506,N_2953,N_4890);
and U7507 (N_7507,N_3128,N_2636);
or U7508 (N_7508,N_4658,N_1038);
xnor U7509 (N_7509,N_3614,N_3724);
or U7510 (N_7510,N_284,N_3344);
nor U7511 (N_7511,N_1096,N_536);
or U7512 (N_7512,N_3897,N_1281);
or U7513 (N_7513,N_3775,N_2930);
nor U7514 (N_7514,N_724,N_2501);
xor U7515 (N_7515,N_1296,N_2184);
nand U7516 (N_7516,N_2890,N_3165);
or U7517 (N_7517,N_4528,N_2671);
xnor U7518 (N_7518,N_3798,N_3033);
or U7519 (N_7519,N_4509,N_3043);
and U7520 (N_7520,N_4296,N_2657);
and U7521 (N_7521,N_3774,N_3395);
nor U7522 (N_7522,N_1508,N_4720);
or U7523 (N_7523,N_3135,N_2549);
or U7524 (N_7524,N_386,N_1303);
xnor U7525 (N_7525,N_3036,N_3412);
nand U7526 (N_7526,N_1522,N_2977);
and U7527 (N_7527,N_1652,N_4733);
xnor U7528 (N_7528,N_2432,N_1902);
nand U7529 (N_7529,N_3431,N_1536);
nand U7530 (N_7530,N_4110,N_4961);
xnor U7531 (N_7531,N_3329,N_2492);
and U7532 (N_7532,N_438,N_1911);
and U7533 (N_7533,N_4586,N_3851);
nand U7534 (N_7534,N_2210,N_2747);
xor U7535 (N_7535,N_3152,N_53);
xnor U7536 (N_7536,N_3965,N_927);
or U7537 (N_7537,N_2535,N_2889);
or U7538 (N_7538,N_3216,N_1660);
and U7539 (N_7539,N_4634,N_854);
nand U7540 (N_7540,N_4775,N_2981);
xor U7541 (N_7541,N_746,N_4967);
and U7542 (N_7542,N_1755,N_2290);
or U7543 (N_7543,N_1232,N_4446);
or U7544 (N_7544,N_3421,N_3090);
and U7545 (N_7545,N_1376,N_3472);
or U7546 (N_7546,N_2691,N_1475);
or U7547 (N_7547,N_277,N_1710);
and U7548 (N_7548,N_3359,N_605);
nand U7549 (N_7549,N_767,N_4405);
nand U7550 (N_7550,N_1387,N_4024);
nand U7551 (N_7551,N_1230,N_2897);
nand U7552 (N_7552,N_3146,N_1871);
nor U7553 (N_7553,N_2049,N_1137);
nand U7554 (N_7554,N_199,N_4144);
and U7555 (N_7555,N_1065,N_4315);
nand U7556 (N_7556,N_2985,N_2688);
nand U7557 (N_7557,N_1799,N_4403);
nor U7558 (N_7558,N_2128,N_3370);
and U7559 (N_7559,N_1393,N_4302);
xor U7560 (N_7560,N_614,N_4469);
or U7561 (N_7561,N_94,N_1497);
or U7562 (N_7562,N_1771,N_2611);
and U7563 (N_7563,N_2232,N_4556);
nor U7564 (N_7564,N_641,N_3661);
xor U7565 (N_7565,N_3100,N_1131);
xor U7566 (N_7566,N_4448,N_2762);
xnor U7567 (N_7567,N_320,N_3150);
xor U7568 (N_7568,N_4140,N_2807);
nor U7569 (N_7569,N_4296,N_3182);
nor U7570 (N_7570,N_319,N_858);
nand U7571 (N_7571,N_1584,N_3581);
nand U7572 (N_7572,N_2142,N_773);
and U7573 (N_7573,N_2544,N_642);
or U7574 (N_7574,N_1251,N_2049);
xnor U7575 (N_7575,N_976,N_3702);
nand U7576 (N_7576,N_3269,N_57);
nor U7577 (N_7577,N_1534,N_4210);
and U7578 (N_7578,N_3763,N_3629);
or U7579 (N_7579,N_1502,N_4637);
nor U7580 (N_7580,N_4851,N_395);
nor U7581 (N_7581,N_216,N_2854);
xor U7582 (N_7582,N_46,N_4336);
nor U7583 (N_7583,N_3624,N_1202);
nand U7584 (N_7584,N_2905,N_4999);
and U7585 (N_7585,N_646,N_549);
or U7586 (N_7586,N_3450,N_2913);
xnor U7587 (N_7587,N_3005,N_1504);
nand U7588 (N_7588,N_1935,N_920);
nor U7589 (N_7589,N_1425,N_2961);
nand U7590 (N_7590,N_1086,N_3654);
nor U7591 (N_7591,N_4600,N_4249);
or U7592 (N_7592,N_2316,N_4679);
or U7593 (N_7593,N_3414,N_4471);
nand U7594 (N_7594,N_4976,N_3177);
or U7595 (N_7595,N_4139,N_3463);
nor U7596 (N_7596,N_4178,N_3874);
nor U7597 (N_7597,N_2106,N_267);
nor U7598 (N_7598,N_1038,N_2581);
and U7599 (N_7599,N_4269,N_822);
or U7600 (N_7600,N_3475,N_2762);
nand U7601 (N_7601,N_2849,N_972);
nor U7602 (N_7602,N_1902,N_1912);
and U7603 (N_7603,N_2098,N_1711);
nor U7604 (N_7604,N_1060,N_1048);
xnor U7605 (N_7605,N_1231,N_2674);
xor U7606 (N_7606,N_3087,N_2812);
or U7607 (N_7607,N_2715,N_2326);
xor U7608 (N_7608,N_261,N_4828);
and U7609 (N_7609,N_2548,N_1544);
nor U7610 (N_7610,N_3927,N_938);
or U7611 (N_7611,N_1304,N_4);
xnor U7612 (N_7612,N_2240,N_4949);
nor U7613 (N_7613,N_4351,N_2130);
or U7614 (N_7614,N_1911,N_2071);
nand U7615 (N_7615,N_2950,N_4963);
nand U7616 (N_7616,N_4913,N_4139);
nand U7617 (N_7617,N_2607,N_1705);
nor U7618 (N_7618,N_3421,N_346);
xnor U7619 (N_7619,N_2822,N_250);
nor U7620 (N_7620,N_2842,N_3815);
nand U7621 (N_7621,N_1453,N_2929);
or U7622 (N_7622,N_3950,N_2963);
nand U7623 (N_7623,N_1123,N_1303);
or U7624 (N_7624,N_4601,N_3714);
xnor U7625 (N_7625,N_3202,N_3973);
nand U7626 (N_7626,N_3109,N_3191);
xor U7627 (N_7627,N_1715,N_962);
or U7628 (N_7628,N_3251,N_3810);
xor U7629 (N_7629,N_1208,N_2052);
xnor U7630 (N_7630,N_3527,N_4780);
xor U7631 (N_7631,N_2073,N_1784);
xor U7632 (N_7632,N_4123,N_4276);
nand U7633 (N_7633,N_1550,N_1001);
and U7634 (N_7634,N_4224,N_3731);
xor U7635 (N_7635,N_2879,N_3745);
and U7636 (N_7636,N_559,N_2855);
xnor U7637 (N_7637,N_4427,N_3551);
nand U7638 (N_7638,N_2512,N_4607);
or U7639 (N_7639,N_1367,N_2717);
nand U7640 (N_7640,N_3024,N_2258);
and U7641 (N_7641,N_3553,N_428);
xor U7642 (N_7642,N_1955,N_1060);
nand U7643 (N_7643,N_3274,N_2004);
nand U7644 (N_7644,N_1664,N_1319);
xnor U7645 (N_7645,N_2158,N_678);
xor U7646 (N_7646,N_2432,N_3791);
nand U7647 (N_7647,N_2007,N_4109);
xor U7648 (N_7648,N_3776,N_4469);
nor U7649 (N_7649,N_2830,N_4556);
and U7650 (N_7650,N_2225,N_2867);
nand U7651 (N_7651,N_775,N_3569);
nand U7652 (N_7652,N_3766,N_3963);
xor U7653 (N_7653,N_4563,N_2268);
or U7654 (N_7654,N_935,N_636);
xnor U7655 (N_7655,N_1836,N_1295);
nand U7656 (N_7656,N_2278,N_1124);
or U7657 (N_7657,N_4327,N_502);
and U7658 (N_7658,N_4138,N_2631);
xnor U7659 (N_7659,N_1220,N_774);
nand U7660 (N_7660,N_3207,N_922);
and U7661 (N_7661,N_3147,N_4834);
and U7662 (N_7662,N_4711,N_471);
and U7663 (N_7663,N_1982,N_1244);
or U7664 (N_7664,N_2078,N_2663);
xnor U7665 (N_7665,N_2595,N_2780);
and U7666 (N_7666,N_2110,N_3784);
xor U7667 (N_7667,N_3901,N_2968);
or U7668 (N_7668,N_3146,N_2648);
nand U7669 (N_7669,N_1807,N_1281);
nand U7670 (N_7670,N_4419,N_382);
xor U7671 (N_7671,N_3396,N_4917);
nand U7672 (N_7672,N_4805,N_2349);
and U7673 (N_7673,N_1249,N_4556);
or U7674 (N_7674,N_4364,N_4062);
nor U7675 (N_7675,N_163,N_1961);
or U7676 (N_7676,N_2175,N_1275);
and U7677 (N_7677,N_3774,N_1442);
xor U7678 (N_7678,N_4329,N_4536);
or U7679 (N_7679,N_4484,N_4296);
nand U7680 (N_7680,N_991,N_4203);
nand U7681 (N_7681,N_297,N_3754);
nand U7682 (N_7682,N_1809,N_374);
or U7683 (N_7683,N_3260,N_2818);
nand U7684 (N_7684,N_3271,N_4087);
nor U7685 (N_7685,N_3331,N_4174);
xor U7686 (N_7686,N_3992,N_4341);
nand U7687 (N_7687,N_2145,N_4953);
or U7688 (N_7688,N_3304,N_4777);
and U7689 (N_7689,N_1418,N_3902);
nor U7690 (N_7690,N_70,N_4873);
and U7691 (N_7691,N_4390,N_3620);
and U7692 (N_7692,N_2143,N_3545);
and U7693 (N_7693,N_3140,N_2295);
nand U7694 (N_7694,N_4113,N_1868);
xnor U7695 (N_7695,N_1888,N_763);
nor U7696 (N_7696,N_1469,N_2224);
nand U7697 (N_7697,N_4778,N_4023);
nand U7698 (N_7698,N_2949,N_4504);
nand U7699 (N_7699,N_3982,N_3129);
nor U7700 (N_7700,N_3863,N_457);
xnor U7701 (N_7701,N_1028,N_4283);
xor U7702 (N_7702,N_2156,N_2124);
and U7703 (N_7703,N_1810,N_407);
xor U7704 (N_7704,N_2222,N_180);
xor U7705 (N_7705,N_1618,N_2181);
nand U7706 (N_7706,N_21,N_1342);
nor U7707 (N_7707,N_60,N_2337);
nor U7708 (N_7708,N_4164,N_924);
or U7709 (N_7709,N_2139,N_3158);
xor U7710 (N_7710,N_2723,N_2943);
nor U7711 (N_7711,N_4920,N_1193);
or U7712 (N_7712,N_2264,N_738);
nand U7713 (N_7713,N_741,N_2744);
nor U7714 (N_7714,N_3496,N_2948);
and U7715 (N_7715,N_3926,N_2399);
xnor U7716 (N_7716,N_4659,N_505);
and U7717 (N_7717,N_3358,N_2178);
nor U7718 (N_7718,N_2206,N_3116);
nor U7719 (N_7719,N_3503,N_593);
and U7720 (N_7720,N_2060,N_3942);
xnor U7721 (N_7721,N_4122,N_1562);
and U7722 (N_7722,N_2544,N_4398);
and U7723 (N_7723,N_2817,N_1747);
nand U7724 (N_7724,N_1881,N_4301);
nor U7725 (N_7725,N_2425,N_3755);
and U7726 (N_7726,N_1882,N_4069);
nand U7727 (N_7727,N_401,N_3696);
or U7728 (N_7728,N_1079,N_93);
nand U7729 (N_7729,N_425,N_894);
and U7730 (N_7730,N_1396,N_198);
and U7731 (N_7731,N_468,N_59);
or U7732 (N_7732,N_1869,N_4772);
and U7733 (N_7733,N_1176,N_3928);
nand U7734 (N_7734,N_2166,N_3894);
or U7735 (N_7735,N_2899,N_1259);
xnor U7736 (N_7736,N_2548,N_319);
or U7737 (N_7737,N_3961,N_303);
xnor U7738 (N_7738,N_3601,N_3221);
nor U7739 (N_7739,N_3026,N_1456);
nor U7740 (N_7740,N_2366,N_4712);
and U7741 (N_7741,N_3614,N_4703);
nor U7742 (N_7742,N_3662,N_2986);
xor U7743 (N_7743,N_3690,N_4663);
or U7744 (N_7744,N_809,N_1632);
nand U7745 (N_7745,N_2031,N_726);
or U7746 (N_7746,N_2631,N_25);
nand U7747 (N_7747,N_4222,N_1396);
or U7748 (N_7748,N_472,N_1934);
and U7749 (N_7749,N_2366,N_3718);
nand U7750 (N_7750,N_1877,N_4551);
or U7751 (N_7751,N_1494,N_2980);
nor U7752 (N_7752,N_256,N_334);
or U7753 (N_7753,N_2454,N_4642);
nor U7754 (N_7754,N_4596,N_2977);
nor U7755 (N_7755,N_1705,N_3680);
nor U7756 (N_7756,N_2126,N_1424);
and U7757 (N_7757,N_3725,N_2733);
or U7758 (N_7758,N_2631,N_516);
nand U7759 (N_7759,N_847,N_152);
and U7760 (N_7760,N_2052,N_3640);
nor U7761 (N_7761,N_86,N_942);
and U7762 (N_7762,N_2695,N_3136);
xnor U7763 (N_7763,N_1789,N_1745);
and U7764 (N_7764,N_66,N_2881);
or U7765 (N_7765,N_1815,N_1348);
nor U7766 (N_7766,N_1601,N_1702);
or U7767 (N_7767,N_86,N_977);
or U7768 (N_7768,N_737,N_2309);
or U7769 (N_7769,N_3201,N_2522);
nor U7770 (N_7770,N_157,N_702);
xor U7771 (N_7771,N_4778,N_314);
nand U7772 (N_7772,N_1668,N_936);
and U7773 (N_7773,N_1328,N_4998);
or U7774 (N_7774,N_3376,N_628);
nor U7775 (N_7775,N_1404,N_1074);
or U7776 (N_7776,N_651,N_4862);
nand U7777 (N_7777,N_883,N_2722);
nand U7778 (N_7778,N_1965,N_92);
and U7779 (N_7779,N_847,N_4239);
nand U7780 (N_7780,N_3247,N_980);
nor U7781 (N_7781,N_652,N_3322);
xnor U7782 (N_7782,N_427,N_3838);
and U7783 (N_7783,N_586,N_233);
xnor U7784 (N_7784,N_4750,N_4074);
nor U7785 (N_7785,N_7,N_1028);
and U7786 (N_7786,N_2717,N_4758);
or U7787 (N_7787,N_4041,N_2653);
or U7788 (N_7788,N_1943,N_2598);
and U7789 (N_7789,N_1808,N_45);
nand U7790 (N_7790,N_1988,N_3228);
nor U7791 (N_7791,N_3362,N_288);
or U7792 (N_7792,N_668,N_1201);
and U7793 (N_7793,N_3282,N_2294);
nor U7794 (N_7794,N_1478,N_2233);
and U7795 (N_7795,N_4281,N_3296);
nand U7796 (N_7796,N_185,N_4358);
nor U7797 (N_7797,N_2414,N_4718);
xor U7798 (N_7798,N_1010,N_3656);
nor U7799 (N_7799,N_2568,N_2268);
or U7800 (N_7800,N_1680,N_2261);
xor U7801 (N_7801,N_877,N_1776);
nand U7802 (N_7802,N_2710,N_4717);
or U7803 (N_7803,N_2641,N_1058);
nand U7804 (N_7804,N_4867,N_1720);
nand U7805 (N_7805,N_329,N_2998);
nor U7806 (N_7806,N_653,N_2290);
and U7807 (N_7807,N_290,N_839);
nand U7808 (N_7808,N_1016,N_1162);
or U7809 (N_7809,N_76,N_3113);
xor U7810 (N_7810,N_3431,N_957);
and U7811 (N_7811,N_3107,N_4210);
nand U7812 (N_7812,N_516,N_4449);
or U7813 (N_7813,N_1309,N_2034);
xor U7814 (N_7814,N_2704,N_1594);
nor U7815 (N_7815,N_1312,N_3564);
or U7816 (N_7816,N_4832,N_1683);
nand U7817 (N_7817,N_1933,N_2416);
or U7818 (N_7818,N_4869,N_368);
nand U7819 (N_7819,N_1644,N_1476);
or U7820 (N_7820,N_1129,N_632);
or U7821 (N_7821,N_720,N_3818);
and U7822 (N_7822,N_1537,N_3932);
or U7823 (N_7823,N_1216,N_2249);
and U7824 (N_7824,N_2825,N_2686);
or U7825 (N_7825,N_2746,N_1808);
and U7826 (N_7826,N_2054,N_533);
and U7827 (N_7827,N_3978,N_3350);
nand U7828 (N_7828,N_2915,N_4969);
or U7829 (N_7829,N_3770,N_4728);
nor U7830 (N_7830,N_3925,N_2836);
nand U7831 (N_7831,N_3149,N_4404);
xor U7832 (N_7832,N_4114,N_1004);
and U7833 (N_7833,N_1045,N_1761);
xor U7834 (N_7834,N_1721,N_4938);
nand U7835 (N_7835,N_2407,N_214);
nand U7836 (N_7836,N_2377,N_388);
xnor U7837 (N_7837,N_2129,N_3752);
xor U7838 (N_7838,N_154,N_1196);
xnor U7839 (N_7839,N_811,N_3436);
nand U7840 (N_7840,N_4542,N_3648);
or U7841 (N_7841,N_4087,N_519);
nand U7842 (N_7842,N_2872,N_1785);
or U7843 (N_7843,N_1367,N_4422);
and U7844 (N_7844,N_4382,N_1794);
and U7845 (N_7845,N_165,N_1814);
nand U7846 (N_7846,N_1344,N_1686);
nor U7847 (N_7847,N_548,N_648);
or U7848 (N_7848,N_993,N_553);
xor U7849 (N_7849,N_2381,N_738);
xor U7850 (N_7850,N_190,N_2524);
nor U7851 (N_7851,N_758,N_4737);
xor U7852 (N_7852,N_1435,N_704);
and U7853 (N_7853,N_1588,N_4832);
or U7854 (N_7854,N_973,N_1345);
xnor U7855 (N_7855,N_676,N_825);
and U7856 (N_7856,N_629,N_2743);
and U7857 (N_7857,N_698,N_2703);
and U7858 (N_7858,N_673,N_2376);
nand U7859 (N_7859,N_3322,N_1175);
nand U7860 (N_7860,N_1227,N_137);
nand U7861 (N_7861,N_2111,N_4172);
nor U7862 (N_7862,N_446,N_518);
nor U7863 (N_7863,N_134,N_3015);
xor U7864 (N_7864,N_715,N_1318);
xor U7865 (N_7865,N_3596,N_879);
and U7866 (N_7866,N_3257,N_3254);
nor U7867 (N_7867,N_4047,N_2913);
or U7868 (N_7868,N_3010,N_2353);
xor U7869 (N_7869,N_1881,N_2612);
and U7870 (N_7870,N_2031,N_1362);
or U7871 (N_7871,N_1164,N_947);
and U7872 (N_7872,N_4360,N_4108);
nand U7873 (N_7873,N_3470,N_3479);
xor U7874 (N_7874,N_4241,N_3148);
xnor U7875 (N_7875,N_1993,N_2471);
or U7876 (N_7876,N_3262,N_1887);
nand U7877 (N_7877,N_1889,N_1185);
xor U7878 (N_7878,N_3540,N_459);
nor U7879 (N_7879,N_3919,N_3679);
and U7880 (N_7880,N_2905,N_3237);
nand U7881 (N_7881,N_72,N_4758);
and U7882 (N_7882,N_1145,N_3931);
and U7883 (N_7883,N_4258,N_2681);
xnor U7884 (N_7884,N_2040,N_539);
and U7885 (N_7885,N_1610,N_1799);
nor U7886 (N_7886,N_4623,N_3561);
nor U7887 (N_7887,N_4910,N_3122);
nand U7888 (N_7888,N_4493,N_2837);
xnor U7889 (N_7889,N_1013,N_1381);
and U7890 (N_7890,N_4360,N_2945);
and U7891 (N_7891,N_3494,N_147);
and U7892 (N_7892,N_4080,N_3578);
and U7893 (N_7893,N_3392,N_2942);
nor U7894 (N_7894,N_4854,N_3660);
xnor U7895 (N_7895,N_3350,N_3239);
xnor U7896 (N_7896,N_3327,N_1557);
xnor U7897 (N_7897,N_4790,N_480);
or U7898 (N_7898,N_859,N_4716);
nand U7899 (N_7899,N_2729,N_3193);
and U7900 (N_7900,N_4403,N_889);
nand U7901 (N_7901,N_1305,N_1573);
xnor U7902 (N_7902,N_3609,N_2867);
or U7903 (N_7903,N_3345,N_81);
xnor U7904 (N_7904,N_2628,N_1949);
and U7905 (N_7905,N_957,N_1508);
or U7906 (N_7906,N_2534,N_4784);
and U7907 (N_7907,N_1313,N_1813);
nand U7908 (N_7908,N_1390,N_2519);
nand U7909 (N_7909,N_4467,N_2776);
or U7910 (N_7910,N_4098,N_2921);
nand U7911 (N_7911,N_1877,N_2504);
nand U7912 (N_7912,N_2052,N_1322);
or U7913 (N_7913,N_2117,N_1806);
nand U7914 (N_7914,N_3977,N_217);
nor U7915 (N_7915,N_1537,N_4095);
nor U7916 (N_7916,N_748,N_4075);
nor U7917 (N_7917,N_2051,N_172);
and U7918 (N_7918,N_238,N_4164);
or U7919 (N_7919,N_3289,N_1710);
xor U7920 (N_7920,N_4556,N_1413);
and U7921 (N_7921,N_227,N_471);
or U7922 (N_7922,N_4424,N_1278);
xnor U7923 (N_7923,N_1264,N_2770);
and U7924 (N_7924,N_4454,N_2054);
and U7925 (N_7925,N_4177,N_234);
or U7926 (N_7926,N_2857,N_1645);
xnor U7927 (N_7927,N_1716,N_3808);
and U7928 (N_7928,N_3193,N_1283);
nand U7929 (N_7929,N_1589,N_2506);
or U7930 (N_7930,N_952,N_4957);
or U7931 (N_7931,N_3513,N_3989);
or U7932 (N_7932,N_3439,N_2450);
and U7933 (N_7933,N_979,N_843);
xnor U7934 (N_7934,N_1631,N_4806);
nand U7935 (N_7935,N_4598,N_4023);
nand U7936 (N_7936,N_3938,N_3307);
and U7937 (N_7937,N_2182,N_2124);
or U7938 (N_7938,N_1693,N_449);
xor U7939 (N_7939,N_1912,N_3832);
nand U7940 (N_7940,N_3549,N_2383);
xnor U7941 (N_7941,N_669,N_2193);
or U7942 (N_7942,N_4406,N_1211);
xor U7943 (N_7943,N_4243,N_4982);
nand U7944 (N_7944,N_3170,N_4935);
nand U7945 (N_7945,N_3137,N_1963);
nand U7946 (N_7946,N_3332,N_3739);
xor U7947 (N_7947,N_4158,N_326);
or U7948 (N_7948,N_4933,N_1039);
and U7949 (N_7949,N_3997,N_2473);
and U7950 (N_7950,N_1642,N_4253);
nor U7951 (N_7951,N_4909,N_3821);
nor U7952 (N_7952,N_4982,N_1408);
and U7953 (N_7953,N_424,N_2422);
and U7954 (N_7954,N_3103,N_2431);
nand U7955 (N_7955,N_2735,N_471);
xnor U7956 (N_7956,N_159,N_1337);
xnor U7957 (N_7957,N_1199,N_1465);
xor U7958 (N_7958,N_3,N_2153);
or U7959 (N_7959,N_3123,N_1176);
xnor U7960 (N_7960,N_3010,N_2604);
nor U7961 (N_7961,N_2207,N_649);
and U7962 (N_7962,N_4486,N_3177);
xnor U7963 (N_7963,N_4718,N_2641);
or U7964 (N_7964,N_1243,N_303);
nor U7965 (N_7965,N_1113,N_1562);
nand U7966 (N_7966,N_3792,N_4404);
xnor U7967 (N_7967,N_4445,N_2566);
nor U7968 (N_7968,N_1760,N_4618);
nand U7969 (N_7969,N_1986,N_525);
or U7970 (N_7970,N_1631,N_3403);
or U7971 (N_7971,N_1577,N_2832);
and U7972 (N_7972,N_2404,N_4877);
nor U7973 (N_7973,N_1106,N_636);
xor U7974 (N_7974,N_4547,N_264);
and U7975 (N_7975,N_1849,N_4244);
or U7976 (N_7976,N_2513,N_3300);
nand U7977 (N_7977,N_128,N_1995);
and U7978 (N_7978,N_17,N_2185);
or U7979 (N_7979,N_685,N_1696);
or U7980 (N_7980,N_2164,N_1345);
nand U7981 (N_7981,N_4082,N_1720);
xnor U7982 (N_7982,N_394,N_4491);
or U7983 (N_7983,N_4917,N_4478);
xnor U7984 (N_7984,N_4405,N_3109);
or U7985 (N_7985,N_3753,N_4086);
xnor U7986 (N_7986,N_2513,N_3112);
nand U7987 (N_7987,N_4246,N_932);
xor U7988 (N_7988,N_4245,N_3889);
nor U7989 (N_7989,N_249,N_354);
nor U7990 (N_7990,N_3598,N_965);
or U7991 (N_7991,N_4974,N_4201);
xnor U7992 (N_7992,N_3862,N_210);
xnor U7993 (N_7993,N_3952,N_4586);
or U7994 (N_7994,N_2834,N_1197);
and U7995 (N_7995,N_3100,N_469);
or U7996 (N_7996,N_1287,N_2534);
nor U7997 (N_7997,N_4643,N_1277);
nand U7998 (N_7998,N_2844,N_4811);
nor U7999 (N_7999,N_3791,N_4195);
and U8000 (N_8000,N_1740,N_2328);
xor U8001 (N_8001,N_4933,N_2668);
xnor U8002 (N_8002,N_3460,N_3028);
xnor U8003 (N_8003,N_1784,N_435);
or U8004 (N_8004,N_4983,N_453);
nand U8005 (N_8005,N_143,N_1318);
nor U8006 (N_8006,N_4246,N_4624);
nor U8007 (N_8007,N_3806,N_1834);
or U8008 (N_8008,N_2064,N_4417);
nor U8009 (N_8009,N_34,N_2999);
nand U8010 (N_8010,N_1019,N_243);
nand U8011 (N_8011,N_2955,N_4572);
or U8012 (N_8012,N_3601,N_1349);
xnor U8013 (N_8013,N_1132,N_1680);
and U8014 (N_8014,N_1456,N_2400);
and U8015 (N_8015,N_3339,N_3047);
xor U8016 (N_8016,N_62,N_916);
nor U8017 (N_8017,N_2679,N_442);
xnor U8018 (N_8018,N_2593,N_3946);
nand U8019 (N_8019,N_4181,N_4045);
xnor U8020 (N_8020,N_376,N_3521);
nand U8021 (N_8021,N_4122,N_3657);
or U8022 (N_8022,N_4588,N_783);
or U8023 (N_8023,N_2187,N_3176);
nor U8024 (N_8024,N_317,N_4772);
or U8025 (N_8025,N_1322,N_1622);
or U8026 (N_8026,N_4248,N_1041);
xnor U8027 (N_8027,N_480,N_4075);
or U8028 (N_8028,N_3825,N_2166);
nor U8029 (N_8029,N_3960,N_3404);
xor U8030 (N_8030,N_1941,N_1609);
or U8031 (N_8031,N_3712,N_1596);
nand U8032 (N_8032,N_249,N_4740);
xnor U8033 (N_8033,N_2501,N_2246);
nand U8034 (N_8034,N_1357,N_1589);
nor U8035 (N_8035,N_1211,N_4215);
nor U8036 (N_8036,N_778,N_4177);
nand U8037 (N_8037,N_211,N_824);
and U8038 (N_8038,N_2852,N_1565);
xor U8039 (N_8039,N_2029,N_4273);
nand U8040 (N_8040,N_3156,N_2896);
xnor U8041 (N_8041,N_841,N_3587);
xnor U8042 (N_8042,N_1192,N_2116);
or U8043 (N_8043,N_4422,N_1116);
xor U8044 (N_8044,N_2594,N_3212);
xnor U8045 (N_8045,N_3158,N_3157);
nand U8046 (N_8046,N_546,N_989);
and U8047 (N_8047,N_4928,N_4107);
nand U8048 (N_8048,N_87,N_1891);
or U8049 (N_8049,N_256,N_4212);
xor U8050 (N_8050,N_1344,N_2399);
nand U8051 (N_8051,N_1923,N_4996);
nor U8052 (N_8052,N_3795,N_4926);
or U8053 (N_8053,N_1842,N_1449);
nor U8054 (N_8054,N_476,N_3689);
nand U8055 (N_8055,N_100,N_4571);
nand U8056 (N_8056,N_2778,N_3040);
or U8057 (N_8057,N_1524,N_1511);
or U8058 (N_8058,N_1388,N_3600);
and U8059 (N_8059,N_1902,N_4043);
nand U8060 (N_8060,N_3113,N_4654);
or U8061 (N_8061,N_1060,N_903);
xor U8062 (N_8062,N_3679,N_3066);
xnor U8063 (N_8063,N_1491,N_2083);
nor U8064 (N_8064,N_217,N_1062);
nand U8065 (N_8065,N_872,N_491);
nor U8066 (N_8066,N_762,N_90);
or U8067 (N_8067,N_800,N_4180);
or U8068 (N_8068,N_837,N_4130);
nand U8069 (N_8069,N_1199,N_2775);
nor U8070 (N_8070,N_4332,N_2523);
xor U8071 (N_8071,N_3743,N_2192);
xnor U8072 (N_8072,N_4091,N_1);
and U8073 (N_8073,N_3572,N_1997);
xnor U8074 (N_8074,N_132,N_3070);
nor U8075 (N_8075,N_4468,N_1554);
nand U8076 (N_8076,N_2145,N_4951);
nand U8077 (N_8077,N_621,N_3291);
nor U8078 (N_8078,N_1330,N_1240);
or U8079 (N_8079,N_345,N_1298);
and U8080 (N_8080,N_1720,N_1379);
and U8081 (N_8081,N_4984,N_3648);
nor U8082 (N_8082,N_55,N_1826);
nand U8083 (N_8083,N_2456,N_2212);
nor U8084 (N_8084,N_4399,N_742);
nand U8085 (N_8085,N_1173,N_2296);
nand U8086 (N_8086,N_1798,N_1369);
nor U8087 (N_8087,N_637,N_4341);
or U8088 (N_8088,N_2639,N_310);
nor U8089 (N_8089,N_4257,N_1865);
and U8090 (N_8090,N_3557,N_4881);
nor U8091 (N_8091,N_1535,N_508);
and U8092 (N_8092,N_568,N_3902);
nor U8093 (N_8093,N_3956,N_514);
nand U8094 (N_8094,N_366,N_4722);
xor U8095 (N_8095,N_1328,N_2184);
and U8096 (N_8096,N_2548,N_4880);
xnor U8097 (N_8097,N_1138,N_4455);
and U8098 (N_8098,N_1847,N_1825);
nand U8099 (N_8099,N_3921,N_1467);
and U8100 (N_8100,N_2696,N_65);
nand U8101 (N_8101,N_3840,N_4756);
nand U8102 (N_8102,N_1770,N_3589);
nor U8103 (N_8103,N_4700,N_3027);
xor U8104 (N_8104,N_2078,N_4144);
xor U8105 (N_8105,N_1990,N_1359);
nor U8106 (N_8106,N_4633,N_4019);
and U8107 (N_8107,N_455,N_245);
and U8108 (N_8108,N_2091,N_1822);
nor U8109 (N_8109,N_368,N_2168);
and U8110 (N_8110,N_3386,N_585);
xor U8111 (N_8111,N_634,N_750);
nor U8112 (N_8112,N_4230,N_2084);
and U8113 (N_8113,N_2015,N_3333);
nor U8114 (N_8114,N_4505,N_4414);
nor U8115 (N_8115,N_586,N_3713);
and U8116 (N_8116,N_4490,N_1097);
nand U8117 (N_8117,N_1537,N_4431);
nand U8118 (N_8118,N_3547,N_2211);
xnor U8119 (N_8119,N_1474,N_1773);
nor U8120 (N_8120,N_3676,N_3662);
nand U8121 (N_8121,N_2351,N_2826);
and U8122 (N_8122,N_3044,N_3297);
and U8123 (N_8123,N_4959,N_1743);
xor U8124 (N_8124,N_2678,N_2366);
nor U8125 (N_8125,N_2096,N_2749);
and U8126 (N_8126,N_4053,N_4227);
or U8127 (N_8127,N_3633,N_4321);
xnor U8128 (N_8128,N_455,N_3638);
xor U8129 (N_8129,N_1641,N_2261);
nand U8130 (N_8130,N_4229,N_1576);
nand U8131 (N_8131,N_132,N_560);
nor U8132 (N_8132,N_4341,N_3147);
or U8133 (N_8133,N_3058,N_3841);
nor U8134 (N_8134,N_4624,N_3540);
nand U8135 (N_8135,N_715,N_1889);
nand U8136 (N_8136,N_1287,N_199);
nor U8137 (N_8137,N_3173,N_3243);
and U8138 (N_8138,N_2064,N_4602);
or U8139 (N_8139,N_2566,N_310);
xnor U8140 (N_8140,N_2474,N_3860);
nor U8141 (N_8141,N_966,N_4);
nor U8142 (N_8142,N_1206,N_4410);
and U8143 (N_8143,N_4644,N_947);
xnor U8144 (N_8144,N_498,N_3428);
nand U8145 (N_8145,N_2335,N_833);
nand U8146 (N_8146,N_2217,N_4087);
nor U8147 (N_8147,N_2710,N_1250);
and U8148 (N_8148,N_3773,N_3071);
nor U8149 (N_8149,N_2097,N_4496);
xor U8150 (N_8150,N_2466,N_3182);
and U8151 (N_8151,N_2905,N_419);
and U8152 (N_8152,N_3675,N_1762);
nand U8153 (N_8153,N_3662,N_3087);
or U8154 (N_8154,N_2987,N_3595);
nand U8155 (N_8155,N_3994,N_2319);
or U8156 (N_8156,N_3111,N_4474);
and U8157 (N_8157,N_738,N_799);
xnor U8158 (N_8158,N_4273,N_290);
nor U8159 (N_8159,N_520,N_670);
or U8160 (N_8160,N_3879,N_2955);
nor U8161 (N_8161,N_3061,N_4031);
and U8162 (N_8162,N_879,N_1104);
or U8163 (N_8163,N_1088,N_1172);
or U8164 (N_8164,N_4558,N_4086);
xor U8165 (N_8165,N_3322,N_207);
or U8166 (N_8166,N_492,N_4309);
nor U8167 (N_8167,N_1109,N_2273);
xnor U8168 (N_8168,N_840,N_1649);
nor U8169 (N_8169,N_3135,N_2711);
nand U8170 (N_8170,N_1801,N_1565);
or U8171 (N_8171,N_4264,N_1990);
and U8172 (N_8172,N_2867,N_631);
nand U8173 (N_8173,N_3726,N_4528);
xnor U8174 (N_8174,N_2366,N_3063);
or U8175 (N_8175,N_663,N_2606);
nand U8176 (N_8176,N_3893,N_4833);
nand U8177 (N_8177,N_619,N_1631);
and U8178 (N_8178,N_4013,N_3775);
nor U8179 (N_8179,N_1123,N_3211);
nor U8180 (N_8180,N_1095,N_3141);
nand U8181 (N_8181,N_180,N_2067);
and U8182 (N_8182,N_4887,N_1095);
nand U8183 (N_8183,N_2350,N_4520);
nor U8184 (N_8184,N_100,N_4586);
xnor U8185 (N_8185,N_1391,N_740);
nand U8186 (N_8186,N_4657,N_3379);
xnor U8187 (N_8187,N_97,N_4025);
and U8188 (N_8188,N_3687,N_1103);
nor U8189 (N_8189,N_766,N_3636);
nand U8190 (N_8190,N_467,N_1911);
nand U8191 (N_8191,N_762,N_2311);
xnor U8192 (N_8192,N_1255,N_1039);
nor U8193 (N_8193,N_1472,N_2191);
nand U8194 (N_8194,N_222,N_307);
or U8195 (N_8195,N_2102,N_1498);
nand U8196 (N_8196,N_353,N_1918);
xor U8197 (N_8197,N_3836,N_3308);
and U8198 (N_8198,N_648,N_1055);
nor U8199 (N_8199,N_1080,N_4757);
or U8200 (N_8200,N_966,N_1724);
and U8201 (N_8201,N_1253,N_711);
xor U8202 (N_8202,N_3881,N_2234);
nor U8203 (N_8203,N_4881,N_307);
nand U8204 (N_8204,N_2590,N_1528);
and U8205 (N_8205,N_2080,N_4304);
nand U8206 (N_8206,N_3364,N_4912);
nor U8207 (N_8207,N_3115,N_348);
nor U8208 (N_8208,N_590,N_244);
and U8209 (N_8209,N_2639,N_2733);
nor U8210 (N_8210,N_3279,N_34);
nand U8211 (N_8211,N_4906,N_2361);
nand U8212 (N_8212,N_2752,N_3022);
or U8213 (N_8213,N_2377,N_3384);
or U8214 (N_8214,N_2921,N_462);
nand U8215 (N_8215,N_4664,N_2301);
and U8216 (N_8216,N_4203,N_562);
xor U8217 (N_8217,N_2408,N_1502);
xnor U8218 (N_8218,N_3273,N_47);
nor U8219 (N_8219,N_4841,N_3336);
or U8220 (N_8220,N_2502,N_1967);
or U8221 (N_8221,N_428,N_1671);
nand U8222 (N_8222,N_414,N_4438);
xor U8223 (N_8223,N_162,N_1645);
nor U8224 (N_8224,N_3902,N_3448);
xor U8225 (N_8225,N_1417,N_1309);
nand U8226 (N_8226,N_795,N_1039);
nand U8227 (N_8227,N_1594,N_444);
or U8228 (N_8228,N_2143,N_1776);
xor U8229 (N_8229,N_4032,N_4953);
nand U8230 (N_8230,N_475,N_1896);
nand U8231 (N_8231,N_2319,N_107);
or U8232 (N_8232,N_2653,N_4204);
xor U8233 (N_8233,N_4613,N_113);
nand U8234 (N_8234,N_2823,N_1194);
or U8235 (N_8235,N_3842,N_3427);
nor U8236 (N_8236,N_3773,N_772);
and U8237 (N_8237,N_178,N_973);
nor U8238 (N_8238,N_2730,N_2396);
or U8239 (N_8239,N_1935,N_3848);
and U8240 (N_8240,N_2854,N_537);
and U8241 (N_8241,N_3738,N_4092);
nor U8242 (N_8242,N_2721,N_2156);
and U8243 (N_8243,N_747,N_1153);
nor U8244 (N_8244,N_2192,N_1993);
xnor U8245 (N_8245,N_4584,N_246);
xor U8246 (N_8246,N_1412,N_4437);
or U8247 (N_8247,N_3228,N_3051);
nor U8248 (N_8248,N_4685,N_2036);
or U8249 (N_8249,N_2116,N_1919);
and U8250 (N_8250,N_4230,N_4713);
and U8251 (N_8251,N_690,N_1978);
xnor U8252 (N_8252,N_2374,N_1588);
and U8253 (N_8253,N_1481,N_3148);
and U8254 (N_8254,N_4250,N_70);
or U8255 (N_8255,N_1902,N_1264);
nor U8256 (N_8256,N_3652,N_69);
xor U8257 (N_8257,N_438,N_85);
and U8258 (N_8258,N_3829,N_4602);
and U8259 (N_8259,N_2626,N_2597);
or U8260 (N_8260,N_1790,N_16);
and U8261 (N_8261,N_431,N_1855);
xnor U8262 (N_8262,N_14,N_2079);
or U8263 (N_8263,N_80,N_333);
and U8264 (N_8264,N_3473,N_3965);
and U8265 (N_8265,N_3237,N_1044);
or U8266 (N_8266,N_3883,N_3810);
xnor U8267 (N_8267,N_1219,N_2396);
nand U8268 (N_8268,N_3984,N_4066);
nand U8269 (N_8269,N_4188,N_3552);
and U8270 (N_8270,N_4434,N_2284);
or U8271 (N_8271,N_1214,N_1909);
and U8272 (N_8272,N_1662,N_4645);
and U8273 (N_8273,N_2165,N_3354);
nor U8274 (N_8274,N_1953,N_3809);
and U8275 (N_8275,N_1800,N_1007);
and U8276 (N_8276,N_4533,N_2523);
xnor U8277 (N_8277,N_2737,N_4676);
or U8278 (N_8278,N_976,N_3914);
nor U8279 (N_8279,N_2276,N_3082);
nand U8280 (N_8280,N_2224,N_1161);
or U8281 (N_8281,N_199,N_2808);
and U8282 (N_8282,N_2714,N_2916);
and U8283 (N_8283,N_647,N_2290);
and U8284 (N_8284,N_3360,N_4937);
nor U8285 (N_8285,N_891,N_673);
and U8286 (N_8286,N_2646,N_2022);
or U8287 (N_8287,N_3945,N_4644);
or U8288 (N_8288,N_4405,N_4755);
or U8289 (N_8289,N_3085,N_4285);
or U8290 (N_8290,N_2505,N_3270);
xnor U8291 (N_8291,N_4817,N_4989);
nor U8292 (N_8292,N_37,N_2648);
and U8293 (N_8293,N_4077,N_4930);
xor U8294 (N_8294,N_1720,N_3497);
and U8295 (N_8295,N_2478,N_949);
or U8296 (N_8296,N_4044,N_1065);
xor U8297 (N_8297,N_298,N_630);
xor U8298 (N_8298,N_1028,N_4726);
nor U8299 (N_8299,N_2476,N_3346);
or U8300 (N_8300,N_4651,N_1174);
nor U8301 (N_8301,N_3280,N_1890);
and U8302 (N_8302,N_752,N_4104);
nand U8303 (N_8303,N_3096,N_4460);
xnor U8304 (N_8304,N_706,N_3584);
nor U8305 (N_8305,N_2552,N_3784);
and U8306 (N_8306,N_201,N_1570);
xnor U8307 (N_8307,N_782,N_4674);
nand U8308 (N_8308,N_3874,N_245);
or U8309 (N_8309,N_337,N_4973);
and U8310 (N_8310,N_4119,N_4092);
nor U8311 (N_8311,N_4423,N_3165);
nor U8312 (N_8312,N_1694,N_3332);
nand U8313 (N_8313,N_2584,N_369);
or U8314 (N_8314,N_4621,N_3631);
and U8315 (N_8315,N_4252,N_3427);
nand U8316 (N_8316,N_2258,N_3801);
or U8317 (N_8317,N_3640,N_4923);
xnor U8318 (N_8318,N_2515,N_3811);
xnor U8319 (N_8319,N_1930,N_2203);
and U8320 (N_8320,N_2091,N_4868);
nand U8321 (N_8321,N_4319,N_9);
or U8322 (N_8322,N_4302,N_2888);
or U8323 (N_8323,N_36,N_943);
xor U8324 (N_8324,N_711,N_446);
or U8325 (N_8325,N_1639,N_375);
or U8326 (N_8326,N_1018,N_2676);
nor U8327 (N_8327,N_435,N_1956);
nor U8328 (N_8328,N_100,N_3128);
and U8329 (N_8329,N_2498,N_3740);
nor U8330 (N_8330,N_4909,N_807);
nor U8331 (N_8331,N_3810,N_399);
nor U8332 (N_8332,N_4961,N_3574);
or U8333 (N_8333,N_2880,N_3517);
and U8334 (N_8334,N_3898,N_293);
xor U8335 (N_8335,N_1468,N_2528);
and U8336 (N_8336,N_4944,N_2478);
nor U8337 (N_8337,N_4798,N_4466);
and U8338 (N_8338,N_2850,N_1508);
nand U8339 (N_8339,N_2234,N_2573);
nand U8340 (N_8340,N_3548,N_526);
nand U8341 (N_8341,N_2838,N_4386);
or U8342 (N_8342,N_4766,N_871);
and U8343 (N_8343,N_2357,N_762);
nor U8344 (N_8344,N_2317,N_1345);
nand U8345 (N_8345,N_2962,N_200);
or U8346 (N_8346,N_281,N_1612);
and U8347 (N_8347,N_1364,N_2133);
and U8348 (N_8348,N_4348,N_4806);
or U8349 (N_8349,N_1116,N_3176);
or U8350 (N_8350,N_3631,N_1845);
xnor U8351 (N_8351,N_4678,N_313);
xor U8352 (N_8352,N_78,N_2646);
nor U8353 (N_8353,N_1470,N_373);
xor U8354 (N_8354,N_4382,N_3850);
or U8355 (N_8355,N_4388,N_4429);
and U8356 (N_8356,N_1217,N_4445);
or U8357 (N_8357,N_1029,N_1360);
nor U8358 (N_8358,N_676,N_3733);
xnor U8359 (N_8359,N_894,N_2369);
xor U8360 (N_8360,N_694,N_2753);
and U8361 (N_8361,N_6,N_4435);
or U8362 (N_8362,N_2569,N_4726);
xor U8363 (N_8363,N_4267,N_2209);
and U8364 (N_8364,N_3324,N_1986);
nor U8365 (N_8365,N_223,N_1981);
nand U8366 (N_8366,N_1855,N_1356);
xor U8367 (N_8367,N_1987,N_2189);
or U8368 (N_8368,N_111,N_2762);
nand U8369 (N_8369,N_2620,N_2006);
nor U8370 (N_8370,N_2971,N_1924);
nor U8371 (N_8371,N_521,N_989);
nor U8372 (N_8372,N_2659,N_1848);
and U8373 (N_8373,N_2583,N_628);
or U8374 (N_8374,N_1891,N_4849);
xor U8375 (N_8375,N_2244,N_2103);
nor U8376 (N_8376,N_247,N_595);
or U8377 (N_8377,N_2675,N_992);
and U8378 (N_8378,N_3372,N_2917);
nand U8379 (N_8379,N_3820,N_1456);
nor U8380 (N_8380,N_3756,N_96);
nor U8381 (N_8381,N_3837,N_3432);
xnor U8382 (N_8382,N_3300,N_3679);
and U8383 (N_8383,N_1577,N_4008);
nand U8384 (N_8384,N_2277,N_2496);
or U8385 (N_8385,N_0,N_4558);
or U8386 (N_8386,N_4172,N_3716);
and U8387 (N_8387,N_4745,N_1099);
and U8388 (N_8388,N_2112,N_1157);
nor U8389 (N_8389,N_1443,N_3770);
nand U8390 (N_8390,N_1553,N_4169);
nand U8391 (N_8391,N_158,N_1739);
or U8392 (N_8392,N_714,N_4423);
and U8393 (N_8393,N_2130,N_3598);
nor U8394 (N_8394,N_1156,N_2814);
xor U8395 (N_8395,N_4616,N_3276);
nor U8396 (N_8396,N_1652,N_951);
and U8397 (N_8397,N_4804,N_537);
nor U8398 (N_8398,N_1620,N_3619);
and U8399 (N_8399,N_193,N_1679);
nand U8400 (N_8400,N_4523,N_3318);
xor U8401 (N_8401,N_1293,N_3693);
xor U8402 (N_8402,N_3383,N_991);
xnor U8403 (N_8403,N_751,N_3732);
or U8404 (N_8404,N_2344,N_1053);
and U8405 (N_8405,N_1210,N_4113);
or U8406 (N_8406,N_907,N_1273);
nor U8407 (N_8407,N_675,N_563);
nand U8408 (N_8408,N_209,N_3201);
xor U8409 (N_8409,N_2375,N_1657);
xor U8410 (N_8410,N_2542,N_3496);
xnor U8411 (N_8411,N_805,N_4141);
and U8412 (N_8412,N_3304,N_1331);
and U8413 (N_8413,N_1832,N_2562);
nand U8414 (N_8414,N_311,N_3048);
or U8415 (N_8415,N_3366,N_4314);
and U8416 (N_8416,N_2678,N_2942);
nor U8417 (N_8417,N_2757,N_2937);
or U8418 (N_8418,N_566,N_63);
or U8419 (N_8419,N_2509,N_501);
xnor U8420 (N_8420,N_1580,N_4870);
or U8421 (N_8421,N_1259,N_4705);
nor U8422 (N_8422,N_2906,N_2186);
and U8423 (N_8423,N_2947,N_926);
xnor U8424 (N_8424,N_2798,N_1129);
xor U8425 (N_8425,N_4378,N_1265);
nand U8426 (N_8426,N_431,N_2793);
or U8427 (N_8427,N_852,N_4716);
nor U8428 (N_8428,N_2970,N_2632);
and U8429 (N_8429,N_2509,N_3983);
nor U8430 (N_8430,N_3624,N_682);
nand U8431 (N_8431,N_2858,N_409);
or U8432 (N_8432,N_2116,N_4337);
and U8433 (N_8433,N_2170,N_3922);
and U8434 (N_8434,N_1939,N_1993);
nand U8435 (N_8435,N_723,N_1330);
nor U8436 (N_8436,N_3970,N_216);
and U8437 (N_8437,N_3118,N_4523);
and U8438 (N_8438,N_1163,N_3725);
and U8439 (N_8439,N_1383,N_3770);
or U8440 (N_8440,N_4845,N_1073);
nand U8441 (N_8441,N_1976,N_2721);
nor U8442 (N_8442,N_2367,N_291);
nand U8443 (N_8443,N_2016,N_626);
xnor U8444 (N_8444,N_3576,N_4703);
xnor U8445 (N_8445,N_4831,N_286);
nor U8446 (N_8446,N_4162,N_1343);
xnor U8447 (N_8447,N_1402,N_2734);
nor U8448 (N_8448,N_271,N_4808);
or U8449 (N_8449,N_1375,N_459);
nand U8450 (N_8450,N_3077,N_1641);
nand U8451 (N_8451,N_194,N_295);
and U8452 (N_8452,N_83,N_4879);
nand U8453 (N_8453,N_3000,N_31);
or U8454 (N_8454,N_2892,N_1285);
nor U8455 (N_8455,N_2753,N_444);
nand U8456 (N_8456,N_4510,N_3054);
and U8457 (N_8457,N_620,N_4386);
and U8458 (N_8458,N_117,N_3663);
nand U8459 (N_8459,N_3514,N_787);
xor U8460 (N_8460,N_3681,N_2820);
or U8461 (N_8461,N_3808,N_2854);
nand U8462 (N_8462,N_1927,N_3168);
xor U8463 (N_8463,N_1960,N_2556);
nand U8464 (N_8464,N_4650,N_2032);
xor U8465 (N_8465,N_2649,N_3870);
nor U8466 (N_8466,N_1009,N_1606);
and U8467 (N_8467,N_3644,N_3850);
xor U8468 (N_8468,N_1976,N_3371);
nor U8469 (N_8469,N_786,N_4747);
and U8470 (N_8470,N_2048,N_1546);
nand U8471 (N_8471,N_2185,N_4614);
nand U8472 (N_8472,N_2548,N_3594);
or U8473 (N_8473,N_3270,N_1736);
nor U8474 (N_8474,N_1743,N_812);
and U8475 (N_8475,N_4609,N_4568);
or U8476 (N_8476,N_833,N_109);
nor U8477 (N_8477,N_992,N_4938);
or U8478 (N_8478,N_308,N_637);
nand U8479 (N_8479,N_4880,N_4088);
nor U8480 (N_8480,N_4438,N_1318);
nor U8481 (N_8481,N_4134,N_1385);
or U8482 (N_8482,N_3734,N_2816);
or U8483 (N_8483,N_440,N_4172);
or U8484 (N_8484,N_3360,N_4017);
xor U8485 (N_8485,N_4290,N_18);
nand U8486 (N_8486,N_2859,N_1696);
nand U8487 (N_8487,N_3257,N_1763);
and U8488 (N_8488,N_1424,N_2741);
and U8489 (N_8489,N_4285,N_4722);
and U8490 (N_8490,N_1279,N_1483);
nand U8491 (N_8491,N_3482,N_4737);
xor U8492 (N_8492,N_3037,N_636);
nor U8493 (N_8493,N_3197,N_471);
nor U8494 (N_8494,N_4352,N_2419);
or U8495 (N_8495,N_1679,N_4764);
or U8496 (N_8496,N_1672,N_3821);
and U8497 (N_8497,N_970,N_3889);
xor U8498 (N_8498,N_19,N_1212);
nor U8499 (N_8499,N_4041,N_3665);
nor U8500 (N_8500,N_1740,N_4056);
or U8501 (N_8501,N_1139,N_1445);
xnor U8502 (N_8502,N_2539,N_728);
and U8503 (N_8503,N_4159,N_916);
and U8504 (N_8504,N_4133,N_2592);
or U8505 (N_8505,N_884,N_3601);
nand U8506 (N_8506,N_2102,N_3196);
and U8507 (N_8507,N_2074,N_1045);
or U8508 (N_8508,N_4702,N_1569);
and U8509 (N_8509,N_4766,N_30);
and U8510 (N_8510,N_2566,N_1751);
or U8511 (N_8511,N_937,N_403);
nand U8512 (N_8512,N_415,N_1588);
and U8513 (N_8513,N_4562,N_4897);
or U8514 (N_8514,N_824,N_1335);
xnor U8515 (N_8515,N_1966,N_1464);
nor U8516 (N_8516,N_3107,N_2214);
nand U8517 (N_8517,N_2384,N_803);
and U8518 (N_8518,N_3716,N_1549);
or U8519 (N_8519,N_2764,N_1604);
nand U8520 (N_8520,N_1360,N_268);
xor U8521 (N_8521,N_2847,N_3214);
xnor U8522 (N_8522,N_2187,N_816);
and U8523 (N_8523,N_2945,N_3117);
nor U8524 (N_8524,N_2046,N_3273);
nand U8525 (N_8525,N_4422,N_1397);
and U8526 (N_8526,N_716,N_3087);
xnor U8527 (N_8527,N_4749,N_4174);
and U8528 (N_8528,N_2530,N_3783);
and U8529 (N_8529,N_1145,N_4201);
or U8530 (N_8530,N_497,N_4999);
nand U8531 (N_8531,N_4586,N_174);
and U8532 (N_8532,N_2788,N_4896);
nor U8533 (N_8533,N_1216,N_4211);
or U8534 (N_8534,N_2945,N_4814);
nor U8535 (N_8535,N_992,N_1200);
nand U8536 (N_8536,N_2059,N_2389);
or U8537 (N_8537,N_182,N_2177);
nor U8538 (N_8538,N_1103,N_257);
xor U8539 (N_8539,N_115,N_1229);
xnor U8540 (N_8540,N_3648,N_3154);
nand U8541 (N_8541,N_3909,N_4295);
xor U8542 (N_8542,N_4518,N_1798);
nand U8543 (N_8543,N_143,N_892);
nand U8544 (N_8544,N_841,N_1854);
nor U8545 (N_8545,N_3133,N_3100);
xnor U8546 (N_8546,N_2368,N_3193);
nand U8547 (N_8547,N_4570,N_1212);
nand U8548 (N_8548,N_1525,N_2511);
nand U8549 (N_8549,N_116,N_2447);
nor U8550 (N_8550,N_399,N_571);
xor U8551 (N_8551,N_4378,N_4187);
xnor U8552 (N_8552,N_2319,N_1614);
nor U8553 (N_8553,N_4694,N_3936);
and U8554 (N_8554,N_615,N_1977);
xor U8555 (N_8555,N_3070,N_1859);
nand U8556 (N_8556,N_3212,N_1991);
nor U8557 (N_8557,N_4904,N_3813);
nand U8558 (N_8558,N_2606,N_3408);
and U8559 (N_8559,N_2418,N_3725);
and U8560 (N_8560,N_3595,N_2948);
or U8561 (N_8561,N_2405,N_3580);
and U8562 (N_8562,N_1403,N_1462);
or U8563 (N_8563,N_3638,N_2593);
or U8564 (N_8564,N_3638,N_3636);
nand U8565 (N_8565,N_4818,N_3597);
or U8566 (N_8566,N_3521,N_3391);
and U8567 (N_8567,N_2366,N_4615);
and U8568 (N_8568,N_4047,N_2324);
nand U8569 (N_8569,N_4921,N_3379);
or U8570 (N_8570,N_939,N_4244);
and U8571 (N_8571,N_273,N_3837);
or U8572 (N_8572,N_701,N_1588);
and U8573 (N_8573,N_317,N_2936);
or U8574 (N_8574,N_3269,N_2424);
or U8575 (N_8575,N_932,N_1294);
nor U8576 (N_8576,N_3221,N_541);
or U8577 (N_8577,N_1924,N_2931);
xnor U8578 (N_8578,N_2344,N_82);
or U8579 (N_8579,N_4440,N_70);
or U8580 (N_8580,N_999,N_3477);
and U8581 (N_8581,N_1625,N_3374);
or U8582 (N_8582,N_2911,N_766);
and U8583 (N_8583,N_3420,N_2353);
nor U8584 (N_8584,N_3951,N_4837);
xnor U8585 (N_8585,N_2417,N_593);
and U8586 (N_8586,N_4572,N_1890);
nand U8587 (N_8587,N_3107,N_2928);
nand U8588 (N_8588,N_4984,N_1559);
nor U8589 (N_8589,N_3700,N_608);
or U8590 (N_8590,N_677,N_2629);
xnor U8591 (N_8591,N_1380,N_471);
nand U8592 (N_8592,N_4329,N_635);
xnor U8593 (N_8593,N_2292,N_6);
xor U8594 (N_8594,N_832,N_4981);
and U8595 (N_8595,N_4319,N_3588);
nor U8596 (N_8596,N_3508,N_3650);
and U8597 (N_8597,N_4189,N_2420);
nor U8598 (N_8598,N_1016,N_2409);
or U8599 (N_8599,N_2718,N_19);
or U8600 (N_8600,N_2092,N_2365);
nand U8601 (N_8601,N_4430,N_3365);
or U8602 (N_8602,N_3432,N_2584);
xnor U8603 (N_8603,N_2281,N_1163);
and U8604 (N_8604,N_3446,N_1033);
xnor U8605 (N_8605,N_3051,N_1535);
xor U8606 (N_8606,N_2873,N_652);
nand U8607 (N_8607,N_1541,N_1179);
nor U8608 (N_8608,N_2513,N_2463);
or U8609 (N_8609,N_1412,N_3634);
or U8610 (N_8610,N_3813,N_2664);
xnor U8611 (N_8611,N_33,N_3247);
nor U8612 (N_8612,N_3515,N_975);
nor U8613 (N_8613,N_389,N_4323);
and U8614 (N_8614,N_112,N_3293);
nor U8615 (N_8615,N_3633,N_4553);
and U8616 (N_8616,N_4049,N_3978);
nand U8617 (N_8617,N_4379,N_740);
and U8618 (N_8618,N_4943,N_552);
or U8619 (N_8619,N_3193,N_4682);
or U8620 (N_8620,N_2073,N_1951);
and U8621 (N_8621,N_3612,N_4853);
and U8622 (N_8622,N_1203,N_4056);
or U8623 (N_8623,N_1881,N_3956);
xor U8624 (N_8624,N_4933,N_4801);
xnor U8625 (N_8625,N_3567,N_2236);
xor U8626 (N_8626,N_2086,N_3775);
nand U8627 (N_8627,N_1602,N_2744);
xnor U8628 (N_8628,N_2540,N_258);
xor U8629 (N_8629,N_1335,N_3529);
nor U8630 (N_8630,N_591,N_4260);
or U8631 (N_8631,N_4549,N_4823);
xnor U8632 (N_8632,N_4326,N_2679);
nand U8633 (N_8633,N_2008,N_3570);
nor U8634 (N_8634,N_1026,N_1541);
nor U8635 (N_8635,N_249,N_1204);
nand U8636 (N_8636,N_1608,N_619);
or U8637 (N_8637,N_3471,N_2076);
and U8638 (N_8638,N_4525,N_256);
and U8639 (N_8639,N_4068,N_925);
or U8640 (N_8640,N_4878,N_296);
xnor U8641 (N_8641,N_1474,N_121);
xor U8642 (N_8642,N_1412,N_1073);
xnor U8643 (N_8643,N_1893,N_4256);
xnor U8644 (N_8644,N_4383,N_2454);
xnor U8645 (N_8645,N_4237,N_2041);
nor U8646 (N_8646,N_3484,N_1581);
nor U8647 (N_8647,N_904,N_1540);
and U8648 (N_8648,N_2021,N_206);
or U8649 (N_8649,N_3132,N_908);
nand U8650 (N_8650,N_3526,N_2304);
or U8651 (N_8651,N_1842,N_459);
nor U8652 (N_8652,N_3165,N_716);
or U8653 (N_8653,N_4521,N_3112);
and U8654 (N_8654,N_3204,N_2723);
or U8655 (N_8655,N_3267,N_2531);
nor U8656 (N_8656,N_2300,N_2188);
nor U8657 (N_8657,N_1784,N_2298);
xnor U8658 (N_8658,N_1574,N_3091);
nor U8659 (N_8659,N_1729,N_2588);
and U8660 (N_8660,N_4387,N_2578);
nand U8661 (N_8661,N_1386,N_3222);
nand U8662 (N_8662,N_4814,N_1400);
or U8663 (N_8663,N_4616,N_4840);
nor U8664 (N_8664,N_2131,N_3094);
or U8665 (N_8665,N_3782,N_4611);
nand U8666 (N_8666,N_438,N_451);
nand U8667 (N_8667,N_3630,N_1618);
xnor U8668 (N_8668,N_3391,N_1177);
and U8669 (N_8669,N_1426,N_792);
and U8670 (N_8670,N_774,N_736);
and U8671 (N_8671,N_2002,N_2702);
or U8672 (N_8672,N_3854,N_2326);
nor U8673 (N_8673,N_4739,N_531);
nand U8674 (N_8674,N_1591,N_2375);
nand U8675 (N_8675,N_2212,N_4050);
nand U8676 (N_8676,N_3161,N_3145);
nand U8677 (N_8677,N_4968,N_1095);
nor U8678 (N_8678,N_1632,N_4598);
nor U8679 (N_8679,N_3638,N_2061);
nor U8680 (N_8680,N_4961,N_2267);
and U8681 (N_8681,N_2900,N_4923);
or U8682 (N_8682,N_633,N_1304);
nand U8683 (N_8683,N_2953,N_1017);
nor U8684 (N_8684,N_395,N_3313);
nor U8685 (N_8685,N_4201,N_1614);
nand U8686 (N_8686,N_654,N_2468);
and U8687 (N_8687,N_1804,N_1260);
nor U8688 (N_8688,N_177,N_1512);
xnor U8689 (N_8689,N_3763,N_709);
or U8690 (N_8690,N_1636,N_2866);
xnor U8691 (N_8691,N_1438,N_3319);
nor U8692 (N_8692,N_2532,N_885);
or U8693 (N_8693,N_211,N_3301);
xnor U8694 (N_8694,N_4490,N_2375);
nand U8695 (N_8695,N_916,N_2744);
or U8696 (N_8696,N_1038,N_2770);
and U8697 (N_8697,N_4976,N_3976);
xnor U8698 (N_8698,N_1753,N_3555);
xnor U8699 (N_8699,N_1912,N_2179);
or U8700 (N_8700,N_4588,N_1586);
and U8701 (N_8701,N_2970,N_2665);
nor U8702 (N_8702,N_4128,N_2805);
nor U8703 (N_8703,N_836,N_3062);
or U8704 (N_8704,N_2407,N_2616);
nand U8705 (N_8705,N_2228,N_1788);
nand U8706 (N_8706,N_1024,N_4666);
and U8707 (N_8707,N_3411,N_2821);
or U8708 (N_8708,N_4683,N_4113);
and U8709 (N_8709,N_2098,N_2517);
xnor U8710 (N_8710,N_214,N_3963);
xor U8711 (N_8711,N_3779,N_364);
nand U8712 (N_8712,N_3932,N_547);
and U8713 (N_8713,N_2589,N_2520);
nand U8714 (N_8714,N_3984,N_1832);
xor U8715 (N_8715,N_565,N_4743);
and U8716 (N_8716,N_602,N_4170);
nor U8717 (N_8717,N_3093,N_4824);
xor U8718 (N_8718,N_4908,N_221);
nand U8719 (N_8719,N_4117,N_4249);
nand U8720 (N_8720,N_4354,N_647);
xnor U8721 (N_8721,N_1171,N_4911);
or U8722 (N_8722,N_3148,N_3137);
nand U8723 (N_8723,N_3819,N_213);
nand U8724 (N_8724,N_3136,N_4629);
or U8725 (N_8725,N_12,N_2919);
nand U8726 (N_8726,N_2803,N_3169);
and U8727 (N_8727,N_2125,N_3269);
or U8728 (N_8728,N_926,N_1710);
nor U8729 (N_8729,N_123,N_3165);
and U8730 (N_8730,N_790,N_4265);
or U8731 (N_8731,N_4953,N_876);
nand U8732 (N_8732,N_3427,N_1404);
and U8733 (N_8733,N_2676,N_1339);
nand U8734 (N_8734,N_4494,N_2091);
and U8735 (N_8735,N_2667,N_102);
nand U8736 (N_8736,N_4470,N_4951);
or U8737 (N_8737,N_766,N_1866);
and U8738 (N_8738,N_1159,N_3405);
nor U8739 (N_8739,N_846,N_4999);
and U8740 (N_8740,N_724,N_339);
and U8741 (N_8741,N_3966,N_1413);
or U8742 (N_8742,N_4065,N_4172);
or U8743 (N_8743,N_2674,N_1619);
nor U8744 (N_8744,N_3264,N_4092);
or U8745 (N_8745,N_907,N_150);
or U8746 (N_8746,N_51,N_3413);
and U8747 (N_8747,N_4252,N_2175);
nor U8748 (N_8748,N_1446,N_2763);
and U8749 (N_8749,N_2932,N_2593);
or U8750 (N_8750,N_3762,N_2629);
or U8751 (N_8751,N_3160,N_3749);
and U8752 (N_8752,N_3248,N_3104);
nand U8753 (N_8753,N_2803,N_2162);
or U8754 (N_8754,N_3707,N_2836);
nand U8755 (N_8755,N_3678,N_3927);
nand U8756 (N_8756,N_2354,N_4061);
and U8757 (N_8757,N_2693,N_2282);
and U8758 (N_8758,N_1083,N_4446);
or U8759 (N_8759,N_1569,N_917);
or U8760 (N_8760,N_1536,N_3353);
xor U8761 (N_8761,N_1943,N_375);
nand U8762 (N_8762,N_1542,N_2907);
and U8763 (N_8763,N_3930,N_822);
or U8764 (N_8764,N_73,N_278);
nand U8765 (N_8765,N_2851,N_3498);
and U8766 (N_8766,N_1507,N_69);
nand U8767 (N_8767,N_4082,N_3345);
xnor U8768 (N_8768,N_2316,N_2285);
and U8769 (N_8769,N_2282,N_4699);
nor U8770 (N_8770,N_239,N_3313);
and U8771 (N_8771,N_2513,N_3887);
or U8772 (N_8772,N_2771,N_893);
xnor U8773 (N_8773,N_1809,N_2458);
xnor U8774 (N_8774,N_369,N_2079);
or U8775 (N_8775,N_4123,N_3716);
or U8776 (N_8776,N_2320,N_4277);
or U8777 (N_8777,N_4680,N_1869);
xor U8778 (N_8778,N_28,N_4300);
nor U8779 (N_8779,N_2790,N_2728);
and U8780 (N_8780,N_4230,N_4939);
and U8781 (N_8781,N_3964,N_4032);
xnor U8782 (N_8782,N_4085,N_649);
nor U8783 (N_8783,N_4408,N_2526);
nand U8784 (N_8784,N_4229,N_4399);
xor U8785 (N_8785,N_1051,N_3193);
nor U8786 (N_8786,N_1537,N_3735);
or U8787 (N_8787,N_2930,N_3497);
xor U8788 (N_8788,N_3170,N_689);
or U8789 (N_8789,N_168,N_692);
and U8790 (N_8790,N_1771,N_1414);
nor U8791 (N_8791,N_125,N_980);
and U8792 (N_8792,N_872,N_56);
xor U8793 (N_8793,N_2795,N_486);
and U8794 (N_8794,N_2511,N_4882);
xor U8795 (N_8795,N_821,N_85);
and U8796 (N_8796,N_3882,N_1462);
nand U8797 (N_8797,N_2301,N_5);
xnor U8798 (N_8798,N_2015,N_4156);
nor U8799 (N_8799,N_4874,N_1333);
nor U8800 (N_8800,N_4653,N_4907);
and U8801 (N_8801,N_2630,N_2894);
or U8802 (N_8802,N_217,N_3892);
xor U8803 (N_8803,N_378,N_1608);
nand U8804 (N_8804,N_122,N_1337);
or U8805 (N_8805,N_3248,N_4480);
nor U8806 (N_8806,N_4372,N_581);
nand U8807 (N_8807,N_1291,N_2894);
nor U8808 (N_8808,N_4075,N_4565);
nand U8809 (N_8809,N_2738,N_3186);
nand U8810 (N_8810,N_99,N_2296);
and U8811 (N_8811,N_3595,N_2365);
and U8812 (N_8812,N_2939,N_4916);
nor U8813 (N_8813,N_2840,N_224);
xor U8814 (N_8814,N_254,N_425);
and U8815 (N_8815,N_3090,N_1480);
and U8816 (N_8816,N_3428,N_530);
and U8817 (N_8817,N_4359,N_3612);
xnor U8818 (N_8818,N_1653,N_509);
nor U8819 (N_8819,N_4887,N_3262);
or U8820 (N_8820,N_1303,N_4140);
nor U8821 (N_8821,N_6,N_1919);
or U8822 (N_8822,N_4983,N_3302);
or U8823 (N_8823,N_2231,N_1287);
xnor U8824 (N_8824,N_4996,N_4218);
or U8825 (N_8825,N_3056,N_1513);
nor U8826 (N_8826,N_680,N_3601);
nand U8827 (N_8827,N_889,N_4760);
nand U8828 (N_8828,N_242,N_1256);
xnor U8829 (N_8829,N_4284,N_57);
or U8830 (N_8830,N_1692,N_3933);
nor U8831 (N_8831,N_846,N_3422);
and U8832 (N_8832,N_4241,N_3485);
nand U8833 (N_8833,N_3990,N_2850);
and U8834 (N_8834,N_4451,N_4737);
xnor U8835 (N_8835,N_4145,N_1723);
or U8836 (N_8836,N_3595,N_3918);
nand U8837 (N_8837,N_4106,N_4756);
nand U8838 (N_8838,N_126,N_3452);
and U8839 (N_8839,N_1240,N_989);
nand U8840 (N_8840,N_3902,N_4180);
and U8841 (N_8841,N_827,N_4569);
nand U8842 (N_8842,N_894,N_1401);
nor U8843 (N_8843,N_1523,N_101);
nor U8844 (N_8844,N_554,N_1758);
xor U8845 (N_8845,N_2543,N_680);
or U8846 (N_8846,N_14,N_1117);
nand U8847 (N_8847,N_15,N_3151);
and U8848 (N_8848,N_1571,N_1005);
and U8849 (N_8849,N_483,N_2017);
xnor U8850 (N_8850,N_2662,N_1623);
nand U8851 (N_8851,N_4714,N_4216);
or U8852 (N_8852,N_4455,N_688);
nand U8853 (N_8853,N_294,N_2870);
or U8854 (N_8854,N_2121,N_3665);
nor U8855 (N_8855,N_161,N_4897);
or U8856 (N_8856,N_4767,N_3403);
and U8857 (N_8857,N_1130,N_1285);
and U8858 (N_8858,N_3381,N_1674);
xor U8859 (N_8859,N_424,N_4412);
nor U8860 (N_8860,N_276,N_4068);
or U8861 (N_8861,N_2051,N_3657);
xnor U8862 (N_8862,N_4880,N_1196);
nor U8863 (N_8863,N_23,N_4238);
and U8864 (N_8864,N_2487,N_3342);
and U8865 (N_8865,N_241,N_2201);
and U8866 (N_8866,N_4829,N_4363);
nor U8867 (N_8867,N_4727,N_4110);
nor U8868 (N_8868,N_1980,N_39);
xor U8869 (N_8869,N_4325,N_4079);
xor U8870 (N_8870,N_1963,N_1501);
xnor U8871 (N_8871,N_311,N_4783);
or U8872 (N_8872,N_333,N_1388);
nand U8873 (N_8873,N_710,N_4003);
nand U8874 (N_8874,N_4087,N_825);
xor U8875 (N_8875,N_1433,N_1446);
or U8876 (N_8876,N_1305,N_4353);
nor U8877 (N_8877,N_3931,N_3224);
and U8878 (N_8878,N_3221,N_29);
nor U8879 (N_8879,N_3211,N_4298);
or U8880 (N_8880,N_2876,N_911);
or U8881 (N_8881,N_1992,N_3673);
or U8882 (N_8882,N_2500,N_3828);
and U8883 (N_8883,N_4440,N_273);
xnor U8884 (N_8884,N_3800,N_1877);
nand U8885 (N_8885,N_508,N_4647);
and U8886 (N_8886,N_2924,N_3082);
nor U8887 (N_8887,N_332,N_1445);
and U8888 (N_8888,N_2292,N_2867);
xnor U8889 (N_8889,N_1635,N_3801);
xor U8890 (N_8890,N_756,N_2975);
nor U8891 (N_8891,N_3034,N_3412);
or U8892 (N_8892,N_4630,N_2137);
and U8893 (N_8893,N_152,N_551);
or U8894 (N_8894,N_1771,N_4211);
xnor U8895 (N_8895,N_1741,N_1370);
nand U8896 (N_8896,N_3484,N_4623);
nor U8897 (N_8897,N_95,N_2987);
or U8898 (N_8898,N_70,N_2196);
nand U8899 (N_8899,N_1109,N_3291);
xnor U8900 (N_8900,N_128,N_3278);
xor U8901 (N_8901,N_128,N_659);
xnor U8902 (N_8902,N_1843,N_3760);
nor U8903 (N_8903,N_3388,N_2900);
or U8904 (N_8904,N_2760,N_4305);
or U8905 (N_8905,N_3682,N_4822);
xnor U8906 (N_8906,N_101,N_2461);
nand U8907 (N_8907,N_1006,N_4795);
or U8908 (N_8908,N_2430,N_3957);
or U8909 (N_8909,N_3659,N_1273);
and U8910 (N_8910,N_4139,N_2754);
xor U8911 (N_8911,N_1842,N_2891);
nand U8912 (N_8912,N_2245,N_1686);
nor U8913 (N_8913,N_1393,N_2335);
or U8914 (N_8914,N_1257,N_3382);
xor U8915 (N_8915,N_4070,N_1617);
and U8916 (N_8916,N_239,N_2915);
and U8917 (N_8917,N_2224,N_4365);
nand U8918 (N_8918,N_2413,N_1701);
nor U8919 (N_8919,N_925,N_1888);
or U8920 (N_8920,N_1699,N_2819);
and U8921 (N_8921,N_1912,N_4229);
nand U8922 (N_8922,N_4478,N_4455);
nand U8923 (N_8923,N_1939,N_638);
or U8924 (N_8924,N_1360,N_4647);
nand U8925 (N_8925,N_1146,N_912);
nor U8926 (N_8926,N_4123,N_4778);
nor U8927 (N_8927,N_60,N_1409);
nor U8928 (N_8928,N_2089,N_3399);
nor U8929 (N_8929,N_208,N_4570);
or U8930 (N_8930,N_4405,N_2378);
nand U8931 (N_8931,N_1041,N_2841);
and U8932 (N_8932,N_2860,N_4740);
xnor U8933 (N_8933,N_559,N_1462);
xor U8934 (N_8934,N_3662,N_402);
or U8935 (N_8935,N_4165,N_4515);
xor U8936 (N_8936,N_556,N_413);
nor U8937 (N_8937,N_101,N_3946);
nor U8938 (N_8938,N_4251,N_289);
nand U8939 (N_8939,N_3011,N_460);
xnor U8940 (N_8940,N_3330,N_1108);
or U8941 (N_8941,N_4395,N_3030);
and U8942 (N_8942,N_190,N_3634);
nor U8943 (N_8943,N_116,N_4724);
nand U8944 (N_8944,N_3671,N_1558);
and U8945 (N_8945,N_98,N_915);
xnor U8946 (N_8946,N_2441,N_3481);
xor U8947 (N_8947,N_911,N_3867);
or U8948 (N_8948,N_688,N_4592);
or U8949 (N_8949,N_1381,N_969);
nor U8950 (N_8950,N_3108,N_2236);
nand U8951 (N_8951,N_2051,N_4434);
and U8952 (N_8952,N_4160,N_4895);
nand U8953 (N_8953,N_1247,N_3535);
nor U8954 (N_8954,N_2432,N_2518);
and U8955 (N_8955,N_2321,N_354);
nor U8956 (N_8956,N_1882,N_1141);
or U8957 (N_8957,N_3102,N_529);
xnor U8958 (N_8958,N_90,N_4177);
nand U8959 (N_8959,N_3965,N_4970);
or U8960 (N_8960,N_4579,N_2413);
and U8961 (N_8961,N_4666,N_4380);
nor U8962 (N_8962,N_1495,N_2961);
nand U8963 (N_8963,N_1136,N_1356);
xor U8964 (N_8964,N_2248,N_1165);
and U8965 (N_8965,N_2413,N_181);
or U8966 (N_8966,N_296,N_4050);
and U8967 (N_8967,N_2028,N_4275);
and U8968 (N_8968,N_4180,N_2759);
nor U8969 (N_8969,N_1510,N_3592);
nor U8970 (N_8970,N_587,N_1206);
nand U8971 (N_8971,N_2493,N_3813);
and U8972 (N_8972,N_1062,N_4893);
nor U8973 (N_8973,N_2912,N_1225);
xor U8974 (N_8974,N_1323,N_3270);
nand U8975 (N_8975,N_3544,N_4267);
nor U8976 (N_8976,N_338,N_3813);
or U8977 (N_8977,N_3707,N_3927);
nand U8978 (N_8978,N_2468,N_4964);
or U8979 (N_8979,N_3212,N_2745);
xor U8980 (N_8980,N_3080,N_1887);
nor U8981 (N_8981,N_2182,N_1202);
nor U8982 (N_8982,N_204,N_23);
nor U8983 (N_8983,N_3330,N_4889);
or U8984 (N_8984,N_594,N_3294);
or U8985 (N_8985,N_228,N_3976);
nor U8986 (N_8986,N_4401,N_98);
or U8987 (N_8987,N_3138,N_4215);
or U8988 (N_8988,N_1001,N_2064);
and U8989 (N_8989,N_691,N_3293);
nand U8990 (N_8990,N_3605,N_1222);
nand U8991 (N_8991,N_4778,N_4202);
xor U8992 (N_8992,N_1026,N_2609);
and U8993 (N_8993,N_4915,N_1858);
xor U8994 (N_8994,N_3684,N_2367);
or U8995 (N_8995,N_1591,N_1147);
or U8996 (N_8996,N_2180,N_4465);
xnor U8997 (N_8997,N_4153,N_2930);
or U8998 (N_8998,N_3169,N_3047);
and U8999 (N_8999,N_2859,N_85);
and U9000 (N_9000,N_785,N_4301);
nand U9001 (N_9001,N_1862,N_4650);
xor U9002 (N_9002,N_43,N_4824);
nand U9003 (N_9003,N_1293,N_3354);
nand U9004 (N_9004,N_169,N_4842);
and U9005 (N_9005,N_2700,N_4481);
or U9006 (N_9006,N_3362,N_4185);
nand U9007 (N_9007,N_185,N_1359);
nand U9008 (N_9008,N_2570,N_2319);
nand U9009 (N_9009,N_3419,N_585);
xnor U9010 (N_9010,N_3719,N_3469);
nor U9011 (N_9011,N_2613,N_4575);
nand U9012 (N_9012,N_2284,N_3087);
nor U9013 (N_9013,N_1142,N_1538);
or U9014 (N_9014,N_1008,N_824);
or U9015 (N_9015,N_577,N_2009);
or U9016 (N_9016,N_2881,N_3994);
nor U9017 (N_9017,N_3767,N_4571);
nor U9018 (N_9018,N_2357,N_1944);
nor U9019 (N_9019,N_403,N_3642);
and U9020 (N_9020,N_3280,N_2277);
and U9021 (N_9021,N_4824,N_86);
or U9022 (N_9022,N_777,N_869);
and U9023 (N_9023,N_200,N_4084);
nand U9024 (N_9024,N_1545,N_647);
xor U9025 (N_9025,N_1208,N_935);
xnor U9026 (N_9026,N_4034,N_4841);
or U9027 (N_9027,N_4082,N_2284);
nand U9028 (N_9028,N_3699,N_926);
nor U9029 (N_9029,N_3205,N_3647);
nor U9030 (N_9030,N_802,N_4462);
or U9031 (N_9031,N_2038,N_2794);
xnor U9032 (N_9032,N_1961,N_2143);
and U9033 (N_9033,N_4088,N_530);
nor U9034 (N_9034,N_20,N_2581);
nand U9035 (N_9035,N_2645,N_3865);
nor U9036 (N_9036,N_273,N_2191);
nor U9037 (N_9037,N_2071,N_3117);
nand U9038 (N_9038,N_409,N_1886);
and U9039 (N_9039,N_4620,N_59);
xnor U9040 (N_9040,N_1251,N_3495);
or U9041 (N_9041,N_839,N_1529);
nand U9042 (N_9042,N_932,N_2702);
or U9043 (N_9043,N_4040,N_2154);
xor U9044 (N_9044,N_2801,N_4735);
or U9045 (N_9045,N_1000,N_4323);
nand U9046 (N_9046,N_4187,N_1712);
xor U9047 (N_9047,N_735,N_1973);
nand U9048 (N_9048,N_1477,N_392);
nor U9049 (N_9049,N_1054,N_4808);
nor U9050 (N_9050,N_4364,N_2647);
nor U9051 (N_9051,N_4642,N_804);
and U9052 (N_9052,N_3732,N_3547);
nor U9053 (N_9053,N_4937,N_918);
or U9054 (N_9054,N_1106,N_4285);
or U9055 (N_9055,N_3054,N_1363);
and U9056 (N_9056,N_4296,N_1318);
nand U9057 (N_9057,N_4313,N_2060);
nand U9058 (N_9058,N_164,N_4399);
and U9059 (N_9059,N_518,N_1927);
or U9060 (N_9060,N_4793,N_844);
xnor U9061 (N_9061,N_1750,N_2119);
nand U9062 (N_9062,N_2885,N_2069);
or U9063 (N_9063,N_4984,N_3562);
and U9064 (N_9064,N_1408,N_1438);
or U9065 (N_9065,N_178,N_4551);
and U9066 (N_9066,N_465,N_3578);
or U9067 (N_9067,N_1575,N_3034);
and U9068 (N_9068,N_2857,N_2322);
nand U9069 (N_9069,N_3737,N_4422);
nor U9070 (N_9070,N_33,N_3334);
nand U9071 (N_9071,N_1794,N_3655);
nand U9072 (N_9072,N_1811,N_701);
or U9073 (N_9073,N_1675,N_1038);
or U9074 (N_9074,N_4713,N_2758);
and U9075 (N_9075,N_77,N_2620);
xnor U9076 (N_9076,N_3235,N_2454);
xor U9077 (N_9077,N_3816,N_4623);
and U9078 (N_9078,N_281,N_3570);
or U9079 (N_9079,N_2634,N_4212);
and U9080 (N_9080,N_4829,N_2040);
nor U9081 (N_9081,N_1355,N_1436);
or U9082 (N_9082,N_3619,N_2593);
xor U9083 (N_9083,N_1475,N_2962);
or U9084 (N_9084,N_3174,N_1569);
or U9085 (N_9085,N_1969,N_3437);
nor U9086 (N_9086,N_2549,N_2277);
or U9087 (N_9087,N_813,N_2059);
or U9088 (N_9088,N_4367,N_964);
xnor U9089 (N_9089,N_1804,N_2012);
xnor U9090 (N_9090,N_3208,N_320);
xor U9091 (N_9091,N_1500,N_1452);
nor U9092 (N_9092,N_4306,N_3035);
and U9093 (N_9093,N_452,N_1072);
or U9094 (N_9094,N_3403,N_2156);
nand U9095 (N_9095,N_1441,N_4690);
nor U9096 (N_9096,N_12,N_4394);
nor U9097 (N_9097,N_95,N_2025);
and U9098 (N_9098,N_2243,N_1690);
nor U9099 (N_9099,N_2941,N_4728);
and U9100 (N_9100,N_1787,N_298);
nor U9101 (N_9101,N_3029,N_3459);
nand U9102 (N_9102,N_3361,N_1087);
nor U9103 (N_9103,N_516,N_4483);
and U9104 (N_9104,N_1725,N_1822);
xor U9105 (N_9105,N_4623,N_1651);
xnor U9106 (N_9106,N_441,N_528);
nand U9107 (N_9107,N_2285,N_2158);
nand U9108 (N_9108,N_1378,N_3511);
nand U9109 (N_9109,N_3231,N_834);
nand U9110 (N_9110,N_2471,N_861);
and U9111 (N_9111,N_342,N_4612);
nand U9112 (N_9112,N_998,N_2241);
nor U9113 (N_9113,N_958,N_3356);
nor U9114 (N_9114,N_170,N_2342);
and U9115 (N_9115,N_2757,N_2383);
and U9116 (N_9116,N_2762,N_934);
nor U9117 (N_9117,N_4411,N_4696);
nor U9118 (N_9118,N_4695,N_1828);
xor U9119 (N_9119,N_1051,N_1189);
and U9120 (N_9120,N_345,N_3462);
or U9121 (N_9121,N_4360,N_3396);
or U9122 (N_9122,N_4304,N_793);
and U9123 (N_9123,N_496,N_3658);
xnor U9124 (N_9124,N_4892,N_3671);
and U9125 (N_9125,N_4296,N_212);
nand U9126 (N_9126,N_4189,N_4172);
nor U9127 (N_9127,N_4035,N_538);
xor U9128 (N_9128,N_1336,N_4267);
nor U9129 (N_9129,N_1551,N_4623);
nand U9130 (N_9130,N_4197,N_3637);
xnor U9131 (N_9131,N_1333,N_1712);
nand U9132 (N_9132,N_2874,N_2851);
and U9133 (N_9133,N_4297,N_3132);
xnor U9134 (N_9134,N_1791,N_2151);
xnor U9135 (N_9135,N_1974,N_1443);
xor U9136 (N_9136,N_3204,N_2053);
and U9137 (N_9137,N_682,N_1820);
nand U9138 (N_9138,N_778,N_2671);
and U9139 (N_9139,N_1328,N_1251);
or U9140 (N_9140,N_2352,N_4051);
nor U9141 (N_9141,N_166,N_2127);
xnor U9142 (N_9142,N_3213,N_728);
and U9143 (N_9143,N_3277,N_1608);
nand U9144 (N_9144,N_575,N_3908);
nor U9145 (N_9145,N_1348,N_4376);
xnor U9146 (N_9146,N_3016,N_714);
and U9147 (N_9147,N_1791,N_949);
nand U9148 (N_9148,N_3902,N_1606);
nor U9149 (N_9149,N_1703,N_3696);
or U9150 (N_9150,N_2145,N_2324);
nand U9151 (N_9151,N_533,N_1708);
or U9152 (N_9152,N_440,N_2651);
xor U9153 (N_9153,N_4976,N_1485);
and U9154 (N_9154,N_941,N_619);
nand U9155 (N_9155,N_1317,N_4122);
nor U9156 (N_9156,N_4804,N_1865);
xor U9157 (N_9157,N_4,N_3342);
nand U9158 (N_9158,N_4803,N_3527);
nand U9159 (N_9159,N_636,N_3410);
or U9160 (N_9160,N_4412,N_1091);
and U9161 (N_9161,N_2848,N_746);
or U9162 (N_9162,N_2281,N_439);
and U9163 (N_9163,N_2472,N_2819);
nor U9164 (N_9164,N_3072,N_2106);
nand U9165 (N_9165,N_3828,N_2048);
or U9166 (N_9166,N_1181,N_4168);
nand U9167 (N_9167,N_438,N_2143);
and U9168 (N_9168,N_696,N_1157);
nand U9169 (N_9169,N_4545,N_1644);
nor U9170 (N_9170,N_4639,N_4564);
nand U9171 (N_9171,N_3640,N_4112);
xor U9172 (N_9172,N_2395,N_4155);
and U9173 (N_9173,N_2697,N_2915);
nand U9174 (N_9174,N_1496,N_4395);
xor U9175 (N_9175,N_2836,N_4681);
xor U9176 (N_9176,N_2771,N_337);
nor U9177 (N_9177,N_1113,N_945);
nand U9178 (N_9178,N_3408,N_2782);
nor U9179 (N_9179,N_4410,N_790);
nand U9180 (N_9180,N_3122,N_4466);
xnor U9181 (N_9181,N_3932,N_2631);
xnor U9182 (N_9182,N_1248,N_599);
nor U9183 (N_9183,N_1977,N_2129);
nand U9184 (N_9184,N_3279,N_376);
and U9185 (N_9185,N_3645,N_3520);
nand U9186 (N_9186,N_2436,N_4177);
or U9187 (N_9187,N_2799,N_926);
nand U9188 (N_9188,N_3506,N_408);
xor U9189 (N_9189,N_360,N_1281);
nor U9190 (N_9190,N_3996,N_4718);
nand U9191 (N_9191,N_425,N_4024);
and U9192 (N_9192,N_128,N_4336);
nor U9193 (N_9193,N_4473,N_1294);
xor U9194 (N_9194,N_4486,N_4693);
or U9195 (N_9195,N_2612,N_1658);
nor U9196 (N_9196,N_822,N_3374);
or U9197 (N_9197,N_3945,N_1476);
nand U9198 (N_9198,N_1253,N_4439);
or U9199 (N_9199,N_251,N_3359);
xor U9200 (N_9200,N_131,N_3566);
xnor U9201 (N_9201,N_1763,N_2383);
nand U9202 (N_9202,N_1450,N_4147);
xnor U9203 (N_9203,N_2665,N_4658);
and U9204 (N_9204,N_3214,N_3597);
or U9205 (N_9205,N_4331,N_1639);
nor U9206 (N_9206,N_4151,N_154);
xor U9207 (N_9207,N_2735,N_1299);
xor U9208 (N_9208,N_352,N_4137);
xor U9209 (N_9209,N_3000,N_2549);
xnor U9210 (N_9210,N_3294,N_926);
or U9211 (N_9211,N_327,N_1369);
nand U9212 (N_9212,N_2855,N_1058);
nor U9213 (N_9213,N_640,N_4379);
nand U9214 (N_9214,N_2034,N_2243);
nand U9215 (N_9215,N_3336,N_3737);
nand U9216 (N_9216,N_3159,N_3318);
xor U9217 (N_9217,N_3968,N_785);
and U9218 (N_9218,N_4438,N_3791);
or U9219 (N_9219,N_3837,N_1329);
nor U9220 (N_9220,N_119,N_3869);
nand U9221 (N_9221,N_2979,N_3484);
nand U9222 (N_9222,N_4249,N_1308);
or U9223 (N_9223,N_3265,N_740);
or U9224 (N_9224,N_436,N_2757);
and U9225 (N_9225,N_1268,N_4470);
or U9226 (N_9226,N_751,N_782);
and U9227 (N_9227,N_4372,N_1677);
or U9228 (N_9228,N_4220,N_4491);
and U9229 (N_9229,N_2143,N_2839);
and U9230 (N_9230,N_4279,N_2676);
nor U9231 (N_9231,N_1217,N_2016);
nand U9232 (N_9232,N_3859,N_2868);
nand U9233 (N_9233,N_4713,N_3324);
and U9234 (N_9234,N_1539,N_840);
nor U9235 (N_9235,N_3570,N_314);
xnor U9236 (N_9236,N_4399,N_1823);
xor U9237 (N_9237,N_588,N_4539);
xnor U9238 (N_9238,N_4490,N_3400);
and U9239 (N_9239,N_1879,N_4685);
or U9240 (N_9240,N_4632,N_560);
xnor U9241 (N_9241,N_2784,N_1263);
nand U9242 (N_9242,N_4417,N_2464);
and U9243 (N_9243,N_3890,N_1452);
xor U9244 (N_9244,N_4144,N_3565);
nor U9245 (N_9245,N_1668,N_4670);
nand U9246 (N_9246,N_2084,N_3714);
xor U9247 (N_9247,N_1474,N_12);
xor U9248 (N_9248,N_1610,N_2528);
or U9249 (N_9249,N_113,N_2047);
and U9250 (N_9250,N_3079,N_4228);
or U9251 (N_9251,N_4453,N_2841);
nand U9252 (N_9252,N_3183,N_3206);
and U9253 (N_9253,N_23,N_59);
nand U9254 (N_9254,N_503,N_2083);
nand U9255 (N_9255,N_1565,N_1693);
or U9256 (N_9256,N_1911,N_3510);
and U9257 (N_9257,N_491,N_1305);
and U9258 (N_9258,N_4629,N_2155);
xnor U9259 (N_9259,N_1699,N_2443);
and U9260 (N_9260,N_668,N_289);
nand U9261 (N_9261,N_2895,N_614);
or U9262 (N_9262,N_4606,N_3579);
and U9263 (N_9263,N_165,N_827);
xor U9264 (N_9264,N_83,N_2528);
nand U9265 (N_9265,N_2167,N_4729);
or U9266 (N_9266,N_4579,N_849);
and U9267 (N_9267,N_3360,N_1205);
nor U9268 (N_9268,N_978,N_3497);
nand U9269 (N_9269,N_3433,N_1157);
or U9270 (N_9270,N_1286,N_1945);
nand U9271 (N_9271,N_1512,N_3158);
and U9272 (N_9272,N_1653,N_1452);
and U9273 (N_9273,N_671,N_2081);
xor U9274 (N_9274,N_3499,N_182);
or U9275 (N_9275,N_1443,N_3543);
or U9276 (N_9276,N_2982,N_1518);
and U9277 (N_9277,N_3692,N_4788);
nand U9278 (N_9278,N_2475,N_2139);
or U9279 (N_9279,N_2287,N_1224);
nand U9280 (N_9280,N_4149,N_2057);
nand U9281 (N_9281,N_1416,N_656);
nor U9282 (N_9282,N_1223,N_576);
nor U9283 (N_9283,N_3032,N_655);
or U9284 (N_9284,N_4585,N_204);
and U9285 (N_9285,N_242,N_665);
or U9286 (N_9286,N_3100,N_652);
xnor U9287 (N_9287,N_263,N_139);
xnor U9288 (N_9288,N_1757,N_2930);
and U9289 (N_9289,N_4723,N_1350);
xnor U9290 (N_9290,N_1055,N_3203);
nand U9291 (N_9291,N_4502,N_4058);
nor U9292 (N_9292,N_1524,N_3821);
xor U9293 (N_9293,N_574,N_396);
nand U9294 (N_9294,N_2839,N_2023);
nor U9295 (N_9295,N_3397,N_1274);
or U9296 (N_9296,N_1916,N_3073);
nand U9297 (N_9297,N_948,N_911);
nor U9298 (N_9298,N_2775,N_4005);
nor U9299 (N_9299,N_1189,N_1485);
and U9300 (N_9300,N_2808,N_3418);
nor U9301 (N_9301,N_2959,N_264);
xnor U9302 (N_9302,N_3014,N_2554);
nor U9303 (N_9303,N_744,N_3337);
xor U9304 (N_9304,N_2449,N_4510);
or U9305 (N_9305,N_4288,N_1884);
nor U9306 (N_9306,N_376,N_3);
nor U9307 (N_9307,N_1630,N_474);
and U9308 (N_9308,N_2032,N_1946);
nor U9309 (N_9309,N_2296,N_1847);
nor U9310 (N_9310,N_1199,N_1263);
xnor U9311 (N_9311,N_4096,N_3029);
xnor U9312 (N_9312,N_2315,N_79);
and U9313 (N_9313,N_1905,N_3690);
nor U9314 (N_9314,N_282,N_1800);
xor U9315 (N_9315,N_2431,N_1063);
nand U9316 (N_9316,N_4535,N_105);
nand U9317 (N_9317,N_3189,N_1866);
nand U9318 (N_9318,N_1556,N_4612);
nand U9319 (N_9319,N_3838,N_2628);
and U9320 (N_9320,N_1292,N_596);
and U9321 (N_9321,N_666,N_651);
or U9322 (N_9322,N_410,N_695);
nor U9323 (N_9323,N_1068,N_2680);
xor U9324 (N_9324,N_3745,N_1548);
and U9325 (N_9325,N_1720,N_917);
xnor U9326 (N_9326,N_2217,N_2632);
and U9327 (N_9327,N_3554,N_1044);
nand U9328 (N_9328,N_3083,N_2772);
xor U9329 (N_9329,N_1927,N_1809);
nor U9330 (N_9330,N_1077,N_4431);
or U9331 (N_9331,N_3948,N_4247);
nor U9332 (N_9332,N_4332,N_1127);
or U9333 (N_9333,N_66,N_1883);
or U9334 (N_9334,N_303,N_3704);
nor U9335 (N_9335,N_3038,N_2576);
and U9336 (N_9336,N_2380,N_2958);
nand U9337 (N_9337,N_4229,N_954);
or U9338 (N_9338,N_854,N_4207);
xnor U9339 (N_9339,N_4333,N_1689);
nand U9340 (N_9340,N_4017,N_3027);
nand U9341 (N_9341,N_4382,N_1591);
or U9342 (N_9342,N_3380,N_3434);
xnor U9343 (N_9343,N_2944,N_2502);
nor U9344 (N_9344,N_4185,N_2309);
xor U9345 (N_9345,N_1161,N_1868);
xnor U9346 (N_9346,N_2182,N_1094);
xor U9347 (N_9347,N_1786,N_1494);
or U9348 (N_9348,N_802,N_4439);
xnor U9349 (N_9349,N_174,N_132);
and U9350 (N_9350,N_3594,N_2266);
or U9351 (N_9351,N_3177,N_3777);
nand U9352 (N_9352,N_4501,N_606);
or U9353 (N_9353,N_426,N_3984);
nor U9354 (N_9354,N_1414,N_2058);
or U9355 (N_9355,N_2880,N_4900);
nand U9356 (N_9356,N_3744,N_3687);
xnor U9357 (N_9357,N_1512,N_1714);
or U9358 (N_9358,N_4906,N_1381);
nand U9359 (N_9359,N_821,N_2271);
nand U9360 (N_9360,N_1967,N_3858);
nor U9361 (N_9361,N_641,N_3533);
nand U9362 (N_9362,N_1097,N_2706);
and U9363 (N_9363,N_1407,N_4426);
xnor U9364 (N_9364,N_564,N_813);
and U9365 (N_9365,N_911,N_4110);
and U9366 (N_9366,N_1332,N_599);
nor U9367 (N_9367,N_3963,N_2185);
xor U9368 (N_9368,N_2034,N_2873);
and U9369 (N_9369,N_3346,N_3267);
or U9370 (N_9370,N_2283,N_1833);
xnor U9371 (N_9371,N_3004,N_1054);
nor U9372 (N_9372,N_280,N_2007);
xor U9373 (N_9373,N_2971,N_303);
or U9374 (N_9374,N_4150,N_1991);
and U9375 (N_9375,N_4183,N_3549);
and U9376 (N_9376,N_1950,N_4262);
nor U9377 (N_9377,N_2068,N_4141);
and U9378 (N_9378,N_734,N_127);
xor U9379 (N_9379,N_83,N_2022);
or U9380 (N_9380,N_3387,N_4702);
nor U9381 (N_9381,N_1954,N_3291);
xnor U9382 (N_9382,N_1815,N_3178);
nor U9383 (N_9383,N_36,N_1561);
or U9384 (N_9384,N_3218,N_2300);
or U9385 (N_9385,N_4529,N_3143);
nand U9386 (N_9386,N_2424,N_1909);
xnor U9387 (N_9387,N_1031,N_3024);
xor U9388 (N_9388,N_4038,N_1293);
and U9389 (N_9389,N_1591,N_2394);
nor U9390 (N_9390,N_1065,N_2089);
nand U9391 (N_9391,N_4809,N_3526);
xor U9392 (N_9392,N_477,N_1169);
or U9393 (N_9393,N_3929,N_4310);
nor U9394 (N_9394,N_3164,N_1150);
xor U9395 (N_9395,N_2578,N_3789);
or U9396 (N_9396,N_1226,N_3341);
or U9397 (N_9397,N_4681,N_4752);
or U9398 (N_9398,N_2984,N_3678);
xnor U9399 (N_9399,N_3565,N_3776);
and U9400 (N_9400,N_2252,N_1519);
nand U9401 (N_9401,N_2619,N_4571);
nand U9402 (N_9402,N_1948,N_2021);
or U9403 (N_9403,N_2345,N_3138);
nor U9404 (N_9404,N_4609,N_151);
or U9405 (N_9405,N_4131,N_2605);
or U9406 (N_9406,N_1940,N_3013);
and U9407 (N_9407,N_396,N_3826);
xnor U9408 (N_9408,N_4458,N_4903);
xor U9409 (N_9409,N_1964,N_1922);
nand U9410 (N_9410,N_2770,N_1093);
and U9411 (N_9411,N_3802,N_3631);
or U9412 (N_9412,N_2574,N_1760);
or U9413 (N_9413,N_3358,N_1395);
nor U9414 (N_9414,N_2224,N_2474);
and U9415 (N_9415,N_2576,N_544);
nand U9416 (N_9416,N_3181,N_2704);
and U9417 (N_9417,N_4791,N_481);
nor U9418 (N_9418,N_2601,N_473);
or U9419 (N_9419,N_3546,N_270);
nor U9420 (N_9420,N_239,N_2600);
nand U9421 (N_9421,N_3630,N_2380);
and U9422 (N_9422,N_3706,N_1840);
nor U9423 (N_9423,N_4185,N_4776);
or U9424 (N_9424,N_4702,N_3887);
nor U9425 (N_9425,N_2171,N_694);
and U9426 (N_9426,N_2609,N_1707);
xnor U9427 (N_9427,N_3669,N_3703);
xnor U9428 (N_9428,N_3155,N_2863);
nand U9429 (N_9429,N_2655,N_4917);
xnor U9430 (N_9430,N_640,N_247);
nor U9431 (N_9431,N_1172,N_3460);
nand U9432 (N_9432,N_3816,N_1868);
or U9433 (N_9433,N_2401,N_3507);
nor U9434 (N_9434,N_1435,N_3503);
or U9435 (N_9435,N_3619,N_2695);
or U9436 (N_9436,N_326,N_3476);
or U9437 (N_9437,N_1287,N_2052);
or U9438 (N_9438,N_2923,N_4756);
or U9439 (N_9439,N_1508,N_4100);
nand U9440 (N_9440,N_4968,N_241);
xnor U9441 (N_9441,N_4637,N_2968);
nor U9442 (N_9442,N_387,N_101);
and U9443 (N_9443,N_163,N_374);
nand U9444 (N_9444,N_2954,N_261);
or U9445 (N_9445,N_3411,N_4407);
or U9446 (N_9446,N_3037,N_2176);
or U9447 (N_9447,N_1748,N_595);
nor U9448 (N_9448,N_267,N_3699);
nor U9449 (N_9449,N_878,N_1733);
and U9450 (N_9450,N_3999,N_4619);
nand U9451 (N_9451,N_1431,N_3033);
nand U9452 (N_9452,N_2775,N_4356);
and U9453 (N_9453,N_1608,N_2231);
or U9454 (N_9454,N_4822,N_3065);
and U9455 (N_9455,N_1639,N_1154);
xnor U9456 (N_9456,N_1213,N_493);
nand U9457 (N_9457,N_3923,N_3452);
nand U9458 (N_9458,N_2783,N_3732);
xnor U9459 (N_9459,N_2701,N_2663);
and U9460 (N_9460,N_4277,N_4841);
nand U9461 (N_9461,N_2329,N_2587);
or U9462 (N_9462,N_3070,N_2752);
nor U9463 (N_9463,N_1084,N_3180);
nor U9464 (N_9464,N_3103,N_4836);
nor U9465 (N_9465,N_2342,N_1910);
nor U9466 (N_9466,N_2601,N_106);
nor U9467 (N_9467,N_3716,N_4721);
and U9468 (N_9468,N_4078,N_4448);
or U9469 (N_9469,N_775,N_1560);
and U9470 (N_9470,N_4576,N_3831);
nor U9471 (N_9471,N_4466,N_2965);
or U9472 (N_9472,N_2649,N_4837);
nor U9473 (N_9473,N_1746,N_3954);
xnor U9474 (N_9474,N_2861,N_3452);
and U9475 (N_9475,N_1912,N_1843);
nor U9476 (N_9476,N_4973,N_2705);
and U9477 (N_9477,N_2674,N_4485);
nand U9478 (N_9478,N_1145,N_3224);
and U9479 (N_9479,N_3865,N_807);
and U9480 (N_9480,N_2192,N_2435);
xnor U9481 (N_9481,N_4314,N_4252);
xnor U9482 (N_9482,N_1684,N_4213);
nor U9483 (N_9483,N_3666,N_1348);
xor U9484 (N_9484,N_2934,N_4603);
nand U9485 (N_9485,N_3363,N_238);
or U9486 (N_9486,N_168,N_3689);
xnor U9487 (N_9487,N_4950,N_2807);
or U9488 (N_9488,N_1610,N_118);
and U9489 (N_9489,N_914,N_493);
and U9490 (N_9490,N_3896,N_3393);
and U9491 (N_9491,N_4002,N_116);
or U9492 (N_9492,N_4241,N_332);
xnor U9493 (N_9493,N_2706,N_858);
nand U9494 (N_9494,N_3722,N_4906);
or U9495 (N_9495,N_3464,N_714);
xor U9496 (N_9496,N_3175,N_65);
or U9497 (N_9497,N_2504,N_456);
or U9498 (N_9498,N_487,N_1815);
nand U9499 (N_9499,N_776,N_2100);
nor U9500 (N_9500,N_3408,N_4500);
nand U9501 (N_9501,N_559,N_4069);
and U9502 (N_9502,N_3216,N_3281);
or U9503 (N_9503,N_117,N_3498);
xnor U9504 (N_9504,N_4079,N_216);
nor U9505 (N_9505,N_1167,N_4103);
nand U9506 (N_9506,N_4421,N_2634);
nand U9507 (N_9507,N_1364,N_2368);
and U9508 (N_9508,N_2714,N_2332);
nor U9509 (N_9509,N_4100,N_163);
nor U9510 (N_9510,N_3746,N_4075);
or U9511 (N_9511,N_3860,N_4806);
and U9512 (N_9512,N_542,N_3690);
or U9513 (N_9513,N_1326,N_2153);
xnor U9514 (N_9514,N_2876,N_4777);
nand U9515 (N_9515,N_4584,N_2926);
and U9516 (N_9516,N_1965,N_4190);
xnor U9517 (N_9517,N_4551,N_1838);
nand U9518 (N_9518,N_3681,N_3215);
xnor U9519 (N_9519,N_452,N_319);
nor U9520 (N_9520,N_4709,N_3189);
and U9521 (N_9521,N_4692,N_3126);
or U9522 (N_9522,N_4592,N_1799);
nor U9523 (N_9523,N_3064,N_2827);
nand U9524 (N_9524,N_3520,N_104);
or U9525 (N_9525,N_4523,N_3035);
xnor U9526 (N_9526,N_3448,N_1203);
and U9527 (N_9527,N_4866,N_2338);
or U9528 (N_9528,N_1512,N_3208);
or U9529 (N_9529,N_2921,N_2818);
nor U9530 (N_9530,N_2755,N_582);
xor U9531 (N_9531,N_2780,N_1694);
xor U9532 (N_9532,N_592,N_4915);
nor U9533 (N_9533,N_3898,N_3515);
nor U9534 (N_9534,N_2135,N_4425);
or U9535 (N_9535,N_2687,N_952);
nand U9536 (N_9536,N_3306,N_316);
and U9537 (N_9537,N_1942,N_1002);
xnor U9538 (N_9538,N_345,N_1121);
nand U9539 (N_9539,N_4282,N_4742);
nor U9540 (N_9540,N_4106,N_4372);
or U9541 (N_9541,N_2937,N_2869);
xnor U9542 (N_9542,N_2936,N_893);
nor U9543 (N_9543,N_673,N_1850);
or U9544 (N_9544,N_3287,N_3858);
xor U9545 (N_9545,N_3188,N_3125);
or U9546 (N_9546,N_91,N_2429);
or U9547 (N_9547,N_3608,N_4525);
and U9548 (N_9548,N_1153,N_839);
and U9549 (N_9549,N_3889,N_3627);
xor U9550 (N_9550,N_1345,N_1110);
nor U9551 (N_9551,N_658,N_1434);
and U9552 (N_9552,N_1394,N_4831);
nor U9553 (N_9553,N_2160,N_4551);
nand U9554 (N_9554,N_2727,N_2920);
or U9555 (N_9555,N_2810,N_516);
nor U9556 (N_9556,N_4637,N_893);
or U9557 (N_9557,N_637,N_2626);
and U9558 (N_9558,N_371,N_3879);
xor U9559 (N_9559,N_740,N_2607);
nor U9560 (N_9560,N_1124,N_2638);
and U9561 (N_9561,N_1202,N_1825);
or U9562 (N_9562,N_2078,N_3834);
and U9563 (N_9563,N_1095,N_3747);
nand U9564 (N_9564,N_357,N_4914);
or U9565 (N_9565,N_694,N_2928);
nor U9566 (N_9566,N_4907,N_343);
and U9567 (N_9567,N_4372,N_1420);
nor U9568 (N_9568,N_2163,N_1526);
xor U9569 (N_9569,N_3793,N_645);
nand U9570 (N_9570,N_2606,N_3259);
nor U9571 (N_9571,N_4210,N_3004);
or U9572 (N_9572,N_3586,N_1943);
nand U9573 (N_9573,N_4802,N_3504);
xor U9574 (N_9574,N_2133,N_1449);
and U9575 (N_9575,N_299,N_2522);
nor U9576 (N_9576,N_3084,N_4904);
nand U9577 (N_9577,N_1781,N_3686);
and U9578 (N_9578,N_348,N_247);
nor U9579 (N_9579,N_92,N_4188);
nand U9580 (N_9580,N_1188,N_4255);
xor U9581 (N_9581,N_3771,N_2338);
nor U9582 (N_9582,N_38,N_519);
and U9583 (N_9583,N_1544,N_462);
nand U9584 (N_9584,N_4823,N_2202);
or U9585 (N_9585,N_425,N_551);
or U9586 (N_9586,N_730,N_1457);
nor U9587 (N_9587,N_1621,N_4860);
and U9588 (N_9588,N_4898,N_2717);
xor U9589 (N_9589,N_969,N_4548);
nor U9590 (N_9590,N_1695,N_904);
or U9591 (N_9591,N_1438,N_1418);
nor U9592 (N_9592,N_1550,N_1342);
nor U9593 (N_9593,N_4413,N_97);
and U9594 (N_9594,N_1372,N_4456);
and U9595 (N_9595,N_2936,N_324);
and U9596 (N_9596,N_1021,N_1019);
nand U9597 (N_9597,N_4207,N_3573);
and U9598 (N_9598,N_150,N_3358);
xor U9599 (N_9599,N_3349,N_3277);
or U9600 (N_9600,N_2661,N_773);
nor U9601 (N_9601,N_4692,N_2682);
xnor U9602 (N_9602,N_4166,N_4870);
xor U9603 (N_9603,N_107,N_3085);
nand U9604 (N_9604,N_2374,N_2089);
nor U9605 (N_9605,N_3980,N_1646);
or U9606 (N_9606,N_4273,N_4171);
nand U9607 (N_9607,N_3674,N_4013);
nand U9608 (N_9608,N_1382,N_3810);
xor U9609 (N_9609,N_3373,N_166);
and U9610 (N_9610,N_3396,N_2246);
and U9611 (N_9611,N_380,N_4847);
and U9612 (N_9612,N_4496,N_2941);
nand U9613 (N_9613,N_247,N_938);
xor U9614 (N_9614,N_437,N_4369);
nor U9615 (N_9615,N_3434,N_1538);
nand U9616 (N_9616,N_2933,N_3998);
or U9617 (N_9617,N_768,N_2073);
nor U9618 (N_9618,N_2482,N_803);
or U9619 (N_9619,N_4310,N_2565);
or U9620 (N_9620,N_2536,N_4435);
nand U9621 (N_9621,N_540,N_3553);
nand U9622 (N_9622,N_4222,N_834);
nor U9623 (N_9623,N_1310,N_3748);
and U9624 (N_9624,N_2192,N_3111);
nand U9625 (N_9625,N_4867,N_4580);
and U9626 (N_9626,N_497,N_3069);
or U9627 (N_9627,N_1408,N_3716);
and U9628 (N_9628,N_2396,N_3733);
nand U9629 (N_9629,N_2969,N_3865);
and U9630 (N_9630,N_4533,N_3512);
xor U9631 (N_9631,N_2133,N_430);
and U9632 (N_9632,N_408,N_3962);
nor U9633 (N_9633,N_1549,N_1047);
nor U9634 (N_9634,N_4964,N_1235);
and U9635 (N_9635,N_1093,N_1840);
or U9636 (N_9636,N_4230,N_2860);
xor U9637 (N_9637,N_4240,N_1174);
and U9638 (N_9638,N_2487,N_1816);
nor U9639 (N_9639,N_189,N_4388);
xor U9640 (N_9640,N_4904,N_3161);
nor U9641 (N_9641,N_3986,N_2903);
nor U9642 (N_9642,N_2625,N_1838);
xor U9643 (N_9643,N_1138,N_3361);
nor U9644 (N_9644,N_2419,N_4718);
and U9645 (N_9645,N_795,N_662);
and U9646 (N_9646,N_1815,N_455);
or U9647 (N_9647,N_2508,N_2967);
or U9648 (N_9648,N_1850,N_4451);
or U9649 (N_9649,N_2770,N_2087);
xnor U9650 (N_9650,N_4351,N_471);
or U9651 (N_9651,N_2151,N_4677);
nor U9652 (N_9652,N_2870,N_2457);
and U9653 (N_9653,N_2315,N_4296);
nand U9654 (N_9654,N_1929,N_3732);
or U9655 (N_9655,N_3116,N_2107);
and U9656 (N_9656,N_303,N_830);
or U9657 (N_9657,N_2109,N_4070);
nor U9658 (N_9658,N_3499,N_3601);
or U9659 (N_9659,N_2414,N_3816);
xor U9660 (N_9660,N_1563,N_1443);
and U9661 (N_9661,N_4146,N_3783);
nor U9662 (N_9662,N_3850,N_4668);
nand U9663 (N_9663,N_4274,N_1731);
and U9664 (N_9664,N_2633,N_2373);
or U9665 (N_9665,N_1951,N_3860);
and U9666 (N_9666,N_4501,N_3157);
nand U9667 (N_9667,N_1711,N_3106);
nor U9668 (N_9668,N_2751,N_4078);
nor U9669 (N_9669,N_889,N_4181);
nor U9670 (N_9670,N_166,N_4825);
nand U9671 (N_9671,N_2563,N_3146);
nand U9672 (N_9672,N_1199,N_2279);
or U9673 (N_9673,N_1170,N_1869);
and U9674 (N_9674,N_3033,N_1642);
and U9675 (N_9675,N_65,N_4541);
nand U9676 (N_9676,N_20,N_656);
and U9677 (N_9677,N_909,N_2911);
nor U9678 (N_9678,N_476,N_2653);
nand U9679 (N_9679,N_195,N_1371);
nand U9680 (N_9680,N_3271,N_4894);
xnor U9681 (N_9681,N_4499,N_447);
nand U9682 (N_9682,N_4116,N_3491);
nor U9683 (N_9683,N_2713,N_1703);
nor U9684 (N_9684,N_3601,N_212);
and U9685 (N_9685,N_2438,N_2702);
or U9686 (N_9686,N_3435,N_676);
nor U9687 (N_9687,N_2579,N_534);
nor U9688 (N_9688,N_657,N_4207);
nand U9689 (N_9689,N_4557,N_3465);
nor U9690 (N_9690,N_2582,N_1660);
nand U9691 (N_9691,N_2725,N_4065);
nand U9692 (N_9692,N_733,N_4117);
nor U9693 (N_9693,N_3270,N_1058);
xor U9694 (N_9694,N_4708,N_2315);
nor U9695 (N_9695,N_4455,N_1419);
xnor U9696 (N_9696,N_746,N_1002);
nand U9697 (N_9697,N_465,N_4502);
nand U9698 (N_9698,N_2983,N_2720);
or U9699 (N_9699,N_4106,N_2922);
and U9700 (N_9700,N_1898,N_65);
nand U9701 (N_9701,N_1310,N_2989);
and U9702 (N_9702,N_2090,N_689);
and U9703 (N_9703,N_1668,N_1275);
xnor U9704 (N_9704,N_1976,N_4617);
and U9705 (N_9705,N_1710,N_1777);
and U9706 (N_9706,N_3495,N_3766);
nor U9707 (N_9707,N_2086,N_3609);
and U9708 (N_9708,N_4018,N_3678);
and U9709 (N_9709,N_3163,N_1433);
or U9710 (N_9710,N_1831,N_2678);
and U9711 (N_9711,N_4959,N_3516);
nor U9712 (N_9712,N_284,N_2232);
nand U9713 (N_9713,N_2635,N_292);
nor U9714 (N_9714,N_1520,N_3711);
nor U9715 (N_9715,N_2429,N_2811);
nor U9716 (N_9716,N_3987,N_2656);
and U9717 (N_9717,N_2696,N_4520);
nor U9718 (N_9718,N_3228,N_4520);
nand U9719 (N_9719,N_1407,N_2014);
nor U9720 (N_9720,N_1219,N_1395);
or U9721 (N_9721,N_2583,N_556);
or U9722 (N_9722,N_4601,N_2837);
nand U9723 (N_9723,N_102,N_96);
and U9724 (N_9724,N_1139,N_3744);
nor U9725 (N_9725,N_137,N_3166);
nor U9726 (N_9726,N_256,N_3861);
xor U9727 (N_9727,N_2516,N_2330);
and U9728 (N_9728,N_3162,N_840);
and U9729 (N_9729,N_3350,N_3417);
or U9730 (N_9730,N_2266,N_1965);
nor U9731 (N_9731,N_4546,N_4850);
nor U9732 (N_9732,N_2515,N_4361);
or U9733 (N_9733,N_3521,N_3974);
or U9734 (N_9734,N_1851,N_1055);
and U9735 (N_9735,N_1527,N_3766);
xnor U9736 (N_9736,N_2290,N_4134);
or U9737 (N_9737,N_3566,N_2406);
and U9738 (N_9738,N_1007,N_1481);
nor U9739 (N_9739,N_826,N_1221);
nor U9740 (N_9740,N_254,N_1156);
and U9741 (N_9741,N_2982,N_2394);
xor U9742 (N_9742,N_1371,N_2472);
or U9743 (N_9743,N_2250,N_3977);
nor U9744 (N_9744,N_3785,N_3677);
nor U9745 (N_9745,N_4105,N_354);
xor U9746 (N_9746,N_3040,N_3598);
xor U9747 (N_9747,N_1353,N_3565);
nand U9748 (N_9748,N_1950,N_513);
or U9749 (N_9749,N_1233,N_172);
and U9750 (N_9750,N_998,N_2051);
nor U9751 (N_9751,N_3728,N_2924);
xnor U9752 (N_9752,N_3239,N_1398);
nand U9753 (N_9753,N_1668,N_2162);
and U9754 (N_9754,N_390,N_4624);
and U9755 (N_9755,N_2923,N_2424);
and U9756 (N_9756,N_2437,N_568);
nand U9757 (N_9757,N_3757,N_4858);
or U9758 (N_9758,N_4308,N_2736);
nand U9759 (N_9759,N_255,N_2052);
nor U9760 (N_9760,N_4628,N_3446);
nand U9761 (N_9761,N_707,N_385);
and U9762 (N_9762,N_518,N_142);
and U9763 (N_9763,N_1702,N_1952);
or U9764 (N_9764,N_3411,N_978);
nand U9765 (N_9765,N_1064,N_800);
nand U9766 (N_9766,N_4109,N_1236);
nand U9767 (N_9767,N_2155,N_3680);
nand U9768 (N_9768,N_490,N_1370);
or U9769 (N_9769,N_3903,N_3834);
or U9770 (N_9770,N_499,N_2307);
nor U9771 (N_9771,N_811,N_4754);
xnor U9772 (N_9772,N_2474,N_638);
and U9773 (N_9773,N_1751,N_2288);
xnor U9774 (N_9774,N_3193,N_4327);
nor U9775 (N_9775,N_4461,N_503);
nand U9776 (N_9776,N_30,N_3204);
nand U9777 (N_9777,N_4448,N_2129);
nor U9778 (N_9778,N_968,N_55);
and U9779 (N_9779,N_3844,N_1996);
xnor U9780 (N_9780,N_4953,N_857);
nor U9781 (N_9781,N_149,N_3082);
xor U9782 (N_9782,N_2766,N_189);
nand U9783 (N_9783,N_4304,N_4423);
nand U9784 (N_9784,N_3045,N_3845);
and U9785 (N_9785,N_3178,N_692);
xnor U9786 (N_9786,N_2508,N_939);
or U9787 (N_9787,N_568,N_3450);
or U9788 (N_9788,N_4951,N_3874);
nor U9789 (N_9789,N_2790,N_3347);
nand U9790 (N_9790,N_767,N_2364);
or U9791 (N_9791,N_198,N_2918);
xor U9792 (N_9792,N_4392,N_4819);
or U9793 (N_9793,N_4915,N_2275);
or U9794 (N_9794,N_2975,N_2232);
xor U9795 (N_9795,N_2042,N_4595);
nor U9796 (N_9796,N_1863,N_4714);
or U9797 (N_9797,N_84,N_308);
and U9798 (N_9798,N_2675,N_161);
or U9799 (N_9799,N_2614,N_520);
or U9800 (N_9800,N_337,N_4635);
xor U9801 (N_9801,N_2371,N_356);
xor U9802 (N_9802,N_4128,N_4406);
nor U9803 (N_9803,N_2927,N_468);
and U9804 (N_9804,N_4727,N_168);
and U9805 (N_9805,N_3007,N_729);
nand U9806 (N_9806,N_2645,N_4476);
xor U9807 (N_9807,N_4859,N_1458);
nor U9808 (N_9808,N_3646,N_2681);
or U9809 (N_9809,N_2903,N_2991);
and U9810 (N_9810,N_2711,N_4000);
or U9811 (N_9811,N_1911,N_4805);
or U9812 (N_9812,N_229,N_1314);
nor U9813 (N_9813,N_4221,N_816);
and U9814 (N_9814,N_1570,N_2769);
or U9815 (N_9815,N_2861,N_1721);
and U9816 (N_9816,N_3175,N_2192);
nor U9817 (N_9817,N_844,N_3722);
nand U9818 (N_9818,N_4156,N_1996);
xnor U9819 (N_9819,N_1232,N_2808);
or U9820 (N_9820,N_1476,N_1243);
or U9821 (N_9821,N_4680,N_2114);
and U9822 (N_9822,N_4727,N_1268);
and U9823 (N_9823,N_4499,N_4343);
nand U9824 (N_9824,N_3364,N_1477);
xnor U9825 (N_9825,N_3468,N_826);
xor U9826 (N_9826,N_1411,N_4976);
nand U9827 (N_9827,N_2612,N_742);
xor U9828 (N_9828,N_4218,N_3192);
xnor U9829 (N_9829,N_495,N_4643);
nand U9830 (N_9830,N_3877,N_3316);
xor U9831 (N_9831,N_458,N_4787);
and U9832 (N_9832,N_640,N_3610);
or U9833 (N_9833,N_3052,N_4012);
and U9834 (N_9834,N_565,N_4834);
xor U9835 (N_9835,N_1001,N_1736);
nand U9836 (N_9836,N_1813,N_2705);
nand U9837 (N_9837,N_3458,N_1213);
nand U9838 (N_9838,N_667,N_859);
and U9839 (N_9839,N_4169,N_3173);
nand U9840 (N_9840,N_2728,N_906);
and U9841 (N_9841,N_1817,N_4375);
and U9842 (N_9842,N_2862,N_4670);
and U9843 (N_9843,N_657,N_1987);
and U9844 (N_9844,N_3444,N_4069);
nand U9845 (N_9845,N_1169,N_4886);
and U9846 (N_9846,N_4304,N_3071);
and U9847 (N_9847,N_3625,N_1096);
nor U9848 (N_9848,N_4779,N_1947);
or U9849 (N_9849,N_1265,N_4124);
xnor U9850 (N_9850,N_1577,N_732);
xnor U9851 (N_9851,N_2336,N_1750);
xor U9852 (N_9852,N_1017,N_4710);
and U9853 (N_9853,N_4836,N_1879);
and U9854 (N_9854,N_3111,N_2746);
nor U9855 (N_9855,N_607,N_4637);
xor U9856 (N_9856,N_919,N_2074);
nand U9857 (N_9857,N_3327,N_4641);
and U9858 (N_9858,N_4330,N_1513);
xor U9859 (N_9859,N_4737,N_2536);
nor U9860 (N_9860,N_4755,N_961);
and U9861 (N_9861,N_4183,N_1973);
nand U9862 (N_9862,N_52,N_219);
or U9863 (N_9863,N_549,N_1880);
or U9864 (N_9864,N_4295,N_3506);
and U9865 (N_9865,N_3754,N_2462);
nor U9866 (N_9866,N_3238,N_2484);
nand U9867 (N_9867,N_1469,N_1841);
xor U9868 (N_9868,N_4490,N_4267);
and U9869 (N_9869,N_2875,N_603);
nor U9870 (N_9870,N_3784,N_974);
or U9871 (N_9871,N_3779,N_112);
or U9872 (N_9872,N_2367,N_1317);
xnor U9873 (N_9873,N_137,N_3086);
nor U9874 (N_9874,N_4632,N_595);
nor U9875 (N_9875,N_4232,N_4193);
xnor U9876 (N_9876,N_4551,N_1833);
nor U9877 (N_9877,N_3798,N_654);
xor U9878 (N_9878,N_4310,N_1776);
or U9879 (N_9879,N_633,N_2444);
or U9880 (N_9880,N_346,N_4191);
nand U9881 (N_9881,N_2159,N_2782);
xor U9882 (N_9882,N_1409,N_1082);
or U9883 (N_9883,N_4941,N_2136);
or U9884 (N_9884,N_2872,N_3709);
or U9885 (N_9885,N_3208,N_2274);
nand U9886 (N_9886,N_2948,N_1434);
and U9887 (N_9887,N_3981,N_2215);
and U9888 (N_9888,N_2816,N_4731);
nand U9889 (N_9889,N_3085,N_2465);
nand U9890 (N_9890,N_3280,N_4660);
nand U9891 (N_9891,N_94,N_81);
xor U9892 (N_9892,N_2063,N_1758);
and U9893 (N_9893,N_120,N_685);
or U9894 (N_9894,N_3633,N_4975);
nor U9895 (N_9895,N_374,N_3525);
nor U9896 (N_9896,N_1163,N_1341);
nand U9897 (N_9897,N_1160,N_2908);
or U9898 (N_9898,N_1924,N_695);
nor U9899 (N_9899,N_3651,N_3659);
and U9900 (N_9900,N_3815,N_1822);
and U9901 (N_9901,N_1873,N_2464);
xnor U9902 (N_9902,N_1592,N_4637);
nand U9903 (N_9903,N_653,N_220);
and U9904 (N_9904,N_3705,N_3114);
or U9905 (N_9905,N_4092,N_2206);
and U9906 (N_9906,N_3718,N_4351);
or U9907 (N_9907,N_1509,N_4289);
nor U9908 (N_9908,N_297,N_4035);
nor U9909 (N_9909,N_4078,N_1446);
or U9910 (N_9910,N_3305,N_1041);
nor U9911 (N_9911,N_2862,N_1529);
and U9912 (N_9912,N_3247,N_2319);
xor U9913 (N_9913,N_1163,N_124);
nor U9914 (N_9914,N_3883,N_885);
and U9915 (N_9915,N_869,N_3820);
nor U9916 (N_9916,N_3070,N_4237);
xnor U9917 (N_9917,N_3439,N_1534);
nor U9918 (N_9918,N_2501,N_4421);
xnor U9919 (N_9919,N_828,N_1470);
or U9920 (N_9920,N_4132,N_627);
or U9921 (N_9921,N_1712,N_5);
nand U9922 (N_9922,N_4999,N_2940);
nor U9923 (N_9923,N_1049,N_2648);
or U9924 (N_9924,N_1759,N_1357);
xor U9925 (N_9925,N_1414,N_2665);
nand U9926 (N_9926,N_4120,N_2439);
and U9927 (N_9927,N_1430,N_347);
or U9928 (N_9928,N_3923,N_3238);
nand U9929 (N_9929,N_4262,N_2296);
and U9930 (N_9930,N_1719,N_2896);
xnor U9931 (N_9931,N_3729,N_1356);
or U9932 (N_9932,N_4163,N_1648);
nor U9933 (N_9933,N_2455,N_4655);
and U9934 (N_9934,N_693,N_4508);
xnor U9935 (N_9935,N_545,N_1529);
nor U9936 (N_9936,N_4709,N_3585);
or U9937 (N_9937,N_1777,N_4202);
xnor U9938 (N_9938,N_724,N_4837);
and U9939 (N_9939,N_493,N_754);
xnor U9940 (N_9940,N_4276,N_2188);
or U9941 (N_9941,N_3701,N_420);
and U9942 (N_9942,N_1475,N_2901);
nand U9943 (N_9943,N_1466,N_4845);
or U9944 (N_9944,N_369,N_2962);
or U9945 (N_9945,N_4830,N_348);
or U9946 (N_9946,N_1390,N_4850);
nand U9947 (N_9947,N_4481,N_3505);
and U9948 (N_9948,N_24,N_2275);
nor U9949 (N_9949,N_4138,N_1853);
nand U9950 (N_9950,N_3483,N_2170);
and U9951 (N_9951,N_4032,N_1484);
nor U9952 (N_9952,N_2757,N_1256);
nand U9953 (N_9953,N_1690,N_2438);
and U9954 (N_9954,N_4895,N_812);
and U9955 (N_9955,N_4278,N_3727);
nand U9956 (N_9956,N_2416,N_4387);
xor U9957 (N_9957,N_414,N_2163);
or U9958 (N_9958,N_1289,N_3578);
xor U9959 (N_9959,N_2753,N_4135);
xor U9960 (N_9960,N_136,N_2023);
xor U9961 (N_9961,N_476,N_881);
nand U9962 (N_9962,N_4055,N_3035);
xnor U9963 (N_9963,N_210,N_992);
or U9964 (N_9964,N_2335,N_755);
and U9965 (N_9965,N_1099,N_4691);
xnor U9966 (N_9966,N_3504,N_4874);
nor U9967 (N_9967,N_2298,N_4799);
and U9968 (N_9968,N_1419,N_2728);
nor U9969 (N_9969,N_3530,N_1266);
nand U9970 (N_9970,N_4174,N_4491);
or U9971 (N_9971,N_3248,N_3331);
xor U9972 (N_9972,N_2751,N_3692);
nor U9973 (N_9973,N_3404,N_3104);
and U9974 (N_9974,N_1679,N_4986);
xor U9975 (N_9975,N_172,N_1476);
or U9976 (N_9976,N_1953,N_4473);
nor U9977 (N_9977,N_2287,N_2344);
nor U9978 (N_9978,N_1174,N_3679);
nor U9979 (N_9979,N_4320,N_128);
nand U9980 (N_9980,N_585,N_1879);
and U9981 (N_9981,N_515,N_2788);
nand U9982 (N_9982,N_1545,N_1221);
and U9983 (N_9983,N_4288,N_660);
nand U9984 (N_9984,N_2538,N_2242);
nand U9985 (N_9985,N_3288,N_56);
xor U9986 (N_9986,N_4171,N_400);
and U9987 (N_9987,N_3656,N_3719);
and U9988 (N_9988,N_1450,N_3333);
and U9989 (N_9989,N_3950,N_880);
and U9990 (N_9990,N_1105,N_1160);
or U9991 (N_9991,N_4698,N_3612);
xor U9992 (N_9992,N_3012,N_1020);
xnor U9993 (N_9993,N_4866,N_2363);
xnor U9994 (N_9994,N_3715,N_1636);
or U9995 (N_9995,N_4697,N_3370);
xnor U9996 (N_9996,N_74,N_4266);
xor U9997 (N_9997,N_2633,N_4788);
or U9998 (N_9998,N_4591,N_858);
xnor U9999 (N_9999,N_62,N_718);
xor U10000 (N_10000,N_9292,N_6136);
xor U10001 (N_10001,N_8308,N_5150);
or U10002 (N_10002,N_6040,N_6051);
and U10003 (N_10003,N_5681,N_7097);
xnor U10004 (N_10004,N_5479,N_7338);
and U10005 (N_10005,N_9061,N_5677);
or U10006 (N_10006,N_6841,N_7614);
nor U10007 (N_10007,N_9725,N_8555);
or U10008 (N_10008,N_6364,N_6579);
or U10009 (N_10009,N_9450,N_5546);
nand U10010 (N_10010,N_6050,N_5971);
or U10011 (N_10011,N_8892,N_9182);
xor U10012 (N_10012,N_8982,N_9038);
xnor U10013 (N_10013,N_7836,N_9935);
nor U10014 (N_10014,N_5032,N_8082);
or U10015 (N_10015,N_8448,N_8239);
nand U10016 (N_10016,N_7281,N_8581);
nor U10017 (N_10017,N_5423,N_8145);
nor U10018 (N_10018,N_6906,N_6299);
or U10019 (N_10019,N_5612,N_9624);
nand U10020 (N_10020,N_5721,N_8821);
and U10021 (N_10021,N_7298,N_6154);
or U10022 (N_10022,N_5236,N_5338);
and U10023 (N_10023,N_6010,N_7823);
and U10024 (N_10024,N_7531,N_7885);
or U10025 (N_10025,N_9246,N_5140);
nor U10026 (N_10026,N_9490,N_7718);
nor U10027 (N_10027,N_9621,N_6560);
xnor U10028 (N_10028,N_8087,N_5081);
and U10029 (N_10029,N_8961,N_5895);
and U10030 (N_10030,N_5038,N_9667);
nand U10031 (N_10031,N_9976,N_5171);
nand U10032 (N_10032,N_5824,N_5389);
nand U10033 (N_10033,N_9794,N_9817);
or U10034 (N_10034,N_7131,N_6362);
nand U10035 (N_10035,N_5607,N_8538);
or U10036 (N_10036,N_6496,N_6721);
nand U10037 (N_10037,N_6619,N_9938);
or U10038 (N_10038,N_9748,N_6885);
xor U10039 (N_10039,N_7840,N_9287);
and U10040 (N_10040,N_9379,N_6416);
nor U10041 (N_10041,N_6336,N_7665);
nand U10042 (N_10042,N_6564,N_6803);
xor U10043 (N_10043,N_7814,N_7103);
or U10044 (N_10044,N_8282,N_5601);
or U10045 (N_10045,N_8384,N_9240);
xor U10046 (N_10046,N_7457,N_8419);
xnor U10047 (N_10047,N_8013,N_5745);
nand U10048 (N_10048,N_7164,N_8460);
nand U10049 (N_10049,N_6012,N_6300);
nand U10050 (N_10050,N_5536,N_8339);
nor U10051 (N_10051,N_7162,N_9630);
nand U10052 (N_10052,N_7036,N_8285);
and U10053 (N_10053,N_5242,N_5420);
xnor U10054 (N_10054,N_6848,N_5221);
and U10055 (N_10055,N_9361,N_7916);
or U10056 (N_10056,N_9496,N_6297);
xnor U10057 (N_10057,N_5588,N_5282);
and U10058 (N_10058,N_6189,N_9284);
nand U10059 (N_10059,N_9632,N_9552);
or U10060 (N_10060,N_8995,N_7236);
and U10061 (N_10061,N_9645,N_8932);
nand U10062 (N_10062,N_5443,N_9278);
or U10063 (N_10063,N_5910,N_6630);
or U10064 (N_10064,N_6174,N_7721);
or U10065 (N_10065,N_9875,N_9074);
or U10066 (N_10066,N_7636,N_8747);
nor U10067 (N_10067,N_5089,N_9824);
nand U10068 (N_10068,N_6184,N_6991);
xnor U10069 (N_10069,N_8700,N_8847);
nand U10070 (N_10070,N_8710,N_7908);
and U10071 (N_10071,N_5117,N_8634);
or U10072 (N_10072,N_9364,N_5432);
nor U10073 (N_10073,N_5245,N_5956);
xor U10074 (N_10074,N_7589,N_9729);
xnor U10075 (N_10075,N_7137,N_6175);
nand U10076 (N_10076,N_7657,N_6891);
xnor U10077 (N_10077,N_5699,N_7535);
nor U10078 (N_10078,N_8449,N_8949);
and U10079 (N_10079,N_6983,N_7556);
and U10080 (N_10080,N_6463,N_5967);
and U10081 (N_10081,N_5813,N_5156);
nand U10082 (N_10082,N_7024,N_8111);
or U10083 (N_10083,N_5115,N_7639);
and U10084 (N_10084,N_9285,N_5944);
xnor U10085 (N_10085,N_9017,N_5387);
or U10086 (N_10086,N_5505,N_5010);
and U10087 (N_10087,N_8766,N_6015);
nand U10088 (N_10088,N_7980,N_9759);
xnor U10089 (N_10089,N_8610,N_9649);
xnor U10090 (N_10090,N_6753,N_5599);
nor U10091 (N_10091,N_7355,N_7749);
nand U10092 (N_10092,N_5110,N_9111);
nor U10093 (N_10093,N_8655,N_5873);
nand U10094 (N_10094,N_7870,N_7524);
nand U10095 (N_10095,N_9333,N_8341);
nor U10096 (N_10096,N_6859,N_7660);
or U10097 (N_10097,N_7929,N_9521);
nor U10098 (N_10098,N_7901,N_5593);
xnor U10099 (N_10099,N_5399,N_6536);
xnor U10100 (N_10100,N_6747,N_6361);
nand U10101 (N_10101,N_9627,N_9427);
or U10102 (N_10102,N_5487,N_9719);
and U10103 (N_10103,N_6858,N_9513);
or U10104 (N_10104,N_9181,N_9788);
or U10105 (N_10105,N_6277,N_6759);
xor U10106 (N_10106,N_6041,N_9110);
nor U10107 (N_10107,N_8957,N_5583);
and U10108 (N_10108,N_8675,N_9377);
xnor U10109 (N_10109,N_9105,N_8180);
and U10110 (N_10110,N_6992,N_9234);
or U10111 (N_10111,N_8377,N_8006);
xor U10112 (N_10112,N_7565,N_8836);
nor U10113 (N_10113,N_7922,N_5059);
xor U10114 (N_10114,N_8148,N_8474);
and U10115 (N_10115,N_8043,N_6679);
xnor U10116 (N_10116,N_7456,N_8576);
and U10117 (N_10117,N_9943,N_7654);
or U10118 (N_10118,N_7742,N_8992);
nor U10119 (N_10119,N_8191,N_9389);
nand U10120 (N_10120,N_6457,N_5142);
and U10121 (N_10121,N_7089,N_6166);
nor U10122 (N_10122,N_6818,N_9332);
nor U10123 (N_10123,N_5569,N_7093);
or U10124 (N_10124,N_6168,N_5416);
or U10125 (N_10125,N_8073,N_9214);
nand U10126 (N_10126,N_9233,N_9149);
xnor U10127 (N_10127,N_6107,N_5698);
or U10128 (N_10128,N_6478,N_6220);
nand U10129 (N_10129,N_7384,N_6898);
xor U10130 (N_10130,N_9020,N_8653);
and U10131 (N_10131,N_9779,N_7612);
nor U10132 (N_10132,N_6837,N_7017);
and U10133 (N_10133,N_5608,N_7078);
and U10134 (N_10134,N_7926,N_9668);
nand U10135 (N_10135,N_8939,N_8107);
nor U10136 (N_10136,N_5957,N_5326);
and U10137 (N_10137,N_9541,N_9777);
nand U10138 (N_10138,N_8228,N_7973);
nor U10139 (N_10139,N_9901,N_5853);
and U10140 (N_10140,N_8058,N_5336);
and U10141 (N_10141,N_5237,N_5587);
nor U10142 (N_10142,N_9544,N_8519);
xnor U10143 (N_10143,N_6755,N_7307);
and U10144 (N_10144,N_7573,N_7308);
or U10145 (N_10145,N_6485,N_8876);
xnor U10146 (N_10146,N_6371,N_7874);
or U10147 (N_10147,N_7372,N_6698);
and U10148 (N_10148,N_8647,N_8959);
nor U10149 (N_10149,N_9067,N_6238);
xnor U10150 (N_10150,N_6521,N_9307);
and U10151 (N_10151,N_7702,N_7163);
nor U10152 (N_10152,N_7149,N_6825);
nand U10153 (N_10153,N_9986,N_8160);
or U10154 (N_10154,N_6352,N_9642);
nor U10155 (N_10155,N_7116,N_8556);
nand U10156 (N_10156,N_9732,N_8866);
or U10157 (N_10157,N_9955,N_9699);
and U10158 (N_10158,N_9727,N_7489);
nor U10159 (N_10159,N_7268,N_8170);
and U10160 (N_10160,N_7506,N_9972);
nor U10161 (N_10161,N_9420,N_8953);
or U10162 (N_10162,N_9706,N_8965);
nor U10163 (N_10163,N_5567,N_5259);
and U10164 (N_10164,N_7509,N_6545);
nand U10165 (N_10165,N_9394,N_6172);
xnor U10166 (N_10166,N_6195,N_9454);
xnor U10167 (N_10167,N_9353,N_6023);
and U10168 (N_10168,N_8758,N_9228);
or U10169 (N_10169,N_6910,N_9126);
and U10170 (N_10170,N_9549,N_8664);
nand U10171 (N_10171,N_6334,N_8832);
nor U10172 (N_10172,N_7054,N_9478);
nor U10173 (N_10173,N_9428,N_6732);
xor U10174 (N_10174,N_8728,N_6231);
or U10175 (N_10175,N_7864,N_5973);
and U10176 (N_10176,N_5785,N_9658);
or U10177 (N_10177,N_6090,N_6607);
or U10178 (N_10178,N_5070,N_9969);
xor U10179 (N_10179,N_5923,N_7817);
nor U10180 (N_10180,N_9674,N_8739);
nand U10181 (N_10181,N_8571,N_5276);
or U10182 (N_10182,N_9147,N_8410);
nand U10183 (N_10183,N_5342,N_6280);
and U10184 (N_10184,N_5535,N_6538);
nor U10185 (N_10185,N_7959,N_7831);
nand U10186 (N_10186,N_7315,N_9470);
nor U10187 (N_10187,N_8184,N_5462);
and U10188 (N_10188,N_9753,N_5120);
nand U10189 (N_10189,N_6053,N_5656);
nand U10190 (N_10190,N_9328,N_5468);
nand U10191 (N_10191,N_6613,N_8105);
and U10192 (N_10192,N_8386,N_6928);
nor U10193 (N_10193,N_8679,N_8331);
nand U10194 (N_10194,N_6286,N_5868);
nand U10195 (N_10195,N_6530,N_9184);
nor U10196 (N_10196,N_8681,N_5606);
or U10197 (N_10197,N_8383,N_9906);
xor U10198 (N_10198,N_6969,N_6420);
nand U10199 (N_10199,N_7580,N_9712);
or U10200 (N_10200,N_9447,N_9888);
and U10201 (N_10201,N_6654,N_9516);
xor U10202 (N_10202,N_7157,N_5643);
nor U10203 (N_10203,N_9601,N_8888);
nand U10204 (N_10204,N_5625,N_9078);
nand U10205 (N_10205,N_5347,N_5794);
nor U10206 (N_10206,N_6594,N_9960);
xor U10207 (N_10207,N_8085,N_7518);
or U10208 (N_10208,N_9306,N_9599);
and U10209 (N_10209,N_9646,N_9019);
nor U10210 (N_10210,N_6513,N_5159);
nand U10211 (N_10211,N_5859,N_7627);
and U10212 (N_10212,N_9188,N_5284);
or U10213 (N_10213,N_5321,N_7354);
nor U10214 (N_10214,N_6633,N_5410);
and U10215 (N_10215,N_8201,N_7205);
nand U10216 (N_10216,N_6216,N_8176);
xnor U10217 (N_10217,N_7300,N_6271);
nand U10218 (N_10218,N_6740,N_6659);
xnor U10219 (N_10219,N_9979,N_8935);
nor U10220 (N_10220,N_6417,N_5015);
and U10221 (N_10221,N_8324,N_6715);
and U10222 (N_10222,N_6735,N_6965);
xnor U10223 (N_10223,N_5368,N_7217);
nand U10224 (N_10224,N_9553,N_9354);
and U10225 (N_10225,N_8607,N_5844);
nand U10226 (N_10226,N_9066,N_7925);
or U10227 (N_10227,N_5870,N_7053);
or U10228 (N_10228,N_6527,N_9302);
nand U10229 (N_10229,N_9161,N_6877);
and U10230 (N_10230,N_8938,N_6274);
and U10231 (N_10231,N_9293,N_8746);
or U10232 (N_10232,N_8596,N_6842);
nor U10233 (N_10233,N_6751,N_6080);
or U10234 (N_10234,N_7529,N_5922);
nand U10235 (N_10235,N_9371,N_6475);
nor U10236 (N_10236,N_7110,N_7195);
nand U10237 (N_10237,N_8485,N_6021);
or U10238 (N_10238,N_6745,N_6767);
nor U10239 (N_10239,N_7108,N_8459);
or U10240 (N_10240,N_6409,N_6451);
or U10241 (N_10241,N_5635,N_5203);
xnor U10242 (N_10242,N_7043,N_6990);
and U10243 (N_10243,N_7343,N_6785);
xnor U10244 (N_10244,N_5497,N_7494);
or U10245 (N_10245,N_6639,N_6318);
xor U10246 (N_10246,N_8335,N_9932);
xor U10247 (N_10247,N_5915,N_7468);
or U10248 (N_10248,N_9772,N_7813);
xor U10249 (N_10249,N_5042,N_6089);
and U10250 (N_10250,N_7486,N_9376);
nand U10251 (N_10251,N_9033,N_7152);
xor U10252 (N_10252,N_6902,N_7821);
or U10253 (N_10253,N_5467,N_6942);
xnor U10254 (N_10254,N_6309,N_6007);
and U10255 (N_10255,N_9408,N_6224);
nand U10256 (N_10256,N_7329,N_7726);
xor U10257 (N_10257,N_5441,N_9143);
or U10258 (N_10258,N_6256,N_6595);
or U10259 (N_10259,N_6319,N_7407);
nor U10260 (N_10260,N_9760,N_6844);
and U10261 (N_10261,N_8985,N_8151);
xor U10262 (N_10262,N_7644,N_9678);
xor U10263 (N_10263,N_6623,N_5207);
xor U10264 (N_10264,N_9030,N_6695);
or U10265 (N_10265,N_6640,N_5706);
and U10266 (N_10266,N_5810,N_9623);
or U10267 (N_10267,N_9119,N_9576);
nor U10268 (N_10268,N_9208,N_8629);
or U10269 (N_10269,N_9031,N_8052);
nand U10270 (N_10270,N_5757,N_9786);
xor U10271 (N_10271,N_7902,N_7290);
or U10272 (N_10272,N_8856,N_7047);
or U10273 (N_10273,N_5506,N_5104);
or U10274 (N_10274,N_6330,N_9296);
xnor U10275 (N_10275,N_8712,N_8908);
and U10276 (N_10276,N_5648,N_8973);
nor U10277 (N_10277,N_8054,N_8473);
and U10278 (N_10278,N_9962,N_6079);
and U10279 (N_10279,N_6047,N_5252);
nor U10280 (N_10280,N_8863,N_5480);
nor U10281 (N_10281,N_5154,N_9254);
nand U10282 (N_10282,N_5437,N_5238);
xnor U10283 (N_10283,N_6285,N_7490);
nand U10284 (N_10284,N_8703,N_8051);
nor U10285 (N_10285,N_8624,N_7410);
or U10286 (N_10286,N_6625,N_9936);
xor U10287 (N_10287,N_6084,N_9224);
and U10288 (N_10288,N_9315,N_8776);
nor U10289 (N_10289,N_8393,N_6348);
nand U10290 (N_10290,N_9403,N_5313);
nand U10291 (N_10291,N_8257,N_5324);
or U10292 (N_10292,N_6452,N_5823);
and U10293 (N_10293,N_8567,N_5921);
and U10294 (N_10294,N_7899,N_8956);
or U10295 (N_10295,N_6028,N_9439);
xnor U10296 (N_10296,N_7561,N_9800);
and U10297 (N_10297,N_6814,N_9052);
nor U10298 (N_10298,N_6546,N_9350);
or U10299 (N_10299,N_8650,N_7398);
or U10300 (N_10300,N_9550,N_5981);
or U10301 (N_10301,N_9511,N_9889);
nand U10302 (N_10302,N_6161,N_5118);
nand U10303 (N_10303,N_8913,N_6367);
or U10304 (N_10304,N_5881,N_5143);
nor U10305 (N_10305,N_5006,N_8027);
nand U10306 (N_10306,N_8352,N_9101);
xnor U10307 (N_10307,N_8903,N_6972);
xnor U10308 (N_10308,N_9839,N_6381);
xor U10309 (N_10309,N_7179,N_7099);
xnor U10310 (N_10310,N_9579,N_7058);
or U10311 (N_10311,N_8875,N_5071);
nand U10312 (N_10312,N_5550,N_7211);
xor U10313 (N_10313,N_6620,N_8857);
and U10314 (N_10314,N_9663,N_7714);
nor U10315 (N_10315,N_8035,N_5948);
xor U10316 (N_10316,N_6544,N_9747);
nand U10317 (N_10317,N_6370,N_8822);
and U10318 (N_10318,N_6415,N_8367);
or U10319 (N_10319,N_7421,N_9483);
nor U10320 (N_10320,N_6569,N_5109);
nand U10321 (N_10321,N_6192,N_8217);
nor U10322 (N_10322,N_9449,N_7231);
and U10323 (N_10323,N_7264,N_5742);
nor U10324 (N_10324,N_5220,N_6374);
nor U10325 (N_10325,N_7632,N_6704);
and U10326 (N_10326,N_9297,N_5703);
nor U10327 (N_10327,N_5604,N_7228);
and U10328 (N_10328,N_9048,N_7375);
nand U10329 (N_10329,N_9411,N_6757);
and U10330 (N_10330,N_6105,N_5894);
xor U10331 (N_10331,N_6567,N_6315);
nor U10332 (N_10332,N_6197,N_8458);
nor U10333 (N_10333,N_7571,N_6480);
xnor U10334 (N_10334,N_5013,N_5575);
or U10335 (N_10335,N_6185,N_7761);
or U10336 (N_10336,N_7363,N_5206);
nand U10337 (N_10337,N_6237,N_5830);
xor U10338 (N_10338,N_9885,N_5210);
nand U10339 (N_10339,N_9073,N_6124);
or U10340 (N_10340,N_7952,N_8838);
or U10341 (N_10341,N_9342,N_7956);
nor U10342 (N_10342,N_9092,N_6295);
or U10343 (N_10343,N_5499,N_9661);
nor U10344 (N_10344,N_7458,N_8967);
or U10345 (N_10345,N_9679,N_9393);
or U10346 (N_10346,N_6155,N_7792);
or U10347 (N_10347,N_8503,N_7334);
xnor U10348 (N_10348,N_8824,N_7880);
or U10349 (N_10349,N_5637,N_5655);
and U10350 (N_10350,N_6213,N_7493);
nand U10351 (N_10351,N_9721,N_7318);
and U10352 (N_10352,N_8560,N_7672);
or U10353 (N_10353,N_9415,N_9963);
and U10354 (N_10354,N_7866,N_7500);
nor U10355 (N_10355,N_5626,N_6181);
or U10356 (N_10356,N_9473,N_8723);
or U10357 (N_10357,N_6997,N_9891);
nor U10358 (N_10358,N_5854,N_7085);
nor U10359 (N_10359,N_8986,N_7275);
or U10360 (N_10360,N_8848,N_8726);
nand U10361 (N_10361,N_9688,N_7664);
or U10362 (N_10362,N_6208,N_6039);
or U10363 (N_10363,N_6046,N_8318);
and U10364 (N_10364,N_9156,N_9993);
and U10365 (N_10365,N_6482,N_8976);
nand U10366 (N_10366,N_8731,N_7904);
xor U10367 (N_10367,N_5050,N_6385);
nand U10368 (N_10368,N_7985,N_6072);
and U10369 (N_10369,N_8493,N_8490);
nor U10370 (N_10370,N_9175,N_5791);
nor U10371 (N_10371,N_8994,N_5363);
or U10372 (N_10372,N_6800,N_8140);
xor U10373 (N_10373,N_6995,N_9499);
or U10374 (N_10374,N_8288,N_8498);
nor U10375 (N_10375,N_6850,N_6832);
nand U10376 (N_10376,N_5543,N_7540);
xor U10377 (N_10377,N_9382,N_8411);
and U10378 (N_10378,N_8934,N_5809);
xor U10379 (N_10379,N_6020,N_9141);
and U10380 (N_10380,N_6383,N_8198);
or U10381 (N_10381,N_6043,N_5357);
or U10382 (N_10382,N_6522,N_9273);
xor U10383 (N_10383,N_6784,N_6982);
nor U10384 (N_10384,N_8488,N_9804);
or U10385 (N_10385,N_8553,N_6943);
nand U10386 (N_10386,N_5179,N_5380);
or U10387 (N_10387,N_5557,N_6100);
or U10388 (N_10388,N_7747,N_8253);
nor U10389 (N_10389,N_8868,N_9247);
nand U10390 (N_10390,N_7400,N_7596);
xor U10391 (N_10391,N_8842,N_5461);
xor U10392 (N_10392,N_5063,N_7434);
and U10393 (N_10393,N_7168,N_8918);
nand U10394 (N_10394,N_5771,N_5585);
and U10395 (N_10395,N_5805,N_9933);
and U10396 (N_10396,N_6118,N_7402);
xor U10397 (N_10397,N_5724,N_9050);
nand U10398 (N_10398,N_9947,N_9456);
nand U10399 (N_10399,N_5934,N_9244);
or U10400 (N_10400,N_9262,N_9977);
and U10401 (N_10401,N_8302,N_6699);
nand U10402 (N_10402,N_7577,N_8867);
or U10403 (N_10403,N_8820,N_9555);
nand U10404 (N_10404,N_6575,N_8770);
or U10405 (N_10405,N_5958,N_5527);
or U10406 (N_10406,N_8778,N_8414);
nand U10407 (N_10407,N_9647,N_6686);
nand U10408 (N_10408,N_5620,N_7087);
nand U10409 (N_10409,N_6874,N_8350);
and U10410 (N_10410,N_6422,N_6988);
or U10411 (N_10411,N_9303,N_5216);
nand U10412 (N_10412,N_7674,N_6541);
xor U10413 (N_10413,N_6535,N_6186);
and U10414 (N_10414,N_5350,N_7301);
nand U10415 (N_10415,N_5086,N_7186);
xor U10416 (N_10416,N_9968,N_7252);
nor U10417 (N_10417,N_9144,N_8855);
and U10418 (N_10418,N_8173,N_9745);
or U10419 (N_10419,N_9185,N_5534);
or U10420 (N_10420,N_9488,N_8455);
and U10421 (N_10421,N_5827,N_6217);
nand U10422 (N_10422,N_6345,N_8181);
xor U10423 (N_10423,N_9311,N_7691);
nand U10424 (N_10424,N_9931,N_9413);
nor U10425 (N_10425,N_7013,N_8740);
nor U10426 (N_10426,N_6221,N_9662);
nor U10427 (N_10427,N_8660,N_6289);
xor U10428 (N_10428,N_9012,N_9225);
nand U10429 (N_10429,N_9929,N_7610);
and U10430 (N_10430,N_9040,N_5214);
and U10431 (N_10431,N_6391,N_7746);
xor U10432 (N_10432,N_5440,N_5586);
xnor U10433 (N_10433,N_7933,N_6616);
nand U10434 (N_10434,N_9220,N_7026);
or U10435 (N_10435,N_9298,N_7125);
xor U10436 (N_10436,N_9299,N_7142);
or U10437 (N_10437,N_7428,N_7616);
nor U10438 (N_10438,N_6812,N_5343);
xnor U10439 (N_10439,N_8428,N_7005);
xor U10440 (N_10440,N_7359,N_7436);
or U10441 (N_10441,N_6250,N_6909);
or U10442 (N_10442,N_8260,N_5163);
nor U10443 (N_10443,N_6888,N_7133);
nor U10444 (N_10444,N_6490,N_5865);
xnor U10445 (N_10445,N_5223,N_8344);
and U10446 (N_10446,N_5621,N_5867);
nand U10447 (N_10447,N_9452,N_9265);
nand U10448 (N_10448,N_5036,N_6102);
or U10449 (N_10449,N_7845,N_6957);
and U10450 (N_10450,N_6660,N_6954);
and U10451 (N_10451,N_6986,N_9819);
or U10452 (N_10452,N_8415,N_5014);
and U10453 (N_10453,N_9118,N_6338);
and U10454 (N_10454,N_5660,N_8423);
xnor U10455 (N_10455,N_7481,N_9603);
nand U10456 (N_10456,N_8036,N_8227);
and U10457 (N_10457,N_9357,N_5933);
and U10458 (N_10458,N_9589,N_6222);
xor U10459 (N_10459,N_8907,N_8835);
nor U10460 (N_10460,N_7101,N_5776);
nand U10461 (N_10461,N_7272,N_8646);
nand U10462 (N_10462,N_9169,N_8117);
or U10463 (N_10463,N_6343,N_8319);
and U10464 (N_10464,N_6789,N_7071);
nor U10465 (N_10465,N_6109,N_7000);
nor U10466 (N_10466,N_6293,N_5168);
xor U10467 (N_10467,N_9372,N_7852);
nand U10468 (N_10468,N_5838,N_7451);
or U10469 (N_10469,N_9942,N_8144);
xor U10470 (N_10470,N_8642,N_7160);
nor U10471 (N_10471,N_5084,N_7304);
nand U10472 (N_10472,N_7470,N_9352);
or U10473 (N_10473,N_5056,N_8923);
or U10474 (N_10474,N_6473,N_8002);
xnor U10475 (N_10475,N_6183,N_5918);
nand U10476 (N_10476,N_9590,N_5365);
or U10477 (N_10477,N_5629,N_6458);
and U10478 (N_10478,N_8549,N_9770);
and U10479 (N_10479,N_5227,N_5714);
xor U10480 (N_10480,N_5307,N_5502);
xor U10481 (N_10481,N_7669,N_8912);
nor U10482 (N_10482,N_9453,N_8153);
nor U10483 (N_10483,N_8042,N_9807);
and U10484 (N_10484,N_6426,N_5875);
or U10485 (N_10485,N_8385,N_5683);
xnor U10486 (N_10486,N_9854,N_6855);
or U10487 (N_10487,N_8944,N_6406);
xor U10488 (N_10488,N_8483,N_9459);
xor U10489 (N_10489,N_5149,N_8958);
or U10490 (N_10490,N_7191,N_5997);
and U10491 (N_10491,N_6069,N_5576);
nand U10492 (N_10492,N_7937,N_6064);
and U10493 (N_10493,N_7215,N_6147);
or U10494 (N_10494,N_9858,N_8438);
nor U10495 (N_10495,N_9381,N_8130);
nand U10496 (N_10496,N_5740,N_8094);
nor U10497 (N_10497,N_8436,N_6796);
nor U10498 (N_10498,N_6266,N_9122);
and U10499 (N_10499,N_8074,N_9565);
nand U10500 (N_10500,N_6158,N_8584);
nor U10501 (N_10501,N_6498,N_6889);
and U10502 (N_10502,N_5391,N_7221);
xor U10503 (N_10503,N_7716,N_8590);
and U10504 (N_10504,N_5419,N_6907);
or U10505 (N_10505,N_7807,N_8790);
xnor U10506 (N_10506,N_9641,N_6897);
nand U10507 (N_10507,N_9847,N_9840);
and U10508 (N_10508,N_8182,N_9384);
xor U10509 (N_10509,N_5209,N_7846);
or U10510 (N_10510,N_6141,N_8696);
nand U10511 (N_10511,N_6746,N_6143);
or U10512 (N_10512,N_9681,N_7176);
and U10513 (N_10513,N_5178,N_8550);
nor U10514 (N_10514,N_9226,N_9675);
xnor U10515 (N_10515,N_6648,N_7537);
nor U10516 (N_10516,N_6781,N_5349);
nor U10517 (N_10517,N_6313,N_8524);
nor U10518 (N_10518,N_7467,N_8089);
and U10519 (N_10519,N_5951,N_9952);
nand U10520 (N_10520,N_8190,N_6156);
and U10521 (N_10521,N_8216,N_7257);
xor U10522 (N_10522,N_5723,N_5067);
and U10523 (N_10523,N_9063,N_6034);
xnor U10524 (N_10524,N_9618,N_7797);
or U10525 (N_10525,N_8463,N_8240);
nor U10526 (N_10526,N_8095,N_5533);
xnor U10527 (N_10527,N_5820,N_9945);
nand U10528 (N_10528,N_7649,N_5968);
or U10529 (N_10529,N_9016,N_8505);
nor U10530 (N_10530,N_5891,N_9577);
and U10531 (N_10531,N_5026,N_6097);
nor U10532 (N_10532,N_7618,N_7733);
and U10533 (N_10533,N_6783,N_5815);
nor U10534 (N_10534,N_6306,N_7136);
xor U10535 (N_10535,N_7905,N_5458);
nand U10536 (N_10536,N_6776,N_7358);
nor U10537 (N_10537,N_7951,N_9008);
nand U10538 (N_10538,N_6244,N_7543);
nor U10539 (N_10539,N_5687,N_6499);
and U10540 (N_10540,N_9150,N_9173);
and U10541 (N_10541,N_7829,N_7027);
nor U10542 (N_10542,N_6934,N_7254);
and U10543 (N_10543,N_7313,N_7939);
and U10544 (N_10544,N_5852,N_7737);
xnor U10545 (N_10545,N_9401,N_6282);
or U10546 (N_10546,N_8312,N_7625);
xor U10547 (N_10547,N_7111,N_7624);
or U10548 (N_10548,N_9317,N_7765);
or U10549 (N_10549,N_7248,N_9857);
nand U10550 (N_10550,N_8001,N_6113);
or U10551 (N_10551,N_8673,N_9596);
xor U10552 (N_10552,N_9004,N_8666);
nor U10553 (N_10553,N_8057,N_5741);
or U10554 (N_10554,N_7302,N_9733);
or U10555 (N_10555,N_7723,N_8812);
or U10556 (N_10556,N_9501,N_7096);
or U10557 (N_10557,N_6828,N_6835);
or U10558 (N_10558,N_8466,N_5900);
or U10559 (N_10559,N_5355,N_5986);
nor U10560 (N_10560,N_9425,N_7551);
nor U10561 (N_10561,N_8387,N_6082);
nand U10562 (N_10562,N_5846,N_8698);
xnor U10563 (N_10563,N_5589,N_8276);
nand U10564 (N_10564,N_7471,N_7764);
and U10565 (N_10565,N_8916,N_5498);
and U10566 (N_10566,N_8254,N_8714);
nand U10567 (N_10567,N_7585,N_5603);
nor U10568 (N_10568,N_6421,N_7562);
nor U10569 (N_10569,N_8159,N_8063);
nand U10570 (N_10570,N_6651,N_5195);
or U10571 (N_10571,N_7201,N_8437);
nand U10572 (N_10572,N_5219,N_7138);
xnor U10573 (N_10573,N_8686,N_8635);
xnor U10574 (N_10574,N_8846,N_5519);
nor U10575 (N_10575,N_6775,N_9290);
nor U10576 (N_10576,N_6628,N_5394);
nor U10577 (N_10577,N_5878,N_9179);
and U10578 (N_10578,N_9421,N_5673);
nand U10579 (N_10579,N_6294,N_9029);
xnor U10580 (N_10580,N_9432,N_6970);
nand U10581 (N_10581,N_5887,N_9438);
nor U10582 (N_10582,N_5406,N_5995);
or U10583 (N_10583,N_7541,N_9165);
or U10584 (N_10584,N_9281,N_7014);
nor U10585 (N_10585,N_9463,N_9978);
nor U10586 (N_10586,N_8984,N_9248);
and U10587 (N_10587,N_9782,N_8542);
nor U10588 (N_10588,N_7059,N_5716);
or U10589 (N_10589,N_9564,N_9853);
xnor U10590 (N_10590,N_7385,N_7064);
nor U10591 (N_10591,N_7241,N_8015);
and U10592 (N_10592,N_6187,N_7390);
or U10593 (N_10593,N_7871,N_8162);
xor U10594 (N_10594,N_7913,N_7403);
xnor U10595 (N_10595,N_8397,N_5275);
nor U10596 (N_10596,N_5330,N_6979);
nand U10597 (N_10597,N_7172,N_5281);
xnor U10598 (N_10598,N_8626,N_9822);
and U10599 (N_10599,N_8129,N_8569);
or U10600 (N_10600,N_7572,N_9082);
nand U10601 (N_10601,N_8286,N_9626);
or U10602 (N_10602,N_7847,N_7414);
or U10603 (N_10603,N_6003,N_7708);
and U10604 (N_10604,N_7943,N_5503);
and U10605 (N_10605,N_5539,N_5613);
xor U10606 (N_10606,N_6937,N_7144);
nor U10607 (N_10607,N_7271,N_9791);
nor U10608 (N_10608,N_7045,N_5334);
nand U10609 (N_10609,N_8563,N_6489);
xor U10610 (N_10610,N_8026,N_7431);
or U10611 (N_10611,N_7763,N_5882);
nor U10612 (N_10612,N_5215,N_7469);
nor U10613 (N_10613,N_5899,N_6194);
xnor U10614 (N_10614,N_7928,N_9696);
or U10615 (N_10615,N_7730,N_7324);
xnor U10616 (N_10616,N_6723,N_7987);
or U10617 (N_10617,N_9625,N_8163);
and U10618 (N_10618,N_5744,N_5835);
xor U10619 (N_10619,N_6703,N_8854);
or U10620 (N_10620,N_9289,N_9838);
or U10621 (N_10621,N_9255,N_6245);
or U10622 (N_10622,N_8247,N_5571);
and U10623 (N_10623,N_9609,N_9862);
or U10624 (N_10624,N_5806,N_8108);
nand U10625 (N_10625,N_9023,N_7748);
nand U10626 (N_10626,N_6846,N_8775);
nand U10627 (N_10627,N_5624,N_5141);
nor U10628 (N_10628,N_9967,N_8734);
nand U10629 (N_10629,N_7311,N_7353);
or U10630 (N_10630,N_6908,N_6836);
xnor U10631 (N_10631,N_9341,N_6344);
xor U10632 (N_10632,N_5068,N_6744);
and U10633 (N_10633,N_9792,N_8224);
and U10634 (N_10634,N_7591,N_6000);
xor U10635 (N_10635,N_6230,N_5578);
or U10636 (N_10636,N_5793,N_7521);
or U10637 (N_10637,N_8098,N_5041);
or U10638 (N_10638,N_5911,N_5136);
xor U10639 (N_10639,N_5789,N_6057);
and U10640 (N_10640,N_8575,N_7296);
or U10641 (N_10641,N_9628,N_7464);
nand U10642 (N_10642,N_7155,N_8265);
xnor U10643 (N_10643,N_7229,N_9575);
nand U10644 (N_10644,N_8283,N_6706);
xnor U10645 (N_10645,N_9041,N_6508);
and U10646 (N_10646,N_5964,N_9974);
or U10647 (N_10647,N_6996,N_8917);
nand U10648 (N_10648,N_7424,N_9908);
xor U10649 (N_10649,N_8439,N_8619);
or U10650 (N_10650,N_9518,N_8891);
xnor U10651 (N_10651,N_5383,N_7575);
or U10652 (N_10652,N_9937,N_5025);
nor U10653 (N_10653,N_9002,N_6547);
or U10654 (N_10654,N_8663,N_5689);
xor U10655 (N_10655,N_7740,N_7588);
xor U10656 (N_10656,N_7212,N_8399);
nor U10657 (N_10657,N_8527,N_7336);
or U10658 (N_10658,N_5329,N_5269);
nand U10659 (N_10659,N_5490,N_9741);
xor U10660 (N_10660,N_5077,N_6608);
nand U10661 (N_10661,N_7923,N_5199);
nor U10662 (N_10662,N_7510,N_7107);
and U10663 (N_10663,N_7485,N_7505);
nand U10664 (N_10664,N_7793,N_5661);
and U10665 (N_10665,N_7222,N_5517);
or U10666 (N_10666,N_6267,N_5783);
and U10667 (N_10667,N_5095,N_7965);
xor U10668 (N_10668,N_5024,N_9525);
xnor U10669 (N_10669,N_9257,N_7197);
xor U10670 (N_10670,N_7619,N_6252);
xor U10671 (N_10671,N_5781,N_7031);
or U10672 (N_10672,N_5617,N_5976);
and U10673 (N_10673,N_7583,N_5384);
xor U10674 (N_10674,N_7717,N_8978);
nor U10675 (N_10675,N_5615,N_6948);
nor U10676 (N_10676,N_8409,N_9291);
or U10677 (N_10677,N_7430,N_5618);
nor U10678 (N_10678,N_6324,N_7200);
or U10679 (N_10679,N_5270,N_9433);
or U10680 (N_10680,N_6281,N_5605);
xnor U10681 (N_10681,N_9683,N_8800);
or U10682 (N_10682,N_9754,N_6333);
or U10683 (N_10683,N_7185,N_5763);
or U10684 (N_10684,N_5476,N_8172);
nor U10685 (N_10685,N_8644,N_7227);
nor U10686 (N_10686,N_9211,N_5414);
xnor U10687 (N_10687,N_9689,N_6402);
or U10688 (N_10688,N_9849,N_9343);
nor U10689 (N_10689,N_9392,N_5359);
xnor U10690 (N_10690,N_5849,N_7507);
xor U10691 (N_10691,N_7736,N_6707);
and U10692 (N_10692,N_9461,N_7883);
nand U10693 (N_10693,N_7564,N_8861);
and U10694 (N_10694,N_7129,N_8322);
nor U10695 (N_10695,N_7843,N_7917);
nand U10696 (N_10696,N_9831,N_8514);
or U10697 (N_10697,N_8738,N_6218);
or U10698 (N_10698,N_6568,N_6550);
nor U10699 (N_10699,N_7487,N_8218);
nand U10700 (N_10700,N_7983,N_5082);
and U10701 (N_10701,N_9409,N_5501);
nand U10702 (N_10702,N_7189,N_9677);
and U10703 (N_10703,N_8597,N_9435);
and U10704 (N_10704,N_8363,N_6525);
or U10705 (N_10705,N_7224,N_5488);
nand U10706 (N_10706,N_5430,N_7406);
or U10707 (N_10707,N_8078,N_5906);
nand U10708 (N_10708,N_7670,N_9108);
xnor U10709 (N_10709,N_8044,N_7759);
xnor U10710 (N_10710,N_5641,N_8467);
nand U10711 (N_10711,N_8772,N_5097);
or U10712 (N_10712,N_7533,N_9390);
or U10713 (N_10713,N_5185,N_6702);
xor U10714 (N_10714,N_8391,N_7879);
or U10715 (N_10715,N_9710,N_7898);
and U10716 (N_10716,N_5966,N_5471);
xor U10717 (N_10717,N_8199,N_7240);
nor U10718 (N_10718,N_6408,N_8705);
or U10719 (N_10719,N_6924,N_8433);
nor U10720 (N_10720,N_9391,N_6626);
or U10721 (N_10721,N_5572,N_8989);
and U10722 (N_10722,N_7938,N_8340);
and U10723 (N_10723,N_5905,N_7440);
or U10724 (N_10724,N_5304,N_9430);
nor U10725 (N_10725,N_7809,N_9167);
and U10726 (N_10726,N_7141,N_9312);
nand U10727 (N_10727,N_5765,N_6140);
or U10728 (N_10728,N_7595,N_5855);
or U10729 (N_10729,N_5508,N_9168);
and U10730 (N_10730,N_7109,N_6273);
nor U10731 (N_10731,N_9789,N_8877);
or U10732 (N_10732,N_5941,N_8375);
nor U10733 (N_10733,N_8905,N_6018);
xor U10734 (N_10734,N_8970,N_9295);
and U10735 (N_10735,N_5524,N_5426);
nand U10736 (N_10736,N_6887,N_6207);
nand U10737 (N_10737,N_6204,N_5392);
or U10738 (N_10738,N_6953,N_6303);
nand U10739 (N_10739,N_7631,N_5902);
nor U10740 (N_10740,N_7559,N_5278);
or U10741 (N_10741,N_6173,N_8930);
or U10742 (N_10742,N_5770,N_6742);
nand U10743 (N_10743,N_7785,N_7539);
nor U10744 (N_10744,N_6094,N_7316);
nor U10745 (N_10745,N_8494,N_7364);
or U10746 (N_10746,N_7940,N_6632);
or U10747 (N_10747,N_5474,N_8298);
xor U10748 (N_10748,N_9337,N_7992);
nand U10749 (N_10749,N_9338,N_6322);
and U10750 (N_10750,N_6912,N_8348);
xor U10751 (N_10751,N_9172,N_5408);
xor U10752 (N_10752,N_5538,N_5268);
or U10753 (N_10753,N_5273,N_9468);
nor U10754 (N_10754,N_9157,N_6514);
nand U10755 (N_10755,N_7601,N_8895);
xnor U10756 (N_10756,N_6398,N_7993);
or U10757 (N_10757,N_8408,N_5644);
xnor U10758 (N_10758,N_6946,N_6975);
and U10759 (N_10759,N_8966,N_9404);
nand U10760 (N_10760,N_7009,N_7713);
nor U10761 (N_10761,N_8789,N_5743);
nand U10762 (N_10762,N_9956,N_6998);
or U10763 (N_10763,N_8220,N_6122);
xnor U10764 (N_10764,N_9212,N_7634);
nand U10765 (N_10765,N_6604,N_5305);
or U10766 (N_10766,N_7854,N_8100);
xor U10767 (N_10767,N_9656,N_6808);
nor U10768 (N_10768,N_6119,N_6961);
nand U10769 (N_10769,N_7453,N_8878);
or U10770 (N_10770,N_9698,N_6433);
nand U10771 (N_10771,N_8398,N_5121);
xnor U10772 (N_10772,N_5301,N_5153);
nand U10773 (N_10773,N_6977,N_8120);
nand U10774 (N_10774,N_8083,N_9402);
nand U10775 (N_10775,N_9653,N_8554);
nor U10776 (N_10776,N_9202,N_8311);
nand U10777 (N_10777,N_5004,N_5845);
nand U10778 (N_10778,N_9314,N_6350);
nor U10779 (N_10779,N_6260,N_7482);
and U10780 (N_10780,N_9724,N_9359);
nand U10781 (N_10781,N_8922,N_5549);
or U10782 (N_10782,N_8255,N_9075);
nor U10783 (N_10783,N_7114,N_6665);
or U10784 (N_10784,N_6693,N_8354);
nand U10785 (N_10785,N_7153,N_7528);
nand U10786 (N_10786,N_6865,N_5386);
nand U10787 (N_10787,N_9763,N_7477);
or U10788 (N_10788,N_9283,N_7999);
or U10789 (N_10789,N_8279,N_5482);
and U10790 (N_10790,N_9990,N_5494);
and U10791 (N_10791,N_6205,N_8713);
or U10792 (N_10792,N_9006,N_6656);
nor U10793 (N_10793,N_7380,N_8515);
and U10794 (N_10794,N_6930,N_8632);
or U10795 (N_10795,N_8782,N_7579);
nand U10796 (N_10796,N_8200,N_5537);
xor U10797 (N_10797,N_6896,N_7273);
xor U10798 (N_10798,N_8358,N_7538);
nor U10799 (N_10799,N_9965,N_5130);
xnor U10800 (N_10800,N_9121,N_6939);
nand U10801 (N_10801,N_7530,N_6901);
nand U10802 (N_10802,N_6359,N_6688);
and U10803 (N_10803,N_7423,N_7796);
or U10804 (N_10804,N_6128,N_8359);
nand U10805 (N_10805,N_8565,N_6869);
and U10806 (N_10806,N_6866,N_7557);
and U10807 (N_10807,N_8007,N_6159);
xor U10808 (N_10808,N_7210,N_8022);
nor U10809 (N_10809,N_8149,N_6883);
xor U10810 (N_10810,N_8602,N_9099);
nor U10811 (N_10811,N_5481,N_8583);
xnor U10812 (N_10812,N_9405,N_5201);
or U10813 (N_10813,N_7743,N_6440);
or U10814 (N_10814,N_9313,N_6733);
xor U10815 (N_10815,N_7868,N_9484);
xnor U10816 (N_10816,N_6246,N_9846);
xnor U10817 (N_10817,N_6922,N_6890);
and U10818 (N_10818,N_5422,N_7062);
nor U10819 (N_10819,N_5552,N_6030);
xor U10820 (N_10820,N_6736,N_6615);
nand U10821 (N_10821,N_5836,N_9123);
and U10822 (N_10822,N_8579,N_8771);
nand U10823 (N_10823,N_9900,N_5295);
nand U10824 (N_10824,N_8744,N_8360);
or U10825 (N_10825,N_8272,N_7637);
nand U10826 (N_10826,N_8192,N_8975);
and U10827 (N_10827,N_5339,N_6209);
nand U10828 (N_10828,N_9114,N_8929);
nor U10829 (N_10829,N_9507,N_9304);
xnor U10830 (N_10830,N_8592,N_5335);
nor U10831 (N_10831,N_6894,N_6795);
or U10832 (N_10832,N_5228,N_6582);
or U10833 (N_10833,N_8683,N_8884);
xor U10834 (N_10834,N_5667,N_6710);
and U10835 (N_10835,N_6672,N_5428);
nand U10836 (N_10836,N_7077,N_6602);
xnor U10837 (N_10837,N_7623,N_8114);
and U10838 (N_10838,N_6752,N_5969);
xor U10839 (N_10839,N_5713,N_5581);
or U10840 (N_10840,N_9487,N_9730);
xnor U10841 (N_10841,N_6650,N_8071);
and U10842 (N_10842,N_6572,N_7166);
nor U10843 (N_10843,N_6180,N_7199);
nand U10844 (N_10844,N_8638,N_7232);
xnor U10845 (N_10845,N_5989,N_9189);
or U10846 (N_10846,N_9829,N_6346);
nand U10847 (N_10847,N_7881,N_5045);
and U10848 (N_10848,N_6351,N_9801);
nand U10849 (N_10849,N_9250,N_9416);
nor U10850 (N_10850,N_9406,N_6876);
nand U10851 (N_10851,N_7859,N_9113);
and U10852 (N_10852,N_7703,N_8418);
nor U10853 (N_10853,N_6627,N_8578);
xor U10854 (N_10854,N_7692,N_7370);
nor U10855 (N_10855,N_6066,N_5319);
nor U10856 (N_10856,N_8127,N_8209);
nor U10857 (N_10857,N_8507,N_7483);
xnor U10858 (N_10858,N_5054,N_5286);
xor U10859 (N_10859,N_5311,N_7484);
xor U10860 (N_10860,N_7261,N_8229);
xor U10861 (N_10861,N_5545,N_5308);
and U10862 (N_10862,N_6585,N_8817);
nand U10863 (N_10863,N_5364,N_9495);
or U10864 (N_10864,N_8389,N_6022);
xor U10865 (N_10865,N_6949,N_8313);
or U10866 (N_10866,N_6236,N_7839);
nand U10867 (N_10867,N_5733,N_8756);
nand U10868 (N_10868,N_8278,N_8701);
nor U10869 (N_10869,N_6247,N_5472);
nand U10870 (N_10870,N_8764,N_6407);
nor U10871 (N_10871,N_6610,N_5208);
nand U10872 (N_10872,N_7659,N_9514);
nand U10873 (N_10873,N_5170,N_7330);
or U10874 (N_10874,N_8309,N_8548);
nand U10875 (N_10875,N_8676,N_6291);
nor U10876 (N_10876,N_7069,N_7006);
nor U10877 (N_10877,N_5671,N_7724);
nand U10878 (N_10878,N_9878,N_6556);
nand U10879 (N_10879,N_5965,N_8513);
and U10880 (N_10880,N_9509,N_5352);
xnor U10881 (N_10881,N_6950,N_9429);
or U10882 (N_10882,N_7277,N_6509);
and U10883 (N_10883,N_7351,N_8572);
nor U10884 (N_10884,N_8910,N_9125);
or U10885 (N_10885,N_5863,N_5772);
nor U10886 (N_10886,N_5840,N_6609);
xor U10887 (N_10887,N_7156,N_8539);
xor U10888 (N_10888,N_7666,N_8222);
xnor U10889 (N_10889,N_5659,N_7080);
or U10890 (N_10890,N_6296,N_7280);
or U10891 (N_10891,N_5345,N_6465);
and U10892 (N_10892,N_9037,N_6624);
nand U10893 (N_10893,N_7279,N_8067);
nor U10894 (N_10894,N_7473,N_7237);
nor U10895 (N_10895,N_5192,N_7790);
or U10896 (N_10896,N_6340,N_5732);
and U10897 (N_10897,N_6813,N_8733);
or U10898 (N_10898,N_8290,N_8141);
nor U10899 (N_10899,N_7954,N_5547);
nand U10900 (N_10900,N_5411,N_6714);
or U10901 (N_10901,N_7603,N_8680);
and U10902 (N_10902,N_8788,N_5931);
nand U10903 (N_10903,N_6311,N_6316);
nor U10904 (N_10904,N_9100,N_8004);
or U10905 (N_10905,N_8749,N_6444);
xnor U10906 (N_10906,N_6474,N_5526);
nor U10907 (N_10907,N_6952,N_7102);
nand U10908 (N_10908,N_7067,N_7783);
or U10909 (N_10909,N_5947,N_5651);
or U10910 (N_10910,N_8296,N_7806);
and U10911 (N_10911,N_7534,N_5514);
nor U10912 (N_10912,N_5847,N_6794);
nand U10913 (N_10913,N_5939,N_8535);
xor U10914 (N_10914,N_6052,N_9680);
or U10915 (N_10915,N_7893,N_9042);
nand U10916 (N_10916,N_6110,N_6577);
and U10917 (N_10917,N_8055,N_8987);
xnor U10918 (N_10918,N_6317,N_9010);
nor U10919 (N_10919,N_6472,N_5057);
nor U10920 (N_10920,N_8532,N_9673);
nor U10921 (N_10921,N_6048,N_8871);
or U10922 (N_10922,N_6798,N_6720);
and U10923 (N_10923,N_5803,N_8049);
or U10924 (N_10924,N_5857,N_9494);
or U10925 (N_10925,N_9467,N_9664);
xor U10926 (N_10926,N_7776,N_9951);
nor U10927 (N_10927,N_8300,N_7777);
nand U10928 (N_10928,N_7668,N_5642);
nor U10929 (N_10929,N_8147,N_9258);
nand U10930 (N_10930,N_8225,N_9320);
xnor U10931 (N_10931,N_7225,N_8648);
nor U10932 (N_10932,N_8661,N_8671);
or U10933 (N_10933,N_8068,N_6144);
or U10934 (N_10934,N_8077,N_8882);
nor U10935 (N_10935,N_7374,N_5949);
nor U10936 (N_10936,N_7432,N_9708);
nand U10937 (N_10937,N_7288,N_9058);
nand U10938 (N_10938,N_7501,N_9112);
nand U10939 (N_10939,N_7711,N_9783);
or U10940 (N_10940,N_9773,N_8444);
and U10941 (N_10941,N_9230,N_6690);
and U10942 (N_10942,N_8598,N_7461);
or U10943 (N_10943,N_7826,N_8215);
nand U10944 (N_10944,N_8783,N_8475);
nor U10945 (N_10945,N_5950,N_7148);
or U10946 (N_10946,N_8595,N_9536);
and U10947 (N_10947,N_6974,N_6459);
and U10948 (N_10948,N_8803,N_5570);
or U10949 (N_10949,N_7550,N_7084);
nand U10950 (N_10950,N_6655,N_5860);
nor U10951 (N_10951,N_9448,N_8931);
or U10952 (N_10952,N_7286,N_5148);
nand U10953 (N_10953,N_6239,N_8587);
or U10954 (N_10954,N_9610,N_6881);
and U10955 (N_10955,N_6911,N_7558);
or U10956 (N_10956,N_7379,N_7862);
and U10957 (N_10957,N_6272,N_8005);
nor U10958 (N_10958,N_5101,N_7250);
nand U10959 (N_10959,N_6524,N_5108);
nand U10960 (N_10960,N_9348,N_9327);
xor U10961 (N_10961,N_6774,N_5294);
xnor U10962 (N_10962,N_8441,N_7673);
nor U10963 (N_10963,N_9915,N_6761);
nand U10964 (N_10964,N_7117,N_6959);
xor U10965 (N_10965,N_6137,N_6684);
nor U10966 (N_10966,N_5800,N_8499);
nor U10967 (N_10967,N_9940,N_6642);
nor U10968 (N_10968,N_6093,N_9903);
nor U10969 (N_10969,N_9758,N_7088);
and U10970 (N_10970,N_9190,N_7658);
and U10971 (N_10971,N_8540,N_5822);
nand U10972 (N_10972,N_9812,N_5099);
and U10973 (N_10973,N_5987,N_5730);
xnor U10974 (N_10974,N_7167,N_6539);
xor U10975 (N_10975,N_5738,N_6071);
and U10976 (N_10976,N_7827,N_6134);
nor U10977 (N_10977,N_5532,N_7177);
xor U10978 (N_10978,N_5728,N_7566);
xor U10979 (N_10979,N_7833,N_7065);
and U10980 (N_10980,N_9643,N_7052);
or U10981 (N_10981,N_9418,N_9153);
xor U10982 (N_10982,N_8787,N_7795);
nor U10983 (N_10983,N_7381,N_7599);
nand U10984 (N_10984,N_6386,N_6854);
nand U10985 (N_10985,N_5255,N_8761);
or U10986 (N_10986,N_7602,N_9098);
and U10987 (N_10987,N_7661,N_6815);
and U10988 (N_10988,N_7563,N_6681);
nand U10989 (N_10989,N_6653,N_7676);
and U10990 (N_10990,N_9859,N_7613);
nand U10991 (N_10991,N_9217,N_5522);
or U10992 (N_10992,N_7945,N_7680);
and U10993 (N_10993,N_8060,N_7707);
or U10994 (N_10994,N_6005,N_8195);
and U10995 (N_10995,N_9769,N_9860);
nand U10996 (N_10996,N_5702,N_8947);
or U10997 (N_10997,N_5066,N_9561);
and U10998 (N_10998,N_7758,N_5048);
nand U10999 (N_10999,N_8954,N_9941);
nand U11000 (N_11000,N_6649,N_6573);
nand U11001 (N_11001,N_7333,N_5760);
and U11002 (N_11002,N_6663,N_5751);
or U11003 (N_11003,N_6634,N_5337);
xor U11004 (N_11004,N_5943,N_6658);
nor U11005 (N_11005,N_8662,N_8134);
nor U11006 (N_11006,N_8521,N_9398);
xnor U11007 (N_11007,N_6713,N_9617);
nand U11008 (N_11008,N_7028,N_9992);
nor U11009 (N_11009,N_5234,N_9363);
xor U11010 (N_11010,N_7314,N_5226);
and U11011 (N_11011,N_7393,N_5230);
nor U11012 (N_11012,N_9309,N_9506);
or U11013 (N_11013,N_6477,N_8118);
xor U11014 (N_11014,N_9001,N_5302);
nand U11015 (N_11015,N_9239,N_9953);
and U11016 (N_11016,N_8523,N_6011);
or U11017 (N_11017,N_6778,N_8076);
nand U11018 (N_11018,N_7319,N_8727);
or U11019 (N_11019,N_8797,N_8872);
nand U11020 (N_11020,N_5649,N_5904);
or U11021 (N_11021,N_7049,N_8769);
xnor U11022 (N_11022,N_8906,N_8684);
xor U11023 (N_11023,N_6645,N_7492);
xor U11024 (N_11024,N_6543,N_8834);
nand U11025 (N_11025,N_5421,N_7520);
nand U11026 (N_11026,N_5028,N_5523);
xnor U11027 (N_11027,N_9442,N_9476);
nor U11028 (N_11028,N_7722,N_8694);
nor U11029 (N_11029,N_7413,N_7397);
and U11030 (N_11030,N_7388,N_7466);
and U11031 (N_11031,N_8447,N_8748);
or U11032 (N_11032,N_6941,N_9802);
nor U11033 (N_11033,N_5229,N_5898);
nand U11034 (N_11034,N_6739,N_6921);
or U11035 (N_11035,N_5759,N_6232);
xor U11036 (N_11036,N_9865,N_9611);
and U11037 (N_11037,N_6133,N_7773);
nor U11038 (N_11038,N_8659,N_6919);
xor U11039 (N_11039,N_9360,N_9957);
and U11040 (N_11040,N_6559,N_9918);
nor U11041 (N_11041,N_8432,N_5920);
and U11042 (N_11042,N_7244,N_8244);
and U11043 (N_11043,N_8370,N_9380);
nor U11044 (N_11044,N_9045,N_7029);
nand U11045 (N_11045,N_6178,N_5405);
and U11046 (N_11046,N_8477,N_6725);
or U11047 (N_11047,N_6253,N_6821);
nand U11048 (N_11048,N_8161,N_9775);
xor U11049 (N_11049,N_9422,N_8711);
nor U11050 (N_11050,N_7633,N_6838);
or U11051 (N_11051,N_6918,N_8235);
or U11052 (N_11052,N_6436,N_6177);
nor U11053 (N_11053,N_7988,N_7850);
nor U11054 (N_11054,N_7341,N_7946);
nand U11055 (N_11055,N_7667,N_7974);
and U11056 (N_11056,N_8757,N_8481);
xor U11057 (N_11057,N_9551,N_6152);
xor U11058 (N_11058,N_7548,N_9375);
and U11059 (N_11059,N_7844,N_7115);
xor U11060 (N_11060,N_7927,N_8066);
xnor U11061 (N_11061,N_9218,N_5072);
nor U11062 (N_11062,N_9922,N_6349);
nor U11063 (N_11063,N_8099,N_8849);
xnor U11064 (N_11064,N_9723,N_7699);
nor U11065 (N_11065,N_7106,N_8295);
or U11066 (N_11066,N_5762,N_9637);
nor U11067 (N_11067,N_7894,N_6534);
and U11068 (N_11068,N_5623,N_8179);
xor U11069 (N_11069,N_7536,N_7638);
nand U11070 (N_11070,N_8355,N_8674);
xor U11071 (N_11071,N_9159,N_8990);
or U11072 (N_11072,N_7960,N_5614);
xnor U11073 (N_11073,N_9106,N_8445);
nand U11074 (N_11074,N_8237,N_8911);
or U11075 (N_11075,N_6269,N_8487);
and U11076 (N_11076,N_7675,N_7499);
and U11077 (N_11077,N_8732,N_7276);
and U11078 (N_11078,N_7989,N_8133);
and U11079 (N_11079,N_5008,N_9345);
nand U11080 (N_11080,N_5390,N_7450);
xor U11081 (N_11081,N_7972,N_7350);
nand U11082 (N_11082,N_9818,N_5158);
and U11083 (N_11083,N_7787,N_7630);
or U11084 (N_11084,N_9369,N_8933);
nand U11085 (N_11085,N_5232,N_5452);
or U11086 (N_11086,N_6824,N_7391);
or U11087 (N_11087,N_5222,N_8707);
or U11088 (N_11088,N_6603,N_6445);
nor U11089 (N_11089,N_7243,N_8755);
xnor U11090 (N_11090,N_7134,N_8640);
and U11091 (N_11091,N_9084,N_5217);
xor U11092 (N_11092,N_5157,N_5622);
nor U11093 (N_11093,N_6980,N_8132);
or U11094 (N_11094,N_9833,N_9080);
nor U11095 (N_11095,N_5448,N_8996);
or U11096 (N_11096,N_9695,N_9062);
nand U11097 (N_11097,N_7782,N_9517);
and U11098 (N_11098,N_5521,N_9757);
nor U11099 (N_11099,N_6114,N_8991);
nor U11100 (N_11100,N_8588,N_6871);
nor U11101 (N_11101,N_7590,N_5942);
and U11102 (N_11102,N_8024,N_9140);
nand U11103 (N_11103,N_7798,N_5718);
or U11104 (N_11104,N_7357,N_9557);
xor U11105 (N_11105,N_8645,N_7170);
nand U11106 (N_11106,N_9640,N_8941);
nor U11107 (N_11107,N_8320,N_5133);
and U11108 (N_11108,N_5260,N_5182);
xor U11109 (N_11109,N_9451,N_6310);
or U11110 (N_11110,N_8695,N_8249);
xnor U11111 (N_11111,N_7435,N_9522);
nand U11112 (N_11112,N_6989,N_9183);
and U11113 (N_11113,N_8558,N_6754);
nand U11114 (N_11114,N_6261,N_9616);
or U11115 (N_11115,N_9538,N_8743);
nand U11116 (N_11116,N_5691,N_6120);
nor U11117 (N_11117,N_6958,N_5690);
or U11118 (N_11118,N_5172,N_9018);
and U11119 (N_11119,N_7293,N_5884);
nor U11120 (N_11120,N_6829,N_7788);
or U11121 (N_11121,N_5784,N_5401);
xor U11122 (N_11122,N_5012,N_7387);
and U11123 (N_11123,N_9083,N_5285);
or U11124 (N_11124,N_5551,N_6337);
nand U11125 (N_11125,N_9021,N_7900);
xnor U11126 (N_11126,N_7073,N_5871);
nand U11127 (N_11127,N_8794,N_9836);
or U11128 (N_11128,N_9636,N_5792);
nand U11129 (N_11129,N_9959,N_5189);
or U11130 (N_11130,N_7100,N_8969);
nor U11131 (N_11131,N_5123,N_9563);
nor U11132 (N_11132,N_9545,N_8221);
xnor U11133 (N_11133,N_5874,N_7967);
and U11134 (N_11134,N_6233,N_9489);
xnor U11135 (N_11135,N_7295,N_9571);
nor U11136 (N_11136,N_9081,N_5496);
nand U11137 (N_11137,N_7181,N_9009);
nor U11138 (N_11138,N_9991,N_6933);
xor U11139 (N_11139,N_8781,N_6734);
and U11140 (N_11140,N_9934,N_5436);
and U11141 (N_11141,N_6517,N_8188);
nand U11142 (N_11142,N_5851,N_6687);
nand U11143 (N_11143,N_5645,N_7516);
nand U11144 (N_11144,N_5137,N_8517);
nor U11145 (N_11145,N_5991,N_6372);
nor U11146 (N_11146,N_7944,N_7145);
nand U11147 (N_11147,N_7082,N_8264);
xnor U11148 (N_11148,N_6060,N_6506);
or U11149 (N_11149,N_7063,N_8018);
nand U11150 (N_11150,N_6685,N_6142);
nand U11151 (N_11151,N_5555,N_5146);
nand U11152 (N_11152,N_9570,N_7855);
or U11153 (N_11153,N_7498,N_6978);
and U11154 (N_11154,N_5630,N_5940);
nor U11155 (N_11155,N_8506,N_7690);
xor U11156 (N_11156,N_5788,N_9705);
xor U11157 (N_11157,N_7417,N_8164);
or U11158 (N_11158,N_8033,N_8586);
nor U11159 (N_11159,N_7694,N_7253);
nand U11160 (N_11160,N_7984,N_7942);
nor U11161 (N_11161,N_7704,N_5073);
or U11162 (N_11162,N_7218,N_8886);
xnor U11163 (N_11163,N_7567,N_5439);
xnor U11164 (N_11164,N_7950,N_7383);
nor U11165 (N_11165,N_9715,N_6387);
nand U11166 (N_11166,N_9534,N_8365);
or U11167 (N_11167,N_5719,N_7386);
or U11168 (N_11168,N_9742,N_6852);
and U11169 (N_11169,N_7433,N_5866);
nor U11170 (N_11170,N_5694,N_5447);
or U11171 (N_11171,N_7964,N_5100);
and U11172 (N_11172,N_7123,N_7542);
and U11173 (N_11173,N_7869,N_6314);
and U11174 (N_11174,N_5712,N_9966);
or U11175 (N_11175,N_6425,N_7878);
xnor U11176 (N_11176,N_9024,N_5160);
and U11177 (N_11177,N_7448,N_8434);
and U11178 (N_11178,N_5291,N_9585);
xor U11179 (N_11179,N_7426,N_9780);
xor U11180 (N_11180,N_9532,N_9355);
xor U11181 (N_11181,N_9911,N_5111);
and U11182 (N_11182,N_9199,N_6923);
and U11183 (N_11183,N_9999,N_7576);
and U11184 (N_11184,N_8112,N_8830);
nor U11185 (N_11185,N_8266,N_5828);
nor U11186 (N_11186,N_9094,N_5795);
and U11187 (N_11187,N_9655,N_6756);
xor U11188 (N_11188,N_7835,N_8028);
nand U11189 (N_11189,N_5764,N_9607);
and U11190 (N_11190,N_5883,N_9948);
and U11191 (N_11191,N_6523,N_8357);
nand U11192 (N_11192,N_5346,N_7310);
and U11193 (N_11193,N_5258,N_6670);
or U11194 (N_11194,N_5735,N_6242);
nor U11195 (N_11195,N_9235,N_5796);
nand U11196 (N_11196,N_5797,N_5459);
nor U11197 (N_11197,N_5382,N_8039);
xor U11198 (N_11198,N_8484,N_8960);
nand U11199 (N_11199,N_8613,N_9480);
nor U11200 (N_11200,N_8725,N_7754);
nand U11201 (N_11201,N_7122,N_7822);
nor U11202 (N_11202,N_5665,N_7180);
xor U11203 (N_11203,N_9117,N_7523);
xor U11204 (N_11204,N_8526,N_5240);
and U11205 (N_11205,N_8702,N_6369);
and U11206 (N_11206,N_7503,N_7475);
nand U11207 (N_11207,N_9895,N_8786);
nand U11208 (N_11208,N_8652,N_6087);
or U11209 (N_11209,N_9434,N_7750);
nor U11210 (N_11210,N_5917,N_5634);
and U11211 (N_11211,N_6357,N_5561);
and U11212 (N_11212,N_8119,N_5378);
or U11213 (N_11213,N_9477,N_7757);
or U11214 (N_11214,N_6729,N_9347);
nor U11215 (N_11215,N_9294,N_9912);
xnor U11216 (N_11216,N_7838,N_9709);
and U11217 (N_11217,N_9252,N_7976);
nand U11218 (N_11218,N_5283,N_9043);
or U11219 (N_11219,N_8349,N_8326);
and U11220 (N_11220,N_6738,N_6611);
nand U11221 (N_11221,N_9586,N_6176);
nor U11222 (N_11222,N_5191,N_5358);
and U11223 (N_11223,N_8413,N_5098);
nand U11224 (N_11224,N_9774,N_8826);
nand U11225 (N_11225,N_7206,N_9798);
nand U11226 (N_11226,N_5047,N_8719);
and U11227 (N_11227,N_7606,N_5510);
or U11228 (N_11228,N_5174,N_7365);
xor U11229 (N_11229,N_7021,N_8431);
or U11230 (N_11230,N_7996,N_6762);
and U11231 (N_11231,N_9588,N_8268);
and U11232 (N_11232,N_9498,N_8116);
or U11233 (N_11233,N_8023,N_7445);
and U11234 (N_11234,N_8405,N_6819);
or U11235 (N_11235,N_9841,N_7415);
and U11236 (N_11236,N_7920,N_6139);
xor U11237 (N_11237,N_7647,N_5080);
xnor U11238 (N_11238,N_8518,N_8371);
nand U11239 (N_11239,N_5725,N_9266);
nand U11240 (N_11240,N_8885,N_7495);
nor U11241 (N_11241,N_7150,N_8245);
nor U11242 (N_11242,N_5650,N_9276);
and U11243 (N_11243,N_5662,N_8730);
nand U11244 (N_11244,N_5049,N_6460);
and U11245 (N_11245,N_8837,N_7193);
xnor U11246 (N_11246,N_6895,N_7184);
nand U11247 (N_11247,N_6925,N_5043);
nor U11248 (N_11248,N_9491,N_8902);
or U11249 (N_11249,N_6160,N_5970);
and U11250 (N_11250,N_8333,N_7812);
nor U11251 (N_11251,N_8537,N_8065);
or U11252 (N_11252,N_9863,N_5924);
and U11253 (N_11253,N_8243,N_5022);
xor U11254 (N_11254,N_7171,N_6399);
or U11255 (N_11255,N_6956,N_6674);
and U11256 (N_11256,N_9766,N_6973);
xor U11257 (N_11257,N_5594,N_5396);
nor U11258 (N_11258,N_6368,N_8426);
nor U11259 (N_11259,N_9566,N_5055);
xor U11260 (N_11260,N_6728,N_9905);
or U11261 (N_11261,N_6491,N_8373);
nand U11262 (N_11262,N_8294,N_6301);
and U11263 (N_11263,N_5990,N_5631);
nor U11264 (N_11264,N_6820,N_7770);
nand U11265 (N_11265,N_8382,N_6581);
nand U11266 (N_11266,N_8840,N_5636);
nand U11267 (N_11267,N_8207,N_9861);
and U11268 (N_11268,N_8643,N_5512);
xor U11269 (N_11269,N_6914,N_7745);
xnor U11270 (N_11270,N_7995,N_8040);
or U11271 (N_11271,N_5982,N_7842);
and U11272 (N_11272,N_7907,N_9323);
nor U11273 (N_11273,N_8605,N_7578);
xnor U11274 (N_11274,N_9548,N_7342);
and U11275 (N_11275,N_9269,N_7192);
nor U11276 (N_11276,N_8667,N_6913);
xnor U11277 (N_11277,N_9064,N_8547);
nor U11278 (N_11278,N_6410,N_7970);
nor U11279 (N_11279,N_8860,N_5034);
nor U11280 (N_11280,N_9573,N_5500);
nand U11281 (N_11281,N_5218,N_8508);
or U11282 (N_11282,N_9440,N_6279);
or U11283 (N_11283,N_7270,N_6182);
and U11284 (N_11284,N_9055,N_9620);
or U11285 (N_11285,N_7147,N_6198);
and U11286 (N_11286,N_8928,N_9274);
or U11287 (N_11287,N_6671,N_9424);
nor U11288 (N_11288,N_6014,N_5980);
nand U11289 (N_11289,N_6356,N_7245);
or U11290 (N_11290,N_7918,N_9520);
and U11291 (N_11291,N_7643,N_5814);
nand U11292 (N_11292,N_6432,N_5296);
or U11293 (N_11293,N_5375,N_8924);
nor U11294 (N_11294,N_8785,N_5695);
and U11295 (N_11295,N_7911,N_9787);
and U11296 (N_11296,N_6801,N_9158);
and U11297 (N_11297,N_8402,N_6116);
and U11298 (N_11298,N_6226,N_9091);
xor U11299 (N_11299,N_5914,N_5872);
or U11300 (N_11300,N_9335,N_7712);
and U11301 (N_11301,N_6597,N_8814);
xor U11302 (N_11302,N_6403,N_7143);
or U11303 (N_11303,N_6968,N_9090);
and U11304 (N_11304,N_6511,N_9560);
xnor U11305 (N_11305,N_6931,N_9954);
nand U11306 (N_11306,N_7463,N_6570);
and U11307 (N_11307,N_8806,N_7012);
xor U11308 (N_11308,N_9330,N_9260);
or U11309 (N_11309,N_9946,N_7604);
nor U11310 (N_11310,N_6927,N_8585);
nor U11311 (N_11311,N_8879,N_8767);
xnor U11312 (N_11312,N_7118,N_9000);
nand U11313 (N_11313,N_6151,N_9855);
and U11314 (N_11314,N_9277,N_8424);
and U11315 (N_11315,N_9595,N_9921);
nor U11316 (N_11316,N_7188,N_5850);
and U11317 (N_11317,N_8754,N_6589);
xnor U11318 (N_11318,N_9015,N_5327);
nand U11319 (N_11319,N_6095,N_9830);
and U11320 (N_11320,N_7256,N_7635);
nor U11321 (N_11321,N_7339,N_8672);
xor U11322 (N_11322,N_5726,N_7857);
or U11323 (N_11323,N_5431,N_5627);
nand U11324 (N_11324,N_8303,N_6437);
or U11325 (N_11325,N_8395,N_6354);
or U11326 (N_11326,N_9065,N_6647);
nand U11327 (N_11327,N_8269,N_7549);
nand U11328 (N_11328,N_6586,N_8937);
or U11329 (N_11329,N_9584,N_8845);
xor U11330 (N_11330,N_6540,N_9378);
nor U11331 (N_11331,N_5106,N_6078);
xnor U11332 (N_11332,N_9572,N_9166);
and U11333 (N_11333,N_8943,N_6418);
nand U11334 (N_11334,N_8811,N_5403);
xor U11335 (N_11335,N_6068,N_6788);
or U11336 (N_11336,N_5841,N_8203);
and U11337 (N_11337,N_9803,N_9734);
or U11338 (N_11338,N_9148,N_7044);
or U11339 (N_11339,N_5113,N_6748);
nand U11340 (N_11340,N_8135,N_9070);
nand U11341 (N_11341,N_8186,N_8617);
xor U11342 (N_11342,N_7719,N_6899);
nand U11343 (N_11343,N_7429,N_8654);
or U11344 (N_11344,N_9909,N_5246);
nand U11345 (N_11345,N_7126,N_7688);
and U11346 (N_11346,N_9170,N_5094);
xor U11347 (N_11347,N_6148,N_5739);
and U11348 (N_11348,N_5188,N_8250);
nor U11349 (N_11349,N_7772,N_5092);
or U11350 (N_11350,N_7592,N_7775);
and U11351 (N_11351,N_6404,N_5829);
nand U11352 (N_11352,N_6905,N_7034);
and U11353 (N_11353,N_8799,N_6467);
xor U11354 (N_11354,N_7008,N_7305);
nor U11355 (N_11355,N_7258,N_5777);
xnor U11356 (N_11356,N_7508,N_8168);
and U11357 (N_11357,N_9280,N_6662);
nor U11358 (N_11358,N_7075,N_6966);
nor U11359 (N_11359,N_9665,N_6131);
nor U11360 (N_11360,N_6312,N_8347);
nor U11361 (N_11361,N_5516,N_7335);
and U11362 (N_11362,N_7811,N_8599);
or U11363 (N_11363,N_5016,N_9423);
and U11364 (N_11364,N_8557,N_8407);
and U11365 (N_11365,N_5107,N_9950);
or U11366 (N_11366,N_9176,N_5666);
and U11367 (N_11367,N_5277,N_7679);
nand U11368 (N_11368,N_5429,N_8353);
or U11369 (N_11369,N_9864,N_9826);
and U11370 (N_11370,N_8138,N_7705);
xor U11371 (N_11371,N_7808,N_8951);
xnor U11372 (N_11372,N_7935,N_5254);
and U11373 (N_11373,N_8204,N_5211);
or U11374 (N_11374,N_7395,N_6132);
nand U11375 (N_11375,N_5271,N_6308);
or U11376 (N_11376,N_9821,N_5445);
or U11377 (N_11377,N_7491,N_9816);
nor U11378 (N_11378,N_7701,N_6764);
or U11379 (N_11379,N_9194,N_8574);
or U11380 (N_11380,N_6593,N_5053);
and U11381 (N_11381,N_5493,N_5579);
and U11382 (N_11382,N_5300,N_8614);
or U11383 (N_11383,N_6127,N_8000);
xnor U11384 (N_11384,N_7048,N_6036);
or U11385 (N_11385,N_9426,N_9205);
and U11386 (N_11386,N_5755,N_9871);
or U11387 (N_11387,N_6532,N_8092);
or U11388 (N_11388,N_9629,N_6395);
or U11389 (N_11389,N_8457,N_9046);
and U11390 (N_11390,N_9417,N_7820);
or U11391 (N_11391,N_5489,N_6378);
nand U11392 (N_11392,N_5530,N_5096);
xor U11393 (N_11393,N_8559,N_7130);
nand U11394 (N_11394,N_9445,N_6962);
and U11395 (N_11395,N_7640,N_8202);
and U11396 (N_11396,N_8137,N_8143);
nor U11397 (N_11397,N_6971,N_5880);
or U11398 (N_11398,N_7016,N_7582);
and U11399 (N_11399,N_9107,N_6400);
xor U11400 (N_11400,N_7735,N_7303);
and U11401 (N_11401,N_7216,N_5616);
or U11402 (N_11402,N_6915,N_5135);
nor U11403 (N_11403,N_9650,N_5685);
or U11404 (N_11404,N_5393,N_7265);
xor U11405 (N_11405,N_5657,N_6677);
nand U11406 (N_11406,N_6392,N_6429);
nor U11407 (N_11407,N_5676,N_6355);
nand U11408 (N_11408,N_6793,N_9152);
and U11409 (N_11409,N_7919,N_5798);
xnor U11410 (N_11410,N_8231,N_7678);
xnor U11411 (N_11411,N_7249,N_8670);
and U11412 (N_11412,N_5400,N_7895);
or U11413 (N_11413,N_9644,N_7178);
and U11414 (N_11414,N_8167,N_5727);
nor U11415 (N_11415,N_9365,N_6805);
nor U11416 (N_11416,N_8378,N_9431);
and U11417 (N_11417,N_6940,N_9060);
or U11418 (N_11418,N_8482,N_6673);
and U11419 (N_11419,N_6170,N_8921);
nand U11420 (N_11420,N_8314,N_5369);
nand U11421 (N_11421,N_7998,N_8825);
nand U11422 (N_11422,N_5144,N_9638);
and U11423 (N_11423,N_8469,N_5961);
nand U11424 (N_11424,N_7728,N_7991);
nor U11425 (N_11425,N_7611,N_7068);
or U11426 (N_11426,N_5197,N_7642);
or U11427 (N_11427,N_6257,N_6709);
nand U11428 (N_11428,N_7003,N_9884);
and U11429 (N_11429,N_6678,N_7405);
or U11430 (N_11430,N_7738,N_7682);
or U11431 (N_11431,N_9288,N_6588);
and U11432 (N_11432,N_8896,N_8773);
xor U11433 (N_11433,N_6254,N_9687);
and U11434 (N_11434,N_6562,N_9093);
and U11435 (N_11435,N_5169,N_5176);
nand U11436 (N_11436,N_9923,N_5065);
and U11437 (N_11437,N_9077,N_9533);
and U11438 (N_11438,N_8156,N_7419);
xnor U11439 (N_11439,N_7323,N_8853);
or U11440 (N_11440,N_7072,N_9805);
or U11441 (N_11441,N_6870,N_7526);
or U11442 (N_11442,N_5138,N_5935);
and U11443 (N_11443,N_8346,N_7609);
nand U11444 (N_11444,N_5858,N_9256);
and U11445 (N_11445,N_9492,N_7947);
xor U11446 (N_11446,N_9203,N_8327);
xnor U11447 (N_11447,N_6860,N_5790);
xor U11448 (N_11448,N_7966,N_9469);
xnor U11449 (N_11449,N_7849,N_9809);
nor U11450 (N_11450,N_7196,N_6486);
nor U11451 (N_11451,N_6013,N_6675);
and U11452 (N_11452,N_9765,N_9368);
and U11453 (N_11453,N_8536,N_5020);
xnor U11454 (N_11454,N_9939,N_7791);
or U11455 (N_11455,N_6366,N_6049);
xor U11456 (N_11456,N_7443,N_9535);
nand U11457 (N_11457,N_9598,N_7779);
nor U11458 (N_11458,N_8561,N_5591);
or U11459 (N_11459,N_8533,N_6393);
xor U11460 (N_11460,N_5492,N_5856);
or U11461 (N_11461,N_8053,N_7626);
and U11462 (N_11462,N_5161,N_6512);
nand U11463 (N_11463,N_9700,N_6103);
and U11464 (N_11464,N_9286,N_7766);
nor U11465 (N_11465,N_6365,N_8573);
xnor U11466 (N_11466,N_5198,N_5078);
nor U11467 (N_11467,N_9515,N_5639);
nor U11468 (N_11468,N_5938,N_5253);
xor U11469 (N_11469,N_5754,N_5062);
and U11470 (N_11470,N_8175,N_8241);
nand U11471 (N_11471,N_8362,N_7169);
or U11472 (N_11472,N_6304,N_8275);
xnor U11473 (N_11473,N_8110,N_5274);
xor U11474 (N_11474,N_6726,N_9707);
and U11475 (N_11475,N_6566,N_7219);
and U11476 (N_11476,N_9085,N_8197);
and U11477 (N_11477,N_8021,N_5609);
or U11478 (N_11478,N_5239,N_7337);
and U11479 (N_11479,N_9339,N_9528);
nor U11480 (N_11480,N_6305,N_5477);
xor U11481 (N_11481,N_6557,N_9155);
xor U11482 (N_11482,N_5746,N_9005);
and U11483 (N_11483,N_6235,N_8946);
nor U11484 (N_11484,N_8315,N_5975);
and U11485 (N_11485,N_8657,N_8823);
and U11486 (N_11486,N_7409,N_9475);
nand U11487 (N_11487,N_7799,N_6056);
xor U11488 (N_11488,N_7367,N_7057);
or U11489 (N_11489,N_7056,N_6439);
or U11490 (N_11490,N_9925,N_5388);
xnor U11491 (N_11491,N_6073,N_8948);
and U11492 (N_11492,N_6135,N_5952);
or U11493 (N_11493,N_7425,N_9686);
nor U11494 (N_11494,N_7677,N_8616);
or U11495 (N_11495,N_8765,N_9232);
or U11496 (N_11496,N_9735,N_9386);
nand U11497 (N_11497,N_7299,N_6032);
xnor U11498 (N_11498,N_9414,N_6981);
nor U11499 (N_11499,N_7371,N_6430);
nand U11500 (N_11500,N_6875,N_7309);
nor U11501 (N_11501,N_6831,N_5693);
nor U11502 (N_11502,N_7574,N_6561);
or U11503 (N_11503,N_8925,N_6248);
or U11504 (N_11504,N_5928,N_5145);
xor U11505 (N_11505,N_8724,N_9731);
or U11506 (N_11506,N_8682,N_6008);
nor U11507 (N_11507,N_9146,N_7628);
nand U11508 (N_11508,N_7234,N_5058);
nor U11509 (N_11509,N_5314,N_5361);
and U11510 (N_11510,N_5817,N_5162);
nor U11511 (N_11511,N_8025,N_9044);
nor U11512 (N_11512,N_8435,N_9137);
xnor U11513 (N_11513,N_5085,N_9701);
or U11514 (N_11514,N_8804,N_5647);
nor U11515 (N_11515,N_6441,N_9071);
nand U11516 (N_11516,N_9970,N_8316);
or U11517 (N_11517,N_7331,N_5680);
nand U11518 (N_11518,N_7086,N_6206);
or U11519 (N_11519,N_8881,N_7587);
xor U11520 (N_11520,N_6083,N_7382);
or U11521 (N_11521,N_8873,N_5580);
and U11522 (N_11522,N_5628,N_6993);
xor U11523 (N_11523,N_5225,N_6830);
xor U11524 (N_11524,N_6461,N_8551);
nand U11525 (N_11525,N_8277,N_6777);
nand U11526 (N_11526,N_7368,N_6600);
or U11527 (N_11527,N_8692,N_8016);
or U11528 (N_11528,N_6984,N_9238);
nand U11529 (N_11529,N_9718,N_7326);
nand U11530 (N_11530,N_9129,N_7327);
and U11531 (N_11531,N_6214,N_9329);
xor U11532 (N_11532,N_5064,N_8716);
nand U11533 (N_11533,N_9872,N_9510);
nand U11534 (N_11534,N_7504,N_9744);
and U11535 (N_11535,N_5303,N_7886);
or U11536 (N_11536,N_5602,N_9558);
xor U11537 (N_11537,N_8258,N_8717);
xor U11538 (N_11538,N_6423,N_7262);
and U11539 (N_11539,N_5926,N_7978);
xor U11540 (N_11540,N_8396,N_6492);
nand U11541 (N_11541,N_7033,N_9633);
xor U11542 (N_11542,N_6823,N_8677);
or U11543 (N_11543,N_9717,N_8476);
or U11544 (N_11544,N_6964,N_6592);
nand U11545 (N_11545,N_9237,N_9351);
or U11546 (N_11546,N_9987,N_6123);
nor U11547 (N_11547,N_8805,N_9308);
and U11548 (N_11548,N_9028,N_5999);
xnor U11549 (N_11549,N_5509,N_5289);
and U11550 (N_11550,N_6027,N_7438);
xnor U11551 (N_11551,N_9088,N_6196);
or U11552 (N_11552,N_6342,N_5577);
and U11553 (N_11553,N_9893,N_7214);
xnor U11554 (N_11554,N_9340,N_9367);
nor U11555 (N_11555,N_8791,N_7553);
and U11556 (N_11556,N_5775,N_5682);
xor U11557 (N_11557,N_8479,N_6379);
nor U11558 (N_11558,N_8865,N_9917);
nand U11559 (N_11559,N_8425,N_8287);
nor U11560 (N_11560,N_5518,N_7554);
or U11561 (N_11561,N_9526,N_9654);
and U11562 (N_11562,N_7328,N_7853);
nand U11563 (N_11563,N_5287,N_9994);
xnor U11564 (N_11564,N_7202,N_5454);
xor U11565 (N_11565,N_8808,N_9441);
or U11566 (N_11566,N_6691,N_6092);
nor U11567 (N_11567,N_7756,N_5563);
xnor U11568 (N_11568,N_5913,N_7650);
and U11569 (N_11569,N_7032,N_5559);
and U11570 (N_11570,N_7344,N_6652);
nor U11571 (N_11571,N_9924,N_5224);
nor U11572 (N_11572,N_9264,N_8267);
nand U11573 (N_11573,N_7858,N_7223);
or U11574 (N_11574,N_8496,N_9346);
nand U11575 (N_11575,N_8704,N_9843);
nor U11576 (N_11576,N_5688,N_9508);
xnor U11577 (N_11577,N_9634,N_9852);
or U11578 (N_11578,N_6455,N_5088);
and U11579 (N_11579,N_8656,N_5864);
xnor U11580 (N_11580,N_7015,N_8020);
nand U11581 (N_11581,N_8142,N_9460);
xnor U11582 (N_11582,N_7607,N_5341);
nand U11583 (N_11583,N_8246,N_9622);
nand U11584 (N_11584,N_7416,N_6179);
or U11585 (N_11585,N_5507,N_9697);
nand U11586 (N_11586,N_8774,N_8829);
or U11587 (N_11587,N_9568,N_5351);
xor U11588 (N_11588,N_6750,N_6327);
nor U11589 (N_11589,N_8019,N_7856);
and U11590 (N_11590,N_7340,N_9178);
and U11591 (N_11591,N_8529,N_5018);
or U11592 (N_11592,N_9200,N_8971);
nand U11593 (N_11593,N_6944,N_8668);
nor U11594 (N_11594,N_9659,N_9397);
nand U11595 (N_11595,N_6612,N_9471);
xnor U11596 (N_11596,N_5247,N_6287);
or U11597 (N_11597,N_9743,N_6076);
nor U11598 (N_11598,N_6596,N_6617);
nand U11599 (N_11599,N_8745,N_7478);
or U11600 (N_11600,N_6229,N_6469);
and U11601 (N_11601,N_9592,N_6947);
xor U11602 (N_11602,N_6129,N_5686);
nand U11603 (N_11603,N_9103,N_7135);
or U11604 (N_11604,N_8032,N_6716);
and U11605 (N_11605,N_9193,N_7004);
and U11606 (N_11606,N_7007,N_5737);
or U11607 (N_11607,N_5565,N_5652);
xnor U11608 (N_11608,N_7349,N_7771);
or U11609 (N_11609,N_5194,N_8718);
nand U11610 (N_11610,N_6037,N_7274);
or U11611 (N_11611,N_9213,N_8510);
xnor U11612 (N_11612,N_6845,N_8259);
xnor U11613 (N_11613,N_9795,N_8795);
and U11614 (N_11614,N_8890,N_7151);
xnor U11615 (N_11615,N_6782,N_6765);
or U11616 (N_11616,N_6804,N_8927);
nor U11617 (N_11617,N_5548,N_6580);
nand U11618 (N_11618,N_7452,N_7022);
nand U11619 (N_11619,N_5919,N_7198);
and U11620 (N_11620,N_8102,N_5139);
xnor U11621 (N_11621,N_8088,N_5711);
or U11622 (N_11622,N_9749,N_7437);
or U11623 (N_11623,N_9605,N_5491);
xnor U11624 (N_11624,N_6019,N_7442);
nor U11625 (N_11625,N_9136,N_6999);
xor U11626 (N_11626,N_8568,N_9145);
and U11627 (N_11627,N_8041,N_6605);
nand U11628 (N_11628,N_6779,N_9790);
xnor U11629 (N_11629,N_7039,N_5102);
or U11630 (N_11630,N_9210,N_5280);
or U11631 (N_11631,N_6727,N_6552);
and U11632 (N_11632,N_8440,N_8639);
nand U11633 (N_11633,N_8495,N_8150);
and U11634 (N_11634,N_8859,N_7345);
xnor U11635 (N_11635,N_5774,N_9671);
xor U11636 (N_11636,N_8446,N_6827);
nor U11637 (N_11637,N_6917,N_9639);
or U11638 (N_11638,N_5190,N_8564);
nand U11639 (N_11639,N_9102,N_6920);
nor U11640 (N_11640,N_7953,N_5449);
and U11641 (N_11641,N_7420,N_9635);
nor U11642 (N_11642,N_7322,N_6339);
xor U11643 (N_11643,N_6631,N_6502);
nand U11644 (N_11644,N_8525,N_9562);
nand U11645 (N_11645,N_7784,N_5360);
nor U11646 (N_11646,N_5816,N_8883);
nor U11647 (N_11647,N_6263,N_8128);
and U11648 (N_11648,N_5119,N_7689);
xnor U11649 (N_11649,N_6276,N_9322);
or U11650 (N_11650,N_8501,N_6618);
xor U11651 (N_11651,N_7396,N_6749);
xor U11652 (N_11652,N_9631,N_6712);
nor U11653 (N_11653,N_5093,N_8914);
and U11654 (N_11654,N_7941,N_6448);
nand U11655 (N_11655,N_7909,N_9241);
nand U11656 (N_11656,N_7496,N_5233);
nand U11657 (N_11657,N_6932,N_6390);
and U11658 (N_11658,N_8815,N_7727);
nor U11659 (N_11659,N_5262,N_6042);
nor U11660 (N_11660,N_9529,N_6323);
and U11661 (N_11661,N_7462,N_8086);
and U11662 (N_11662,N_6904,N_9834);
nand U11663 (N_11663,N_7656,N_6689);
xnor U11664 (N_11664,N_8183,N_6985);
and U11665 (N_11665,N_7362,N_5243);
or U11666 (N_11666,N_8011,N_7949);
nand U11667 (N_11667,N_5415,N_8392);
xnor U11668 (N_11668,N_8850,N_6017);
and U11669 (N_11669,N_6833,N_7502);
nor U11670 (N_11670,N_7018,N_5520);
nor U11671 (N_11671,N_9465,N_8452);
and U11672 (N_11672,N_7497,N_6571);
nor U11673 (N_11673,N_8940,N_8611);
or U11674 (N_11674,N_9022,N_7930);
nand U11675 (N_11675,N_7139,N_5413);
xnor U11676 (N_11676,N_7810,N_9996);
nand U11677 (N_11677,N_6200,N_6636);
xor U11678 (N_11678,N_8131,N_7292);
and U11679 (N_11679,N_7278,N_5362);
or U11680 (N_11680,N_5122,N_6851);
xor U11681 (N_11681,N_6157,N_7287);
nand U11682 (N_11682,N_5478,N_9896);
xnor U11683 (N_11683,N_5200,N_8735);
or U11684 (N_11684,N_9881,N_5184);
xor U11685 (N_11685,N_5984,N_5560);
or U11686 (N_11686,N_8270,N_9958);
and U11687 (N_11687,N_6171,N_7104);
nand U11688 (N_11688,N_5261,N_7863);
nand U11689 (N_11689,N_6817,N_5366);
nand U11690 (N_11690,N_8376,N_8406);
and U11691 (N_11691,N_5640,N_5435);
and U11692 (N_11692,N_8813,N_8291);
nand U11693 (N_11693,N_8113,N_6797);
or U11694 (N_11694,N_5960,N_9612);
xnor U11695 (N_11695,N_7404,N_7159);
and U11696 (N_11696,N_9670,N_8582);
nor U11697 (N_11697,N_9530,N_5039);
nand U11698 (N_11698,N_8736,N_5061);
and U11699 (N_11699,N_7872,N_8899);
or U11700 (N_11700,N_6241,N_8504);
xnor U11701 (N_11701,N_6298,N_8633);
or U11702 (N_11702,N_5558,N_5125);
nand U11703 (N_11703,N_7729,N_9272);
nor U11704 (N_11704,N_7751,N_7710);
or U11705 (N_11705,N_7906,N_7932);
nor U11706 (N_11706,N_5427,N_8187);
nand U11707 (N_11707,N_6495,N_5839);
or U11708 (N_11708,N_9187,N_7046);
nor U11709 (N_11709,N_5442,N_6061);
nand U11710 (N_11710,N_5731,N_5251);
and U11711 (N_11711,N_8374,N_8210);
nand U11712 (N_11712,N_8456,N_9385);
and U11713 (N_11713,N_9497,N_7011);
and U11714 (N_11714,N_8465,N_6528);
xor U11715 (N_11715,N_9319,N_6963);
and U11716 (N_11716,N_9316,N_6711);
nand U11717 (N_11717,N_9869,N_5573);
and U11718 (N_11718,N_5885,N_8915);
nor U11719 (N_11719,N_6766,N_6225);
or U11720 (N_11720,N_8687,N_8621);
or U11721 (N_11721,N_5484,N_7986);
xor U11722 (N_11722,N_5753,N_8403);
xor U11723 (N_11723,N_5315,N_6033);
and U11724 (N_11724,N_7546,N_5653);
or U11725 (N_11725,N_6255,N_5597);
or U11726 (N_11726,N_9868,N_5320);
xor U11727 (N_11727,N_7597,N_7023);
xor U11728 (N_11728,N_8366,N_5486);
or U11729 (N_11729,N_8516,N_8509);
nor U11730 (N_11730,N_7753,N_6884);
or U11731 (N_11731,N_5709,N_8061);
or U11732 (N_11732,N_8792,N_8169);
and U11733 (N_11733,N_8261,N_9691);
nor U11734 (N_11734,N_6554,N_6697);
xor U11735 (N_11735,N_5804,N_7066);
xnor U11736 (N_11736,N_7819,N_8037);
nor U11737 (N_11737,N_7512,N_6892);
nor U11738 (N_11738,N_6413,N_6537);
and U11739 (N_11739,N_6661,N_9672);
nand U11740 (N_11740,N_8577,N_7235);
nor U11741 (N_11741,N_9407,N_5424);
xnor U11742 (N_11742,N_9845,N_5235);
nor U11743 (N_11743,N_7803,N_9613);
and U11744 (N_11744,N_8936,N_9761);
and U11745 (N_11745,N_7158,N_8234);
and U11746 (N_11746,N_7860,N_8827);
or U11747 (N_11747,N_6644,N_9720);
nand U11748 (N_11748,N_6696,N_6622);
nor U11749 (N_11749,N_5893,N_9581);
nor U11750 (N_11750,N_6772,N_9593);
nor U11751 (N_11751,N_5114,N_7693);
or U11752 (N_11752,N_8534,N_8541);
and U11753 (N_11753,N_8649,N_5831);
nand U11754 (N_11754,N_8862,N_5264);
or U11755 (N_11755,N_9301,N_7459);
xor U11756 (N_11756,N_8779,N_7552);
and U11757 (N_11757,N_8689,N_9738);
or U11758 (N_11758,N_5638,N_6976);
nor U11759 (N_11759,N_9171,N_6657);
or U11760 (N_11760,N_5903,N_5808);
or U11761 (N_11761,N_9652,N_9666);
or U11762 (N_11762,N_8289,N_8236);
and U11763 (N_11763,N_7686,N_6606);
xor U11764 (N_11764,N_5574,N_6038);
xor U11765 (N_11765,N_6935,N_6446);
and U11766 (N_11766,N_9781,N_9325);
nand U11767 (N_11767,N_6533,N_7569);
xnor U11768 (N_11768,N_9395,N_5456);
nand U11769 (N_11769,N_7896,N_7242);
nand U11770 (N_11770,N_7165,N_9808);
nand U11771 (N_11771,N_5129,N_6471);
nand U11772 (N_11772,N_5288,N_5715);
and U11773 (N_11773,N_6700,N_7038);
xnor U11774 (N_11774,N_8325,N_8858);
xor U11775 (N_11775,N_5463,N_8136);
nand U11776 (N_11776,N_5299,N_9882);
nand U11777 (N_11777,N_7025,N_8889);
or U11778 (N_11778,N_6210,N_5372);
nor U11779 (N_11779,N_7098,N_5370);
and U11780 (N_11780,N_8317,N_8874);
nand U11781 (N_11781,N_7648,N_5052);
nor U11782 (N_11782,N_5708,N_6162);
or U11783 (N_11783,N_8274,N_7695);
and U11784 (N_11784,N_9201,N_6555);
xnor U11785 (N_11785,N_8093,N_7092);
or U11786 (N_11786,N_5483,N_8669);
xnor U11787 (N_11787,N_5654,N_7525);
nand U11788 (N_11788,N_9995,N_6878);
and U11789 (N_11789,N_5633,N_8977);
xor U11790 (N_11790,N_9713,N_8942);
xor U11791 (N_11791,N_9186,N_6325);
xor U11792 (N_11792,N_8688,N_6125);
xnor U11793 (N_11793,N_5091,N_9174);
or U11794 (N_11794,N_8768,N_9358);
nor U11795 (N_11795,N_7769,N_5465);
nand U11796 (N_11796,N_9660,N_6228);
and U11797 (N_11797,N_7968,N_9887);
and U11798 (N_11798,N_8031,N_8230);
nor U11799 (N_11799,N_5937,N_6434);
xor U11800 (N_11800,N_9242,N_7961);
or U11801 (N_11801,N_5173,N_5409);
and U11802 (N_11802,N_7778,N_5678);
and U11803 (N_11803,N_7971,N_9574);
or U11804 (N_11804,N_6411,N_8453);
or U11805 (N_11805,N_9980,N_9975);
xor U11806 (N_11806,N_8115,N_8096);
nor U11807 (N_11807,N_5155,N_5376);
or U11808 (N_11808,N_9279,N_7255);
nand U11809 (N_11809,N_5886,N_5180);
or U11810 (N_11810,N_7990,N_9785);
nor U11811 (N_11811,N_9537,N_7394);
nand U11812 (N_11812,N_6401,N_9268);
nor U11813 (N_11813,N_7522,N_6212);
or U11814 (N_11814,N_7828,N_5087);
nand U11815 (N_11815,N_8898,N_7060);
nand U11816 (N_11816,N_5729,N_6099);
xor U11817 (N_11817,N_5381,N_9949);
xor U11818 (N_11818,N_9047,N_7605);
or U11819 (N_11819,N_8762,N_8332);
nor U11820 (N_11820,N_8763,N_5310);
nor U11821 (N_11821,N_7399,N_7105);
and U11822 (N_11822,N_9479,N_5434);
and U11823 (N_11823,N_9251,N_6360);
nand U11824 (N_11824,N_8894,N_9690);
nand U11825 (N_11825,N_6519,N_7681);
or U11826 (N_11826,N_7655,N_8570);
nor U11827 (N_11827,N_8658,N_9115);
nor U11828 (N_11828,N_7910,N_8034);
nor U11829 (N_11829,N_7207,N_5825);
nand U11830 (N_11830,N_5658,N_6270);
xnor U11831 (N_11831,N_9531,N_6578);
or U11832 (N_11832,N_9740,N_9594);
xor U11833 (N_11833,N_6510,N_5040);
or U11834 (N_11834,N_7568,N_8337);
nand U11835 (N_11835,N_9784,N_7994);
and U11836 (N_11836,N_5417,N_9305);
xnor U11837 (N_11837,N_5127,N_5932);
or U11838 (N_11838,N_7912,N_9866);
or U11839 (N_11839,N_8993,N_9944);
xnor U11840 (N_11840,N_6449,N_5112);
nor U11841 (N_11841,N_8887,N_7294);
and U11842 (N_11842,N_6864,N_5710);
xnor U11843 (N_11843,N_7890,N_9089);
nand U11844 (N_11844,N_9462,N_6435);
xor U11845 (N_11845,N_8589,N_8968);
and U11846 (N_11846,N_5241,N_7474);
and U11847 (N_11847,N_8427,N_8816);
and U11848 (N_11848,N_5037,N_6405);
or U11849 (N_11849,N_8753,N_6442);
nor U11850 (N_11850,N_9810,N_5554);
and U11851 (N_11851,N_8531,N_5475);
and U11852 (N_11852,N_5888,N_9602);
xor U11853 (N_11853,N_6847,N_6431);
nor U11854 (N_11854,N_5027,N_5779);
xnor U11855 (N_11855,N_5193,N_9275);
or U11856 (N_11856,N_8472,N_7476);
nand U11857 (N_11857,N_8972,N_7187);
or U11858 (N_11858,N_8299,N_5132);
and U11859 (N_11859,N_5600,N_7544);
nand U11860 (N_11860,N_6666,N_7805);
or U11861 (N_11861,N_6587,N_7297);
and U11862 (N_11862,N_9825,N_9216);
and U11863 (N_11863,N_5167,N_6856);
xnor U11864 (N_11864,N_6065,N_6741);
or U11865 (N_11865,N_7781,N_6101);
or U11866 (N_11866,N_5402,N_8486);
nand U11867 (N_11867,N_7802,N_5927);
xor U11868 (N_11868,N_5266,N_9894);
and U11869 (N_11869,N_8511,N_9437);
or U11870 (N_11870,N_9591,N_9997);
xnor U11871 (N_11871,N_6382,N_5962);
or U11872 (N_11872,N_5672,N_6026);
or U11873 (N_11873,N_7183,N_5485);
nor U11874 (N_11874,N_6692,N_8722);
and U11875 (N_11875,N_6790,N_9130);
and U11876 (N_11876,N_6067,N_6583);
nand U11877 (N_11877,N_7685,N_8964);
nand U11878 (N_11878,N_7955,N_6165);
and U11879 (N_11879,N_9436,N_7460);
and U11880 (N_11880,N_9886,N_8307);
xor U11881 (N_11881,N_8489,N_5748);
nor U11882 (N_11882,N_7418,N_5152);
nor U11883 (N_11883,N_8893,N_8809);
or U11884 (N_11884,N_5131,N_9068);
nor U11885 (N_11885,N_7291,N_6520);
or U11886 (N_11886,N_9221,N_9913);
nor U11887 (N_11887,N_9356,N_6810);
and U11888 (N_11888,N_9842,N_8394);
xnor U11889 (N_11889,N_8742,N_5811);
nand U11890 (N_11890,N_6149,N_5632);
and U11891 (N_11891,N_9133,N_9764);
or U11892 (N_11892,N_9752,N_9087);
xnor U11893 (N_11893,N_7204,N_6307);
and U11894 (N_11894,N_5786,N_9387);
or U11895 (N_11895,N_6493,N_6994);
xor U11896 (N_11896,N_6786,N_8046);
nor U11897 (N_11897,N_8003,N_6724);
xnor U11898 (N_11898,N_8342,N_5889);
nor U11899 (N_11899,N_9767,N_6667);
xnor U11900 (N_11900,N_6412,N_8233);
and U11901 (N_11901,N_8390,N_8566);
nor U11902 (N_11902,N_7762,N_8252);
nand U11903 (N_11903,N_7837,N_7312);
nand U11904 (N_11904,N_9366,N_9458);
nor U11905 (N_11905,N_5861,N_5819);
nor U11906 (N_11906,N_7709,N_7584);
and U11907 (N_11907,N_7794,N_9981);
and U11908 (N_11908,N_5090,N_7289);
and U11909 (N_11909,N_9198,N_9615);
nand U11910 (N_11910,N_6900,N_7801);
or U11911 (N_11911,N_8369,N_9209);
and U11912 (N_11912,N_9902,N_9196);
or U11913 (N_11913,N_6234,N_9162);
and U11914 (N_11914,N_9567,N_6731);
nor U11915 (N_11915,N_6290,N_9814);
or U11916 (N_11916,N_6394,N_6454);
nor U11917 (N_11917,N_9120,N_7124);
or U11918 (N_11918,N_9222,N_6773);
nor U11919 (N_11919,N_5126,N_6494);
xor U11920 (N_11920,N_6464,N_9124);
nand U11921 (N_11921,N_7083,N_9502);
or U11922 (N_11922,N_8345,N_8280);
nor U11923 (N_11923,N_8623,N_5769);
nor U11924 (N_11924,N_5750,N_7934);
nor U11925 (N_11925,N_9739,N_5244);
or U11926 (N_11926,N_8196,N_9003);
or U11927 (N_11927,N_7969,N_6563);
nand U11928 (N_11928,N_6730,N_5177);
or U11929 (N_11929,N_8125,N_9919);
xnor U11930 (N_11930,N_6737,N_6070);
nor U11931 (N_11931,N_9259,N_6009);
xor U11932 (N_11932,N_5309,N_9474);
nand U11933 (N_11933,N_9988,N_9493);
nor U11934 (N_11934,N_9485,N_9049);
xor U11935 (N_11935,N_9180,N_8729);
or U11936 (N_11936,N_6377,N_9892);
and U11937 (N_11937,N_7861,N_8232);
nor U11938 (N_11938,N_6886,N_7651);
nand U11939 (N_11939,N_8292,N_9076);
xor U11940 (N_11940,N_6284,N_7449);
nand U11941 (N_11941,N_9778,N_7641);
nor U11942 (N_11942,N_6096,N_9504);
nand U11943 (N_11943,N_8123,N_8152);
or U11944 (N_11944,N_7731,N_6278);
nor U11945 (N_11945,N_8796,N_8451);
nor U11946 (N_11946,N_8637,N_5353);
and U11947 (N_11947,N_5993,N_5019);
or U11948 (N_11948,N_5267,N_5704);
nand U11949 (N_11949,N_5998,N_8329);
xnor U11950 (N_11950,N_5312,N_6839);
nor U11951 (N_11951,N_8075,N_7472);
nand U11952 (N_11952,N_9056,N_7422);
nand U11953 (N_11953,N_6668,N_5455);
nor U11954 (N_11954,N_8750,N_7074);
and U11955 (N_11955,N_8974,N_5446);
or U11956 (N_11956,N_6326,N_6077);
nor U11957 (N_11957,N_7348,N_9486);
or U11958 (N_11958,N_8454,N_5469);
and U11959 (N_11959,N_6518,N_7511);
and U11960 (N_11960,N_6375,N_9215);
xnor U11961 (N_11961,N_5356,N_8492);
nand U11962 (N_11962,N_6075,N_8012);
xnor U11963 (N_11963,N_9034,N_8997);
nand U11964 (N_11964,N_8752,N_7545);
or U11965 (N_11965,N_5929,N_8600);
and U11966 (N_11966,N_7208,N_7752);
and U11967 (N_11967,N_5869,N_6111);
nor U11968 (N_11968,N_5778,N_7360);
or U11969 (N_11969,N_9231,N_6054);
nand U11970 (N_11970,N_5955,N_8461);
nand U11971 (N_11971,N_9482,N_5540);
and U11972 (N_11972,N_8062,N_6347);
nor U11973 (N_11973,N_5317,N_5407);
nor U11974 (N_11974,N_9737,N_7284);
nand U11975 (N_11975,N_8368,N_6879);
nand U11976 (N_11976,N_5598,N_9191);
xnor U11977 (N_11977,N_5134,N_9059);
nand U11978 (N_11978,N_9815,N_7816);
and U11979 (N_11979,N_8330,N_6466);
and U11980 (N_11980,N_8522,N_9027);
xnor U11981 (N_11981,N_5818,N_9396);
or U11982 (N_11982,N_8226,N_8609);
nand U11983 (N_11983,N_9985,N_5473);
xnor U11984 (N_11984,N_5562,N_5385);
nand U11985 (N_11985,N_7936,N_7010);
xnor U11986 (N_11986,N_5544,N_5196);
or U11987 (N_11987,N_6169,N_8165);
and U11988 (N_11988,N_9383,N_9580);
or U11989 (N_11989,N_9127,N_9973);
nand U11990 (N_11990,N_5202,N_8281);
nor U11991 (N_11991,N_6549,N_9569);
or U11992 (N_11992,N_9547,N_6262);
and U11993 (N_11993,N_6117,N_5821);
nor U11994 (N_11994,N_6770,N_7132);
and U11995 (N_11995,N_7128,N_6091);
nor U11996 (N_11996,N_8106,N_5801);
xor U11997 (N_11997,N_5011,N_6130);
nand U11998 (N_11998,N_6916,N_7824);
xnor U11999 (N_11999,N_9910,N_7306);
and U12000 (N_12000,N_9961,N_8591);
and U12001 (N_12001,N_7220,N_9026);
xnor U12002 (N_12002,N_9243,N_8784);
and U12003 (N_12003,N_9703,N_7441);
xnor U12004 (N_12004,N_6211,N_9692);
and U12005 (N_12005,N_7408,N_8047);
and U12006 (N_12006,N_8699,N_6867);
nor U12007 (N_12007,N_8185,N_8963);
nand U12008 (N_12008,N_6792,N_6006);
nor U12009 (N_12009,N_7725,N_5340);
nand U12010 (N_12010,N_5007,N_6335);
xor U12011 (N_12011,N_7615,N_5331);
and U12012 (N_12012,N_6488,N_7527);
nand U12013 (N_12013,N_9736,N_8193);
and U12014 (N_12014,N_6576,N_8139);
xor U12015 (N_12015,N_9466,N_7621);
nand U12016 (N_12016,N_6505,N_8841);
nand U12017 (N_12017,N_6163,N_6694);
xnor U12018 (N_12018,N_9223,N_8999);
nand U12019 (N_12019,N_6938,N_8851);
xor U12020 (N_12020,N_9512,N_9751);
or U12021 (N_12021,N_6758,N_8158);
xnor U12022 (N_12022,N_7401,N_5584);
xnor U12023 (N_12023,N_9728,N_7547);
nor U12024 (N_12024,N_7325,N_9086);
nand U12025 (N_12025,N_5963,N_6565);
nor U12026 (N_12026,N_8998,N_5023);
nand U12027 (N_12027,N_8627,N_7055);
xnor U12028 (N_12028,N_5619,N_5075);
and U12029 (N_12029,N_9245,N_6388);
and U12030 (N_12030,N_9920,N_9229);
nor U12031 (N_12031,N_6574,N_7683);
xor U12032 (N_12032,N_6112,N_6363);
or U12033 (N_12033,N_6614,N_7377);
nand U12034 (N_12034,N_8685,N_7175);
or U12035 (N_12035,N_5747,N_7091);
and U12036 (N_12036,N_5466,N_6321);
or U12037 (N_12037,N_5912,N_6516);
xnor U12038 (N_12038,N_6153,N_5596);
nand U12039 (N_12039,N_5707,N_5780);
nor U12040 (N_12040,N_6638,N_9771);
nand U12041 (N_12041,N_6029,N_8818);
nor U12042 (N_12042,N_8777,N_5031);
nor U12043 (N_12043,N_7020,N_9876);
and U12044 (N_12044,N_6243,N_7019);
and U12045 (N_12045,N_6849,N_7251);
nor U12046 (N_12046,N_8056,N_6676);
nand U12047 (N_12047,N_6868,N_7392);
and U12048 (N_12048,N_5901,N_7140);
and U12049 (N_12049,N_9374,N_8500);
nand U12050 (N_12050,N_5318,N_8952);
nor U12051 (N_12051,N_5328,N_9318);
and U12052 (N_12052,N_7127,N_9914);
nand U12053 (N_12053,N_5003,N_5470);
nor U12054 (N_12054,N_8328,N_7260);
or U12055 (N_12055,N_6219,N_6945);
nor U12056 (N_12056,N_8601,N_5453);
xor U12057 (N_12057,N_9971,N_5761);
or U12058 (N_12058,N_5862,N_6987);
nor U12059 (N_12059,N_8919,N_6055);
and U12060 (N_12060,N_6427,N_9326);
xnor U12061 (N_12061,N_5700,N_5128);
nor U12062 (N_12062,N_6811,N_7815);
and U12063 (N_12063,N_7884,N_5257);
nand U12064 (N_12064,N_6857,N_9399);
and U12065 (N_12065,N_7706,N_8442);
nand U12066 (N_12066,N_7146,N_9813);
nand U12067 (N_12067,N_8090,N_9873);
and U12068 (N_12068,N_9300,N_8828);
and U12069 (N_12069,N_9554,N_8900);
or U12070 (N_12070,N_9503,N_5322);
and U12071 (N_12071,N_9608,N_8464);
and U12072 (N_12072,N_6834,N_8693);
xnor U12073 (N_12073,N_9267,N_6193);
nor U12074 (N_12074,N_6414,N_7818);
xor U12075 (N_12075,N_7997,N_5105);
or U12076 (N_12076,N_6529,N_9848);
xnor U12077 (N_12077,N_9236,N_9930);
nand U12078 (N_12078,N_6088,N_6484);
xnor U12079 (N_12079,N_5837,N_6373);
nand U12080 (N_12080,N_8706,N_8072);
nand U12081 (N_12081,N_6771,N_7361);
and U12082 (N_12082,N_9711,N_9684);
nor U12083 (N_12083,N_6873,N_6288);
or U12084 (N_12084,N_5325,N_7903);
nor U12085 (N_12085,N_6138,N_6501);
nand U12086 (N_12086,N_5954,N_5166);
nor U12087 (N_12087,N_6558,N_8544);
and U12088 (N_12088,N_6292,N_7233);
or U12089 (N_12089,N_6063,N_6669);
nand U12090 (N_12090,N_6504,N_7532);
or U12091 (N_12091,N_9109,N_6320);
xor U12092 (N_12092,N_7593,N_9904);
xnor U12093 (N_12093,N_5936,N_8530);
nor U12094 (N_12094,N_8372,N_8121);
nand U12095 (N_12095,N_7446,N_7230);
nand U12096 (N_12096,N_8780,N_6936);
or U12097 (N_12097,N_5767,N_6438);
xnor U12098 (N_12098,N_7427,N_6104);
nor U12099 (N_12099,N_7239,N_6203);
nand U12100 (N_12100,N_5582,N_8155);
and U12101 (N_12101,N_5033,N_8470);
nand U12102 (N_12102,N_5879,N_8880);
and U12103 (N_12103,N_7517,N_5165);
nand U12104 (N_12104,N_9142,N_6031);
and U12105 (N_12105,N_9192,N_6106);
nor U12106 (N_12106,N_5332,N_7581);
xor U12107 (N_12107,N_8404,N_6769);
nand U12108 (N_12108,N_9054,N_9898);
nand U12109 (N_12109,N_7739,N_7465);
xnor U12110 (N_12110,N_8429,N_8008);
nor U12111 (N_12111,N_5758,N_9132);
nand U12112 (N_12112,N_8219,N_8546);
nor U12113 (N_12113,N_5186,N_6397);
xor U12114 (N_12114,N_5592,N_9669);
nor U12115 (N_12115,N_8297,N_8014);
nor U12116 (N_12116,N_5890,N_9540);
nand U12117 (N_12117,N_9702,N_7981);
nand U12118 (N_12118,N_5985,N_5001);
nand U12119 (N_12119,N_7266,N_8798);
or U12120 (N_12120,N_9793,N_7887);
nand U12121 (N_12121,N_9519,N_5272);
nor U12122 (N_12122,N_5994,N_6240);
xor U12123 (N_12123,N_7979,N_8381);
nand U12124 (N_12124,N_8109,N_5675);
nor U12125 (N_12125,N_6396,N_9983);
nand U12126 (N_12126,N_7332,N_8810);
nand U12127 (N_12127,N_8864,N_6807);
or U12128 (N_12128,N_8843,N_7076);
or U12129 (N_12129,N_9270,N_6590);
nor U12130 (N_12130,N_9851,N_7378);
nand U12131 (N_12131,N_7373,N_9685);
xnor U12132 (N_12132,N_7875,N_8029);
nand U12133 (N_12133,N_7439,N_7035);
or U12134 (N_12134,N_5734,N_9344);
nand U12135 (N_12135,N_9578,N_5768);
nor U12136 (N_12136,N_6719,N_6621);
or U12137 (N_12137,N_6328,N_9388);
nor U12138 (N_12138,N_9163,N_5525);
xnor U12139 (N_12139,N_8793,N_9768);
nand U12140 (N_12140,N_7514,N_7697);
xor U12141 (N_12141,N_5664,N_9204);
nor U12142 (N_12142,N_5293,N_9261);
nor U12143 (N_12143,N_8691,N_6074);
nor U12144 (N_12144,N_6880,N_6249);
xor U12145 (N_12145,N_6121,N_8336);
nand U12146 (N_12146,N_5000,N_5610);
nand U12147 (N_12147,N_9007,N_5983);
or U12148 (N_12148,N_8901,N_8620);
and U12149 (N_12149,N_5749,N_5848);
nand U12150 (N_12150,N_9880,N_7687);
xnor U12151 (N_12151,N_8361,N_6470);
nand U12152 (N_12152,N_7834,N_8471);
and U12153 (N_12153,N_8430,N_6717);
xor U12154 (N_12154,N_5279,N_6840);
or U12155 (N_12155,N_5877,N_6780);
and U12156 (N_12156,N_8981,N_7914);
nand U12157 (N_12157,N_7629,N_8048);
nor U12158 (N_12158,N_5802,N_9104);
xor U12159 (N_12159,N_6258,N_9820);
nor U12160 (N_12160,N_7832,N_7889);
nor U12161 (N_12161,N_8491,N_7050);
and U12162 (N_12162,N_9890,N_6081);
nor U12163 (N_12163,N_9776,N_9331);
nor U12164 (N_12164,N_5705,N_5916);
or U12165 (N_12165,N_7804,N_6341);
and U12166 (N_12166,N_7962,N_5298);
or U12167 (N_12167,N_8831,N_5812);
nand U12168 (N_12168,N_8010,N_7741);
or U12169 (N_12169,N_7081,N_9139);
nor U12170 (N_12170,N_8103,N_8400);
nand U12171 (N_12171,N_5250,N_9053);
xnor U12172 (N_12172,N_5595,N_6722);
xnor U12173 (N_12173,N_8697,N_6456);
or U12174 (N_12174,N_7161,N_6384);
nor U12175 (N_12175,N_8512,N_5457);
xor U12176 (N_12176,N_7090,N_8079);
or U12177 (N_12177,N_6584,N_8101);
and U12178 (N_12178,N_7376,N_7317);
or U12179 (N_12179,N_8751,N_5843);
nor U12180 (N_12180,N_5256,N_5373);
xnor U12181 (N_12181,N_7002,N_8263);
nor U12182 (N_12182,N_6058,N_7455);
xor U12183 (N_12183,N_9926,N_9505);
and U12184 (N_12184,N_8844,N_9867);
or U12185 (N_12185,N_5265,N_8628);
xnor U12186 (N_12186,N_8306,N_9128);
nand U12187 (N_12187,N_5896,N_8126);
nand U12188 (N_12188,N_8962,N_7369);
xor U12189 (N_12189,N_8416,N_5029);
xor U12190 (N_12190,N_6487,N_6802);
nand U12191 (N_12191,N_5752,N_9928);
xnor U12192 (N_12192,N_9750,N_7780);
nor U12193 (N_12193,N_7663,N_7174);
xor U12194 (N_12194,N_9539,N_9362);
nand U12195 (N_12195,N_7190,N_9600);
nand U12196 (N_12196,N_6164,N_7041);
nor U12197 (N_12197,N_5444,N_9207);
xnor U12198 (N_12198,N_8926,N_5736);
xor U12199 (N_12199,N_8980,N_7095);
xnor U12200 (N_12200,N_7586,N_5354);
xor U12201 (N_12201,N_9443,N_5248);
nand U12202 (N_12202,N_6843,N_7051);
nor U12203 (N_12203,N_6259,N_9799);
nor U12204 (N_12204,N_9011,N_7555);
nor U12205 (N_12205,N_6787,N_9310);
and U12206 (N_12206,N_5908,N_8124);
xnor U12207 (N_12207,N_5213,N_5807);
nor U12208 (N_12208,N_8091,N_7515);
xnor U12209 (N_12209,N_6002,N_5021);
xor U12210 (N_12210,N_6108,N_5766);
nor U12211 (N_12211,N_7513,N_5464);
xnor U12212 (N_12212,N_5002,N_9850);
nor U12213 (N_12213,N_8625,N_5826);
xnor U12214 (N_12214,N_8678,N_7001);
xnor U12215 (N_12215,N_5529,N_9151);
xnor U12216 (N_12216,N_5892,N_5344);
or U12217 (N_12217,N_5834,N_9321);
and U12218 (N_12218,N_6826,N_5249);
and U12219 (N_12219,N_9334,N_8356);
nand U12220 (N_12220,N_8709,N_7209);
and U12221 (N_12221,N_5611,N_9823);
xor U12222 (N_12222,N_5663,N_9879);
and U12223 (N_12223,N_8064,N_8759);
or U12224 (N_12224,N_8819,N_7119);
nor U12225 (N_12225,N_5679,N_9481);
nor U12226 (N_12226,N_7617,N_9349);
and U12227 (N_12227,N_5124,N_6358);
and U12228 (N_12228,N_9227,N_8497);
or U12229 (N_12229,N_5692,N_8084);
nor U12230 (N_12230,N_5756,N_9219);
and U12231 (N_12231,N_5397,N_5333);
or U12232 (N_12232,N_6531,N_9057);
and U12233 (N_12233,N_9870,N_5030);
nor U12234 (N_12234,N_7921,N_9877);
nor U12235 (N_12235,N_9899,N_7113);
nand U12236 (N_12236,N_7444,N_5996);
and U12237 (N_12237,N_6799,N_9025);
nand U12238 (N_12238,N_8251,N_7411);
nor U12239 (N_12239,N_5460,N_7891);
and U12240 (N_12240,N_6468,N_9035);
nand U12241 (N_12241,N_5348,N_6190);
xnor U12242 (N_12242,N_7269,N_6500);
and U12243 (N_12243,N_5832,N_6450);
and U12244 (N_12244,N_9036,N_8009);
xor U12245 (N_12245,N_6951,N_5897);
xor U12246 (N_12246,N_6862,N_7356);
nor U12247 (N_12247,N_8690,N_5946);
and U12248 (N_12248,N_8604,N_5720);
xnor U12249 (N_12249,N_7830,N_7283);
and U12250 (N_12250,N_8636,N_6872);
nor U12251 (N_12251,N_9373,N_7734);
xor U12252 (N_12252,N_9582,N_5568);
and U12253 (N_12253,N_9806,N_6167);
or U12254 (N_12254,N_7646,N_9837);
nand U12255 (N_12255,N_8242,N_5959);
xor U12256 (N_12256,N_9907,N_7030);
nor U12257 (N_12257,N_6763,N_8284);
or U12258 (N_12258,N_7320,N_9446);
nor U12259 (N_12259,N_7040,N_6227);
nand U12260 (N_12260,N_8651,N_6223);
and U12261 (N_12261,N_9253,N_6551);
or U12262 (N_12262,N_8194,N_7662);
nor U12263 (N_12263,N_8594,N_5553);
or U12264 (N_12264,N_6718,N_8178);
nand U12265 (N_12265,N_7121,N_8741);
nor U12266 (N_12266,N_7848,N_5103);
nand U12267 (N_12267,N_8904,N_8562);
nand U12268 (N_12268,N_6443,N_8050);
nor U12269 (N_12269,N_6453,N_6822);
nand U12270 (N_12270,N_9856,N_5978);
nor U12271 (N_12271,N_6146,N_8608);
nand U12272 (N_12272,N_5701,N_7285);
or U12273 (N_12273,N_5513,N_8081);
and U12274 (N_12274,N_9556,N_9998);
and U12275 (N_12275,N_6929,N_9472);
nand U12276 (N_12276,N_6476,N_8543);
nor U12277 (N_12277,N_7841,N_6016);
and U12278 (N_12278,N_9648,N_5377);
or U12279 (N_12279,N_9704,N_7744);
and U12280 (N_12280,N_7851,N_5204);
or U12281 (N_12281,N_7594,N_6126);
and U12282 (N_12282,N_6629,N_8720);
or U12283 (N_12283,N_6024,N_5009);
nor U12284 (N_12284,N_7958,N_6302);
nor U12285 (N_12285,N_6264,N_9013);
or U12286 (N_12286,N_9796,N_8038);
xnor U12287 (N_12287,N_9069,N_5187);
and U12288 (N_12288,N_5646,N_6202);
xor U12289 (N_12289,N_9657,N_9164);
or U12290 (N_12290,N_6332,N_9916);
xnor U12291 (N_12291,N_9197,N_8618);
nand U12292 (N_12292,N_9651,N_5511);
or U12293 (N_12293,N_9897,N_9324);
xnor U12294 (N_12294,N_5418,N_9756);
or U12295 (N_12295,N_8343,N_8945);
xnor U12296 (N_12296,N_9597,N_7570);
nand U12297 (N_12297,N_7488,N_6188);
or U12298 (N_12298,N_7698,N_9587);
xor U12299 (N_12299,N_8615,N_8310);
nand U12300 (N_12300,N_5684,N_6283);
nor U12301 (N_12301,N_5051,N_9606);
xnor U12302 (N_12302,N_6553,N_6701);
or U12303 (N_12303,N_9138,N_5833);
nor U12304 (N_12304,N_5988,N_8412);
or U12305 (N_12305,N_6275,N_9982);
or U12306 (N_12306,N_7786,N_7226);
or U12307 (N_12307,N_8502,N_8256);
and U12308 (N_12308,N_5379,N_5404);
nor U12309 (N_12309,N_6637,N_7963);
or U12310 (N_12310,N_8443,N_8380);
xnor U12311 (N_12311,N_5787,N_7447);
or U12312 (N_12312,N_6646,N_7454);
nand U12313 (N_12313,N_6816,N_6806);
or U12314 (N_12314,N_5541,N_5046);
nor U12315 (N_12315,N_9797,N_7888);
nand U12316 (N_12316,N_5979,N_8983);
xor U12317 (N_12317,N_6599,N_5069);
xor U12318 (N_12318,N_7774,N_7975);
nor U12319 (N_12319,N_6960,N_5017);
nor U12320 (N_12320,N_6483,N_5669);
nand U12321 (N_12321,N_7897,N_8630);
nor U12322 (N_12322,N_9989,N_7347);
xor U12323 (N_12323,N_8248,N_7282);
nor U12324 (N_12324,N_9079,N_6768);
or U12325 (N_12325,N_5907,N_7120);
xnor U12326 (N_12326,N_9523,N_8622);
nand U12327 (N_12327,N_9726,N_6641);
or U12328 (N_12328,N_7194,N_8097);
and U12329 (N_12329,N_6863,N_6548);
xnor U12330 (N_12330,N_6682,N_6268);
nor U12331 (N_12331,N_8321,N_5515);
and U12332 (N_12332,N_8909,N_8080);
nand U12333 (N_12333,N_7768,N_5183);
xor U12334 (N_12334,N_7867,N_7767);
and U12335 (N_12335,N_7389,N_7203);
and U12336 (N_12336,N_6601,N_7877);
nand U12337 (N_12337,N_5451,N_9116);
nor U12338 (N_12338,N_5205,N_6150);
and U12339 (N_12339,N_8580,N_6098);
and U12340 (N_12340,N_9160,N_7924);
xnor U12341 (N_12341,N_9614,N_6059);
and U12342 (N_12342,N_8422,N_8017);
nand U12343 (N_12343,N_7760,N_7671);
nand U12344 (N_12344,N_5495,N_8520);
nand U12345 (N_12345,N_5876,N_7653);
xnor U12346 (N_12346,N_5542,N_9583);
or U12347 (N_12347,N_9249,N_5083);
nand U12348 (N_12348,N_6045,N_9412);
or U12349 (N_12349,N_8552,N_8641);
or U12350 (N_12350,N_8214,N_6025);
nor U12351 (N_12351,N_9457,N_6967);
or U12352 (N_12352,N_5842,N_9714);
nor U12353 (N_12353,N_6791,N_8154);
xor U12354 (N_12354,N_5231,N_6380);
nor U12355 (N_12355,N_6353,N_6191);
or U12356 (N_12356,N_5297,N_8401);
or U12357 (N_12357,N_9014,N_8030);
xnor U12358 (N_12358,N_9370,N_5395);
xnor U12359 (N_12359,N_5674,N_8593);
nor U12360 (N_12360,N_7684,N_6507);
or U12361 (N_12361,N_6086,N_8420);
xnor U12362 (N_12362,N_5972,N_9844);
nand U12363 (N_12363,N_5977,N_8480);
xor U12364 (N_12364,N_7112,N_5076);
nor U12365 (N_12365,N_8988,N_9419);
or U12366 (N_12366,N_5005,N_9828);
and U12367 (N_12367,N_9177,N_9619);
nand U12368 (N_12368,N_8122,N_8955);
nor U12369 (N_12369,N_8462,N_6145);
xor U12370 (N_12370,N_8631,N_5799);
nor U12371 (N_12371,N_7182,N_7977);
nand U12372 (N_12372,N_7876,N_8223);
or U12373 (N_12373,N_6705,N_6515);
xnor U12374 (N_12374,N_7800,N_8146);
nor U12375 (N_12375,N_7931,N_9072);
nand U12376 (N_12376,N_7352,N_9835);
or U12377 (N_12377,N_8545,N_5035);
nor U12378 (N_12378,N_5060,N_6462);
nor U12379 (N_12379,N_6004,N_7267);
or U12380 (N_12380,N_8528,N_8920);
nand U12381 (N_12381,N_5953,N_6643);
nand U12382 (N_12382,N_6447,N_6419);
nand U12383 (N_12383,N_9542,N_7480);
nand U12384 (N_12384,N_8238,N_7560);
xnor U12385 (N_12385,N_9032,N_8211);
nand U12386 (N_12386,N_9527,N_8603);
and U12387 (N_12387,N_6389,N_8189);
nand U12388 (N_12388,N_5717,N_9693);
or U12389 (N_12389,N_8606,N_8157);
and U12390 (N_12390,N_8807,N_5367);
xor U12391 (N_12391,N_5292,N_9444);
and U12392 (N_12392,N_7366,N_5925);
nand U12393 (N_12393,N_6201,N_8293);
nor U12394 (N_12394,N_7079,N_8323);
nor U12395 (N_12395,N_6085,N_7247);
and U12396 (N_12396,N_7479,N_9604);
or U12397 (N_12397,N_9134,N_9716);
nor U12398 (N_12398,N_5697,N_8379);
and U12399 (N_12399,N_6542,N_5909);
nor U12400 (N_12400,N_7789,N_7213);
or U12401 (N_12401,N_6598,N_8166);
xnor U12402 (N_12402,N_5212,N_5181);
xor U12403 (N_12403,N_6044,N_8174);
or U12404 (N_12404,N_9464,N_9039);
or U12405 (N_12405,N_7042,N_7238);
and U12406 (N_12406,N_5290,N_8665);
or U12407 (N_12407,N_6035,N_7652);
or U12408 (N_12408,N_8421,N_5164);
and U12409 (N_12409,N_7154,N_8271);
or U12410 (N_12410,N_7696,N_9927);
or U12411 (N_12411,N_8870,N_8262);
xnor U12412 (N_12412,N_6331,N_6664);
nor U12413 (N_12413,N_8612,N_8213);
nor U12414 (N_12414,N_8059,N_9154);
xor U12415 (N_12415,N_9097,N_8802);
xnor U12416 (N_12416,N_6503,N_9095);
and U12417 (N_12417,N_7246,N_9543);
nand U12418 (N_12418,N_8721,N_6251);
nor U12419 (N_12419,N_8212,N_8852);
nor U12420 (N_12420,N_5531,N_9263);
nor U12421 (N_12421,N_7259,N_5074);
nand U12422 (N_12422,N_6115,N_8304);
and U12423 (N_12423,N_9676,N_8205);
and U12424 (N_12424,N_6635,N_9755);
nor U12425 (N_12425,N_7037,N_9827);
nand U12426 (N_12426,N_9546,N_6428);
and U12427 (N_12427,N_5670,N_7600);
xor U12428 (N_12428,N_8478,N_6743);
xor U12429 (N_12429,N_7094,N_7892);
nor U12430 (N_12430,N_7755,N_9051);
xor U12431 (N_12431,N_7622,N_6376);
nand U12432 (N_12432,N_9559,N_8869);
nand U12433 (N_12433,N_8273,N_8364);
or U12434 (N_12434,N_6882,N_9195);
nand U12435 (N_12435,N_6680,N_7825);
and U12436 (N_12436,N_5306,N_5151);
or U12437 (N_12437,N_9336,N_6199);
nor U12438 (N_12438,N_9500,N_5945);
xor U12439 (N_12439,N_5564,N_9762);
nor U12440 (N_12440,N_5504,N_6497);
xnor U12441 (N_12441,N_6062,N_8839);
or U12442 (N_12442,N_9271,N_7346);
nor U12443 (N_12443,N_5773,N_7519);
or U12444 (N_12444,N_5116,N_5316);
xnor U12445 (N_12445,N_7915,N_6893);
xnor U12446 (N_12446,N_8833,N_7263);
nor U12447 (N_12447,N_9874,N_5147);
and U12448 (N_12448,N_6683,N_9964);
xnor U12449 (N_12449,N_5528,N_5450);
nor U12450 (N_12450,N_5590,N_5782);
nor U12451 (N_12451,N_8417,N_6861);
or U12452 (N_12452,N_9096,N_7620);
or U12453 (N_12453,N_5696,N_6903);
nor U12454 (N_12454,N_5722,N_7865);
or U12455 (N_12455,N_9206,N_6955);
xnor U12456 (N_12456,N_5566,N_5425);
or U12457 (N_12457,N_7061,N_5412);
xnor U12458 (N_12458,N_6708,N_9131);
xor U12459 (N_12459,N_5556,N_6526);
and U12460 (N_12460,N_5263,N_6215);
xor U12461 (N_12461,N_8334,N_8708);
xnor U12462 (N_12462,N_8305,N_8737);
or U12463 (N_12463,N_9883,N_6481);
nor U12464 (N_12464,N_9282,N_5974);
nor U12465 (N_12465,N_7173,N_7412);
or U12466 (N_12466,N_8069,N_8338);
nor U12467 (N_12467,N_7732,N_7321);
and U12468 (N_12468,N_9832,N_8468);
nor U12469 (N_12469,N_8979,N_7720);
and U12470 (N_12470,N_7645,N_5079);
or U12471 (N_12471,N_8801,N_5438);
or U12472 (N_12472,N_5398,N_5433);
or U12473 (N_12473,N_9746,N_8045);
or U12474 (N_12474,N_8715,N_9694);
or U12475 (N_12475,N_9682,N_8070);
or U12476 (N_12476,N_8104,N_6424);
and U12477 (N_12477,N_9811,N_8351);
nand U12478 (N_12478,N_9984,N_5668);
and U12479 (N_12479,N_8450,N_7608);
and U12480 (N_12480,N_6591,N_5044);
nand U12481 (N_12481,N_6760,N_7882);
or U12482 (N_12482,N_8950,N_6001);
and U12483 (N_12483,N_9135,N_6926);
or U12484 (N_12484,N_7598,N_5930);
nor U12485 (N_12485,N_5323,N_7873);
and U12486 (N_12486,N_7715,N_5374);
nand U12487 (N_12487,N_6479,N_6809);
xnor U12488 (N_12488,N_6265,N_8171);
and U12489 (N_12489,N_8897,N_5175);
and U12490 (N_12490,N_8208,N_8206);
xnor U12491 (N_12491,N_7982,N_5992);
or U12492 (N_12492,N_9722,N_9410);
xor U12493 (N_12493,N_7070,N_8388);
nor U12494 (N_12494,N_6853,N_8301);
xor U12495 (N_12495,N_8177,N_9524);
nor U12496 (N_12496,N_5371,N_7700);
nand U12497 (N_12497,N_7957,N_9455);
or U12498 (N_12498,N_7948,N_8760);
and U12499 (N_12499,N_9400,N_6329);
or U12500 (N_12500,N_6332,N_5064);
nand U12501 (N_12501,N_9968,N_6635);
nor U12502 (N_12502,N_8590,N_5110);
nand U12503 (N_12503,N_9318,N_7780);
and U12504 (N_12504,N_8320,N_6733);
nor U12505 (N_12505,N_8768,N_6160);
xor U12506 (N_12506,N_9809,N_7081);
nand U12507 (N_12507,N_8107,N_6150);
and U12508 (N_12508,N_8728,N_5842);
and U12509 (N_12509,N_7449,N_9984);
nand U12510 (N_12510,N_7485,N_6739);
and U12511 (N_12511,N_5698,N_7739);
nor U12512 (N_12512,N_6323,N_9997);
and U12513 (N_12513,N_8484,N_6969);
or U12514 (N_12514,N_5386,N_9877);
xor U12515 (N_12515,N_7863,N_9108);
nor U12516 (N_12516,N_6709,N_9478);
nor U12517 (N_12517,N_6384,N_7279);
xnor U12518 (N_12518,N_8415,N_7972);
or U12519 (N_12519,N_7245,N_8696);
and U12520 (N_12520,N_9434,N_5782);
nand U12521 (N_12521,N_8605,N_8522);
nor U12522 (N_12522,N_8510,N_7419);
and U12523 (N_12523,N_6292,N_8517);
or U12524 (N_12524,N_7849,N_5469);
nor U12525 (N_12525,N_8587,N_8254);
and U12526 (N_12526,N_6061,N_9364);
or U12527 (N_12527,N_9522,N_6804);
nand U12528 (N_12528,N_5758,N_7367);
or U12529 (N_12529,N_7974,N_5321);
nand U12530 (N_12530,N_9372,N_9476);
or U12531 (N_12531,N_8039,N_7499);
or U12532 (N_12532,N_6670,N_7346);
nor U12533 (N_12533,N_8847,N_9850);
xnor U12534 (N_12534,N_9341,N_8877);
and U12535 (N_12535,N_7794,N_8948);
or U12536 (N_12536,N_5685,N_5790);
and U12537 (N_12537,N_7372,N_9295);
or U12538 (N_12538,N_8692,N_7307);
or U12539 (N_12539,N_6752,N_7994);
and U12540 (N_12540,N_9375,N_6360);
xnor U12541 (N_12541,N_6188,N_7987);
or U12542 (N_12542,N_8100,N_7671);
xnor U12543 (N_12543,N_9960,N_5228);
xnor U12544 (N_12544,N_8462,N_5166);
nand U12545 (N_12545,N_5071,N_8433);
nor U12546 (N_12546,N_7707,N_7693);
xor U12547 (N_12547,N_8917,N_9901);
nand U12548 (N_12548,N_9407,N_9726);
nand U12549 (N_12549,N_7837,N_6049);
nor U12550 (N_12550,N_8477,N_9482);
nand U12551 (N_12551,N_9005,N_7057);
xor U12552 (N_12552,N_8477,N_5261);
xor U12553 (N_12553,N_8493,N_9940);
or U12554 (N_12554,N_8205,N_5710);
nor U12555 (N_12555,N_9735,N_5166);
or U12556 (N_12556,N_8507,N_8140);
nand U12557 (N_12557,N_5430,N_9369);
nor U12558 (N_12558,N_5089,N_6509);
xor U12559 (N_12559,N_6248,N_9590);
and U12560 (N_12560,N_9854,N_6630);
nand U12561 (N_12561,N_5663,N_7300);
or U12562 (N_12562,N_5914,N_6862);
xor U12563 (N_12563,N_6131,N_7841);
and U12564 (N_12564,N_9723,N_7501);
and U12565 (N_12565,N_6832,N_6028);
xor U12566 (N_12566,N_6757,N_9796);
or U12567 (N_12567,N_6419,N_6514);
or U12568 (N_12568,N_9077,N_9050);
nand U12569 (N_12569,N_5978,N_9032);
nand U12570 (N_12570,N_5635,N_8004);
nor U12571 (N_12571,N_5314,N_9868);
nor U12572 (N_12572,N_5254,N_6708);
xnor U12573 (N_12573,N_5891,N_8651);
nor U12574 (N_12574,N_7250,N_7441);
nor U12575 (N_12575,N_5348,N_7777);
nor U12576 (N_12576,N_8401,N_6213);
and U12577 (N_12577,N_9933,N_9287);
and U12578 (N_12578,N_7293,N_8069);
xor U12579 (N_12579,N_7383,N_7534);
and U12580 (N_12580,N_9581,N_7879);
or U12581 (N_12581,N_5724,N_5497);
and U12582 (N_12582,N_8873,N_5464);
and U12583 (N_12583,N_6256,N_7787);
and U12584 (N_12584,N_8348,N_7122);
or U12585 (N_12585,N_7442,N_9249);
and U12586 (N_12586,N_8467,N_6937);
xor U12587 (N_12587,N_5468,N_6970);
or U12588 (N_12588,N_9729,N_9786);
or U12589 (N_12589,N_7437,N_9170);
nand U12590 (N_12590,N_5480,N_8406);
and U12591 (N_12591,N_6092,N_9862);
nand U12592 (N_12592,N_6412,N_9943);
nor U12593 (N_12593,N_7206,N_9084);
nor U12594 (N_12594,N_7054,N_5738);
xor U12595 (N_12595,N_9783,N_9782);
nor U12596 (N_12596,N_5110,N_7105);
nand U12597 (N_12597,N_9763,N_6634);
xor U12598 (N_12598,N_5517,N_5251);
or U12599 (N_12599,N_7530,N_6518);
nand U12600 (N_12600,N_5867,N_9581);
and U12601 (N_12601,N_5237,N_8614);
and U12602 (N_12602,N_9054,N_6744);
xor U12603 (N_12603,N_7917,N_9469);
or U12604 (N_12604,N_6929,N_8411);
or U12605 (N_12605,N_5329,N_8415);
nand U12606 (N_12606,N_9571,N_7044);
xnor U12607 (N_12607,N_7274,N_6027);
or U12608 (N_12608,N_7875,N_5380);
xor U12609 (N_12609,N_9576,N_5881);
nand U12610 (N_12610,N_5094,N_9089);
xor U12611 (N_12611,N_9009,N_8877);
or U12612 (N_12612,N_6304,N_6499);
xor U12613 (N_12613,N_5834,N_5190);
xnor U12614 (N_12614,N_9292,N_8135);
nor U12615 (N_12615,N_9649,N_9257);
nor U12616 (N_12616,N_5634,N_8577);
nand U12617 (N_12617,N_5757,N_6781);
nand U12618 (N_12618,N_9666,N_5707);
nor U12619 (N_12619,N_9723,N_7134);
nand U12620 (N_12620,N_8160,N_7321);
nor U12621 (N_12621,N_7395,N_7360);
or U12622 (N_12622,N_6637,N_8015);
nand U12623 (N_12623,N_8865,N_5059);
nor U12624 (N_12624,N_7775,N_6115);
and U12625 (N_12625,N_8926,N_7290);
nor U12626 (N_12626,N_8488,N_6029);
and U12627 (N_12627,N_6241,N_9725);
nand U12628 (N_12628,N_9966,N_7412);
nor U12629 (N_12629,N_5547,N_7928);
and U12630 (N_12630,N_8158,N_5840);
nor U12631 (N_12631,N_9624,N_5145);
and U12632 (N_12632,N_5983,N_9508);
and U12633 (N_12633,N_9964,N_8517);
nor U12634 (N_12634,N_9641,N_8736);
nand U12635 (N_12635,N_7853,N_5671);
nor U12636 (N_12636,N_6551,N_6507);
xnor U12637 (N_12637,N_6587,N_6815);
or U12638 (N_12638,N_8441,N_8003);
xnor U12639 (N_12639,N_6656,N_9463);
and U12640 (N_12640,N_7841,N_8508);
and U12641 (N_12641,N_9598,N_8680);
xor U12642 (N_12642,N_5188,N_6557);
nor U12643 (N_12643,N_9272,N_6607);
or U12644 (N_12644,N_7122,N_7113);
xor U12645 (N_12645,N_9757,N_6422);
nand U12646 (N_12646,N_7000,N_7606);
or U12647 (N_12647,N_5510,N_5485);
xor U12648 (N_12648,N_8638,N_8073);
or U12649 (N_12649,N_6377,N_7520);
or U12650 (N_12650,N_5952,N_9137);
xnor U12651 (N_12651,N_6361,N_7774);
or U12652 (N_12652,N_7131,N_5746);
and U12653 (N_12653,N_5620,N_7864);
and U12654 (N_12654,N_6277,N_9099);
or U12655 (N_12655,N_9864,N_5568);
xnor U12656 (N_12656,N_8879,N_9151);
nor U12657 (N_12657,N_9789,N_5276);
nor U12658 (N_12658,N_9197,N_8868);
nor U12659 (N_12659,N_5273,N_6582);
nand U12660 (N_12660,N_7232,N_7556);
or U12661 (N_12661,N_5333,N_8911);
nand U12662 (N_12662,N_5877,N_9725);
xor U12663 (N_12663,N_8694,N_8681);
or U12664 (N_12664,N_7077,N_5673);
and U12665 (N_12665,N_9584,N_9659);
xnor U12666 (N_12666,N_7536,N_6399);
xor U12667 (N_12667,N_8155,N_9606);
and U12668 (N_12668,N_7716,N_6978);
and U12669 (N_12669,N_6471,N_9941);
and U12670 (N_12670,N_5858,N_7087);
xor U12671 (N_12671,N_7216,N_6337);
xnor U12672 (N_12672,N_5670,N_8794);
nand U12673 (N_12673,N_6740,N_6144);
or U12674 (N_12674,N_5072,N_5858);
xnor U12675 (N_12675,N_6531,N_6525);
or U12676 (N_12676,N_7896,N_8794);
xnor U12677 (N_12677,N_8412,N_8494);
nor U12678 (N_12678,N_9893,N_9859);
nand U12679 (N_12679,N_9233,N_6843);
xor U12680 (N_12680,N_9684,N_7192);
nand U12681 (N_12681,N_6375,N_9799);
or U12682 (N_12682,N_9818,N_9039);
nor U12683 (N_12683,N_9084,N_6492);
nand U12684 (N_12684,N_9271,N_5613);
nor U12685 (N_12685,N_7791,N_7427);
nand U12686 (N_12686,N_7159,N_7345);
nor U12687 (N_12687,N_9391,N_7630);
and U12688 (N_12688,N_6223,N_9838);
nor U12689 (N_12689,N_6056,N_6000);
nor U12690 (N_12690,N_6651,N_7651);
and U12691 (N_12691,N_7633,N_5946);
nor U12692 (N_12692,N_7141,N_9204);
nor U12693 (N_12693,N_8331,N_8918);
nand U12694 (N_12694,N_5119,N_7079);
xnor U12695 (N_12695,N_6156,N_5412);
nand U12696 (N_12696,N_7226,N_7686);
nand U12697 (N_12697,N_9196,N_7632);
xnor U12698 (N_12698,N_5542,N_7421);
nand U12699 (N_12699,N_7110,N_9356);
nor U12700 (N_12700,N_7114,N_5687);
nand U12701 (N_12701,N_9734,N_6537);
nor U12702 (N_12702,N_6981,N_5672);
nor U12703 (N_12703,N_6452,N_9085);
nor U12704 (N_12704,N_6189,N_9692);
xnor U12705 (N_12705,N_8544,N_6412);
or U12706 (N_12706,N_8887,N_7845);
nand U12707 (N_12707,N_9148,N_6874);
nor U12708 (N_12708,N_5224,N_5624);
or U12709 (N_12709,N_5730,N_8334);
or U12710 (N_12710,N_7592,N_5167);
and U12711 (N_12711,N_9564,N_9331);
nand U12712 (N_12712,N_8081,N_7494);
and U12713 (N_12713,N_9040,N_5765);
nand U12714 (N_12714,N_5730,N_5164);
nand U12715 (N_12715,N_6007,N_6816);
and U12716 (N_12716,N_5913,N_8585);
and U12717 (N_12717,N_6234,N_6548);
nor U12718 (N_12718,N_8635,N_7770);
nand U12719 (N_12719,N_8856,N_6302);
or U12720 (N_12720,N_8294,N_5668);
nand U12721 (N_12721,N_5274,N_6359);
nor U12722 (N_12722,N_6362,N_6724);
nor U12723 (N_12723,N_8073,N_6116);
nor U12724 (N_12724,N_5420,N_7011);
nor U12725 (N_12725,N_6191,N_7010);
xnor U12726 (N_12726,N_8536,N_8930);
nand U12727 (N_12727,N_7911,N_8258);
nand U12728 (N_12728,N_9053,N_9525);
nand U12729 (N_12729,N_8396,N_8296);
nor U12730 (N_12730,N_6871,N_6527);
or U12731 (N_12731,N_6004,N_9759);
xor U12732 (N_12732,N_7124,N_9597);
nand U12733 (N_12733,N_6553,N_8370);
nand U12734 (N_12734,N_8871,N_8517);
and U12735 (N_12735,N_6220,N_7162);
nor U12736 (N_12736,N_6070,N_6270);
or U12737 (N_12737,N_7186,N_6426);
nand U12738 (N_12738,N_9079,N_9043);
or U12739 (N_12739,N_8947,N_7747);
and U12740 (N_12740,N_5260,N_6596);
xor U12741 (N_12741,N_6569,N_7388);
or U12742 (N_12742,N_7433,N_8546);
xor U12743 (N_12743,N_8055,N_8040);
and U12744 (N_12744,N_8706,N_9687);
nand U12745 (N_12745,N_8796,N_9401);
and U12746 (N_12746,N_7432,N_7848);
nor U12747 (N_12747,N_6336,N_5554);
or U12748 (N_12748,N_9872,N_5947);
xor U12749 (N_12749,N_9252,N_7729);
xnor U12750 (N_12750,N_8810,N_7111);
or U12751 (N_12751,N_9211,N_8031);
nor U12752 (N_12752,N_5485,N_8051);
nand U12753 (N_12753,N_9483,N_6568);
nand U12754 (N_12754,N_5250,N_7393);
or U12755 (N_12755,N_9088,N_9392);
nor U12756 (N_12756,N_5912,N_9891);
xor U12757 (N_12757,N_8960,N_5569);
and U12758 (N_12758,N_8639,N_7913);
and U12759 (N_12759,N_8137,N_8083);
and U12760 (N_12760,N_9899,N_5935);
or U12761 (N_12761,N_7098,N_9097);
xor U12762 (N_12762,N_8253,N_9113);
and U12763 (N_12763,N_7807,N_6589);
and U12764 (N_12764,N_7432,N_8544);
or U12765 (N_12765,N_9900,N_9145);
and U12766 (N_12766,N_5062,N_5007);
nand U12767 (N_12767,N_6072,N_7775);
xor U12768 (N_12768,N_9895,N_8218);
or U12769 (N_12769,N_5176,N_5065);
nand U12770 (N_12770,N_8160,N_6405);
and U12771 (N_12771,N_8285,N_5009);
nor U12772 (N_12772,N_6180,N_5433);
xnor U12773 (N_12773,N_9417,N_8831);
xor U12774 (N_12774,N_7074,N_6500);
or U12775 (N_12775,N_7300,N_7035);
xor U12776 (N_12776,N_7977,N_5126);
nand U12777 (N_12777,N_9982,N_8738);
nand U12778 (N_12778,N_6857,N_7586);
and U12779 (N_12779,N_5364,N_8690);
or U12780 (N_12780,N_9539,N_6720);
and U12781 (N_12781,N_8563,N_5828);
or U12782 (N_12782,N_5302,N_7314);
or U12783 (N_12783,N_7701,N_6883);
xnor U12784 (N_12784,N_8639,N_5262);
xor U12785 (N_12785,N_5886,N_5306);
or U12786 (N_12786,N_7007,N_9896);
nand U12787 (N_12787,N_6247,N_5438);
nand U12788 (N_12788,N_6089,N_8827);
nor U12789 (N_12789,N_8419,N_6924);
or U12790 (N_12790,N_7479,N_9465);
xnor U12791 (N_12791,N_6816,N_7751);
nand U12792 (N_12792,N_7972,N_5792);
nand U12793 (N_12793,N_6675,N_9349);
xnor U12794 (N_12794,N_6648,N_5668);
nor U12795 (N_12795,N_9101,N_5722);
nand U12796 (N_12796,N_6097,N_9222);
or U12797 (N_12797,N_6279,N_9834);
nand U12798 (N_12798,N_7566,N_6315);
or U12799 (N_12799,N_9962,N_7292);
or U12800 (N_12800,N_9293,N_6056);
nand U12801 (N_12801,N_7556,N_7664);
nand U12802 (N_12802,N_5781,N_8400);
nor U12803 (N_12803,N_6240,N_7313);
nand U12804 (N_12804,N_9484,N_9157);
or U12805 (N_12805,N_9616,N_5130);
or U12806 (N_12806,N_8825,N_6889);
or U12807 (N_12807,N_5667,N_7172);
nand U12808 (N_12808,N_8508,N_9951);
nor U12809 (N_12809,N_5041,N_9463);
nand U12810 (N_12810,N_5248,N_5752);
nor U12811 (N_12811,N_8569,N_5932);
xnor U12812 (N_12812,N_9338,N_7105);
and U12813 (N_12813,N_9787,N_9591);
and U12814 (N_12814,N_8372,N_7961);
xor U12815 (N_12815,N_9997,N_9645);
xor U12816 (N_12816,N_8579,N_9385);
nor U12817 (N_12817,N_9975,N_6641);
nor U12818 (N_12818,N_7947,N_8377);
nor U12819 (N_12819,N_5427,N_8952);
or U12820 (N_12820,N_5934,N_8713);
nor U12821 (N_12821,N_7302,N_9401);
nand U12822 (N_12822,N_8984,N_9521);
nand U12823 (N_12823,N_5480,N_6959);
xnor U12824 (N_12824,N_6138,N_8035);
or U12825 (N_12825,N_6118,N_7803);
xor U12826 (N_12826,N_9983,N_7390);
and U12827 (N_12827,N_8385,N_6916);
xor U12828 (N_12828,N_8986,N_8197);
or U12829 (N_12829,N_8530,N_5509);
nor U12830 (N_12830,N_5286,N_9756);
and U12831 (N_12831,N_9276,N_7042);
nor U12832 (N_12832,N_9680,N_6491);
nand U12833 (N_12833,N_8174,N_7314);
nand U12834 (N_12834,N_7645,N_7410);
nor U12835 (N_12835,N_9660,N_6225);
xor U12836 (N_12836,N_9041,N_6909);
or U12837 (N_12837,N_9994,N_5090);
or U12838 (N_12838,N_7862,N_7863);
and U12839 (N_12839,N_7518,N_7382);
nor U12840 (N_12840,N_8786,N_5681);
nor U12841 (N_12841,N_7168,N_6396);
xnor U12842 (N_12842,N_7780,N_8798);
xnor U12843 (N_12843,N_5274,N_9050);
nor U12844 (N_12844,N_5264,N_6309);
and U12845 (N_12845,N_7855,N_8566);
nor U12846 (N_12846,N_5489,N_8926);
nand U12847 (N_12847,N_9049,N_9620);
xnor U12848 (N_12848,N_8167,N_5579);
and U12849 (N_12849,N_7522,N_9459);
nor U12850 (N_12850,N_8965,N_7961);
and U12851 (N_12851,N_7906,N_8321);
nor U12852 (N_12852,N_5584,N_7417);
nand U12853 (N_12853,N_9133,N_8875);
nand U12854 (N_12854,N_5321,N_8341);
and U12855 (N_12855,N_7373,N_6094);
and U12856 (N_12856,N_9824,N_8406);
and U12857 (N_12857,N_5224,N_8892);
or U12858 (N_12858,N_9672,N_8135);
nor U12859 (N_12859,N_9813,N_5120);
nor U12860 (N_12860,N_6318,N_6492);
or U12861 (N_12861,N_6359,N_5884);
and U12862 (N_12862,N_8368,N_8742);
or U12863 (N_12863,N_7159,N_5168);
and U12864 (N_12864,N_6570,N_7439);
xnor U12865 (N_12865,N_6908,N_5404);
or U12866 (N_12866,N_5762,N_8166);
xnor U12867 (N_12867,N_8005,N_7049);
or U12868 (N_12868,N_5919,N_7354);
xor U12869 (N_12869,N_6956,N_7649);
xnor U12870 (N_12870,N_8403,N_7004);
nand U12871 (N_12871,N_7546,N_8313);
nand U12872 (N_12872,N_6473,N_8759);
or U12873 (N_12873,N_5509,N_7887);
nand U12874 (N_12874,N_9922,N_7999);
xor U12875 (N_12875,N_6736,N_7265);
nand U12876 (N_12876,N_8013,N_7582);
and U12877 (N_12877,N_8088,N_8049);
or U12878 (N_12878,N_9051,N_7655);
xor U12879 (N_12879,N_6538,N_6055);
nor U12880 (N_12880,N_5933,N_6189);
nand U12881 (N_12881,N_8942,N_5051);
or U12882 (N_12882,N_8691,N_5491);
xnor U12883 (N_12883,N_9018,N_7375);
and U12884 (N_12884,N_6710,N_6659);
or U12885 (N_12885,N_5182,N_6672);
nand U12886 (N_12886,N_6533,N_8062);
or U12887 (N_12887,N_8993,N_7808);
nor U12888 (N_12888,N_7274,N_9393);
and U12889 (N_12889,N_9061,N_6021);
and U12890 (N_12890,N_7998,N_8764);
nand U12891 (N_12891,N_9267,N_6928);
nand U12892 (N_12892,N_5779,N_9753);
nand U12893 (N_12893,N_6207,N_6436);
nand U12894 (N_12894,N_7049,N_6242);
or U12895 (N_12895,N_9565,N_8840);
nor U12896 (N_12896,N_9454,N_7351);
nor U12897 (N_12897,N_8798,N_5382);
xnor U12898 (N_12898,N_9075,N_9803);
or U12899 (N_12899,N_7971,N_8212);
or U12900 (N_12900,N_8941,N_6108);
nand U12901 (N_12901,N_5956,N_9790);
xnor U12902 (N_12902,N_5002,N_7398);
and U12903 (N_12903,N_8748,N_6729);
nor U12904 (N_12904,N_9999,N_9688);
or U12905 (N_12905,N_7156,N_9684);
and U12906 (N_12906,N_9159,N_6462);
and U12907 (N_12907,N_7717,N_8186);
and U12908 (N_12908,N_9886,N_7769);
and U12909 (N_12909,N_7971,N_8383);
nor U12910 (N_12910,N_5268,N_8366);
nand U12911 (N_12911,N_8879,N_8743);
nand U12912 (N_12912,N_7600,N_6481);
nor U12913 (N_12913,N_7814,N_6707);
or U12914 (N_12914,N_9164,N_8188);
or U12915 (N_12915,N_5632,N_9849);
xnor U12916 (N_12916,N_9981,N_6646);
nand U12917 (N_12917,N_6350,N_9935);
nor U12918 (N_12918,N_7219,N_9445);
or U12919 (N_12919,N_6794,N_9513);
or U12920 (N_12920,N_8946,N_8216);
nor U12921 (N_12921,N_6838,N_6849);
and U12922 (N_12922,N_9019,N_9602);
and U12923 (N_12923,N_5687,N_9613);
and U12924 (N_12924,N_6890,N_7242);
xor U12925 (N_12925,N_8606,N_7851);
or U12926 (N_12926,N_6082,N_6971);
and U12927 (N_12927,N_9480,N_6212);
xor U12928 (N_12928,N_5705,N_8819);
nand U12929 (N_12929,N_8402,N_5271);
and U12930 (N_12930,N_6581,N_8567);
nand U12931 (N_12931,N_7996,N_9952);
xnor U12932 (N_12932,N_5679,N_5334);
nand U12933 (N_12933,N_5323,N_7229);
nand U12934 (N_12934,N_9125,N_5493);
xnor U12935 (N_12935,N_5092,N_5706);
and U12936 (N_12936,N_5693,N_6142);
and U12937 (N_12937,N_9663,N_6137);
and U12938 (N_12938,N_6791,N_5000);
xnor U12939 (N_12939,N_7891,N_7300);
or U12940 (N_12940,N_9964,N_9330);
nand U12941 (N_12941,N_8321,N_6029);
or U12942 (N_12942,N_9601,N_9599);
xnor U12943 (N_12943,N_9441,N_9687);
and U12944 (N_12944,N_6317,N_8963);
nand U12945 (N_12945,N_6068,N_7229);
xor U12946 (N_12946,N_6790,N_9267);
and U12947 (N_12947,N_6960,N_5977);
or U12948 (N_12948,N_6989,N_9930);
and U12949 (N_12949,N_9754,N_6890);
nor U12950 (N_12950,N_8926,N_6183);
or U12951 (N_12951,N_7539,N_7018);
xor U12952 (N_12952,N_7669,N_9349);
xor U12953 (N_12953,N_6264,N_9687);
xor U12954 (N_12954,N_5346,N_9919);
nand U12955 (N_12955,N_7122,N_5772);
and U12956 (N_12956,N_7746,N_5798);
and U12957 (N_12957,N_6298,N_7801);
nand U12958 (N_12958,N_8187,N_7255);
or U12959 (N_12959,N_5040,N_7640);
xnor U12960 (N_12960,N_8881,N_5679);
and U12961 (N_12961,N_9999,N_9076);
xnor U12962 (N_12962,N_8512,N_6239);
nand U12963 (N_12963,N_5477,N_7171);
or U12964 (N_12964,N_6240,N_8069);
xnor U12965 (N_12965,N_9782,N_6940);
and U12966 (N_12966,N_8330,N_6907);
nand U12967 (N_12967,N_5306,N_6221);
nand U12968 (N_12968,N_9986,N_7995);
xor U12969 (N_12969,N_8483,N_7748);
or U12970 (N_12970,N_8580,N_8942);
and U12971 (N_12971,N_7917,N_9565);
or U12972 (N_12972,N_8789,N_9199);
nor U12973 (N_12973,N_9084,N_6293);
nor U12974 (N_12974,N_9655,N_6130);
nor U12975 (N_12975,N_9133,N_8410);
xnor U12976 (N_12976,N_6259,N_5644);
nor U12977 (N_12977,N_5789,N_8157);
nand U12978 (N_12978,N_5084,N_8576);
and U12979 (N_12979,N_6367,N_9860);
nor U12980 (N_12980,N_5578,N_5770);
nand U12981 (N_12981,N_6636,N_6920);
or U12982 (N_12982,N_8019,N_5782);
nand U12983 (N_12983,N_5144,N_7273);
xor U12984 (N_12984,N_8326,N_7350);
and U12985 (N_12985,N_6362,N_8725);
nor U12986 (N_12986,N_6594,N_7768);
nand U12987 (N_12987,N_6490,N_8106);
nand U12988 (N_12988,N_9989,N_8842);
nor U12989 (N_12989,N_6380,N_8634);
xor U12990 (N_12990,N_5506,N_5685);
nand U12991 (N_12991,N_9105,N_9988);
or U12992 (N_12992,N_9891,N_8726);
or U12993 (N_12993,N_5743,N_8375);
or U12994 (N_12994,N_5023,N_9547);
xnor U12995 (N_12995,N_6435,N_8817);
and U12996 (N_12996,N_7543,N_7667);
or U12997 (N_12997,N_6091,N_6101);
nor U12998 (N_12998,N_9562,N_6689);
xor U12999 (N_12999,N_9298,N_6053);
and U13000 (N_13000,N_9096,N_7788);
nor U13001 (N_13001,N_5870,N_5663);
nand U13002 (N_13002,N_9164,N_9424);
xor U13003 (N_13003,N_8770,N_8501);
nor U13004 (N_13004,N_5986,N_5866);
and U13005 (N_13005,N_5649,N_8351);
or U13006 (N_13006,N_8598,N_5484);
and U13007 (N_13007,N_5966,N_7703);
nor U13008 (N_13008,N_9256,N_6500);
or U13009 (N_13009,N_7026,N_9328);
and U13010 (N_13010,N_7193,N_6883);
nand U13011 (N_13011,N_7321,N_5991);
and U13012 (N_13012,N_5423,N_8296);
or U13013 (N_13013,N_8498,N_6170);
nor U13014 (N_13014,N_9363,N_6347);
or U13015 (N_13015,N_9676,N_6959);
nor U13016 (N_13016,N_6156,N_6219);
and U13017 (N_13017,N_9724,N_5080);
nand U13018 (N_13018,N_5194,N_6061);
or U13019 (N_13019,N_5398,N_9219);
nor U13020 (N_13020,N_7127,N_5325);
xnor U13021 (N_13021,N_5848,N_8525);
xor U13022 (N_13022,N_6538,N_7869);
or U13023 (N_13023,N_6939,N_5747);
xnor U13024 (N_13024,N_7564,N_9517);
or U13025 (N_13025,N_9340,N_8164);
xor U13026 (N_13026,N_9463,N_7282);
and U13027 (N_13027,N_9609,N_6074);
or U13028 (N_13028,N_9007,N_8155);
nand U13029 (N_13029,N_9645,N_9923);
nand U13030 (N_13030,N_9341,N_8255);
xor U13031 (N_13031,N_9325,N_7238);
and U13032 (N_13032,N_6277,N_5270);
xor U13033 (N_13033,N_7107,N_9952);
and U13034 (N_13034,N_9098,N_6740);
and U13035 (N_13035,N_7381,N_8155);
nand U13036 (N_13036,N_9881,N_5781);
and U13037 (N_13037,N_8207,N_8273);
and U13038 (N_13038,N_6030,N_5431);
or U13039 (N_13039,N_9534,N_7961);
and U13040 (N_13040,N_6763,N_9218);
nor U13041 (N_13041,N_9162,N_9614);
or U13042 (N_13042,N_7720,N_5194);
nand U13043 (N_13043,N_7489,N_6267);
xor U13044 (N_13044,N_5293,N_6362);
nor U13045 (N_13045,N_7515,N_8950);
nand U13046 (N_13046,N_5307,N_5884);
xnor U13047 (N_13047,N_5033,N_5713);
nand U13048 (N_13048,N_9576,N_6861);
or U13049 (N_13049,N_9862,N_7464);
and U13050 (N_13050,N_5507,N_9371);
nand U13051 (N_13051,N_7772,N_5153);
nor U13052 (N_13052,N_6557,N_9458);
nand U13053 (N_13053,N_8943,N_7740);
xnor U13054 (N_13054,N_6884,N_5803);
nor U13055 (N_13055,N_6967,N_7390);
xnor U13056 (N_13056,N_5149,N_5745);
nor U13057 (N_13057,N_5085,N_9804);
nand U13058 (N_13058,N_9033,N_9912);
nor U13059 (N_13059,N_5290,N_7903);
or U13060 (N_13060,N_8995,N_5186);
xor U13061 (N_13061,N_6929,N_7481);
and U13062 (N_13062,N_7299,N_9323);
or U13063 (N_13063,N_7443,N_6567);
nand U13064 (N_13064,N_6822,N_5041);
nor U13065 (N_13065,N_9897,N_6166);
xnor U13066 (N_13066,N_5618,N_8446);
and U13067 (N_13067,N_8628,N_8934);
xor U13068 (N_13068,N_9169,N_7985);
nand U13069 (N_13069,N_9986,N_5594);
and U13070 (N_13070,N_6273,N_7405);
or U13071 (N_13071,N_7646,N_6319);
xor U13072 (N_13072,N_7462,N_9082);
xor U13073 (N_13073,N_9790,N_9871);
or U13074 (N_13074,N_6353,N_8658);
nand U13075 (N_13075,N_5174,N_8591);
nor U13076 (N_13076,N_7798,N_9800);
nor U13077 (N_13077,N_9977,N_8723);
and U13078 (N_13078,N_9505,N_8256);
or U13079 (N_13079,N_7290,N_8217);
and U13080 (N_13080,N_8837,N_7227);
and U13081 (N_13081,N_6844,N_5801);
nand U13082 (N_13082,N_7835,N_6387);
or U13083 (N_13083,N_8828,N_9362);
or U13084 (N_13084,N_8472,N_5354);
xnor U13085 (N_13085,N_7931,N_7958);
or U13086 (N_13086,N_7777,N_6783);
and U13087 (N_13087,N_6285,N_6551);
xnor U13088 (N_13088,N_8066,N_9698);
nand U13089 (N_13089,N_7236,N_5566);
and U13090 (N_13090,N_5640,N_8077);
nor U13091 (N_13091,N_9222,N_7895);
nor U13092 (N_13092,N_7431,N_6407);
nor U13093 (N_13093,N_7248,N_5032);
and U13094 (N_13094,N_6872,N_7093);
nor U13095 (N_13095,N_7716,N_8448);
and U13096 (N_13096,N_9081,N_6475);
and U13097 (N_13097,N_9242,N_8042);
xnor U13098 (N_13098,N_9886,N_8835);
and U13099 (N_13099,N_5393,N_6525);
nor U13100 (N_13100,N_5671,N_5130);
nor U13101 (N_13101,N_7770,N_7521);
nand U13102 (N_13102,N_9615,N_9656);
nand U13103 (N_13103,N_6074,N_8471);
nor U13104 (N_13104,N_9059,N_5321);
xnor U13105 (N_13105,N_8581,N_5696);
and U13106 (N_13106,N_9824,N_5781);
xor U13107 (N_13107,N_9706,N_6517);
nor U13108 (N_13108,N_9228,N_8225);
and U13109 (N_13109,N_8203,N_9988);
nand U13110 (N_13110,N_7111,N_8894);
or U13111 (N_13111,N_7652,N_9622);
or U13112 (N_13112,N_5994,N_5012);
or U13113 (N_13113,N_8494,N_7140);
nor U13114 (N_13114,N_9764,N_6649);
and U13115 (N_13115,N_7937,N_9020);
xnor U13116 (N_13116,N_6108,N_7720);
and U13117 (N_13117,N_6311,N_8655);
xor U13118 (N_13118,N_8798,N_7302);
and U13119 (N_13119,N_6051,N_8146);
or U13120 (N_13120,N_5914,N_7429);
nand U13121 (N_13121,N_6407,N_9831);
or U13122 (N_13122,N_7815,N_6957);
xor U13123 (N_13123,N_6466,N_7465);
or U13124 (N_13124,N_7043,N_9325);
and U13125 (N_13125,N_8840,N_5527);
or U13126 (N_13126,N_6896,N_7839);
or U13127 (N_13127,N_6341,N_5265);
xnor U13128 (N_13128,N_6823,N_8456);
nand U13129 (N_13129,N_6245,N_5194);
and U13130 (N_13130,N_9445,N_7036);
xnor U13131 (N_13131,N_9374,N_9207);
xnor U13132 (N_13132,N_8882,N_5928);
xnor U13133 (N_13133,N_6818,N_7124);
xor U13134 (N_13134,N_6541,N_5096);
and U13135 (N_13135,N_5567,N_9490);
and U13136 (N_13136,N_9652,N_6329);
xnor U13137 (N_13137,N_8915,N_9090);
xor U13138 (N_13138,N_5682,N_9774);
nand U13139 (N_13139,N_6444,N_8339);
or U13140 (N_13140,N_9786,N_5370);
xor U13141 (N_13141,N_7973,N_7764);
and U13142 (N_13142,N_5853,N_7319);
nor U13143 (N_13143,N_8800,N_5602);
xor U13144 (N_13144,N_7480,N_6037);
xor U13145 (N_13145,N_7128,N_7186);
nand U13146 (N_13146,N_8268,N_9798);
and U13147 (N_13147,N_8653,N_8992);
nor U13148 (N_13148,N_5083,N_5325);
nor U13149 (N_13149,N_5140,N_6792);
and U13150 (N_13150,N_7843,N_9849);
and U13151 (N_13151,N_7242,N_5264);
xor U13152 (N_13152,N_7691,N_5037);
or U13153 (N_13153,N_5519,N_8367);
and U13154 (N_13154,N_7230,N_6782);
nand U13155 (N_13155,N_5485,N_8891);
nand U13156 (N_13156,N_6666,N_8289);
nor U13157 (N_13157,N_8745,N_8754);
nand U13158 (N_13158,N_7058,N_6692);
and U13159 (N_13159,N_7744,N_9792);
xor U13160 (N_13160,N_6251,N_9718);
nand U13161 (N_13161,N_7466,N_8963);
and U13162 (N_13162,N_5558,N_5568);
xor U13163 (N_13163,N_7590,N_8137);
nor U13164 (N_13164,N_8029,N_7747);
nor U13165 (N_13165,N_9332,N_8267);
or U13166 (N_13166,N_5946,N_8641);
nor U13167 (N_13167,N_8514,N_5475);
or U13168 (N_13168,N_6872,N_7855);
xor U13169 (N_13169,N_9489,N_7845);
nand U13170 (N_13170,N_6400,N_6030);
and U13171 (N_13171,N_6306,N_8148);
or U13172 (N_13172,N_9588,N_8563);
or U13173 (N_13173,N_7020,N_6497);
and U13174 (N_13174,N_9606,N_8095);
nor U13175 (N_13175,N_5574,N_7090);
xor U13176 (N_13176,N_9461,N_9840);
and U13177 (N_13177,N_5208,N_6120);
or U13178 (N_13178,N_5180,N_5208);
and U13179 (N_13179,N_6760,N_7447);
nor U13180 (N_13180,N_6252,N_6739);
and U13181 (N_13181,N_7194,N_8884);
and U13182 (N_13182,N_9284,N_8900);
or U13183 (N_13183,N_8032,N_7676);
nand U13184 (N_13184,N_7638,N_7079);
nand U13185 (N_13185,N_9965,N_6579);
xor U13186 (N_13186,N_7052,N_9318);
and U13187 (N_13187,N_6247,N_9850);
and U13188 (N_13188,N_9780,N_5783);
and U13189 (N_13189,N_7379,N_6932);
nand U13190 (N_13190,N_7374,N_6105);
xor U13191 (N_13191,N_8950,N_9054);
and U13192 (N_13192,N_8498,N_8960);
xnor U13193 (N_13193,N_6408,N_6530);
and U13194 (N_13194,N_7348,N_7759);
or U13195 (N_13195,N_5246,N_7832);
nand U13196 (N_13196,N_5526,N_5035);
xnor U13197 (N_13197,N_5315,N_8744);
nand U13198 (N_13198,N_8787,N_9360);
nand U13199 (N_13199,N_7211,N_9996);
nand U13200 (N_13200,N_7583,N_7833);
or U13201 (N_13201,N_9935,N_5021);
nor U13202 (N_13202,N_5384,N_6057);
or U13203 (N_13203,N_8497,N_6546);
nand U13204 (N_13204,N_5917,N_8678);
nand U13205 (N_13205,N_8870,N_5232);
xor U13206 (N_13206,N_5108,N_6786);
and U13207 (N_13207,N_5499,N_9530);
xnor U13208 (N_13208,N_7577,N_5208);
xnor U13209 (N_13209,N_9563,N_7773);
and U13210 (N_13210,N_5967,N_9633);
or U13211 (N_13211,N_7384,N_5787);
and U13212 (N_13212,N_6260,N_9355);
xnor U13213 (N_13213,N_5051,N_6693);
nor U13214 (N_13214,N_5958,N_6707);
or U13215 (N_13215,N_8251,N_5549);
and U13216 (N_13216,N_8109,N_6543);
or U13217 (N_13217,N_6645,N_7559);
and U13218 (N_13218,N_6669,N_9573);
or U13219 (N_13219,N_5995,N_5906);
nor U13220 (N_13220,N_6526,N_6928);
nand U13221 (N_13221,N_8236,N_9891);
or U13222 (N_13222,N_9351,N_7196);
nor U13223 (N_13223,N_5950,N_9252);
nor U13224 (N_13224,N_5444,N_7824);
nand U13225 (N_13225,N_9295,N_6525);
or U13226 (N_13226,N_7664,N_6446);
xor U13227 (N_13227,N_8453,N_8375);
xor U13228 (N_13228,N_8364,N_7957);
nand U13229 (N_13229,N_7725,N_7338);
and U13230 (N_13230,N_5937,N_7700);
and U13231 (N_13231,N_8825,N_6235);
xnor U13232 (N_13232,N_9861,N_9678);
or U13233 (N_13233,N_7945,N_8727);
nand U13234 (N_13234,N_8691,N_8719);
nor U13235 (N_13235,N_8907,N_9520);
and U13236 (N_13236,N_7540,N_9697);
nor U13237 (N_13237,N_5020,N_5473);
or U13238 (N_13238,N_6509,N_7565);
and U13239 (N_13239,N_8498,N_6265);
nand U13240 (N_13240,N_6852,N_9944);
or U13241 (N_13241,N_7779,N_8901);
xnor U13242 (N_13242,N_6709,N_8070);
nand U13243 (N_13243,N_5727,N_6532);
xnor U13244 (N_13244,N_7369,N_7165);
nand U13245 (N_13245,N_7670,N_6279);
xor U13246 (N_13246,N_9985,N_5324);
nor U13247 (N_13247,N_8814,N_8458);
nor U13248 (N_13248,N_5929,N_7430);
or U13249 (N_13249,N_9178,N_6217);
nor U13250 (N_13250,N_6276,N_9715);
xor U13251 (N_13251,N_5383,N_9304);
nor U13252 (N_13252,N_8857,N_8466);
or U13253 (N_13253,N_8108,N_9059);
xor U13254 (N_13254,N_9968,N_7109);
and U13255 (N_13255,N_8603,N_5086);
nor U13256 (N_13256,N_6663,N_7396);
or U13257 (N_13257,N_6606,N_7568);
and U13258 (N_13258,N_6243,N_6111);
xnor U13259 (N_13259,N_5935,N_9850);
nor U13260 (N_13260,N_8692,N_7633);
nand U13261 (N_13261,N_8737,N_6636);
xnor U13262 (N_13262,N_9083,N_8857);
or U13263 (N_13263,N_6420,N_5213);
nor U13264 (N_13264,N_7061,N_9729);
xor U13265 (N_13265,N_6098,N_6922);
nand U13266 (N_13266,N_5109,N_8185);
and U13267 (N_13267,N_6110,N_8379);
xnor U13268 (N_13268,N_8555,N_5099);
nor U13269 (N_13269,N_6563,N_7465);
xnor U13270 (N_13270,N_9570,N_9912);
and U13271 (N_13271,N_7395,N_5825);
or U13272 (N_13272,N_6463,N_8985);
or U13273 (N_13273,N_5084,N_5216);
nor U13274 (N_13274,N_8412,N_7022);
and U13275 (N_13275,N_6720,N_7899);
xor U13276 (N_13276,N_8912,N_9250);
xor U13277 (N_13277,N_7151,N_9114);
nand U13278 (N_13278,N_9759,N_9456);
nand U13279 (N_13279,N_8122,N_8154);
nand U13280 (N_13280,N_6249,N_9174);
or U13281 (N_13281,N_8688,N_8087);
or U13282 (N_13282,N_9939,N_8123);
or U13283 (N_13283,N_7499,N_6078);
nor U13284 (N_13284,N_8326,N_9775);
or U13285 (N_13285,N_5510,N_7711);
xnor U13286 (N_13286,N_5704,N_9947);
or U13287 (N_13287,N_8101,N_6508);
and U13288 (N_13288,N_8215,N_6902);
xor U13289 (N_13289,N_9756,N_7755);
xnor U13290 (N_13290,N_5262,N_6430);
xnor U13291 (N_13291,N_9015,N_7057);
xor U13292 (N_13292,N_9507,N_6744);
and U13293 (N_13293,N_5126,N_9594);
nand U13294 (N_13294,N_5242,N_7144);
nor U13295 (N_13295,N_7389,N_8684);
or U13296 (N_13296,N_5624,N_9080);
or U13297 (N_13297,N_8885,N_7587);
nor U13298 (N_13298,N_9865,N_7101);
xnor U13299 (N_13299,N_7803,N_7929);
nand U13300 (N_13300,N_6577,N_9081);
nor U13301 (N_13301,N_7819,N_7729);
nand U13302 (N_13302,N_9032,N_9884);
xnor U13303 (N_13303,N_6414,N_7468);
xor U13304 (N_13304,N_6463,N_7022);
nor U13305 (N_13305,N_9646,N_8962);
nor U13306 (N_13306,N_6495,N_5732);
and U13307 (N_13307,N_5604,N_8390);
nor U13308 (N_13308,N_6014,N_5820);
xnor U13309 (N_13309,N_5786,N_5370);
or U13310 (N_13310,N_6675,N_8675);
nand U13311 (N_13311,N_7056,N_6725);
nor U13312 (N_13312,N_6484,N_7682);
and U13313 (N_13313,N_5846,N_5718);
xnor U13314 (N_13314,N_6416,N_5833);
nand U13315 (N_13315,N_8020,N_5248);
xor U13316 (N_13316,N_6918,N_9221);
nor U13317 (N_13317,N_8416,N_5227);
and U13318 (N_13318,N_6321,N_7919);
xor U13319 (N_13319,N_5582,N_9729);
and U13320 (N_13320,N_8862,N_5601);
xor U13321 (N_13321,N_5748,N_7377);
or U13322 (N_13322,N_9828,N_7000);
nand U13323 (N_13323,N_9492,N_6320);
nor U13324 (N_13324,N_9556,N_9467);
nand U13325 (N_13325,N_9916,N_7122);
nand U13326 (N_13326,N_5648,N_6972);
or U13327 (N_13327,N_6566,N_7954);
nand U13328 (N_13328,N_8629,N_8676);
nor U13329 (N_13329,N_8715,N_6382);
and U13330 (N_13330,N_7172,N_5527);
or U13331 (N_13331,N_8002,N_7164);
nand U13332 (N_13332,N_6450,N_9965);
nor U13333 (N_13333,N_7098,N_9055);
xnor U13334 (N_13334,N_7951,N_9603);
or U13335 (N_13335,N_6920,N_6753);
xnor U13336 (N_13336,N_5457,N_9401);
nand U13337 (N_13337,N_5537,N_5944);
nand U13338 (N_13338,N_7453,N_6381);
nor U13339 (N_13339,N_6620,N_7945);
nor U13340 (N_13340,N_9202,N_5238);
and U13341 (N_13341,N_7484,N_8189);
nor U13342 (N_13342,N_6252,N_8919);
nand U13343 (N_13343,N_8489,N_9537);
and U13344 (N_13344,N_7554,N_8554);
nand U13345 (N_13345,N_6252,N_7385);
or U13346 (N_13346,N_9127,N_5595);
nand U13347 (N_13347,N_9663,N_9132);
or U13348 (N_13348,N_8348,N_8418);
nand U13349 (N_13349,N_6658,N_5874);
nor U13350 (N_13350,N_5544,N_5717);
and U13351 (N_13351,N_6466,N_9351);
xor U13352 (N_13352,N_8679,N_6117);
and U13353 (N_13353,N_8155,N_6568);
or U13354 (N_13354,N_9699,N_6155);
nand U13355 (N_13355,N_7918,N_6200);
nor U13356 (N_13356,N_7331,N_9288);
or U13357 (N_13357,N_6948,N_5874);
xor U13358 (N_13358,N_7277,N_8859);
or U13359 (N_13359,N_8408,N_8012);
xnor U13360 (N_13360,N_6142,N_9991);
and U13361 (N_13361,N_6102,N_5195);
nand U13362 (N_13362,N_8564,N_6485);
nand U13363 (N_13363,N_9378,N_5761);
or U13364 (N_13364,N_5731,N_6599);
and U13365 (N_13365,N_7868,N_5354);
nor U13366 (N_13366,N_5580,N_5401);
nand U13367 (N_13367,N_5094,N_5425);
nor U13368 (N_13368,N_5452,N_8693);
xnor U13369 (N_13369,N_6504,N_7716);
xnor U13370 (N_13370,N_6256,N_6056);
xor U13371 (N_13371,N_9332,N_9033);
or U13372 (N_13372,N_7638,N_8279);
xnor U13373 (N_13373,N_5033,N_9813);
xor U13374 (N_13374,N_8936,N_9835);
xnor U13375 (N_13375,N_8124,N_5930);
xnor U13376 (N_13376,N_6247,N_5650);
and U13377 (N_13377,N_9057,N_6344);
and U13378 (N_13378,N_8822,N_5245);
nand U13379 (N_13379,N_7685,N_8854);
nand U13380 (N_13380,N_7380,N_8982);
or U13381 (N_13381,N_6802,N_6714);
xnor U13382 (N_13382,N_7285,N_6290);
or U13383 (N_13383,N_9065,N_6747);
and U13384 (N_13384,N_5419,N_6217);
nor U13385 (N_13385,N_6534,N_6656);
xnor U13386 (N_13386,N_6489,N_5348);
or U13387 (N_13387,N_5513,N_6168);
xor U13388 (N_13388,N_6169,N_7784);
nand U13389 (N_13389,N_9938,N_7299);
nor U13390 (N_13390,N_9212,N_7157);
nor U13391 (N_13391,N_5356,N_6254);
or U13392 (N_13392,N_7267,N_9954);
and U13393 (N_13393,N_7218,N_6136);
or U13394 (N_13394,N_8404,N_5455);
xnor U13395 (N_13395,N_5049,N_9441);
nand U13396 (N_13396,N_7945,N_5962);
or U13397 (N_13397,N_6807,N_6757);
nand U13398 (N_13398,N_5517,N_8953);
xor U13399 (N_13399,N_9252,N_5772);
or U13400 (N_13400,N_9345,N_7752);
nor U13401 (N_13401,N_5488,N_9418);
nand U13402 (N_13402,N_9459,N_6520);
and U13403 (N_13403,N_9575,N_5244);
and U13404 (N_13404,N_5978,N_6666);
and U13405 (N_13405,N_9170,N_7295);
or U13406 (N_13406,N_5101,N_5274);
nand U13407 (N_13407,N_9595,N_6851);
nor U13408 (N_13408,N_5917,N_8302);
nand U13409 (N_13409,N_6209,N_9775);
and U13410 (N_13410,N_7598,N_5421);
or U13411 (N_13411,N_8335,N_6002);
nor U13412 (N_13412,N_5103,N_8024);
nand U13413 (N_13413,N_7359,N_6744);
nor U13414 (N_13414,N_5728,N_5516);
and U13415 (N_13415,N_5338,N_5014);
and U13416 (N_13416,N_5866,N_5141);
nor U13417 (N_13417,N_6813,N_5497);
nand U13418 (N_13418,N_7398,N_8472);
or U13419 (N_13419,N_7336,N_5301);
and U13420 (N_13420,N_5421,N_6977);
or U13421 (N_13421,N_9432,N_5886);
nand U13422 (N_13422,N_7419,N_8067);
and U13423 (N_13423,N_6503,N_5826);
and U13424 (N_13424,N_9084,N_8489);
nor U13425 (N_13425,N_5157,N_5890);
and U13426 (N_13426,N_5027,N_9704);
nand U13427 (N_13427,N_7586,N_8100);
nand U13428 (N_13428,N_9784,N_6797);
nor U13429 (N_13429,N_8539,N_5045);
xnor U13430 (N_13430,N_8612,N_8923);
or U13431 (N_13431,N_8717,N_6395);
or U13432 (N_13432,N_8814,N_7845);
nand U13433 (N_13433,N_5011,N_8802);
nand U13434 (N_13434,N_5192,N_8652);
or U13435 (N_13435,N_7860,N_6730);
or U13436 (N_13436,N_7370,N_8332);
and U13437 (N_13437,N_8814,N_5873);
xnor U13438 (N_13438,N_9156,N_7788);
nand U13439 (N_13439,N_8753,N_7749);
nand U13440 (N_13440,N_5824,N_8732);
xor U13441 (N_13441,N_6413,N_9017);
or U13442 (N_13442,N_6403,N_5984);
xor U13443 (N_13443,N_9318,N_5848);
xor U13444 (N_13444,N_6149,N_5169);
and U13445 (N_13445,N_8327,N_8101);
xor U13446 (N_13446,N_5986,N_9790);
nor U13447 (N_13447,N_6208,N_8622);
xnor U13448 (N_13448,N_6362,N_9055);
nor U13449 (N_13449,N_7073,N_5997);
xnor U13450 (N_13450,N_6184,N_7039);
xor U13451 (N_13451,N_5421,N_8836);
nor U13452 (N_13452,N_7487,N_7897);
nor U13453 (N_13453,N_8758,N_8900);
nand U13454 (N_13454,N_9668,N_6660);
and U13455 (N_13455,N_8524,N_7341);
nor U13456 (N_13456,N_5822,N_7474);
nor U13457 (N_13457,N_8938,N_8215);
xnor U13458 (N_13458,N_8808,N_7934);
xor U13459 (N_13459,N_9493,N_7396);
and U13460 (N_13460,N_6481,N_5406);
or U13461 (N_13461,N_7117,N_7135);
or U13462 (N_13462,N_8525,N_7241);
nor U13463 (N_13463,N_5953,N_7041);
or U13464 (N_13464,N_9830,N_9608);
and U13465 (N_13465,N_8167,N_5020);
nor U13466 (N_13466,N_8985,N_6271);
nand U13467 (N_13467,N_6306,N_5661);
nand U13468 (N_13468,N_5354,N_6080);
nand U13469 (N_13469,N_7915,N_6561);
nor U13470 (N_13470,N_8955,N_8818);
and U13471 (N_13471,N_9361,N_7798);
nand U13472 (N_13472,N_5870,N_6239);
xor U13473 (N_13473,N_8975,N_9715);
nor U13474 (N_13474,N_7018,N_7363);
nor U13475 (N_13475,N_7659,N_7159);
or U13476 (N_13476,N_9129,N_7054);
or U13477 (N_13477,N_9040,N_7154);
nand U13478 (N_13478,N_5096,N_7436);
nand U13479 (N_13479,N_9156,N_9118);
and U13480 (N_13480,N_8337,N_6843);
or U13481 (N_13481,N_7142,N_9906);
nand U13482 (N_13482,N_7059,N_7713);
xnor U13483 (N_13483,N_7252,N_8082);
or U13484 (N_13484,N_7165,N_7924);
and U13485 (N_13485,N_8655,N_8673);
or U13486 (N_13486,N_6709,N_9995);
nor U13487 (N_13487,N_7404,N_8922);
nand U13488 (N_13488,N_5022,N_7888);
nor U13489 (N_13489,N_8964,N_6252);
nand U13490 (N_13490,N_8332,N_8983);
nand U13491 (N_13491,N_6244,N_9656);
nand U13492 (N_13492,N_9508,N_5458);
and U13493 (N_13493,N_8217,N_8507);
nand U13494 (N_13494,N_5927,N_6472);
nand U13495 (N_13495,N_6582,N_6425);
or U13496 (N_13496,N_5312,N_9511);
nor U13497 (N_13497,N_6577,N_7357);
or U13498 (N_13498,N_5137,N_8544);
and U13499 (N_13499,N_9824,N_6348);
or U13500 (N_13500,N_9124,N_9354);
and U13501 (N_13501,N_5610,N_8576);
nand U13502 (N_13502,N_9131,N_6936);
nand U13503 (N_13503,N_6802,N_9810);
xnor U13504 (N_13504,N_5279,N_6337);
nand U13505 (N_13505,N_5556,N_6367);
nand U13506 (N_13506,N_8052,N_5891);
and U13507 (N_13507,N_5522,N_5697);
or U13508 (N_13508,N_5996,N_6268);
xor U13509 (N_13509,N_6763,N_9145);
xnor U13510 (N_13510,N_9180,N_9333);
and U13511 (N_13511,N_9314,N_7029);
xnor U13512 (N_13512,N_8120,N_5913);
and U13513 (N_13513,N_5641,N_9739);
nand U13514 (N_13514,N_9831,N_8427);
xnor U13515 (N_13515,N_9270,N_5867);
or U13516 (N_13516,N_9486,N_7368);
xor U13517 (N_13517,N_8370,N_5404);
nand U13518 (N_13518,N_8238,N_8850);
nand U13519 (N_13519,N_8311,N_5772);
nor U13520 (N_13520,N_8037,N_8438);
or U13521 (N_13521,N_8958,N_9649);
nand U13522 (N_13522,N_9615,N_6038);
or U13523 (N_13523,N_9372,N_5505);
xor U13524 (N_13524,N_6782,N_8630);
nor U13525 (N_13525,N_9150,N_6772);
and U13526 (N_13526,N_8791,N_5578);
and U13527 (N_13527,N_6409,N_9698);
nor U13528 (N_13528,N_5699,N_9432);
nand U13529 (N_13529,N_7147,N_8264);
or U13530 (N_13530,N_8787,N_5581);
nor U13531 (N_13531,N_6863,N_5502);
nand U13532 (N_13532,N_5734,N_9738);
or U13533 (N_13533,N_9971,N_5775);
nand U13534 (N_13534,N_5008,N_5297);
xor U13535 (N_13535,N_8453,N_7824);
or U13536 (N_13536,N_9583,N_5056);
and U13537 (N_13537,N_8675,N_7015);
nor U13538 (N_13538,N_7983,N_5832);
and U13539 (N_13539,N_6106,N_8603);
nand U13540 (N_13540,N_6727,N_7972);
xor U13541 (N_13541,N_9006,N_7098);
nor U13542 (N_13542,N_7897,N_7064);
nor U13543 (N_13543,N_7193,N_7241);
or U13544 (N_13544,N_7872,N_9894);
xnor U13545 (N_13545,N_7424,N_7578);
nor U13546 (N_13546,N_7029,N_9651);
and U13547 (N_13547,N_8021,N_9925);
and U13548 (N_13548,N_5982,N_7601);
nor U13549 (N_13549,N_6950,N_7408);
and U13550 (N_13550,N_7744,N_9759);
xnor U13551 (N_13551,N_9259,N_6568);
nand U13552 (N_13552,N_6307,N_7055);
and U13553 (N_13553,N_6231,N_9022);
or U13554 (N_13554,N_8991,N_6555);
nor U13555 (N_13555,N_5048,N_9044);
nand U13556 (N_13556,N_5474,N_9296);
xnor U13557 (N_13557,N_7545,N_8685);
xnor U13558 (N_13558,N_5962,N_6942);
xor U13559 (N_13559,N_9119,N_6576);
or U13560 (N_13560,N_5803,N_6702);
nand U13561 (N_13561,N_9531,N_6122);
xor U13562 (N_13562,N_7942,N_8468);
nor U13563 (N_13563,N_5109,N_6373);
nor U13564 (N_13564,N_8489,N_6050);
nor U13565 (N_13565,N_9250,N_5373);
nand U13566 (N_13566,N_7849,N_7047);
xor U13567 (N_13567,N_5731,N_9469);
xor U13568 (N_13568,N_7873,N_7732);
nand U13569 (N_13569,N_8658,N_8360);
xnor U13570 (N_13570,N_8118,N_8145);
and U13571 (N_13571,N_8917,N_7693);
or U13572 (N_13572,N_6248,N_9384);
and U13573 (N_13573,N_5707,N_6079);
or U13574 (N_13574,N_6523,N_9489);
or U13575 (N_13575,N_9913,N_9610);
or U13576 (N_13576,N_5521,N_5199);
nand U13577 (N_13577,N_9902,N_6106);
xor U13578 (N_13578,N_9181,N_8788);
and U13579 (N_13579,N_5436,N_8362);
or U13580 (N_13580,N_5506,N_8349);
nand U13581 (N_13581,N_8737,N_6768);
or U13582 (N_13582,N_9877,N_7552);
or U13583 (N_13583,N_6167,N_6871);
and U13584 (N_13584,N_7355,N_9217);
xor U13585 (N_13585,N_7892,N_5302);
nand U13586 (N_13586,N_8514,N_7415);
and U13587 (N_13587,N_9855,N_5911);
xnor U13588 (N_13588,N_8556,N_9598);
nor U13589 (N_13589,N_5962,N_7689);
and U13590 (N_13590,N_7683,N_8988);
and U13591 (N_13591,N_8929,N_7677);
nand U13592 (N_13592,N_7419,N_6797);
xor U13593 (N_13593,N_7435,N_7464);
xor U13594 (N_13594,N_8782,N_5348);
or U13595 (N_13595,N_7191,N_8119);
and U13596 (N_13596,N_7649,N_5001);
nor U13597 (N_13597,N_7602,N_8817);
xnor U13598 (N_13598,N_9131,N_9947);
or U13599 (N_13599,N_6990,N_7525);
and U13600 (N_13600,N_8915,N_9709);
and U13601 (N_13601,N_5660,N_5245);
nor U13602 (N_13602,N_6427,N_5444);
xnor U13603 (N_13603,N_9326,N_8482);
or U13604 (N_13604,N_7212,N_7940);
and U13605 (N_13605,N_9242,N_8798);
nand U13606 (N_13606,N_6490,N_9300);
or U13607 (N_13607,N_6513,N_5941);
nor U13608 (N_13608,N_7621,N_8412);
xnor U13609 (N_13609,N_8702,N_7749);
nor U13610 (N_13610,N_9234,N_5258);
and U13611 (N_13611,N_8002,N_8513);
and U13612 (N_13612,N_7449,N_7847);
nor U13613 (N_13613,N_7217,N_6446);
and U13614 (N_13614,N_5202,N_9336);
xnor U13615 (N_13615,N_6723,N_8666);
or U13616 (N_13616,N_7458,N_5282);
nand U13617 (N_13617,N_5706,N_9330);
xnor U13618 (N_13618,N_5354,N_8436);
xor U13619 (N_13619,N_9804,N_5795);
xnor U13620 (N_13620,N_7823,N_6681);
xnor U13621 (N_13621,N_5423,N_8598);
xnor U13622 (N_13622,N_5714,N_8135);
and U13623 (N_13623,N_8365,N_9468);
or U13624 (N_13624,N_8915,N_6069);
xnor U13625 (N_13625,N_7366,N_9021);
nand U13626 (N_13626,N_9862,N_7342);
or U13627 (N_13627,N_7738,N_9991);
nand U13628 (N_13628,N_8914,N_9510);
or U13629 (N_13629,N_9559,N_8581);
and U13630 (N_13630,N_8864,N_7643);
or U13631 (N_13631,N_8368,N_7041);
or U13632 (N_13632,N_8416,N_8143);
or U13633 (N_13633,N_7969,N_5590);
nand U13634 (N_13634,N_7719,N_9998);
or U13635 (N_13635,N_8268,N_5079);
xor U13636 (N_13636,N_6266,N_6187);
nor U13637 (N_13637,N_7484,N_7892);
or U13638 (N_13638,N_8579,N_9668);
nand U13639 (N_13639,N_9676,N_6043);
nand U13640 (N_13640,N_5606,N_5478);
nor U13641 (N_13641,N_6208,N_8982);
and U13642 (N_13642,N_8948,N_7169);
nor U13643 (N_13643,N_6528,N_9335);
nand U13644 (N_13644,N_9020,N_7052);
or U13645 (N_13645,N_9095,N_8096);
nor U13646 (N_13646,N_7085,N_8902);
or U13647 (N_13647,N_6534,N_9764);
or U13648 (N_13648,N_7606,N_6489);
and U13649 (N_13649,N_9395,N_8472);
or U13650 (N_13650,N_9214,N_8895);
nor U13651 (N_13651,N_5681,N_9586);
xnor U13652 (N_13652,N_6720,N_6428);
and U13653 (N_13653,N_9466,N_5149);
nor U13654 (N_13654,N_6011,N_7751);
nor U13655 (N_13655,N_7375,N_8206);
and U13656 (N_13656,N_6928,N_9412);
and U13657 (N_13657,N_7048,N_9286);
or U13658 (N_13658,N_7930,N_9282);
and U13659 (N_13659,N_8370,N_5714);
and U13660 (N_13660,N_7220,N_9716);
xnor U13661 (N_13661,N_7247,N_5267);
or U13662 (N_13662,N_5251,N_5598);
nor U13663 (N_13663,N_5797,N_5478);
xnor U13664 (N_13664,N_5878,N_9346);
nor U13665 (N_13665,N_6659,N_5755);
xnor U13666 (N_13666,N_5671,N_7299);
or U13667 (N_13667,N_5966,N_9890);
or U13668 (N_13668,N_5107,N_6200);
nand U13669 (N_13669,N_6569,N_7721);
nand U13670 (N_13670,N_9865,N_5229);
nor U13671 (N_13671,N_6487,N_8289);
xnor U13672 (N_13672,N_5054,N_6999);
nor U13673 (N_13673,N_6448,N_9335);
nand U13674 (N_13674,N_5897,N_6916);
or U13675 (N_13675,N_6664,N_8805);
xnor U13676 (N_13676,N_9990,N_8859);
and U13677 (N_13677,N_5675,N_6173);
nand U13678 (N_13678,N_6657,N_6632);
and U13679 (N_13679,N_7505,N_7219);
nand U13680 (N_13680,N_7553,N_9026);
nand U13681 (N_13681,N_9541,N_5918);
nor U13682 (N_13682,N_7756,N_8823);
or U13683 (N_13683,N_7259,N_5206);
nor U13684 (N_13684,N_5826,N_9102);
or U13685 (N_13685,N_7408,N_7580);
nor U13686 (N_13686,N_6460,N_6703);
xor U13687 (N_13687,N_9423,N_7581);
nor U13688 (N_13688,N_7913,N_5550);
xnor U13689 (N_13689,N_5935,N_7367);
xnor U13690 (N_13690,N_7620,N_9197);
and U13691 (N_13691,N_9728,N_9264);
or U13692 (N_13692,N_5855,N_5355);
nor U13693 (N_13693,N_6293,N_6417);
nor U13694 (N_13694,N_6291,N_8753);
and U13695 (N_13695,N_7563,N_8983);
nor U13696 (N_13696,N_7869,N_7347);
and U13697 (N_13697,N_5276,N_8425);
nand U13698 (N_13698,N_5785,N_6538);
or U13699 (N_13699,N_6824,N_8460);
and U13700 (N_13700,N_8552,N_8601);
nor U13701 (N_13701,N_9586,N_5794);
xnor U13702 (N_13702,N_7448,N_7652);
and U13703 (N_13703,N_5109,N_5250);
nor U13704 (N_13704,N_8354,N_8278);
xor U13705 (N_13705,N_8316,N_9813);
or U13706 (N_13706,N_8657,N_5605);
xor U13707 (N_13707,N_6545,N_5334);
nand U13708 (N_13708,N_6721,N_6673);
xnor U13709 (N_13709,N_7072,N_6846);
xor U13710 (N_13710,N_9883,N_8157);
and U13711 (N_13711,N_6862,N_6740);
nand U13712 (N_13712,N_7395,N_7820);
and U13713 (N_13713,N_6668,N_5594);
and U13714 (N_13714,N_8959,N_6916);
nor U13715 (N_13715,N_6224,N_7231);
xnor U13716 (N_13716,N_9366,N_8243);
nor U13717 (N_13717,N_7742,N_8442);
and U13718 (N_13718,N_6927,N_5283);
and U13719 (N_13719,N_9127,N_5768);
xnor U13720 (N_13720,N_8365,N_9740);
and U13721 (N_13721,N_7823,N_5682);
nor U13722 (N_13722,N_9982,N_8901);
nand U13723 (N_13723,N_6087,N_5420);
nand U13724 (N_13724,N_6168,N_5252);
or U13725 (N_13725,N_9510,N_9460);
and U13726 (N_13726,N_7930,N_9244);
nor U13727 (N_13727,N_9899,N_7935);
or U13728 (N_13728,N_7425,N_8558);
nand U13729 (N_13729,N_8525,N_7167);
or U13730 (N_13730,N_6280,N_9951);
nor U13731 (N_13731,N_7855,N_7762);
nor U13732 (N_13732,N_7224,N_5592);
or U13733 (N_13733,N_8913,N_8645);
or U13734 (N_13734,N_8480,N_6158);
or U13735 (N_13735,N_7196,N_5435);
nor U13736 (N_13736,N_8721,N_9796);
and U13737 (N_13737,N_8791,N_5870);
xor U13738 (N_13738,N_9003,N_8728);
nor U13739 (N_13739,N_8129,N_7001);
nor U13740 (N_13740,N_8640,N_6524);
nand U13741 (N_13741,N_6638,N_6454);
and U13742 (N_13742,N_6352,N_5393);
or U13743 (N_13743,N_9130,N_7196);
xor U13744 (N_13744,N_5542,N_8363);
nor U13745 (N_13745,N_9341,N_6749);
nor U13746 (N_13746,N_7674,N_9162);
nor U13747 (N_13747,N_5325,N_5078);
or U13748 (N_13748,N_8893,N_9196);
nand U13749 (N_13749,N_8022,N_5207);
nor U13750 (N_13750,N_5266,N_8118);
nand U13751 (N_13751,N_8906,N_8626);
xor U13752 (N_13752,N_9339,N_9178);
xnor U13753 (N_13753,N_6917,N_7597);
or U13754 (N_13754,N_5828,N_5024);
xnor U13755 (N_13755,N_6844,N_8589);
xnor U13756 (N_13756,N_6356,N_6894);
nor U13757 (N_13757,N_8894,N_8193);
xnor U13758 (N_13758,N_8122,N_9518);
or U13759 (N_13759,N_9234,N_5395);
nor U13760 (N_13760,N_7465,N_6628);
xnor U13761 (N_13761,N_5944,N_8931);
xnor U13762 (N_13762,N_7323,N_8592);
nor U13763 (N_13763,N_9822,N_7136);
or U13764 (N_13764,N_9998,N_9997);
and U13765 (N_13765,N_5752,N_6901);
and U13766 (N_13766,N_8089,N_8460);
nand U13767 (N_13767,N_8757,N_9592);
and U13768 (N_13768,N_6590,N_5468);
nand U13769 (N_13769,N_9815,N_5987);
or U13770 (N_13770,N_5943,N_7513);
nand U13771 (N_13771,N_7427,N_6638);
and U13772 (N_13772,N_9353,N_7084);
or U13773 (N_13773,N_8724,N_8923);
nand U13774 (N_13774,N_7273,N_8324);
or U13775 (N_13775,N_8593,N_6187);
or U13776 (N_13776,N_7170,N_7735);
and U13777 (N_13777,N_7121,N_5065);
xor U13778 (N_13778,N_8623,N_5583);
nand U13779 (N_13779,N_9363,N_8387);
or U13780 (N_13780,N_5324,N_9280);
or U13781 (N_13781,N_5326,N_5301);
xnor U13782 (N_13782,N_7617,N_9874);
xor U13783 (N_13783,N_5561,N_7388);
or U13784 (N_13784,N_8525,N_9096);
xnor U13785 (N_13785,N_6127,N_8103);
xnor U13786 (N_13786,N_9979,N_5758);
xnor U13787 (N_13787,N_7299,N_6336);
xnor U13788 (N_13788,N_7085,N_7198);
nand U13789 (N_13789,N_9015,N_5894);
or U13790 (N_13790,N_5571,N_6896);
xor U13791 (N_13791,N_8373,N_6187);
xnor U13792 (N_13792,N_7808,N_6819);
nand U13793 (N_13793,N_9762,N_7120);
xnor U13794 (N_13794,N_9936,N_8857);
xnor U13795 (N_13795,N_5620,N_6293);
and U13796 (N_13796,N_6549,N_6755);
and U13797 (N_13797,N_7264,N_8089);
or U13798 (N_13798,N_5552,N_7479);
and U13799 (N_13799,N_9376,N_8020);
or U13800 (N_13800,N_7750,N_5704);
xor U13801 (N_13801,N_7944,N_8148);
and U13802 (N_13802,N_9395,N_9941);
and U13803 (N_13803,N_7356,N_6286);
xnor U13804 (N_13804,N_9373,N_7970);
and U13805 (N_13805,N_5948,N_7408);
xnor U13806 (N_13806,N_6066,N_7626);
nand U13807 (N_13807,N_8191,N_7384);
nor U13808 (N_13808,N_7412,N_6649);
xnor U13809 (N_13809,N_5016,N_9223);
and U13810 (N_13810,N_6850,N_5674);
nand U13811 (N_13811,N_9799,N_7012);
nor U13812 (N_13812,N_6517,N_7933);
and U13813 (N_13813,N_8610,N_8952);
nor U13814 (N_13814,N_5541,N_7765);
or U13815 (N_13815,N_9020,N_8416);
nor U13816 (N_13816,N_8261,N_8872);
nor U13817 (N_13817,N_8223,N_7950);
and U13818 (N_13818,N_8047,N_8500);
nor U13819 (N_13819,N_5025,N_7322);
xnor U13820 (N_13820,N_9547,N_8366);
xnor U13821 (N_13821,N_5609,N_8896);
nand U13822 (N_13822,N_9297,N_9526);
and U13823 (N_13823,N_7158,N_7956);
nor U13824 (N_13824,N_8657,N_7589);
xor U13825 (N_13825,N_6996,N_7089);
xor U13826 (N_13826,N_7032,N_6955);
nor U13827 (N_13827,N_8925,N_8452);
nor U13828 (N_13828,N_9916,N_6060);
nor U13829 (N_13829,N_8357,N_9408);
nor U13830 (N_13830,N_6375,N_9426);
nand U13831 (N_13831,N_7463,N_9985);
nor U13832 (N_13832,N_5485,N_5283);
nand U13833 (N_13833,N_7055,N_7408);
or U13834 (N_13834,N_6045,N_6178);
xor U13835 (N_13835,N_8393,N_8353);
nor U13836 (N_13836,N_8776,N_7210);
and U13837 (N_13837,N_5312,N_8553);
nand U13838 (N_13838,N_9326,N_5383);
xnor U13839 (N_13839,N_5661,N_8844);
xnor U13840 (N_13840,N_6893,N_7427);
nand U13841 (N_13841,N_9683,N_7265);
nand U13842 (N_13842,N_5987,N_6959);
nor U13843 (N_13843,N_5442,N_5081);
nand U13844 (N_13844,N_6754,N_9501);
or U13845 (N_13845,N_5448,N_7006);
or U13846 (N_13846,N_9717,N_8607);
nor U13847 (N_13847,N_9663,N_6539);
nor U13848 (N_13848,N_9505,N_7286);
or U13849 (N_13849,N_7394,N_9539);
nor U13850 (N_13850,N_9505,N_6995);
or U13851 (N_13851,N_8086,N_7420);
nand U13852 (N_13852,N_8793,N_8498);
xnor U13853 (N_13853,N_9318,N_8616);
nor U13854 (N_13854,N_8607,N_9000);
xor U13855 (N_13855,N_8551,N_5180);
xnor U13856 (N_13856,N_7117,N_9577);
or U13857 (N_13857,N_5247,N_5917);
and U13858 (N_13858,N_7746,N_5336);
or U13859 (N_13859,N_7314,N_5657);
nor U13860 (N_13860,N_7878,N_5232);
nand U13861 (N_13861,N_8301,N_7957);
and U13862 (N_13862,N_6153,N_5513);
nor U13863 (N_13863,N_5244,N_9566);
or U13864 (N_13864,N_8245,N_5196);
or U13865 (N_13865,N_6081,N_6124);
nor U13866 (N_13866,N_5784,N_8722);
or U13867 (N_13867,N_5143,N_9840);
nor U13868 (N_13868,N_8031,N_9371);
and U13869 (N_13869,N_9002,N_6777);
nor U13870 (N_13870,N_8609,N_8385);
nand U13871 (N_13871,N_5554,N_5890);
nand U13872 (N_13872,N_9019,N_6009);
nor U13873 (N_13873,N_9412,N_5022);
or U13874 (N_13874,N_9024,N_9393);
or U13875 (N_13875,N_5303,N_6214);
xnor U13876 (N_13876,N_6826,N_6396);
and U13877 (N_13877,N_5506,N_5944);
nor U13878 (N_13878,N_7993,N_7916);
and U13879 (N_13879,N_7264,N_6319);
or U13880 (N_13880,N_5543,N_6135);
nor U13881 (N_13881,N_9427,N_7587);
xor U13882 (N_13882,N_5302,N_7482);
xnor U13883 (N_13883,N_6912,N_7117);
nand U13884 (N_13884,N_7859,N_8375);
nand U13885 (N_13885,N_8856,N_7020);
nor U13886 (N_13886,N_6484,N_8913);
or U13887 (N_13887,N_9657,N_7438);
nor U13888 (N_13888,N_5267,N_6059);
nand U13889 (N_13889,N_5025,N_6856);
nor U13890 (N_13890,N_5272,N_6465);
or U13891 (N_13891,N_5629,N_8903);
or U13892 (N_13892,N_9516,N_8821);
xor U13893 (N_13893,N_8895,N_5504);
or U13894 (N_13894,N_9268,N_6862);
or U13895 (N_13895,N_6172,N_5523);
xnor U13896 (N_13896,N_6421,N_9862);
or U13897 (N_13897,N_9113,N_9615);
or U13898 (N_13898,N_9920,N_5985);
nor U13899 (N_13899,N_6587,N_8379);
xor U13900 (N_13900,N_7065,N_9803);
or U13901 (N_13901,N_8157,N_8190);
and U13902 (N_13902,N_8476,N_5698);
and U13903 (N_13903,N_9652,N_7075);
and U13904 (N_13904,N_9081,N_5552);
and U13905 (N_13905,N_8012,N_5400);
nor U13906 (N_13906,N_8723,N_8471);
xnor U13907 (N_13907,N_8569,N_6555);
nor U13908 (N_13908,N_9075,N_7523);
xnor U13909 (N_13909,N_6943,N_9128);
or U13910 (N_13910,N_9959,N_8124);
xnor U13911 (N_13911,N_8759,N_7006);
nand U13912 (N_13912,N_8654,N_5384);
nor U13913 (N_13913,N_5763,N_9523);
or U13914 (N_13914,N_9777,N_7597);
and U13915 (N_13915,N_7035,N_8565);
xor U13916 (N_13916,N_5302,N_9991);
nor U13917 (N_13917,N_6768,N_8607);
nand U13918 (N_13918,N_9414,N_5274);
or U13919 (N_13919,N_5416,N_9038);
and U13920 (N_13920,N_6095,N_7531);
nor U13921 (N_13921,N_7812,N_6567);
or U13922 (N_13922,N_9408,N_6773);
or U13923 (N_13923,N_5823,N_9703);
xnor U13924 (N_13924,N_5652,N_7892);
xor U13925 (N_13925,N_8904,N_5850);
nand U13926 (N_13926,N_8229,N_9363);
xor U13927 (N_13927,N_9403,N_6783);
nor U13928 (N_13928,N_7780,N_9270);
or U13929 (N_13929,N_5661,N_6318);
nand U13930 (N_13930,N_7490,N_7563);
or U13931 (N_13931,N_7302,N_5124);
and U13932 (N_13932,N_5104,N_5411);
xor U13933 (N_13933,N_9016,N_6736);
nor U13934 (N_13934,N_7265,N_7773);
xor U13935 (N_13935,N_6770,N_6013);
nor U13936 (N_13936,N_9473,N_8530);
xnor U13937 (N_13937,N_5574,N_6993);
nor U13938 (N_13938,N_7000,N_7393);
or U13939 (N_13939,N_9661,N_6669);
nor U13940 (N_13940,N_5636,N_5094);
xnor U13941 (N_13941,N_5750,N_8857);
xor U13942 (N_13942,N_5816,N_6936);
xor U13943 (N_13943,N_8252,N_7919);
xor U13944 (N_13944,N_5382,N_6731);
nand U13945 (N_13945,N_5817,N_7193);
xor U13946 (N_13946,N_6885,N_6732);
or U13947 (N_13947,N_8874,N_9785);
xor U13948 (N_13948,N_5343,N_7239);
nand U13949 (N_13949,N_7426,N_7109);
nor U13950 (N_13950,N_8903,N_5591);
nand U13951 (N_13951,N_9755,N_5230);
nor U13952 (N_13952,N_9918,N_8305);
nor U13953 (N_13953,N_7900,N_7058);
and U13954 (N_13954,N_6779,N_7422);
xor U13955 (N_13955,N_5468,N_9897);
xnor U13956 (N_13956,N_9730,N_5147);
xor U13957 (N_13957,N_8902,N_8955);
nand U13958 (N_13958,N_9218,N_8084);
nor U13959 (N_13959,N_5697,N_6488);
and U13960 (N_13960,N_9295,N_6158);
xnor U13961 (N_13961,N_5477,N_6642);
and U13962 (N_13962,N_9279,N_6263);
xor U13963 (N_13963,N_8124,N_8036);
and U13964 (N_13964,N_9339,N_8358);
xor U13965 (N_13965,N_8138,N_8998);
nand U13966 (N_13966,N_9376,N_9595);
nand U13967 (N_13967,N_7920,N_8963);
or U13968 (N_13968,N_8174,N_9355);
xnor U13969 (N_13969,N_5265,N_5301);
and U13970 (N_13970,N_7775,N_8358);
and U13971 (N_13971,N_7356,N_6178);
or U13972 (N_13972,N_5725,N_9151);
or U13973 (N_13973,N_5848,N_7950);
nand U13974 (N_13974,N_9733,N_9671);
or U13975 (N_13975,N_8010,N_5431);
or U13976 (N_13976,N_8126,N_9200);
nor U13977 (N_13977,N_6308,N_8039);
nand U13978 (N_13978,N_6558,N_8184);
or U13979 (N_13979,N_6172,N_7148);
nand U13980 (N_13980,N_6192,N_9983);
or U13981 (N_13981,N_8556,N_8903);
nor U13982 (N_13982,N_5204,N_7650);
or U13983 (N_13983,N_5130,N_5060);
or U13984 (N_13984,N_7585,N_5794);
and U13985 (N_13985,N_8619,N_7973);
nor U13986 (N_13986,N_5980,N_8467);
and U13987 (N_13987,N_8678,N_5396);
and U13988 (N_13988,N_9796,N_8141);
and U13989 (N_13989,N_6402,N_6610);
nor U13990 (N_13990,N_6544,N_5699);
nand U13991 (N_13991,N_6854,N_5028);
and U13992 (N_13992,N_8076,N_6607);
or U13993 (N_13993,N_8604,N_8731);
and U13994 (N_13994,N_6652,N_8716);
or U13995 (N_13995,N_5493,N_5429);
nand U13996 (N_13996,N_6074,N_7008);
or U13997 (N_13997,N_8510,N_5837);
xnor U13998 (N_13998,N_8548,N_5962);
nor U13999 (N_13999,N_7446,N_8268);
or U14000 (N_14000,N_8471,N_7944);
xnor U14001 (N_14001,N_9680,N_8600);
xnor U14002 (N_14002,N_8450,N_6452);
or U14003 (N_14003,N_6226,N_8019);
or U14004 (N_14004,N_8256,N_6933);
and U14005 (N_14005,N_5145,N_5000);
nor U14006 (N_14006,N_9889,N_5562);
xnor U14007 (N_14007,N_7102,N_9918);
nand U14008 (N_14008,N_9655,N_8575);
and U14009 (N_14009,N_8981,N_8458);
nand U14010 (N_14010,N_6279,N_9721);
nor U14011 (N_14011,N_8705,N_9428);
xnor U14012 (N_14012,N_8073,N_6113);
or U14013 (N_14013,N_9172,N_9946);
or U14014 (N_14014,N_7248,N_9438);
or U14015 (N_14015,N_6918,N_9974);
xor U14016 (N_14016,N_8313,N_7839);
xor U14017 (N_14017,N_8437,N_7869);
nand U14018 (N_14018,N_9701,N_6847);
or U14019 (N_14019,N_9851,N_9808);
nor U14020 (N_14020,N_5846,N_6317);
nor U14021 (N_14021,N_5554,N_9076);
nor U14022 (N_14022,N_6391,N_7602);
xor U14023 (N_14023,N_9510,N_5417);
or U14024 (N_14024,N_5488,N_9067);
xor U14025 (N_14025,N_5969,N_8823);
nor U14026 (N_14026,N_8284,N_8797);
xnor U14027 (N_14027,N_5085,N_7808);
and U14028 (N_14028,N_5562,N_8235);
nand U14029 (N_14029,N_6057,N_6118);
nor U14030 (N_14030,N_9693,N_9466);
nand U14031 (N_14031,N_7289,N_5318);
xor U14032 (N_14032,N_7505,N_7723);
nand U14033 (N_14033,N_5088,N_5008);
or U14034 (N_14034,N_6979,N_5641);
nor U14035 (N_14035,N_8265,N_9648);
and U14036 (N_14036,N_8270,N_9087);
or U14037 (N_14037,N_7399,N_7116);
nand U14038 (N_14038,N_5169,N_7132);
or U14039 (N_14039,N_6042,N_8715);
or U14040 (N_14040,N_6752,N_5201);
nor U14041 (N_14041,N_9262,N_9080);
xnor U14042 (N_14042,N_5233,N_6037);
and U14043 (N_14043,N_5802,N_7430);
nor U14044 (N_14044,N_6736,N_6533);
xor U14045 (N_14045,N_7237,N_7632);
nor U14046 (N_14046,N_5652,N_7811);
or U14047 (N_14047,N_7904,N_5417);
xnor U14048 (N_14048,N_9075,N_5832);
or U14049 (N_14049,N_5283,N_8753);
xnor U14050 (N_14050,N_5805,N_6629);
nand U14051 (N_14051,N_8568,N_7056);
xor U14052 (N_14052,N_6293,N_5972);
or U14053 (N_14053,N_9191,N_9577);
and U14054 (N_14054,N_6460,N_7535);
nand U14055 (N_14055,N_9445,N_5389);
or U14056 (N_14056,N_8246,N_7350);
nand U14057 (N_14057,N_6059,N_7584);
nor U14058 (N_14058,N_6254,N_7126);
nor U14059 (N_14059,N_8142,N_8555);
xor U14060 (N_14060,N_6145,N_5963);
or U14061 (N_14061,N_5335,N_8612);
and U14062 (N_14062,N_5861,N_9965);
or U14063 (N_14063,N_6003,N_8441);
or U14064 (N_14064,N_6891,N_5363);
or U14065 (N_14065,N_7131,N_6860);
or U14066 (N_14066,N_7392,N_5089);
xnor U14067 (N_14067,N_5534,N_6594);
nor U14068 (N_14068,N_6367,N_7911);
nand U14069 (N_14069,N_8055,N_7289);
nand U14070 (N_14070,N_8428,N_9303);
and U14071 (N_14071,N_8415,N_9564);
xnor U14072 (N_14072,N_6991,N_7751);
or U14073 (N_14073,N_5790,N_8308);
or U14074 (N_14074,N_5865,N_5593);
nand U14075 (N_14075,N_7268,N_6419);
nand U14076 (N_14076,N_5061,N_7043);
nor U14077 (N_14077,N_9408,N_6852);
nor U14078 (N_14078,N_6055,N_5891);
xnor U14079 (N_14079,N_7390,N_9907);
xor U14080 (N_14080,N_6445,N_5537);
nand U14081 (N_14081,N_6250,N_5663);
and U14082 (N_14082,N_7188,N_8155);
xnor U14083 (N_14083,N_9105,N_5049);
nor U14084 (N_14084,N_9215,N_6242);
nor U14085 (N_14085,N_7089,N_7245);
and U14086 (N_14086,N_8660,N_9919);
and U14087 (N_14087,N_8328,N_5398);
and U14088 (N_14088,N_9023,N_6915);
xnor U14089 (N_14089,N_5434,N_7225);
or U14090 (N_14090,N_8060,N_8421);
and U14091 (N_14091,N_8681,N_9566);
nor U14092 (N_14092,N_5335,N_8448);
nand U14093 (N_14093,N_6110,N_8347);
nor U14094 (N_14094,N_7773,N_6724);
and U14095 (N_14095,N_6707,N_5581);
and U14096 (N_14096,N_8980,N_8880);
and U14097 (N_14097,N_9952,N_6132);
nor U14098 (N_14098,N_7663,N_9304);
or U14099 (N_14099,N_8860,N_7700);
and U14100 (N_14100,N_9873,N_6107);
and U14101 (N_14101,N_9353,N_9538);
xnor U14102 (N_14102,N_6476,N_8922);
nand U14103 (N_14103,N_8104,N_5127);
nand U14104 (N_14104,N_8984,N_8263);
nand U14105 (N_14105,N_9422,N_5384);
nand U14106 (N_14106,N_5528,N_9913);
and U14107 (N_14107,N_5307,N_7324);
xnor U14108 (N_14108,N_9516,N_9791);
nand U14109 (N_14109,N_6325,N_9099);
and U14110 (N_14110,N_8467,N_5435);
and U14111 (N_14111,N_9025,N_6562);
nor U14112 (N_14112,N_6172,N_8629);
nor U14113 (N_14113,N_9349,N_9117);
nor U14114 (N_14114,N_7261,N_7490);
or U14115 (N_14115,N_7780,N_9805);
nor U14116 (N_14116,N_8660,N_6427);
and U14117 (N_14117,N_5358,N_6507);
or U14118 (N_14118,N_7051,N_7055);
and U14119 (N_14119,N_8655,N_7501);
or U14120 (N_14120,N_9898,N_6286);
and U14121 (N_14121,N_6039,N_7536);
nand U14122 (N_14122,N_6049,N_6642);
and U14123 (N_14123,N_5618,N_9957);
xor U14124 (N_14124,N_9196,N_7907);
nor U14125 (N_14125,N_8817,N_7835);
nand U14126 (N_14126,N_8810,N_5018);
nor U14127 (N_14127,N_7078,N_7754);
or U14128 (N_14128,N_8479,N_5044);
and U14129 (N_14129,N_7313,N_9179);
and U14130 (N_14130,N_8411,N_7230);
nand U14131 (N_14131,N_7110,N_6004);
or U14132 (N_14132,N_9652,N_9005);
or U14133 (N_14133,N_9173,N_6803);
and U14134 (N_14134,N_7155,N_9502);
xnor U14135 (N_14135,N_6657,N_7578);
or U14136 (N_14136,N_5865,N_6489);
or U14137 (N_14137,N_5097,N_5920);
xor U14138 (N_14138,N_6057,N_9990);
nand U14139 (N_14139,N_5857,N_9197);
nor U14140 (N_14140,N_6630,N_8441);
nand U14141 (N_14141,N_6370,N_8861);
and U14142 (N_14142,N_5473,N_6550);
nand U14143 (N_14143,N_7459,N_9605);
and U14144 (N_14144,N_5556,N_5624);
nand U14145 (N_14145,N_8978,N_5355);
or U14146 (N_14146,N_5442,N_7694);
nor U14147 (N_14147,N_5681,N_5780);
nand U14148 (N_14148,N_9426,N_7865);
nand U14149 (N_14149,N_7890,N_7774);
xor U14150 (N_14150,N_9180,N_5045);
or U14151 (N_14151,N_5124,N_8605);
nand U14152 (N_14152,N_7674,N_8544);
nor U14153 (N_14153,N_6966,N_6216);
and U14154 (N_14154,N_8115,N_5774);
nand U14155 (N_14155,N_6075,N_6222);
and U14156 (N_14156,N_6356,N_6033);
nor U14157 (N_14157,N_6344,N_6156);
nor U14158 (N_14158,N_5889,N_6593);
or U14159 (N_14159,N_7893,N_6184);
or U14160 (N_14160,N_8231,N_7613);
xor U14161 (N_14161,N_7968,N_9544);
or U14162 (N_14162,N_6638,N_9296);
or U14163 (N_14163,N_7864,N_7390);
xor U14164 (N_14164,N_8155,N_6608);
xnor U14165 (N_14165,N_5587,N_8031);
and U14166 (N_14166,N_7410,N_8661);
nor U14167 (N_14167,N_5424,N_9638);
nand U14168 (N_14168,N_5587,N_9673);
nand U14169 (N_14169,N_9170,N_8081);
xor U14170 (N_14170,N_5937,N_7192);
xor U14171 (N_14171,N_6953,N_5409);
and U14172 (N_14172,N_7169,N_9057);
nor U14173 (N_14173,N_6888,N_7187);
nor U14174 (N_14174,N_7699,N_8380);
nand U14175 (N_14175,N_5940,N_7483);
nor U14176 (N_14176,N_5323,N_5478);
nand U14177 (N_14177,N_9980,N_9790);
xor U14178 (N_14178,N_8472,N_7711);
or U14179 (N_14179,N_8538,N_8568);
and U14180 (N_14180,N_7078,N_6622);
or U14181 (N_14181,N_5551,N_9270);
xor U14182 (N_14182,N_9003,N_8599);
nand U14183 (N_14183,N_9416,N_9780);
nand U14184 (N_14184,N_6564,N_7014);
or U14185 (N_14185,N_5155,N_6221);
nand U14186 (N_14186,N_6674,N_5042);
and U14187 (N_14187,N_7455,N_8890);
nand U14188 (N_14188,N_5046,N_6572);
nand U14189 (N_14189,N_8361,N_7980);
nand U14190 (N_14190,N_8834,N_5335);
or U14191 (N_14191,N_9170,N_9482);
xnor U14192 (N_14192,N_6220,N_6849);
xnor U14193 (N_14193,N_6826,N_5478);
xnor U14194 (N_14194,N_8528,N_8123);
nand U14195 (N_14195,N_9239,N_7394);
nor U14196 (N_14196,N_5764,N_7553);
and U14197 (N_14197,N_9024,N_7589);
or U14198 (N_14198,N_9417,N_8151);
nor U14199 (N_14199,N_9383,N_9930);
nor U14200 (N_14200,N_7691,N_6060);
and U14201 (N_14201,N_7486,N_6276);
and U14202 (N_14202,N_8642,N_6208);
nand U14203 (N_14203,N_9100,N_6878);
nand U14204 (N_14204,N_5605,N_7564);
or U14205 (N_14205,N_9772,N_7244);
xnor U14206 (N_14206,N_8205,N_5505);
and U14207 (N_14207,N_5881,N_5676);
or U14208 (N_14208,N_5922,N_6141);
nor U14209 (N_14209,N_5267,N_9284);
or U14210 (N_14210,N_9305,N_8030);
xnor U14211 (N_14211,N_9382,N_6981);
or U14212 (N_14212,N_7704,N_5162);
or U14213 (N_14213,N_5964,N_7365);
nor U14214 (N_14214,N_7245,N_5534);
xnor U14215 (N_14215,N_8377,N_8773);
and U14216 (N_14216,N_6517,N_7203);
and U14217 (N_14217,N_6651,N_7184);
nand U14218 (N_14218,N_6296,N_8246);
and U14219 (N_14219,N_9666,N_6424);
nor U14220 (N_14220,N_5218,N_6769);
xor U14221 (N_14221,N_9144,N_6156);
and U14222 (N_14222,N_6757,N_9576);
nor U14223 (N_14223,N_6726,N_9157);
or U14224 (N_14224,N_8172,N_7789);
nand U14225 (N_14225,N_6539,N_9987);
xor U14226 (N_14226,N_8561,N_9500);
and U14227 (N_14227,N_8173,N_6355);
nand U14228 (N_14228,N_9701,N_5674);
nand U14229 (N_14229,N_5498,N_5716);
xor U14230 (N_14230,N_7154,N_7066);
nand U14231 (N_14231,N_8237,N_7630);
or U14232 (N_14232,N_9980,N_5687);
xor U14233 (N_14233,N_5658,N_9921);
and U14234 (N_14234,N_5948,N_5483);
nor U14235 (N_14235,N_8826,N_9144);
xor U14236 (N_14236,N_6700,N_6766);
nand U14237 (N_14237,N_9011,N_9460);
nor U14238 (N_14238,N_6690,N_8811);
and U14239 (N_14239,N_8368,N_6630);
or U14240 (N_14240,N_8591,N_5598);
nand U14241 (N_14241,N_9576,N_7386);
nand U14242 (N_14242,N_6241,N_7196);
and U14243 (N_14243,N_5591,N_8657);
or U14244 (N_14244,N_6079,N_9294);
and U14245 (N_14245,N_7118,N_6563);
or U14246 (N_14246,N_5431,N_5481);
or U14247 (N_14247,N_7791,N_6568);
or U14248 (N_14248,N_6555,N_6359);
nand U14249 (N_14249,N_5329,N_9572);
and U14250 (N_14250,N_6870,N_5684);
nor U14251 (N_14251,N_8775,N_5229);
nand U14252 (N_14252,N_5765,N_7474);
or U14253 (N_14253,N_9357,N_5284);
or U14254 (N_14254,N_9637,N_8953);
nor U14255 (N_14255,N_7835,N_8236);
nor U14256 (N_14256,N_6925,N_6263);
xor U14257 (N_14257,N_5659,N_7236);
and U14258 (N_14258,N_5145,N_9622);
xor U14259 (N_14259,N_5607,N_8390);
nor U14260 (N_14260,N_9973,N_6380);
or U14261 (N_14261,N_8093,N_6577);
or U14262 (N_14262,N_7728,N_8156);
and U14263 (N_14263,N_9287,N_5411);
nor U14264 (N_14264,N_6946,N_6594);
xor U14265 (N_14265,N_6936,N_9339);
nand U14266 (N_14266,N_6226,N_5003);
or U14267 (N_14267,N_5541,N_5817);
and U14268 (N_14268,N_7281,N_9037);
xor U14269 (N_14269,N_9960,N_7613);
nor U14270 (N_14270,N_6955,N_8843);
nand U14271 (N_14271,N_9769,N_5784);
xor U14272 (N_14272,N_6249,N_8479);
nand U14273 (N_14273,N_8883,N_9539);
nor U14274 (N_14274,N_5309,N_6901);
xnor U14275 (N_14275,N_7473,N_7321);
and U14276 (N_14276,N_9496,N_7506);
and U14277 (N_14277,N_8637,N_5793);
nor U14278 (N_14278,N_6889,N_8947);
and U14279 (N_14279,N_6314,N_5060);
nor U14280 (N_14280,N_8203,N_9599);
and U14281 (N_14281,N_8122,N_6094);
xnor U14282 (N_14282,N_6547,N_8793);
and U14283 (N_14283,N_8647,N_9334);
xor U14284 (N_14284,N_6782,N_5024);
and U14285 (N_14285,N_9996,N_7856);
nor U14286 (N_14286,N_5057,N_6686);
and U14287 (N_14287,N_6291,N_9146);
xnor U14288 (N_14288,N_7717,N_7312);
and U14289 (N_14289,N_8182,N_6916);
or U14290 (N_14290,N_9518,N_8034);
xor U14291 (N_14291,N_7703,N_6337);
and U14292 (N_14292,N_8607,N_7700);
and U14293 (N_14293,N_5080,N_5949);
nor U14294 (N_14294,N_6393,N_6415);
nand U14295 (N_14295,N_6468,N_9893);
and U14296 (N_14296,N_9949,N_6747);
and U14297 (N_14297,N_7524,N_9250);
or U14298 (N_14298,N_9267,N_9332);
xnor U14299 (N_14299,N_8918,N_5403);
nor U14300 (N_14300,N_7553,N_5480);
and U14301 (N_14301,N_6286,N_5010);
or U14302 (N_14302,N_9564,N_5259);
nor U14303 (N_14303,N_5341,N_6389);
nor U14304 (N_14304,N_8028,N_6282);
or U14305 (N_14305,N_7264,N_9332);
or U14306 (N_14306,N_7555,N_8304);
xor U14307 (N_14307,N_8235,N_7070);
and U14308 (N_14308,N_9915,N_9602);
or U14309 (N_14309,N_9042,N_6100);
nand U14310 (N_14310,N_6245,N_9871);
xor U14311 (N_14311,N_7986,N_7480);
and U14312 (N_14312,N_9080,N_9118);
and U14313 (N_14313,N_5144,N_7655);
and U14314 (N_14314,N_5231,N_8679);
xnor U14315 (N_14315,N_5286,N_9445);
and U14316 (N_14316,N_8737,N_5394);
nor U14317 (N_14317,N_5418,N_5987);
and U14318 (N_14318,N_5532,N_5451);
and U14319 (N_14319,N_8306,N_5835);
nor U14320 (N_14320,N_6061,N_6428);
nand U14321 (N_14321,N_8165,N_5518);
nand U14322 (N_14322,N_7550,N_6631);
xor U14323 (N_14323,N_7905,N_9418);
or U14324 (N_14324,N_7900,N_5825);
or U14325 (N_14325,N_9657,N_6778);
nor U14326 (N_14326,N_9246,N_7660);
nand U14327 (N_14327,N_7716,N_9594);
and U14328 (N_14328,N_9605,N_8738);
xnor U14329 (N_14329,N_9084,N_7151);
xnor U14330 (N_14330,N_8892,N_5323);
or U14331 (N_14331,N_5517,N_8998);
xor U14332 (N_14332,N_5839,N_6639);
nor U14333 (N_14333,N_5350,N_7853);
nor U14334 (N_14334,N_5042,N_8390);
xor U14335 (N_14335,N_8743,N_6522);
nor U14336 (N_14336,N_9464,N_8320);
xnor U14337 (N_14337,N_7988,N_8205);
xor U14338 (N_14338,N_6895,N_6491);
or U14339 (N_14339,N_8393,N_5709);
nor U14340 (N_14340,N_7814,N_8402);
nor U14341 (N_14341,N_5202,N_5580);
or U14342 (N_14342,N_5614,N_6161);
or U14343 (N_14343,N_7545,N_8996);
and U14344 (N_14344,N_8959,N_9108);
and U14345 (N_14345,N_8744,N_8225);
xor U14346 (N_14346,N_6718,N_7150);
xnor U14347 (N_14347,N_6902,N_6667);
nand U14348 (N_14348,N_7200,N_7230);
or U14349 (N_14349,N_8295,N_7801);
and U14350 (N_14350,N_5106,N_9561);
nand U14351 (N_14351,N_7842,N_6973);
nor U14352 (N_14352,N_8679,N_7065);
nor U14353 (N_14353,N_6820,N_7812);
nor U14354 (N_14354,N_8245,N_9260);
xor U14355 (N_14355,N_5838,N_8757);
xor U14356 (N_14356,N_7693,N_6790);
or U14357 (N_14357,N_9531,N_5474);
xor U14358 (N_14358,N_5711,N_8911);
xnor U14359 (N_14359,N_6776,N_9331);
and U14360 (N_14360,N_6461,N_8297);
nor U14361 (N_14361,N_7763,N_5145);
xor U14362 (N_14362,N_7369,N_6760);
nor U14363 (N_14363,N_6460,N_6911);
nor U14364 (N_14364,N_5932,N_5281);
or U14365 (N_14365,N_5682,N_9814);
nor U14366 (N_14366,N_7418,N_6442);
or U14367 (N_14367,N_9037,N_7667);
and U14368 (N_14368,N_8854,N_7558);
nor U14369 (N_14369,N_9985,N_5424);
or U14370 (N_14370,N_5699,N_6908);
xor U14371 (N_14371,N_7025,N_5698);
nor U14372 (N_14372,N_7335,N_6530);
or U14373 (N_14373,N_9011,N_7844);
nand U14374 (N_14374,N_7758,N_9333);
or U14375 (N_14375,N_6404,N_5974);
nand U14376 (N_14376,N_7493,N_6214);
or U14377 (N_14377,N_8622,N_9753);
and U14378 (N_14378,N_7792,N_6099);
xnor U14379 (N_14379,N_5019,N_7123);
nor U14380 (N_14380,N_9201,N_5997);
nor U14381 (N_14381,N_6646,N_5218);
or U14382 (N_14382,N_9007,N_7853);
and U14383 (N_14383,N_5996,N_5559);
nand U14384 (N_14384,N_9405,N_5699);
xnor U14385 (N_14385,N_5628,N_5715);
and U14386 (N_14386,N_7650,N_7603);
nor U14387 (N_14387,N_8979,N_6680);
and U14388 (N_14388,N_6505,N_5659);
or U14389 (N_14389,N_8656,N_6554);
xor U14390 (N_14390,N_9265,N_5526);
or U14391 (N_14391,N_7209,N_5529);
and U14392 (N_14392,N_9181,N_6189);
or U14393 (N_14393,N_8140,N_7576);
nor U14394 (N_14394,N_6702,N_7947);
and U14395 (N_14395,N_7985,N_8940);
nor U14396 (N_14396,N_6562,N_8620);
and U14397 (N_14397,N_5018,N_7226);
nor U14398 (N_14398,N_5001,N_7792);
nor U14399 (N_14399,N_7530,N_8838);
and U14400 (N_14400,N_6434,N_9230);
nor U14401 (N_14401,N_9665,N_9845);
and U14402 (N_14402,N_9525,N_9636);
or U14403 (N_14403,N_5563,N_6457);
nor U14404 (N_14404,N_7341,N_8395);
nor U14405 (N_14405,N_9403,N_7392);
xnor U14406 (N_14406,N_5293,N_8309);
nand U14407 (N_14407,N_8104,N_6877);
or U14408 (N_14408,N_6184,N_9800);
and U14409 (N_14409,N_5431,N_6866);
nor U14410 (N_14410,N_7605,N_8151);
nand U14411 (N_14411,N_5381,N_8895);
nand U14412 (N_14412,N_9200,N_6719);
xor U14413 (N_14413,N_9647,N_9022);
nor U14414 (N_14414,N_9112,N_7892);
nor U14415 (N_14415,N_8022,N_8953);
and U14416 (N_14416,N_9040,N_7210);
xor U14417 (N_14417,N_8925,N_8951);
or U14418 (N_14418,N_5535,N_6362);
and U14419 (N_14419,N_7539,N_7161);
and U14420 (N_14420,N_7134,N_7458);
or U14421 (N_14421,N_8350,N_6859);
and U14422 (N_14422,N_8011,N_8689);
xnor U14423 (N_14423,N_9261,N_7119);
nor U14424 (N_14424,N_7109,N_6166);
and U14425 (N_14425,N_5522,N_7935);
or U14426 (N_14426,N_9305,N_8923);
and U14427 (N_14427,N_6145,N_8880);
nor U14428 (N_14428,N_5448,N_5035);
nand U14429 (N_14429,N_6841,N_9566);
nand U14430 (N_14430,N_7458,N_9853);
nand U14431 (N_14431,N_6395,N_7345);
or U14432 (N_14432,N_6107,N_8017);
nand U14433 (N_14433,N_6374,N_6884);
nand U14434 (N_14434,N_7528,N_9142);
or U14435 (N_14435,N_9350,N_6012);
nand U14436 (N_14436,N_9338,N_7465);
or U14437 (N_14437,N_8128,N_5453);
xnor U14438 (N_14438,N_5373,N_7631);
nand U14439 (N_14439,N_8978,N_5560);
and U14440 (N_14440,N_6110,N_9384);
nand U14441 (N_14441,N_7559,N_9678);
and U14442 (N_14442,N_5447,N_9479);
nand U14443 (N_14443,N_9966,N_6940);
and U14444 (N_14444,N_6659,N_7935);
nor U14445 (N_14445,N_6013,N_8079);
nor U14446 (N_14446,N_5073,N_9079);
or U14447 (N_14447,N_7671,N_6874);
nor U14448 (N_14448,N_9816,N_5511);
or U14449 (N_14449,N_7628,N_7387);
and U14450 (N_14450,N_6430,N_9959);
or U14451 (N_14451,N_6678,N_7094);
or U14452 (N_14452,N_7679,N_8693);
and U14453 (N_14453,N_8458,N_5000);
nand U14454 (N_14454,N_8478,N_6438);
or U14455 (N_14455,N_9121,N_7239);
nor U14456 (N_14456,N_9037,N_7664);
and U14457 (N_14457,N_9105,N_8908);
or U14458 (N_14458,N_7195,N_5685);
or U14459 (N_14459,N_5654,N_9455);
or U14460 (N_14460,N_8808,N_6024);
xor U14461 (N_14461,N_7631,N_5238);
nand U14462 (N_14462,N_8218,N_9037);
nor U14463 (N_14463,N_9043,N_6628);
and U14464 (N_14464,N_5602,N_9527);
and U14465 (N_14465,N_7182,N_9677);
nor U14466 (N_14466,N_6757,N_8109);
and U14467 (N_14467,N_7196,N_9488);
and U14468 (N_14468,N_8067,N_7463);
and U14469 (N_14469,N_5307,N_9057);
nor U14470 (N_14470,N_7142,N_6614);
and U14471 (N_14471,N_6872,N_6149);
nand U14472 (N_14472,N_9631,N_8787);
or U14473 (N_14473,N_5603,N_8160);
nor U14474 (N_14474,N_7524,N_7261);
and U14475 (N_14475,N_6235,N_6173);
nor U14476 (N_14476,N_6951,N_7867);
nor U14477 (N_14477,N_5054,N_7451);
and U14478 (N_14478,N_7313,N_9259);
nand U14479 (N_14479,N_8181,N_5516);
nor U14480 (N_14480,N_5973,N_6526);
and U14481 (N_14481,N_8066,N_8407);
or U14482 (N_14482,N_7090,N_6076);
xor U14483 (N_14483,N_9019,N_5487);
or U14484 (N_14484,N_7832,N_5171);
nor U14485 (N_14485,N_8977,N_8789);
xor U14486 (N_14486,N_5083,N_9948);
and U14487 (N_14487,N_5894,N_6692);
and U14488 (N_14488,N_9444,N_6468);
nor U14489 (N_14489,N_9798,N_9308);
nor U14490 (N_14490,N_7401,N_5889);
and U14491 (N_14491,N_5741,N_9781);
nand U14492 (N_14492,N_6017,N_9038);
nor U14493 (N_14493,N_9107,N_6065);
or U14494 (N_14494,N_7625,N_8188);
nor U14495 (N_14495,N_6657,N_8812);
nand U14496 (N_14496,N_9860,N_8760);
and U14497 (N_14497,N_8210,N_6354);
nand U14498 (N_14498,N_5040,N_6112);
xnor U14499 (N_14499,N_5979,N_7045);
or U14500 (N_14500,N_5069,N_6192);
xor U14501 (N_14501,N_6363,N_9547);
xnor U14502 (N_14502,N_6157,N_7631);
nor U14503 (N_14503,N_9542,N_9079);
and U14504 (N_14504,N_6089,N_5174);
nand U14505 (N_14505,N_8758,N_9389);
nand U14506 (N_14506,N_9726,N_6594);
or U14507 (N_14507,N_9879,N_6406);
nor U14508 (N_14508,N_5378,N_9093);
nor U14509 (N_14509,N_9079,N_8032);
xnor U14510 (N_14510,N_8128,N_7954);
and U14511 (N_14511,N_8256,N_7179);
nor U14512 (N_14512,N_8068,N_6745);
nor U14513 (N_14513,N_6024,N_9480);
and U14514 (N_14514,N_7701,N_9632);
nor U14515 (N_14515,N_9596,N_5078);
and U14516 (N_14516,N_9260,N_5838);
xor U14517 (N_14517,N_6803,N_6732);
and U14518 (N_14518,N_9349,N_6079);
and U14519 (N_14519,N_8958,N_6359);
xnor U14520 (N_14520,N_6193,N_9320);
or U14521 (N_14521,N_9502,N_8752);
nor U14522 (N_14522,N_9820,N_7838);
or U14523 (N_14523,N_6080,N_5426);
and U14524 (N_14524,N_9595,N_7592);
nand U14525 (N_14525,N_8977,N_6067);
and U14526 (N_14526,N_7509,N_7081);
xor U14527 (N_14527,N_9135,N_6578);
nand U14528 (N_14528,N_9260,N_8023);
and U14529 (N_14529,N_5945,N_9727);
nand U14530 (N_14530,N_5163,N_6068);
or U14531 (N_14531,N_7145,N_9396);
nand U14532 (N_14532,N_6022,N_9244);
nand U14533 (N_14533,N_9928,N_6603);
nand U14534 (N_14534,N_9462,N_8870);
xor U14535 (N_14535,N_5116,N_6650);
or U14536 (N_14536,N_5994,N_5272);
nand U14537 (N_14537,N_5939,N_7794);
nor U14538 (N_14538,N_8882,N_5465);
nand U14539 (N_14539,N_5835,N_5790);
nand U14540 (N_14540,N_5630,N_8115);
and U14541 (N_14541,N_8763,N_6636);
nor U14542 (N_14542,N_6776,N_5258);
or U14543 (N_14543,N_6062,N_9584);
xor U14544 (N_14544,N_6038,N_7584);
or U14545 (N_14545,N_9242,N_5117);
nor U14546 (N_14546,N_7028,N_9838);
nand U14547 (N_14547,N_9071,N_8428);
xor U14548 (N_14548,N_9162,N_7012);
nand U14549 (N_14549,N_5458,N_8568);
xnor U14550 (N_14550,N_5322,N_8109);
and U14551 (N_14551,N_8426,N_7964);
and U14552 (N_14552,N_8869,N_6425);
and U14553 (N_14553,N_6977,N_8538);
or U14554 (N_14554,N_6683,N_5728);
xor U14555 (N_14555,N_9432,N_9171);
nor U14556 (N_14556,N_8999,N_7407);
nor U14557 (N_14557,N_7267,N_5407);
nor U14558 (N_14558,N_6490,N_6143);
xor U14559 (N_14559,N_8888,N_7902);
and U14560 (N_14560,N_7929,N_9624);
nand U14561 (N_14561,N_5155,N_5295);
xnor U14562 (N_14562,N_5451,N_5439);
nand U14563 (N_14563,N_5939,N_5987);
xnor U14564 (N_14564,N_5021,N_6182);
xnor U14565 (N_14565,N_7169,N_6688);
or U14566 (N_14566,N_9063,N_9660);
nand U14567 (N_14567,N_8356,N_7195);
or U14568 (N_14568,N_7273,N_6592);
and U14569 (N_14569,N_9886,N_5432);
nand U14570 (N_14570,N_9964,N_9862);
nor U14571 (N_14571,N_8486,N_5076);
xnor U14572 (N_14572,N_8248,N_8651);
xnor U14573 (N_14573,N_8215,N_5674);
nor U14574 (N_14574,N_8014,N_8627);
nand U14575 (N_14575,N_5470,N_8989);
xor U14576 (N_14576,N_9594,N_8975);
xnor U14577 (N_14577,N_7682,N_6902);
and U14578 (N_14578,N_7965,N_6230);
or U14579 (N_14579,N_8058,N_9899);
xnor U14580 (N_14580,N_8924,N_5255);
xnor U14581 (N_14581,N_8479,N_5475);
xor U14582 (N_14582,N_5232,N_7567);
nand U14583 (N_14583,N_9439,N_7443);
xnor U14584 (N_14584,N_5591,N_6115);
nand U14585 (N_14585,N_8664,N_5448);
xnor U14586 (N_14586,N_7105,N_8656);
nand U14587 (N_14587,N_5416,N_5820);
xnor U14588 (N_14588,N_8465,N_6559);
and U14589 (N_14589,N_6030,N_5670);
xnor U14590 (N_14590,N_7539,N_6284);
xor U14591 (N_14591,N_6427,N_9774);
or U14592 (N_14592,N_8296,N_6098);
nor U14593 (N_14593,N_8241,N_6396);
nand U14594 (N_14594,N_8514,N_9647);
and U14595 (N_14595,N_6914,N_5481);
and U14596 (N_14596,N_8200,N_8066);
xor U14597 (N_14597,N_6988,N_9671);
and U14598 (N_14598,N_8611,N_8721);
xnor U14599 (N_14599,N_8553,N_9003);
nand U14600 (N_14600,N_7703,N_8843);
nand U14601 (N_14601,N_9798,N_8194);
and U14602 (N_14602,N_8599,N_7007);
and U14603 (N_14603,N_8133,N_9970);
nor U14604 (N_14604,N_9968,N_9556);
or U14605 (N_14605,N_5682,N_7735);
nor U14606 (N_14606,N_5212,N_5372);
or U14607 (N_14607,N_5414,N_7422);
or U14608 (N_14608,N_6845,N_5313);
xor U14609 (N_14609,N_5709,N_8001);
or U14610 (N_14610,N_8431,N_6163);
nor U14611 (N_14611,N_9748,N_9438);
xnor U14612 (N_14612,N_5461,N_7210);
and U14613 (N_14613,N_9984,N_7621);
and U14614 (N_14614,N_7893,N_9003);
or U14615 (N_14615,N_7159,N_9075);
xnor U14616 (N_14616,N_5166,N_7810);
or U14617 (N_14617,N_6337,N_9552);
xnor U14618 (N_14618,N_7329,N_5855);
nor U14619 (N_14619,N_6190,N_8016);
nor U14620 (N_14620,N_5379,N_8237);
and U14621 (N_14621,N_6600,N_6196);
nand U14622 (N_14622,N_9010,N_5309);
nor U14623 (N_14623,N_8630,N_7795);
and U14624 (N_14624,N_8410,N_6558);
nor U14625 (N_14625,N_7292,N_7286);
and U14626 (N_14626,N_8793,N_8916);
nand U14627 (N_14627,N_9396,N_7707);
nand U14628 (N_14628,N_8182,N_8979);
or U14629 (N_14629,N_9995,N_6581);
xor U14630 (N_14630,N_9671,N_7099);
or U14631 (N_14631,N_7518,N_7106);
or U14632 (N_14632,N_5975,N_8447);
nand U14633 (N_14633,N_8792,N_8989);
nor U14634 (N_14634,N_7844,N_9711);
nor U14635 (N_14635,N_8483,N_9228);
xor U14636 (N_14636,N_9414,N_6119);
nand U14637 (N_14637,N_8118,N_7537);
or U14638 (N_14638,N_6472,N_5036);
xor U14639 (N_14639,N_9278,N_7241);
nor U14640 (N_14640,N_7168,N_6459);
nor U14641 (N_14641,N_7657,N_8629);
xor U14642 (N_14642,N_8204,N_8049);
or U14643 (N_14643,N_9560,N_5013);
and U14644 (N_14644,N_7193,N_8661);
and U14645 (N_14645,N_9489,N_7579);
xnor U14646 (N_14646,N_9334,N_9893);
nand U14647 (N_14647,N_7535,N_7522);
xnor U14648 (N_14648,N_8542,N_9203);
or U14649 (N_14649,N_8624,N_7648);
or U14650 (N_14650,N_6874,N_8271);
and U14651 (N_14651,N_7066,N_8343);
nand U14652 (N_14652,N_6887,N_9941);
and U14653 (N_14653,N_9600,N_6023);
nor U14654 (N_14654,N_6106,N_9539);
xnor U14655 (N_14655,N_7532,N_6475);
nor U14656 (N_14656,N_9724,N_5087);
xor U14657 (N_14657,N_6496,N_9153);
and U14658 (N_14658,N_9437,N_5097);
or U14659 (N_14659,N_5957,N_5939);
and U14660 (N_14660,N_9155,N_6966);
nand U14661 (N_14661,N_8052,N_9335);
xor U14662 (N_14662,N_5607,N_9561);
nand U14663 (N_14663,N_6890,N_6467);
nand U14664 (N_14664,N_9725,N_9321);
and U14665 (N_14665,N_6447,N_7381);
nand U14666 (N_14666,N_8336,N_7077);
xor U14667 (N_14667,N_6638,N_9345);
or U14668 (N_14668,N_7541,N_8443);
xor U14669 (N_14669,N_9008,N_7755);
xor U14670 (N_14670,N_9313,N_6065);
or U14671 (N_14671,N_7262,N_7496);
or U14672 (N_14672,N_9623,N_8853);
or U14673 (N_14673,N_8232,N_6940);
and U14674 (N_14674,N_7845,N_8187);
and U14675 (N_14675,N_9670,N_6130);
or U14676 (N_14676,N_6166,N_5639);
and U14677 (N_14677,N_5500,N_5553);
nor U14678 (N_14678,N_6722,N_6791);
and U14679 (N_14679,N_5970,N_9629);
or U14680 (N_14680,N_5973,N_7735);
and U14681 (N_14681,N_7057,N_5850);
nor U14682 (N_14682,N_9922,N_8736);
xor U14683 (N_14683,N_7764,N_5951);
and U14684 (N_14684,N_9258,N_5225);
and U14685 (N_14685,N_7769,N_6352);
nor U14686 (N_14686,N_7234,N_6579);
and U14687 (N_14687,N_6433,N_6731);
and U14688 (N_14688,N_8005,N_7933);
and U14689 (N_14689,N_5249,N_8951);
nor U14690 (N_14690,N_6440,N_5729);
xor U14691 (N_14691,N_5581,N_8375);
nor U14692 (N_14692,N_7895,N_7293);
and U14693 (N_14693,N_5583,N_9491);
nor U14694 (N_14694,N_8719,N_5604);
and U14695 (N_14695,N_8959,N_9316);
xnor U14696 (N_14696,N_6601,N_8505);
and U14697 (N_14697,N_8615,N_6219);
nor U14698 (N_14698,N_6549,N_9099);
nand U14699 (N_14699,N_8202,N_5327);
xor U14700 (N_14700,N_9286,N_5336);
or U14701 (N_14701,N_7723,N_6490);
nor U14702 (N_14702,N_8129,N_7881);
and U14703 (N_14703,N_5692,N_7626);
or U14704 (N_14704,N_5853,N_6945);
xnor U14705 (N_14705,N_5364,N_9249);
or U14706 (N_14706,N_9573,N_5744);
nor U14707 (N_14707,N_8192,N_7159);
xor U14708 (N_14708,N_8860,N_5072);
or U14709 (N_14709,N_5115,N_9564);
or U14710 (N_14710,N_6355,N_6773);
and U14711 (N_14711,N_9818,N_7168);
nor U14712 (N_14712,N_5035,N_9028);
xor U14713 (N_14713,N_7297,N_6293);
nand U14714 (N_14714,N_7622,N_8188);
nor U14715 (N_14715,N_5911,N_7679);
nor U14716 (N_14716,N_7095,N_8049);
or U14717 (N_14717,N_9694,N_9930);
xor U14718 (N_14718,N_5292,N_7989);
nor U14719 (N_14719,N_5800,N_5644);
nand U14720 (N_14720,N_6925,N_5356);
and U14721 (N_14721,N_9234,N_8074);
and U14722 (N_14722,N_7827,N_7980);
or U14723 (N_14723,N_7407,N_6185);
nor U14724 (N_14724,N_7293,N_5774);
and U14725 (N_14725,N_6505,N_8935);
xnor U14726 (N_14726,N_7156,N_8978);
and U14727 (N_14727,N_8394,N_7891);
or U14728 (N_14728,N_7540,N_8980);
and U14729 (N_14729,N_9343,N_9883);
nand U14730 (N_14730,N_6458,N_8534);
or U14731 (N_14731,N_8369,N_5613);
xor U14732 (N_14732,N_6374,N_8138);
and U14733 (N_14733,N_6369,N_9560);
or U14734 (N_14734,N_7327,N_6932);
nor U14735 (N_14735,N_5626,N_5593);
xnor U14736 (N_14736,N_9042,N_6442);
or U14737 (N_14737,N_5903,N_6841);
nor U14738 (N_14738,N_8837,N_9956);
or U14739 (N_14739,N_9312,N_5397);
nand U14740 (N_14740,N_8343,N_7341);
nand U14741 (N_14741,N_8478,N_8611);
xnor U14742 (N_14742,N_9439,N_7489);
nor U14743 (N_14743,N_9265,N_9312);
and U14744 (N_14744,N_5178,N_8961);
and U14745 (N_14745,N_9775,N_5086);
xor U14746 (N_14746,N_6566,N_9761);
nand U14747 (N_14747,N_7817,N_8119);
and U14748 (N_14748,N_7435,N_7820);
or U14749 (N_14749,N_7024,N_7919);
or U14750 (N_14750,N_9770,N_6019);
nand U14751 (N_14751,N_5829,N_5218);
xnor U14752 (N_14752,N_7464,N_7866);
or U14753 (N_14753,N_8001,N_8370);
nand U14754 (N_14754,N_7609,N_7696);
nor U14755 (N_14755,N_8305,N_9386);
and U14756 (N_14756,N_5944,N_8462);
xnor U14757 (N_14757,N_7651,N_5323);
xnor U14758 (N_14758,N_9346,N_6934);
nor U14759 (N_14759,N_8365,N_9774);
nor U14760 (N_14760,N_9685,N_7013);
xor U14761 (N_14761,N_5839,N_8174);
and U14762 (N_14762,N_8797,N_9003);
and U14763 (N_14763,N_5193,N_7581);
xor U14764 (N_14764,N_9175,N_6094);
nand U14765 (N_14765,N_9159,N_5812);
xnor U14766 (N_14766,N_7857,N_8631);
nand U14767 (N_14767,N_5193,N_9638);
nor U14768 (N_14768,N_7326,N_5904);
and U14769 (N_14769,N_5772,N_7687);
and U14770 (N_14770,N_7844,N_7580);
and U14771 (N_14771,N_9417,N_9099);
nor U14772 (N_14772,N_9531,N_7405);
xnor U14773 (N_14773,N_5689,N_7805);
and U14774 (N_14774,N_5012,N_9911);
xnor U14775 (N_14775,N_9897,N_5584);
nand U14776 (N_14776,N_6709,N_7989);
or U14777 (N_14777,N_5247,N_5021);
nor U14778 (N_14778,N_9095,N_8383);
nand U14779 (N_14779,N_9709,N_9428);
and U14780 (N_14780,N_7179,N_8885);
nor U14781 (N_14781,N_7595,N_6248);
nor U14782 (N_14782,N_7887,N_6265);
nor U14783 (N_14783,N_8689,N_9636);
xor U14784 (N_14784,N_5473,N_8959);
xor U14785 (N_14785,N_5236,N_9852);
nand U14786 (N_14786,N_7359,N_6740);
xnor U14787 (N_14787,N_8492,N_8845);
or U14788 (N_14788,N_5841,N_8020);
nor U14789 (N_14789,N_6710,N_7461);
xor U14790 (N_14790,N_7532,N_6202);
nand U14791 (N_14791,N_6045,N_9245);
and U14792 (N_14792,N_5412,N_8300);
nand U14793 (N_14793,N_8011,N_7017);
or U14794 (N_14794,N_9258,N_7914);
xor U14795 (N_14795,N_8273,N_6460);
xor U14796 (N_14796,N_6194,N_5658);
nor U14797 (N_14797,N_8950,N_5690);
nor U14798 (N_14798,N_5237,N_6238);
or U14799 (N_14799,N_9062,N_6559);
nor U14800 (N_14800,N_8456,N_9269);
or U14801 (N_14801,N_8238,N_9694);
nor U14802 (N_14802,N_5620,N_7252);
or U14803 (N_14803,N_5807,N_6569);
or U14804 (N_14804,N_6269,N_8884);
or U14805 (N_14805,N_9753,N_8656);
xnor U14806 (N_14806,N_7270,N_8800);
or U14807 (N_14807,N_6133,N_6298);
xor U14808 (N_14808,N_6385,N_8289);
and U14809 (N_14809,N_5684,N_7010);
xor U14810 (N_14810,N_6960,N_8460);
or U14811 (N_14811,N_5063,N_8769);
xnor U14812 (N_14812,N_8767,N_6877);
and U14813 (N_14813,N_7269,N_7384);
nand U14814 (N_14814,N_7725,N_8108);
xor U14815 (N_14815,N_8320,N_9991);
nand U14816 (N_14816,N_6393,N_7950);
xor U14817 (N_14817,N_5446,N_7851);
and U14818 (N_14818,N_9745,N_8477);
and U14819 (N_14819,N_5719,N_9568);
or U14820 (N_14820,N_7608,N_6712);
xnor U14821 (N_14821,N_5875,N_8320);
and U14822 (N_14822,N_6561,N_7188);
xor U14823 (N_14823,N_8131,N_7376);
and U14824 (N_14824,N_8531,N_8670);
nor U14825 (N_14825,N_8929,N_7091);
xnor U14826 (N_14826,N_8242,N_7192);
xor U14827 (N_14827,N_6190,N_7522);
nand U14828 (N_14828,N_6934,N_5467);
xor U14829 (N_14829,N_6934,N_7625);
xor U14830 (N_14830,N_6125,N_9096);
or U14831 (N_14831,N_5533,N_8335);
and U14832 (N_14832,N_5051,N_8258);
nand U14833 (N_14833,N_8953,N_8587);
xnor U14834 (N_14834,N_7382,N_8419);
xor U14835 (N_14835,N_9033,N_6227);
and U14836 (N_14836,N_7826,N_9486);
and U14837 (N_14837,N_6388,N_6853);
and U14838 (N_14838,N_8071,N_9347);
and U14839 (N_14839,N_5364,N_9845);
nor U14840 (N_14840,N_6504,N_8166);
nor U14841 (N_14841,N_9634,N_5563);
or U14842 (N_14842,N_7648,N_9487);
xor U14843 (N_14843,N_7154,N_5624);
nor U14844 (N_14844,N_8819,N_6654);
nor U14845 (N_14845,N_7675,N_9915);
nor U14846 (N_14846,N_8210,N_6901);
nor U14847 (N_14847,N_5294,N_9847);
xor U14848 (N_14848,N_8020,N_8504);
nand U14849 (N_14849,N_6368,N_6512);
nand U14850 (N_14850,N_8741,N_7721);
nand U14851 (N_14851,N_9326,N_6762);
nand U14852 (N_14852,N_6374,N_5552);
and U14853 (N_14853,N_5301,N_9666);
nand U14854 (N_14854,N_8633,N_7386);
or U14855 (N_14855,N_6734,N_5270);
or U14856 (N_14856,N_6265,N_7012);
xor U14857 (N_14857,N_8833,N_5564);
xnor U14858 (N_14858,N_7250,N_7832);
or U14859 (N_14859,N_6523,N_5927);
and U14860 (N_14860,N_7068,N_7828);
and U14861 (N_14861,N_9532,N_9458);
or U14862 (N_14862,N_7111,N_9830);
and U14863 (N_14863,N_6341,N_7193);
or U14864 (N_14864,N_7769,N_5325);
nand U14865 (N_14865,N_9916,N_9918);
or U14866 (N_14866,N_6925,N_5269);
or U14867 (N_14867,N_7126,N_9892);
and U14868 (N_14868,N_6383,N_9257);
nand U14869 (N_14869,N_7167,N_5681);
nand U14870 (N_14870,N_6941,N_8528);
and U14871 (N_14871,N_7408,N_8371);
nor U14872 (N_14872,N_9392,N_7432);
and U14873 (N_14873,N_5053,N_5563);
and U14874 (N_14874,N_5327,N_8529);
xor U14875 (N_14875,N_6579,N_9073);
or U14876 (N_14876,N_7176,N_6458);
nand U14877 (N_14877,N_5020,N_6155);
nor U14878 (N_14878,N_5174,N_7670);
nor U14879 (N_14879,N_6458,N_6586);
or U14880 (N_14880,N_7173,N_5815);
or U14881 (N_14881,N_9171,N_7376);
nor U14882 (N_14882,N_5728,N_6150);
nor U14883 (N_14883,N_5062,N_9881);
or U14884 (N_14884,N_9990,N_8828);
nor U14885 (N_14885,N_5862,N_6566);
xor U14886 (N_14886,N_6920,N_5917);
and U14887 (N_14887,N_8780,N_9274);
nor U14888 (N_14888,N_7255,N_5147);
or U14889 (N_14889,N_8983,N_7549);
nand U14890 (N_14890,N_6690,N_8522);
nor U14891 (N_14891,N_7659,N_5153);
nor U14892 (N_14892,N_9040,N_6748);
or U14893 (N_14893,N_6430,N_8207);
nand U14894 (N_14894,N_7151,N_9875);
or U14895 (N_14895,N_5042,N_8356);
nand U14896 (N_14896,N_5208,N_7045);
nand U14897 (N_14897,N_8565,N_8364);
or U14898 (N_14898,N_8313,N_5316);
nand U14899 (N_14899,N_6847,N_8220);
or U14900 (N_14900,N_7235,N_7432);
xor U14901 (N_14901,N_6747,N_7436);
and U14902 (N_14902,N_6242,N_9122);
nor U14903 (N_14903,N_5149,N_8849);
or U14904 (N_14904,N_5632,N_5052);
nor U14905 (N_14905,N_6796,N_8588);
or U14906 (N_14906,N_8984,N_7767);
xor U14907 (N_14907,N_6364,N_9552);
or U14908 (N_14908,N_5274,N_9053);
xor U14909 (N_14909,N_5245,N_9989);
nand U14910 (N_14910,N_9351,N_6203);
and U14911 (N_14911,N_7183,N_8787);
and U14912 (N_14912,N_8644,N_8411);
or U14913 (N_14913,N_5872,N_9967);
and U14914 (N_14914,N_8021,N_9467);
or U14915 (N_14915,N_7351,N_8127);
nor U14916 (N_14916,N_8843,N_8577);
nor U14917 (N_14917,N_6416,N_9429);
and U14918 (N_14918,N_5139,N_5839);
and U14919 (N_14919,N_6079,N_8493);
nor U14920 (N_14920,N_5075,N_6878);
and U14921 (N_14921,N_7698,N_9772);
nor U14922 (N_14922,N_9556,N_7703);
or U14923 (N_14923,N_6819,N_5891);
nor U14924 (N_14924,N_9574,N_7273);
nand U14925 (N_14925,N_9086,N_8885);
nor U14926 (N_14926,N_6006,N_6523);
or U14927 (N_14927,N_9932,N_8263);
xnor U14928 (N_14928,N_8675,N_7192);
nor U14929 (N_14929,N_5477,N_6220);
nor U14930 (N_14930,N_5197,N_9504);
xor U14931 (N_14931,N_8586,N_6487);
and U14932 (N_14932,N_7553,N_8483);
nand U14933 (N_14933,N_5091,N_7595);
nand U14934 (N_14934,N_6648,N_5397);
and U14935 (N_14935,N_6475,N_6130);
nor U14936 (N_14936,N_5554,N_6567);
or U14937 (N_14937,N_5586,N_7860);
nand U14938 (N_14938,N_8117,N_8005);
xor U14939 (N_14939,N_8930,N_6465);
or U14940 (N_14940,N_6482,N_8328);
or U14941 (N_14941,N_9018,N_5282);
nor U14942 (N_14942,N_6883,N_6502);
nand U14943 (N_14943,N_7198,N_8273);
nand U14944 (N_14944,N_8798,N_7638);
nand U14945 (N_14945,N_7324,N_7335);
nand U14946 (N_14946,N_8161,N_7596);
nor U14947 (N_14947,N_8136,N_6993);
nor U14948 (N_14948,N_7844,N_9959);
or U14949 (N_14949,N_5536,N_8473);
and U14950 (N_14950,N_8092,N_6302);
nor U14951 (N_14951,N_7934,N_5585);
xnor U14952 (N_14952,N_9216,N_8531);
xnor U14953 (N_14953,N_8830,N_8022);
nand U14954 (N_14954,N_9924,N_8026);
xor U14955 (N_14955,N_7766,N_7535);
nor U14956 (N_14956,N_7558,N_6248);
nand U14957 (N_14957,N_9251,N_7762);
or U14958 (N_14958,N_8522,N_6977);
nand U14959 (N_14959,N_5956,N_7148);
nor U14960 (N_14960,N_5634,N_5313);
nand U14961 (N_14961,N_5474,N_7692);
nor U14962 (N_14962,N_6478,N_7013);
nand U14963 (N_14963,N_7740,N_8887);
or U14964 (N_14964,N_5469,N_7371);
nand U14965 (N_14965,N_8165,N_7540);
nand U14966 (N_14966,N_9050,N_5437);
xnor U14967 (N_14967,N_5764,N_5821);
xor U14968 (N_14968,N_8602,N_6281);
nand U14969 (N_14969,N_6550,N_6211);
nand U14970 (N_14970,N_5818,N_5504);
xor U14971 (N_14971,N_5228,N_5859);
nor U14972 (N_14972,N_7188,N_9480);
and U14973 (N_14973,N_8775,N_5187);
or U14974 (N_14974,N_5280,N_6745);
and U14975 (N_14975,N_8950,N_9584);
xnor U14976 (N_14976,N_7419,N_7930);
nand U14977 (N_14977,N_8362,N_6918);
nand U14978 (N_14978,N_8698,N_5475);
or U14979 (N_14979,N_8823,N_6451);
nand U14980 (N_14980,N_5838,N_9162);
nor U14981 (N_14981,N_9520,N_7215);
and U14982 (N_14982,N_5060,N_8497);
nor U14983 (N_14983,N_6703,N_7567);
and U14984 (N_14984,N_7442,N_7087);
and U14985 (N_14985,N_8128,N_9685);
xor U14986 (N_14986,N_9090,N_6127);
nand U14987 (N_14987,N_6910,N_9332);
xor U14988 (N_14988,N_5948,N_7916);
nor U14989 (N_14989,N_8788,N_8752);
nand U14990 (N_14990,N_7762,N_5775);
nand U14991 (N_14991,N_7424,N_5714);
nor U14992 (N_14992,N_7791,N_8229);
nor U14993 (N_14993,N_6034,N_5171);
or U14994 (N_14994,N_9246,N_6010);
or U14995 (N_14995,N_6436,N_5230);
or U14996 (N_14996,N_9206,N_5640);
nor U14997 (N_14997,N_8139,N_9203);
or U14998 (N_14998,N_8489,N_7182);
nor U14999 (N_14999,N_5533,N_8441);
nand UO_0 (O_0,N_11892,N_14532);
nor UO_1 (O_1,N_11500,N_11705);
nand UO_2 (O_2,N_12769,N_10847);
or UO_3 (O_3,N_10288,N_11030);
or UO_4 (O_4,N_12228,N_13223);
or UO_5 (O_5,N_14838,N_10873);
nand UO_6 (O_6,N_10826,N_14656);
nor UO_7 (O_7,N_13026,N_14659);
and UO_8 (O_8,N_10033,N_12134);
xor UO_9 (O_9,N_13775,N_11515);
or UO_10 (O_10,N_11548,N_13648);
and UO_11 (O_11,N_12291,N_11420);
nor UO_12 (O_12,N_12252,N_11182);
nor UO_13 (O_13,N_10749,N_12112);
and UO_14 (O_14,N_13524,N_12524);
nand UO_15 (O_15,N_11772,N_11434);
nor UO_16 (O_16,N_12118,N_12827);
and UO_17 (O_17,N_11588,N_13328);
and UO_18 (O_18,N_12785,N_11701);
nor UO_19 (O_19,N_14001,N_13763);
nor UO_20 (O_20,N_12175,N_11468);
xnor UO_21 (O_21,N_12616,N_10010);
nand UO_22 (O_22,N_10709,N_13426);
and UO_23 (O_23,N_14196,N_11081);
or UO_24 (O_24,N_10652,N_13950);
nor UO_25 (O_25,N_10778,N_11095);
nand UO_26 (O_26,N_12028,N_14377);
or UO_27 (O_27,N_12916,N_12305);
nor UO_28 (O_28,N_10861,N_10818);
and UO_29 (O_29,N_12387,N_12347);
nand UO_30 (O_30,N_12946,N_10273);
or UO_31 (O_31,N_11855,N_11417);
nand UO_32 (O_32,N_13310,N_10933);
and UO_33 (O_33,N_14418,N_12718);
xnor UO_34 (O_34,N_11990,N_10874);
xnor UO_35 (O_35,N_14831,N_11384);
and UO_36 (O_36,N_12503,N_13850);
nand UO_37 (O_37,N_10843,N_10993);
nand UO_38 (O_38,N_13810,N_14421);
nor UO_39 (O_39,N_14882,N_12979);
xnor UO_40 (O_40,N_12928,N_14976);
xnor UO_41 (O_41,N_14751,N_14425);
nand UO_42 (O_42,N_10880,N_13510);
and UO_43 (O_43,N_14175,N_12336);
or UO_44 (O_44,N_13423,N_14410);
nor UO_45 (O_45,N_13452,N_10581);
xnor UO_46 (O_46,N_12831,N_13351);
and UO_47 (O_47,N_13016,N_14840);
nand UO_48 (O_48,N_11489,N_10676);
or UO_49 (O_49,N_11714,N_13534);
or UO_50 (O_50,N_11414,N_10090);
nor UO_51 (O_51,N_14512,N_13318);
xnor UO_52 (O_52,N_10468,N_14665);
or UO_53 (O_53,N_11785,N_12915);
or UO_54 (O_54,N_12147,N_13902);
or UO_55 (O_55,N_12110,N_13401);
nand UO_56 (O_56,N_14288,N_12376);
and UO_57 (O_57,N_10975,N_12453);
nand UO_58 (O_58,N_13133,N_10139);
nor UO_59 (O_59,N_10669,N_10465);
xnor UO_60 (O_60,N_11371,N_14587);
nand UO_61 (O_61,N_14752,N_11786);
or UO_62 (O_62,N_13150,N_11383);
xor UO_63 (O_63,N_10599,N_11914);
xor UO_64 (O_64,N_12274,N_14322);
xnor UO_65 (O_65,N_10456,N_10216);
nor UO_66 (O_66,N_11569,N_11689);
nand UO_67 (O_67,N_10539,N_14977);
or UO_68 (O_68,N_12299,N_10004);
or UO_69 (O_69,N_11720,N_14195);
nand UO_70 (O_70,N_13792,N_13306);
nand UO_71 (O_71,N_11265,N_10824);
xnor UO_72 (O_72,N_11181,N_13008);
xor UO_73 (O_73,N_10729,N_14231);
nand UO_74 (O_74,N_14803,N_10814);
and UO_75 (O_75,N_12036,N_13254);
nor UO_76 (O_76,N_12295,N_12481);
xor UO_77 (O_77,N_11243,N_13547);
or UO_78 (O_78,N_11726,N_11213);
and UO_79 (O_79,N_12180,N_14958);
xor UO_80 (O_80,N_11851,N_14079);
and UO_81 (O_81,N_12158,N_10694);
and UO_82 (O_82,N_14750,N_11742);
or UO_83 (O_83,N_13007,N_11062);
nor UO_84 (O_84,N_12354,N_11345);
or UO_85 (O_85,N_14061,N_10274);
nand UO_86 (O_86,N_13335,N_11018);
or UO_87 (O_87,N_11130,N_11981);
nor UO_88 (O_88,N_10124,N_10497);
and UO_89 (O_89,N_12476,N_10422);
nand UO_90 (O_90,N_11973,N_13461);
xnor UO_91 (O_91,N_11799,N_14192);
and UO_92 (O_92,N_13906,N_10209);
or UO_93 (O_93,N_10157,N_14179);
nor UO_94 (O_94,N_12137,N_11970);
nand UO_95 (O_95,N_11312,N_12407);
xor UO_96 (O_96,N_11526,N_13447);
and UO_97 (O_97,N_12455,N_11511);
nand UO_98 (O_98,N_12715,N_13113);
nor UO_99 (O_99,N_12547,N_10828);
or UO_100 (O_100,N_10785,N_10430);
or UO_101 (O_101,N_12938,N_14155);
nand UO_102 (O_102,N_10347,N_13859);
or UO_103 (O_103,N_10807,N_12699);
nor UO_104 (O_104,N_10394,N_10875);
or UO_105 (O_105,N_12952,N_11996);
and UO_106 (O_106,N_10726,N_12320);
nand UO_107 (O_107,N_13023,N_14523);
or UO_108 (O_108,N_14117,N_10120);
or UO_109 (O_109,N_11169,N_11814);
nor UO_110 (O_110,N_10131,N_12678);
or UO_111 (O_111,N_13761,N_11200);
nor UO_112 (O_112,N_11784,N_10223);
nor UO_113 (O_113,N_11887,N_12267);
and UO_114 (O_114,N_14862,N_13301);
nor UO_115 (O_115,N_13390,N_11029);
and UO_116 (O_116,N_14296,N_13292);
and UO_117 (O_117,N_12196,N_11863);
nand UO_118 (O_118,N_12622,N_12604);
xnor UO_119 (O_119,N_14794,N_14841);
nand UO_120 (O_120,N_11930,N_14860);
nand UO_121 (O_121,N_13341,N_14073);
xor UO_122 (O_122,N_10424,N_13414);
nand UO_123 (O_123,N_10498,N_13498);
or UO_124 (O_124,N_14006,N_11398);
and UO_125 (O_125,N_12969,N_11443);
xor UO_126 (O_126,N_10197,N_11798);
or UO_127 (O_127,N_13471,N_12873);
or UO_128 (O_128,N_14373,N_11359);
nand UO_129 (O_129,N_10162,N_14581);
nor UO_130 (O_130,N_10458,N_12934);
and UO_131 (O_131,N_12595,N_10686);
nand UO_132 (O_132,N_13721,N_14283);
and UO_133 (O_133,N_11674,N_13272);
nand UO_134 (O_134,N_11945,N_10077);
xor UO_135 (O_135,N_12582,N_14800);
or UO_136 (O_136,N_10587,N_14570);
or UO_137 (O_137,N_10622,N_12828);
nor UO_138 (O_138,N_12596,N_13595);
or UO_139 (O_139,N_13168,N_14509);
xnor UO_140 (O_140,N_10845,N_13497);
nor UO_141 (O_141,N_10298,N_13374);
xnor UO_142 (O_142,N_13093,N_10115);
or UO_143 (O_143,N_14692,N_12013);
nand UO_144 (O_144,N_12860,N_13283);
or UO_145 (O_145,N_12812,N_13560);
and UO_146 (O_146,N_11488,N_10434);
nand UO_147 (O_147,N_13312,N_10326);
nor UO_148 (O_148,N_14669,N_14878);
and UO_149 (O_149,N_14236,N_12429);
nand UO_150 (O_150,N_14622,N_10038);
nor UO_151 (O_151,N_14045,N_11059);
or UO_152 (O_152,N_10220,N_10883);
or UO_153 (O_153,N_13194,N_12247);
nor UO_154 (O_154,N_13081,N_14607);
and UO_155 (O_155,N_10574,N_11058);
and UO_156 (O_156,N_11953,N_14489);
or UO_157 (O_157,N_13893,N_12723);
nand UO_158 (O_158,N_12039,N_10059);
nor UO_159 (O_159,N_14475,N_13587);
or UO_160 (O_160,N_10588,N_13765);
nand UO_161 (O_161,N_12380,N_13465);
or UO_162 (O_162,N_12141,N_11827);
nand UO_163 (O_163,N_10537,N_10635);
nor UO_164 (O_164,N_10525,N_13702);
nand UO_165 (O_165,N_10436,N_14617);
nand UO_166 (O_166,N_14295,N_13406);
and UO_167 (O_167,N_10538,N_11547);
or UO_168 (O_168,N_10119,N_13323);
and UO_169 (O_169,N_11168,N_14234);
and UO_170 (O_170,N_10986,N_14932);
nor UO_171 (O_171,N_11316,N_13901);
and UO_172 (O_172,N_12691,N_10001);
nand UO_173 (O_173,N_14389,N_11293);
nor UO_174 (O_174,N_11721,N_14020);
xor UO_175 (O_175,N_11937,N_10564);
xnor UO_176 (O_176,N_11803,N_12774);
nor UO_177 (O_177,N_14731,N_11460);
and UO_178 (O_178,N_14388,N_14370);
xor UO_179 (O_179,N_12303,N_13490);
nand UO_180 (O_180,N_14582,N_10406);
nor UO_181 (O_181,N_11551,N_14531);
xor UO_182 (O_182,N_14613,N_12941);
xor UO_183 (O_183,N_13482,N_12795);
xor UO_184 (O_184,N_14398,N_14600);
or UO_185 (O_185,N_14160,N_12197);
nor UO_186 (O_186,N_12572,N_10490);
xnor UO_187 (O_187,N_12760,N_14686);
nand UO_188 (O_188,N_14002,N_12676);
and UO_189 (O_189,N_11745,N_14528);
xnor UO_190 (O_190,N_14652,N_13514);
xor UO_191 (O_191,N_13443,N_14371);
and UO_192 (O_192,N_13910,N_12800);
nand UO_193 (O_193,N_14149,N_14487);
or UO_194 (O_194,N_10397,N_10627);
xnor UO_195 (O_195,N_12082,N_13034);
nor UO_196 (O_196,N_11076,N_11940);
and UO_197 (O_197,N_11894,N_11241);
or UO_198 (O_198,N_14875,N_13554);
xnor UO_199 (O_199,N_10502,N_10585);
and UO_200 (O_200,N_12057,N_13467);
xnor UO_201 (O_201,N_13941,N_14657);
nand UO_202 (O_202,N_11049,N_14836);
or UO_203 (O_203,N_14998,N_10478);
nand UO_204 (O_204,N_10204,N_14627);
and UO_205 (O_205,N_13803,N_10745);
xnor UO_206 (O_206,N_12264,N_10928);
nor UO_207 (O_207,N_10572,N_13118);
or UO_208 (O_208,N_12880,N_10988);
nor UO_209 (O_209,N_13894,N_13974);
nor UO_210 (O_210,N_12312,N_10999);
nor UO_211 (O_211,N_13831,N_14265);
and UO_212 (O_212,N_11439,N_10247);
xor UO_213 (O_213,N_10783,N_14062);
nor UO_214 (O_214,N_10614,N_12738);
or UO_215 (O_215,N_12218,N_11157);
or UO_216 (O_216,N_10487,N_13979);
nand UO_217 (O_217,N_13229,N_10428);
nor UO_218 (O_218,N_11246,N_13486);
xnor UO_219 (O_219,N_11257,N_14473);
or UO_220 (O_220,N_14807,N_14161);
nand UO_221 (O_221,N_10452,N_13431);
and UO_222 (O_222,N_10776,N_14635);
nor UO_223 (O_223,N_10523,N_13170);
nand UO_224 (O_224,N_10018,N_14895);
or UO_225 (O_225,N_11052,N_10407);
nor UO_226 (O_226,N_12050,N_11430);
xnor UO_227 (O_227,N_13046,N_10552);
nor UO_228 (O_228,N_14811,N_12846);
and UO_229 (O_229,N_12975,N_13287);
and UO_230 (O_230,N_11704,N_13891);
and UO_231 (O_231,N_14864,N_13183);
nand UO_232 (O_232,N_13337,N_10336);
or UO_233 (O_233,N_12927,N_14797);
and UO_234 (O_234,N_13260,N_10835);
nor UO_235 (O_235,N_11563,N_12308);
nor UO_236 (O_236,N_13762,N_10291);
nand UO_237 (O_237,N_14099,N_12101);
xor UO_238 (O_238,N_12100,N_10267);
nor UO_239 (O_239,N_14019,N_13152);
nand UO_240 (O_240,N_13493,N_14695);
xor UO_241 (O_241,N_11918,N_14592);
or UO_242 (O_242,N_10196,N_11820);
and UO_243 (O_243,N_13321,N_12468);
xnor UO_244 (O_244,N_10604,N_11882);
nand UO_245 (O_245,N_11131,N_11091);
nand UO_246 (O_246,N_10429,N_10113);
nand UO_247 (O_247,N_13644,N_11365);
and UO_248 (O_248,N_10377,N_12710);
nor UO_249 (O_249,N_11764,N_10736);
and UO_250 (O_250,N_13161,N_11777);
nor UO_251 (O_251,N_11678,N_10659);
or UO_252 (O_252,N_14849,N_11821);
and UO_253 (O_253,N_13109,N_12388);
and UO_254 (O_254,N_13285,N_12398);
xnor UO_255 (O_255,N_14917,N_14955);
nand UO_256 (O_256,N_10868,N_14369);
xor UO_257 (O_257,N_11774,N_10706);
xnor UO_258 (O_258,N_13151,N_13288);
and UO_259 (O_259,N_14818,N_12480);
or UO_260 (O_260,N_14064,N_10270);
or UO_261 (O_261,N_14482,N_13091);
or UO_262 (O_262,N_10127,N_13256);
nand UO_263 (O_263,N_10888,N_13649);
nand UO_264 (O_264,N_11544,N_14804);
and UO_265 (O_265,N_10685,N_12890);
or UO_266 (O_266,N_13243,N_12717);
and UO_267 (O_267,N_14334,N_13782);
or UO_268 (O_268,N_13837,N_14344);
nor UO_269 (O_269,N_13848,N_10961);
nor UO_270 (O_270,N_12750,N_10165);
nand UO_271 (O_271,N_14697,N_10161);
or UO_272 (O_272,N_14813,N_14346);
or UO_273 (O_273,N_12495,N_11612);
nor UO_274 (O_274,N_12607,N_13024);
xnor UO_275 (O_275,N_12744,N_10911);
and UO_276 (O_276,N_11839,N_14121);
nand UO_277 (O_277,N_11687,N_13958);
or UO_278 (O_278,N_14897,N_13821);
or UO_279 (O_279,N_11239,N_11147);
nor UO_280 (O_280,N_11484,N_11218);
nor UO_281 (O_281,N_11270,N_14098);
nor UO_282 (O_282,N_11713,N_14034);
xnor UO_283 (O_283,N_14021,N_10811);
or UO_284 (O_284,N_10333,N_13772);
nor UO_285 (O_285,N_13539,N_11138);
xor UO_286 (O_286,N_11880,N_11260);
xor UO_287 (O_287,N_10766,N_12452);
xor UO_288 (O_288,N_10922,N_10725);
nor UO_289 (O_289,N_10592,N_14088);
nand UO_290 (O_290,N_10373,N_12128);
or UO_291 (O_291,N_12632,N_12432);
xnor UO_292 (O_292,N_10855,N_12319);
and UO_293 (O_293,N_13888,N_12272);
and UO_294 (O_294,N_13061,N_12018);
nor UO_295 (O_295,N_13375,N_14615);
nand UO_296 (O_296,N_12143,N_13867);
xor UO_297 (O_297,N_10962,N_11220);
or UO_298 (O_298,N_12865,N_12426);
nor UO_299 (O_299,N_12681,N_13715);
or UO_300 (O_300,N_12643,N_11259);
and UO_301 (O_301,N_14237,N_14861);
and UO_302 (O_302,N_10664,N_11822);
xnor UO_303 (O_303,N_12912,N_12208);
xnor UO_304 (O_304,N_12569,N_14046);
and UO_305 (O_305,N_12292,N_12701);
xnor UO_306 (O_306,N_13535,N_14423);
nand UO_307 (O_307,N_14145,N_10110);
and UO_308 (O_308,N_13652,N_14967);
or UO_309 (O_309,N_12730,N_13135);
and UO_310 (O_310,N_10050,N_13235);
and UO_311 (O_311,N_10948,N_10385);
nand UO_312 (O_312,N_13005,N_12788);
nor UO_313 (O_313,N_13833,N_13296);
nand UO_314 (O_314,N_12552,N_13824);
or UO_315 (O_315,N_12528,N_10914);
or UO_316 (O_316,N_14380,N_13770);
xor UO_317 (O_317,N_14275,N_13521);
xor UO_318 (O_318,N_13186,N_14116);
and UO_319 (O_319,N_13370,N_13578);
and UO_320 (O_320,N_14515,N_13816);
nand UO_321 (O_321,N_14992,N_13862);
nor UO_322 (O_322,N_14783,N_12450);
xnor UO_323 (O_323,N_10823,N_11919);
nand UO_324 (O_324,N_12649,N_13609);
or UO_325 (O_325,N_10132,N_11116);
or UO_326 (O_326,N_14709,N_13097);
and UO_327 (O_327,N_12527,N_14299);
xnor UO_328 (O_328,N_12116,N_13955);
nand UO_329 (O_329,N_14252,N_11999);
xnor UO_330 (O_330,N_12787,N_14997);
or UO_331 (O_331,N_13620,N_13128);
nand UO_332 (O_332,N_11082,N_13628);
xnor UO_333 (O_333,N_13495,N_12020);
nand UO_334 (O_334,N_12438,N_10268);
or UO_335 (O_335,N_12133,N_14565);
nor UO_336 (O_336,N_10717,N_13156);
nand UO_337 (O_337,N_11173,N_13064);
xor UO_338 (O_338,N_11856,N_10203);
xor UO_339 (O_339,N_10413,N_12583);
and UO_340 (O_340,N_11343,N_11905);
nor UO_341 (O_341,N_12839,N_13018);
xor UO_342 (O_342,N_13975,N_14235);
or UO_343 (O_343,N_12638,N_11989);
and UO_344 (O_344,N_10882,N_13219);
xor UO_345 (O_345,N_13373,N_13206);
and UO_346 (O_346,N_14994,N_11065);
and UO_347 (O_347,N_14363,N_13585);
nand UO_348 (O_348,N_11474,N_10009);
nand UO_349 (O_349,N_14915,N_12745);
nand UO_350 (O_350,N_12215,N_14282);
nand UO_351 (O_351,N_10248,N_11344);
and UO_352 (O_352,N_14248,N_10578);
or UO_353 (O_353,N_13999,N_14760);
or UO_354 (O_354,N_10784,N_10951);
xnor UO_355 (O_355,N_13819,N_14210);
xor UO_356 (O_356,N_11195,N_12820);
nor UO_357 (O_357,N_13866,N_10083);
and UO_358 (O_358,N_14979,N_14082);
nor UO_359 (O_359,N_13531,N_14406);
or UO_360 (O_360,N_11572,N_10054);
and UO_361 (O_361,N_12386,N_11453);
nor UO_362 (O_362,N_13804,N_11516);
nand UO_363 (O_363,N_14345,N_13224);
xnor UO_364 (O_364,N_14229,N_10952);
nand UO_365 (O_365,N_10003,N_13475);
and UO_366 (O_366,N_11824,N_12471);
nand UO_367 (O_367,N_14706,N_14326);
nor UO_368 (O_368,N_14842,N_12870);
nor UO_369 (O_369,N_14758,N_14430);
nand UO_370 (O_370,N_10739,N_13202);
nor UO_371 (O_371,N_12195,N_11373);
or UO_372 (O_372,N_11706,N_13541);
xnor UO_373 (O_373,N_10445,N_10691);
nor UO_374 (O_374,N_12592,N_11001);
and UO_375 (O_375,N_14876,N_14341);
or UO_376 (O_376,N_14514,N_10589);
xor UO_377 (O_377,N_14550,N_10057);
or UO_378 (O_378,N_12921,N_11469);
and UO_379 (O_379,N_12004,N_12086);
and UO_380 (O_380,N_13730,N_11944);
xor UO_381 (O_381,N_12269,N_10972);
nor UO_382 (O_382,N_10226,N_12474);
nor UO_383 (O_383,N_12737,N_14926);
or UO_384 (O_384,N_10047,N_12577);
nand UO_385 (O_385,N_14884,N_14147);
nor UO_386 (O_386,N_11699,N_13174);
xor UO_387 (O_387,N_10315,N_12142);
nand UO_388 (O_388,N_11426,N_10367);
xnor UO_389 (O_389,N_14291,N_13967);
xnor UO_390 (O_390,N_14902,N_13909);
xnor UO_391 (O_391,N_11133,N_13448);
or UO_392 (O_392,N_14017,N_10117);
and UO_393 (O_393,N_11751,N_14859);
or UO_394 (O_394,N_10170,N_14399);
nand UO_395 (O_395,N_12277,N_12329);
nor UO_396 (O_396,N_14232,N_12515);
and UO_397 (O_397,N_12253,N_11664);
nor UO_398 (O_398,N_10927,N_10096);
or UO_399 (O_399,N_12111,N_14596);
nand UO_400 (O_400,N_12856,N_10302);
xor UO_401 (O_401,N_10319,N_14624);
and UO_402 (O_402,N_13073,N_10360);
nand UO_403 (O_403,N_14176,N_12868);
xnor UO_404 (O_404,N_11712,N_11535);
xnor UO_405 (O_405,N_14644,N_11811);
or UO_406 (O_406,N_14721,N_12052);
xnor UO_407 (O_407,N_14662,N_13752);
and UO_408 (O_408,N_11557,N_14153);
nand UO_409 (O_409,N_10402,N_12791);
xnor UO_410 (O_410,N_13264,N_12917);
nand UO_411 (O_411,N_12227,N_12540);
nand UO_412 (O_412,N_14526,N_10476);
nor UO_413 (O_413,N_12982,N_10929);
nor UO_414 (O_414,N_13217,N_12044);
xnor UO_415 (O_415,N_12107,N_12669);
xor UO_416 (O_416,N_14567,N_13897);
and UO_417 (O_417,N_12605,N_11895);
nor UO_418 (O_418,N_12103,N_10337);
nor UO_419 (O_419,N_12685,N_13695);
or UO_420 (O_420,N_14465,N_13853);
nor UO_421 (O_421,N_13342,N_13863);
and UO_422 (O_422,N_13670,N_11767);
nor UO_423 (O_423,N_10485,N_13538);
nand UO_424 (O_424,N_11779,N_13080);
and UO_425 (O_425,N_12830,N_10853);
and UO_426 (O_426,N_12854,N_12712);
nor UO_427 (O_427,N_14560,N_14556);
nand UO_428 (O_428,N_10982,N_12893);
nor UO_429 (O_429,N_14638,N_13949);
and UO_430 (O_430,N_13079,N_13057);
xnor UO_431 (O_431,N_13550,N_13028);
nor UO_432 (O_432,N_10583,N_10125);
or UO_433 (O_433,N_12819,N_14779);
and UO_434 (O_434,N_12011,N_13978);
xnor UO_435 (O_435,N_11553,N_12358);
xnor UO_436 (O_436,N_14786,N_13892);
nor UO_437 (O_437,N_13020,N_11321);
and UO_438 (O_438,N_14133,N_13696);
and UO_439 (O_439,N_11655,N_10792);
or UO_440 (O_440,N_11925,N_11967);
xor UO_441 (O_441,N_11630,N_13719);
and UO_442 (O_442,N_13433,N_14948);
and UO_443 (O_443,N_10177,N_11167);
nor UO_444 (O_444,N_12493,N_13245);
or UO_445 (O_445,N_12853,N_12816);
and UO_446 (O_446,N_12802,N_11229);
and UO_447 (O_447,N_11555,N_11752);
and UO_448 (O_448,N_10568,N_10813);
xnor UO_449 (O_449,N_14287,N_11730);
or UO_450 (O_450,N_13693,N_10256);
xnor UO_451 (O_451,N_14103,N_14402);
and UO_452 (O_452,N_11978,N_11695);
xnor UO_453 (O_453,N_13605,N_12074);
nor UO_454 (O_454,N_10060,N_14879);
xor UO_455 (O_455,N_11838,N_12351);
xor UO_456 (O_456,N_11665,N_10731);
or UO_457 (O_457,N_11425,N_11738);
nor UO_458 (O_458,N_13875,N_13799);
nor UO_459 (O_459,N_13755,N_11593);
and UO_460 (O_460,N_14415,N_11140);
and UO_461 (O_461,N_14700,N_12821);
nor UO_462 (O_462,N_11487,N_14543);
xnor UO_463 (O_463,N_14737,N_13276);
nand UO_464 (O_464,N_12328,N_11028);
xor UO_465 (O_465,N_11235,N_11224);
nor UO_466 (O_466,N_12798,N_13247);
xor UO_467 (O_467,N_13384,N_10168);
or UO_468 (O_468,N_12489,N_11845);
and UO_469 (O_469,N_11875,N_13056);
nor UO_470 (O_470,N_14546,N_11765);
xor UO_471 (O_471,N_13464,N_11888);
and UO_472 (O_472,N_13376,N_11458);
or UO_473 (O_473,N_13385,N_10654);
nor UO_474 (O_474,N_14140,N_10153);
nor UO_475 (O_475,N_12061,N_11295);
and UO_476 (O_476,N_14853,N_11509);
and UO_477 (O_477,N_10656,N_12048);
xnor UO_478 (O_478,N_10591,N_14355);
nor UO_479 (O_479,N_11074,N_10734);
xor UO_480 (O_480,N_14292,N_14660);
nand UO_481 (O_481,N_11891,N_12586);
nor UO_482 (O_482,N_11543,N_13055);
or UO_483 (O_483,N_11690,N_10830);
xor UO_484 (O_484,N_14540,N_11109);
nand UO_485 (O_485,N_13557,N_11727);
xor UO_486 (O_486,N_11204,N_14612);
xnor UO_487 (O_487,N_10839,N_11561);
nor UO_488 (O_488,N_11413,N_10335);
and UO_489 (O_489,N_11203,N_11141);
and UO_490 (O_490,N_14886,N_11326);
or UO_491 (O_491,N_11067,N_10344);
xnor UO_492 (O_492,N_14190,N_11666);
nor UO_493 (O_493,N_12926,N_10954);
and UO_494 (O_494,N_13732,N_14982);
nand UO_495 (O_495,N_10894,N_10594);
xor UO_496 (O_496,N_14379,N_13094);
nand UO_497 (O_497,N_13754,N_13218);
or UO_498 (O_498,N_11486,N_11222);
or UO_499 (O_499,N_10313,N_13001);
nor UO_500 (O_500,N_13751,N_12168);
nand UO_501 (O_501,N_11421,N_12808);
and UO_502 (O_502,N_12516,N_12790);
nand UO_503 (O_503,N_12370,N_13734);
and UO_504 (O_504,N_10881,N_13424);
nor UO_505 (O_505,N_12709,N_12740);
xor UO_506 (O_506,N_14490,N_14026);
nor UO_507 (O_507,N_13293,N_12205);
and UO_508 (O_508,N_10990,N_14674);
nand UO_509 (O_509,N_13813,N_12647);
nand UO_510 (O_510,N_11886,N_13895);
and UO_511 (O_511,N_14313,N_12301);
nand UO_512 (O_512,N_12742,N_12159);
or UO_513 (O_513,N_14314,N_14701);
or UO_514 (O_514,N_11290,N_13717);
nand UO_515 (O_515,N_13656,N_10964);
or UO_516 (O_516,N_10444,N_14722);
xor UO_517 (O_517,N_10376,N_11198);
nand UO_518 (O_518,N_13885,N_10738);
nand UO_519 (O_519,N_10380,N_11211);
nand UO_520 (O_520,N_11399,N_11936);
or UO_521 (O_521,N_12731,N_12207);
xor UO_522 (O_522,N_13569,N_14940);
nand UO_523 (O_523,N_13124,N_11707);
xor UO_524 (O_524,N_12942,N_14636);
xnor UO_525 (O_525,N_11477,N_12814);
nor UO_526 (O_526,N_14664,N_13954);
or UO_527 (O_527,N_14185,N_13795);
nand UO_528 (O_528,N_12535,N_10832);
or UO_529 (O_529,N_10512,N_14197);
and UO_530 (O_530,N_14602,N_12815);
xnor UO_531 (O_531,N_14010,N_11227);
xnor UO_532 (O_532,N_11804,N_11369);
nor UO_533 (O_533,N_11530,N_14485);
xor UO_534 (O_534,N_11935,N_11975);
or UO_535 (O_535,N_10944,N_14130);
nand UO_536 (O_536,N_13905,N_11533);
nand UO_537 (O_537,N_13265,N_11812);
xor UO_538 (O_538,N_14572,N_12985);
nand UO_539 (O_539,N_10339,N_13913);
or UO_540 (O_540,N_11452,N_11170);
nand UO_541 (O_541,N_14041,N_12418);
nand UO_542 (O_542,N_13200,N_13402);
nand UO_543 (O_543,N_14094,N_14869);
xor UO_544 (O_544,N_13491,N_14078);
and UO_545 (O_545,N_14290,N_12722);
xnor UO_546 (O_546,N_12046,N_10351);
nand UO_547 (O_547,N_10860,N_10661);
and UO_548 (O_548,N_11756,N_12561);
nand UO_549 (O_549,N_14454,N_11657);
xor UO_550 (O_550,N_13017,N_11571);
or UO_551 (O_551,N_14688,N_11191);
and UO_552 (O_552,N_12931,N_13230);
nand UO_553 (O_553,N_11951,N_14337);
xnor UO_554 (O_554,N_10850,N_14396);
and UO_555 (O_555,N_11586,N_12241);
nand UO_556 (O_556,N_10229,N_11325);
nand UO_557 (O_557,N_14188,N_14529);
nand UO_558 (O_558,N_13926,N_11470);
nor UO_559 (O_559,N_12629,N_11759);
nor UO_560 (O_560,N_13830,N_10405);
xnor UO_561 (O_561,N_10896,N_13268);
nor UO_562 (O_562,N_13651,N_12573);
or UO_563 (O_563,N_11776,N_13736);
nor UO_564 (O_564,N_11903,N_12414);
nor UO_565 (O_565,N_12874,N_14825);
xor UO_566 (O_566,N_11931,N_13584);
xor UO_567 (O_567,N_11451,N_11959);
or UO_568 (O_568,N_14460,N_14850);
or UO_569 (O_569,N_12879,N_14983);
and UO_570 (O_570,N_11749,N_13936);
or UO_571 (O_571,N_12244,N_10903);
nand UO_572 (O_572,N_13886,N_14468);
xor UO_573 (O_573,N_10398,N_13991);
nand UO_574 (O_574,N_13372,N_14716);
and UO_575 (O_575,N_12682,N_12919);
xnor UO_576 (O_576,N_10909,N_12677);
xor UO_577 (O_577,N_10865,N_12986);
nand UO_578 (O_578,N_11679,N_10940);
and UO_579 (O_579,N_10827,N_14595);
nand UO_580 (O_580,N_10943,N_11817);
nor UO_581 (O_581,N_14632,N_10688);
xor UO_582 (O_582,N_13921,N_13835);
nor UO_583 (O_583,N_12968,N_11292);
or UO_584 (O_584,N_13279,N_14655);
nand UO_585 (O_585,N_13769,N_13136);
nor UO_586 (O_586,N_11615,N_13441);
nor UO_587 (O_587,N_14057,N_13344);
xor UO_588 (O_588,N_11899,N_13549);
nand UO_589 (O_589,N_11405,N_12733);
or UO_590 (O_590,N_10415,N_11394);
nand UO_591 (O_591,N_13241,N_10087);
nor UO_592 (O_592,N_14011,N_14780);
nor UO_593 (O_593,N_12858,N_12339);
and UO_594 (O_594,N_12178,N_11605);
xor UO_595 (O_595,N_11734,N_12887);
nand UO_596 (O_596,N_11427,N_14535);
nor UO_597 (O_597,N_12179,N_11475);
and UO_598 (O_598,N_11036,N_13607);
xor UO_599 (O_599,N_12436,N_13794);
nor UO_600 (O_600,N_12500,N_13654);
nand UO_601 (O_601,N_13100,N_11285);
or UO_602 (O_602,N_14593,N_11370);
or UO_603 (O_603,N_12841,N_12181);
xnor UO_604 (O_604,N_13723,N_14898);
and UO_605 (O_605,N_13166,N_12262);
and UO_606 (O_606,N_13577,N_12679);
nand UO_607 (O_607,N_13332,N_10858);
nand UO_608 (O_608,N_10126,N_11787);
xor UO_609 (O_609,N_12021,N_14198);
xor UO_610 (O_610,N_14776,N_10379);
nor UO_611 (O_611,N_14675,N_13890);
and UO_612 (O_612,N_11731,N_14184);
nand UO_613 (O_613,N_10513,N_13545);
nor UO_614 (O_614,N_11294,N_14154);
nor UO_615 (O_615,N_10837,N_10763);
xor UO_616 (O_616,N_13971,N_10106);
and UO_617 (O_617,N_12825,N_12444);
or UO_618 (O_618,N_14511,N_14450);
and UO_619 (O_619,N_13718,N_14409);
nand UO_620 (O_620,N_11648,N_10704);
nand UO_621 (O_621,N_11920,N_14777);
and UO_622 (O_622,N_14281,N_11296);
xnor UO_623 (O_623,N_10535,N_14357);
nand UO_624 (O_624,N_13044,N_11139);
and UO_625 (O_625,N_10607,N_10227);
and UO_626 (O_626,N_13275,N_10570);
nor UO_627 (O_627,N_12614,N_13589);
nor UO_628 (O_628,N_10494,N_14141);
and UO_629 (O_629,N_12383,N_11185);
nand UO_630 (O_630,N_14851,N_14392);
nor UO_631 (O_631,N_10985,N_14647);
and UO_632 (O_632,N_12543,N_11954);
xor UO_633 (O_633,N_11153,N_13199);
or UO_634 (O_634,N_13038,N_13690);
or UO_635 (O_635,N_13019,N_14727);
and UO_636 (O_636,N_13291,N_14455);
and UO_637 (O_637,N_10515,N_10793);
and UO_638 (O_638,N_13571,N_14193);
nand UO_639 (O_639,N_10802,N_13568);
nand UO_640 (O_640,N_14887,N_11685);
nand UO_641 (O_641,N_11362,N_12891);
nand UO_642 (O_642,N_13544,N_13436);
nand UO_643 (O_643,N_12877,N_12002);
nand UO_644 (O_644,N_14214,N_12322);
nand UO_645 (O_645,N_12555,N_10035);
nand UO_646 (O_646,N_10810,N_12442);
nand UO_647 (O_647,N_14863,N_14328);
nand UO_648 (O_648,N_10055,N_11390);
nand UO_649 (O_649,N_14245,N_10869);
xnor UO_650 (O_650,N_12421,N_14877);
nand UO_651 (O_651,N_14995,N_13391);
and UO_652 (O_652,N_10791,N_12600);
nor UO_653 (O_653,N_13735,N_13961);
or UO_654 (O_654,N_13553,N_10013);
and UO_655 (O_655,N_13858,N_13561);
xor UO_656 (O_656,N_13108,N_11201);
xnor UO_657 (O_657,N_10966,N_14120);
or UO_658 (O_658,N_14336,N_10201);
xnor UO_659 (O_659,N_10673,N_12741);
nor UO_660 (O_660,N_12309,N_13635);
xnor UO_661 (O_661,N_14268,N_14907);
xnor UO_662 (O_662,N_10984,N_11921);
or UO_663 (O_663,N_14986,N_10005);
and UO_664 (O_664,N_12857,N_13052);
and UO_665 (O_665,N_13315,N_14238);
nor UO_666 (O_666,N_13071,N_12078);
nand UO_667 (O_667,N_12041,N_14016);
xor UO_668 (O_668,N_14169,N_13685);
xnor UO_669 (O_669,N_12300,N_12156);
nand UO_670 (O_670,N_14741,N_12040);
xor UO_671 (O_671,N_14014,N_12892);
and UO_672 (O_672,N_10683,N_14186);
nor UO_673 (O_673,N_12509,N_10421);
xnor UO_674 (O_674,N_12249,N_10593);
xnor UO_675 (O_675,N_12780,N_14785);
xor UO_676 (O_676,N_11302,N_12823);
xor UO_677 (O_677,N_11828,N_13294);
xnor UO_678 (O_678,N_10816,N_12302);
nor UO_679 (O_679,N_10871,N_12861);
or UO_680 (O_680,N_11570,N_10042);
xnor UO_681 (O_681,N_14394,N_12959);
nand UO_682 (O_682,N_11034,N_11423);
nand UO_683 (O_683,N_10926,N_14870);
xnor UO_684 (O_684,N_11156,N_13350);
and UO_685 (O_685,N_14484,N_14505);
or UO_686 (O_686,N_10257,N_12005);
xnor UO_687 (O_687,N_13706,N_11314);
xnor UO_688 (O_688,N_11176,N_14909);
nor UO_689 (O_689,N_14348,N_10028);
nor UO_690 (O_690,N_12224,N_14166);
nor UO_691 (O_691,N_12704,N_12807);
and UO_692 (O_692,N_10046,N_13478);
nand UO_693 (O_693,N_13879,N_10775);
nand UO_694 (O_694,N_12034,N_10450);
xnor UO_695 (O_695,N_13697,N_10453);
xnor UO_696 (O_696,N_14561,N_11374);
nand UO_697 (O_697,N_10304,N_12772);
nand UO_698 (O_698,N_13570,N_10979);
xnor UO_699 (O_699,N_13773,N_10343);
nand UO_700 (O_700,N_12496,N_10680);
xnor UO_701 (O_701,N_14824,N_12394);
nor UO_702 (O_702,N_10560,N_12165);
or UO_703 (O_703,N_10278,N_14814);
nand UO_704 (O_704,N_12898,N_12035);
and UO_705 (O_705,N_13249,N_14847);
nor UO_706 (O_706,N_10123,N_11410);
or UO_707 (O_707,N_13882,N_13148);
and UO_708 (O_708,N_13789,N_13209);
nand UO_709 (O_709,N_14381,N_12463);
nand UO_710 (O_710,N_11743,N_14312);
xor UO_711 (O_711,N_10076,N_12449);
and UO_712 (O_712,N_12477,N_13631);
xor UO_713 (O_713,N_10987,N_13601);
nand UO_714 (O_714,N_11275,N_10085);
xor UO_715 (O_715,N_13051,N_10511);
nor UO_716 (O_716,N_13394,N_11221);
and UO_717 (O_717,N_11054,N_12829);
xnor UO_718 (O_718,N_12146,N_12956);
nand UO_719 (O_719,N_13576,N_14023);
xnor UO_720 (O_720,N_11581,N_11667);
nand UO_721 (O_721,N_11806,N_12661);
or UO_722 (O_722,N_11843,N_12067);
or UO_723 (O_723,N_12289,N_12424);
and UO_724 (O_724,N_10743,N_14244);
and UO_725 (O_725,N_10130,N_14440);
xnor UO_726 (O_726,N_14642,N_10255);
or UO_727 (O_727,N_14092,N_14510);
nand UO_728 (O_728,N_13425,N_12186);
or UO_729 (O_729,N_14650,N_12361);
or UO_730 (O_730,N_11741,N_10104);
and UO_731 (O_731,N_11022,N_12526);
xor UO_732 (O_732,N_14331,N_11656);
or UO_733 (O_733,N_14178,N_10259);
nand UO_734 (O_734,N_12381,N_13089);
nand UO_735 (O_735,N_14412,N_12357);
nand UO_736 (O_736,N_12624,N_14488);
or UO_737 (O_737,N_10140,N_13743);
nor UO_738 (O_738,N_14429,N_11075);
and UO_739 (O_739,N_13234,N_14845);
nand UO_740 (O_740,N_13639,N_12633);
nand UO_741 (O_741,N_11696,N_13758);
nor UO_742 (O_742,N_12690,N_14690);
nand UO_743 (O_743,N_11654,N_11092);
and UO_744 (O_744,N_11829,N_13334);
xnor UO_745 (O_745,N_10668,N_13998);
nand UO_746 (O_746,N_11233,N_14927);
nor UO_747 (O_747,N_12311,N_13415);
xnor UO_748 (O_748,N_14439,N_10086);
and UO_749 (O_749,N_13780,N_11305);
xnor UO_750 (O_750,N_13849,N_14359);
nand UO_751 (O_751,N_10974,N_14712);
nor UO_752 (O_752,N_12746,N_14131);
and UO_753 (O_753,N_11651,N_11783);
and UO_754 (O_754,N_14300,N_13800);
and UO_755 (O_755,N_13320,N_13366);
or UO_756 (O_756,N_13588,N_12625);
nand UO_757 (O_757,N_12571,N_11266);
and UO_758 (O_758,N_14766,N_13522);
nor UO_759 (O_759,N_13945,N_10626);
nand UO_760 (O_760,N_10624,N_11818);
nor UO_761 (O_761,N_13257,N_10744);
xnor UO_762 (O_762,N_12127,N_14213);
and UO_763 (O_763,N_14246,N_13070);
nor UO_764 (O_764,N_14521,N_13744);
nand UO_765 (O_765,N_14207,N_13119);
nand UO_766 (O_766,N_11893,N_13013);
or UO_767 (O_767,N_11448,N_14476);
xor UO_768 (O_768,N_13413,N_13793);
or UO_769 (O_769,N_14044,N_11640);
xnor UO_770 (O_770,N_10608,N_10352);
xor UO_771 (O_771,N_10058,N_13040);
xnor UO_772 (O_772,N_10006,N_12824);
and UO_773 (O_773,N_14466,N_10027);
and UO_774 (O_774,N_14228,N_12619);
xnor UO_775 (O_775,N_14754,N_14306);
nor UO_776 (O_776,N_11024,N_13707);
and UO_777 (O_777,N_11789,N_10391);
nor UO_778 (O_778,N_11980,N_12822);
xor UO_779 (O_779,N_14264,N_10671);
nand UO_780 (O_780,N_11653,N_13043);
and UO_781 (O_781,N_11748,N_14933);
nor UO_782 (O_782,N_14968,N_12187);
nor UO_783 (O_783,N_13339,N_14135);
xor UO_784 (O_784,N_14384,N_12170);
nor UO_785 (O_785,N_13917,N_14493);
and UO_786 (O_786,N_14685,N_11591);
nand UO_787 (O_787,N_13144,N_13748);
or UO_788 (O_788,N_13201,N_13621);
or UO_789 (O_789,N_14732,N_14069);
nor UO_790 (O_790,N_11346,N_12659);
and UO_791 (O_791,N_10887,N_13927);
nor UO_792 (O_792,N_12169,N_14205);
and UO_793 (O_793,N_14681,N_14963);
or UO_794 (O_794,N_12538,N_12448);
or UO_795 (O_795,N_11068,N_11733);
nor UO_796 (O_796,N_14260,N_10030);
nor UO_797 (O_797,N_11014,N_10508);
nor UO_798 (O_798,N_10950,N_10089);
and UO_799 (O_799,N_11379,N_14072);
nand UO_800 (O_800,N_12777,N_12226);
and UO_801 (O_801,N_14124,N_10088);
xnor UO_802 (O_802,N_14218,N_13543);
and UO_803 (O_803,N_13360,N_14970);
or UO_804 (O_804,N_13904,N_12562);
and UO_805 (O_805,N_13855,N_11125);
nor UO_806 (O_806,N_14134,N_10710);
and UO_807 (O_807,N_10399,N_10625);
nor UO_808 (O_808,N_13555,N_13783);
nor UO_809 (O_809,N_10084,N_11879);
and UO_810 (O_810,N_10797,N_11622);
and UO_811 (O_811,N_11441,N_11083);
or UO_812 (O_812,N_14435,N_13629);
nor UO_813 (O_813,N_10199,N_13127);
or UO_814 (O_814,N_13326,N_11108);
or UO_815 (O_815,N_14113,N_14874);
and UO_816 (O_816,N_13367,N_10401);
xnor UO_817 (O_817,N_10945,N_11154);
nor UO_818 (O_818,N_10782,N_10427);
or UO_819 (O_819,N_10455,N_13509);
xnor UO_820 (O_820,N_11684,N_12539);
xnor UO_821 (O_821,N_13041,N_12989);
nor UO_822 (O_822,N_12055,N_14993);
xor UO_823 (O_823,N_11528,N_12063);
nor UO_824 (O_824,N_12729,N_12779);
xnor UO_825 (O_825,N_11237,N_10416);
or UO_826 (O_826,N_10438,N_11248);
xnor UO_827 (O_827,N_13253,N_14431);
and UO_828 (O_828,N_13171,N_10579);
nand UO_829 (O_829,N_13232,N_12306);
nor UO_830 (O_830,N_14799,N_12920);
or UO_831 (O_831,N_10277,N_13428);
xnor UO_832 (O_832,N_12770,N_11313);
nand UO_833 (O_833,N_14164,N_10675);
xnor UO_834 (O_834,N_11897,N_12160);
nor UO_835 (O_835,N_12431,N_12797);
nand UO_836 (O_836,N_11585,N_11077);
nor UO_837 (O_837,N_11700,N_11368);
nor UO_838 (O_838,N_13062,N_12786);
nor UO_839 (O_839,N_12978,N_11409);
nor UO_840 (O_840,N_12479,N_14551);
xnor UO_841 (O_841,N_11513,N_14945);
and UO_842 (O_842,N_14952,N_12095);
nor UO_843 (O_843,N_13298,N_12768);
and UO_844 (O_844,N_12219,N_11178);
and UO_845 (O_845,N_12852,N_10279);
nand UO_846 (O_846,N_13887,N_14463);
nand UO_847 (O_847,N_14890,N_11909);
nor UO_848 (O_848,N_11311,N_14227);
nor UO_849 (O_849,N_13606,N_10849);
and UO_850 (O_850,N_14835,N_14321);
xor UO_851 (O_851,N_10527,N_10939);
nor UO_852 (O_852,N_13248,N_11337);
or UO_853 (O_853,N_10469,N_14937);
nor UO_854 (O_854,N_11660,N_12944);
and UO_855 (O_855,N_12428,N_10682);
xor UO_856 (O_856,N_14385,N_12131);
or UO_857 (O_857,N_10462,N_11910);
and UO_858 (O_858,N_14137,N_11473);
xor UO_859 (O_859,N_10634,N_13102);
and UO_860 (O_860,N_12288,N_14942);
nor UO_861 (O_861,N_10386,N_12384);
nor UO_862 (O_862,N_13873,N_10166);
or UO_863 (O_863,N_10590,N_13021);
nand UO_864 (O_864,N_11440,N_11805);
xor UO_865 (O_865,N_13412,N_10056);
xor UO_866 (O_866,N_11300,N_13225);
and UO_867 (O_867,N_12403,N_10052);
nor UO_868 (O_868,N_12060,N_12617);
or UO_869 (O_869,N_14668,N_13766);
or UO_870 (O_870,N_13411,N_11432);
xnor UO_871 (O_871,N_14427,N_14930);
xnor UO_872 (O_872,N_11626,N_14990);
or UO_873 (O_873,N_10864,N_12545);
nand UO_874 (O_874,N_12102,N_10960);
nor UO_875 (O_875,N_14318,N_13922);
and UO_876 (O_876,N_11979,N_13145);
and UO_877 (O_877,N_10156,N_14910);
nand UO_878 (O_878,N_12099,N_12091);
nor UO_879 (O_879,N_12557,N_14966);
xor UO_880 (O_880,N_12245,N_10449);
xnor UO_881 (O_881,N_13208,N_13517);
nor UO_882 (O_882,N_12026,N_12375);
and UO_883 (O_883,N_11043,N_13933);
and UO_884 (O_884,N_12957,N_11580);
nor UO_885 (O_885,N_13307,N_13623);
nand UO_886 (O_886,N_11263,N_13768);
and UO_887 (O_887,N_11255,N_11836);
and UO_888 (O_888,N_10474,N_14503);
nand UO_889 (O_889,N_12123,N_13378);
or UO_890 (O_890,N_14478,N_13671);
nand UO_891 (O_891,N_10019,N_11934);
xor UO_892 (O_892,N_12517,N_14559);
nand UO_893 (O_893,N_10600,N_10872);
xor UO_894 (O_894,N_11524,N_11000);
and UO_895 (O_895,N_12747,N_12732);
nor UO_896 (O_896,N_12088,N_12894);
xnor UO_897 (O_897,N_14191,N_13724);
and UO_898 (O_898,N_14486,N_13434);
nor UO_899 (O_899,N_11624,N_12234);
nor UO_900 (O_900,N_12924,N_12121);
xor UO_901 (O_901,N_11984,N_14212);
and UO_902 (O_902,N_11792,N_14714);
nand UO_903 (O_903,N_10024,N_10510);
nor UO_904 (O_904,N_10917,N_12189);
nand UO_905 (O_905,N_13672,N_13042);
or UO_906 (O_906,N_10187,N_10544);
nor UO_907 (O_907,N_12645,N_10546);
nor UO_908 (O_908,N_11631,N_11438);
and UO_909 (O_909,N_11923,N_12446);
xnor UO_910 (O_910,N_13393,N_11002);
or UO_911 (O_911,N_10697,N_12216);
xor UO_912 (O_912,N_12588,N_13586);
or UO_913 (O_913,N_11119,N_14395);
and UO_914 (O_914,N_10708,N_10532);
or UO_915 (O_915,N_10750,N_14972);
and UO_916 (O_916,N_11341,N_11320);
and UO_917 (O_917,N_12009,N_11702);
xor UO_918 (O_918,N_13346,N_11519);
and UO_919 (O_919,N_12027,N_11889);
nor UO_920 (O_920,N_12014,N_12120);
or UO_921 (O_921,N_12939,N_11913);
nand UO_922 (O_922,N_10597,N_11261);
nand UO_923 (O_923,N_11575,N_12655);
nand UO_924 (O_924,N_13611,N_13329);
nor UO_925 (O_925,N_11864,N_10724);
xor UO_926 (O_926,N_14152,N_10540);
or UO_927 (O_927,N_10804,N_10262);
nor UO_928 (O_928,N_10773,N_14578);
or UO_929 (O_929,N_13637,N_14699);
nand UO_930 (O_930,N_12419,N_11272);
nand UO_931 (O_931,N_10000,N_14987);
xnor UO_932 (O_932,N_11431,N_11046);
nor UO_933 (O_933,N_13986,N_10439);
nand UO_934 (O_934,N_10374,N_10551);
or UO_935 (O_935,N_11032,N_14165);
nor UO_936 (O_936,N_12353,N_10795);
nor UO_937 (O_937,N_10149,N_14277);
xor UO_938 (O_938,N_12610,N_11573);
or UO_939 (O_939,N_13000,N_11286);
nor UO_940 (O_940,N_12345,N_12458);
and UO_941 (O_941,N_13430,N_10573);
nor UO_942 (O_942,N_14743,N_13924);
and UO_943 (O_943,N_11577,N_13112);
or UO_944 (O_944,N_10992,N_13829);
and UO_945 (O_945,N_13454,N_14599);
or UO_946 (O_946,N_14839,N_12611);
or UO_947 (O_947,N_10670,N_10892);
xnor UO_948 (O_948,N_10495,N_10417);
nor UO_949 (O_949,N_12544,N_13067);
nand UO_950 (O_950,N_11600,N_12721);
and UO_951 (O_951,N_14060,N_11791);
nor UO_952 (O_952,N_14215,N_13304);
nor UO_953 (O_953,N_11401,N_10996);
or UO_954 (O_954,N_12209,N_13343);
nor UO_955 (O_955,N_13220,N_14102);
xor UO_956 (O_956,N_10239,N_11604);
nor UO_957 (O_957,N_14136,N_11055);
and UO_958 (O_958,N_14547,N_14031);
and UO_959 (O_959,N_10293,N_13636);
nor UO_960 (O_960,N_14342,N_10375);
or UO_961 (O_961,N_10210,N_14748);
nand UO_962 (O_962,N_11192,N_10014);
nor UO_963 (O_963,N_10488,N_12578);
nor UO_964 (O_964,N_14725,N_10520);
or UO_965 (O_965,N_12631,N_11725);
and UO_966 (O_966,N_11835,N_11985);
and UO_967 (O_967,N_14802,N_13322);
xor UO_968 (O_968,N_14368,N_10765);
xnor UO_969 (O_969,N_11596,N_11737);
xor UO_970 (O_970,N_13286,N_11873);
xnor UO_971 (O_971,N_13727,N_14170);
nor UO_972 (O_972,N_14383,N_11349);
nand UO_973 (O_973,N_14095,N_14555);
and UO_974 (O_974,N_10753,N_14631);
and UO_975 (O_975,N_13037,N_12867);
and UO_976 (O_976,N_13969,N_11736);
or UO_977 (O_977,N_11911,N_14457);
xnor UO_978 (O_978,N_13274,N_14254);
nand UO_979 (O_979,N_14319,N_13439);
xnor UO_980 (O_980,N_14703,N_13579);
and UO_981 (O_981,N_14183,N_10755);
or UO_982 (O_982,N_10957,N_13211);
nor UO_983 (O_983,N_10409,N_11051);
xor UO_984 (O_984,N_13952,N_12434);
nor UO_985 (O_985,N_13036,N_14871);
and UO_986 (O_986,N_12720,N_12714);
nand UO_987 (O_987,N_10418,N_10164);
and UO_988 (O_988,N_10666,N_11926);
nand UO_989 (O_989,N_10312,N_14679);
xnor UO_990 (O_990,N_13982,N_13540);
and UO_991 (O_991,N_12298,N_13870);
nand UO_992 (O_992,N_14445,N_13523);
nor UO_993 (O_993,N_12996,N_11522);
nor UO_994 (O_994,N_14025,N_13946);
or UO_995 (O_995,N_11844,N_12587);
and UO_996 (O_996,N_13348,N_11186);
nand UO_997 (O_997,N_14067,N_11610);
xnor UO_998 (O_998,N_10910,N_13506);
or UO_999 (O_999,N_14654,N_11550);
and UO_1000 (O_1000,N_13914,N_12971);
xnor UO_1001 (O_1001,N_14285,N_13625);
nor UO_1002 (O_1002,N_14956,N_14944);
and UO_1003 (O_1003,N_14637,N_13242);
nor UO_1004 (O_1004,N_12064,N_10679);
nor UO_1005 (O_1005,N_13617,N_14199);
and UO_1006 (O_1006,N_14464,N_13368);
and UO_1007 (O_1007,N_14491,N_13494);
or UO_1008 (O_1008,N_12542,N_14387);
nand UO_1009 (O_1009,N_13563,N_13187);
or UO_1010 (O_1010,N_11537,N_10821);
or UO_1011 (O_1011,N_10859,N_13942);
nand UO_1012 (O_1012,N_10938,N_10491);
and UO_1013 (O_1013,N_10768,N_10234);
xor UO_1014 (O_1014,N_14639,N_13002);
or UO_1015 (O_1015,N_10472,N_14989);
and UO_1016 (O_1016,N_14817,N_13785);
xor UO_1017 (O_1017,N_13386,N_11771);
xor UO_1018 (O_1018,N_11006,N_12935);
nand UO_1019 (O_1019,N_13212,N_12413);
nand UO_1020 (O_1020,N_10191,N_14250);
and UO_1021 (O_1021,N_10531,N_11813);
nand UO_1022 (O_1022,N_13657,N_11115);
and UO_1023 (O_1023,N_11896,N_10321);
or UO_1024 (O_1024,N_11683,N_12203);
and UO_1025 (O_1025,N_13903,N_14343);
or UO_1026 (O_1026,N_11625,N_11740);
or UO_1027 (O_1027,N_12443,N_12826);
and UO_1028 (O_1028,N_11766,N_13684);
and UO_1029 (O_1029,N_12783,N_13289);
xnor UO_1030 (O_1030,N_12490,N_14070);
and UO_1031 (O_1031,N_14894,N_10808);
and UO_1032 (O_1032,N_12364,N_13198);
xor UO_1033 (O_1033,N_12420,N_11193);
xnor UO_1034 (O_1034,N_12232,N_10460);
nand UO_1035 (O_1035,N_13869,N_10245);
xnor UO_1036 (O_1036,N_11271,N_10610);
nor UO_1037 (O_1037,N_14747,N_12568);
xor UO_1038 (O_1038,N_10081,N_10475);
xnor UO_1039 (O_1039,N_13937,N_13594);
nand UO_1040 (O_1040,N_10748,N_14784);
xnor UO_1041 (O_1041,N_14516,N_14071);
xnor UO_1042 (O_1042,N_14083,N_13059);
nand UO_1043 (O_1043,N_14557,N_14677);
nand UO_1044 (O_1044,N_12532,N_12278);
nor UO_1045 (O_1045,N_10236,N_12466);
xor UO_1046 (O_1046,N_13900,N_10163);
nand UO_1047 (O_1047,N_10545,N_10252);
or UO_1048 (O_1048,N_10393,N_11621);
nand UO_1049 (O_1049,N_11329,N_11111);
and UO_1050 (O_1050,N_14620,N_10719);
xor UO_1051 (O_1051,N_12907,N_12073);
nand UO_1052 (O_1052,N_14759,N_10015);
or UO_1053 (O_1053,N_12514,N_13966);
or UO_1054 (O_1054,N_13355,N_11523);
xnor UO_1055 (O_1055,N_11151,N_14507);
or UO_1056 (O_1056,N_13559,N_11869);
nand UO_1057 (O_1057,N_11823,N_13364);
nor UO_1058 (O_1058,N_13058,N_10507);
and UO_1059 (O_1059,N_14413,N_12748);
nand UO_1060 (O_1060,N_11658,N_13261);
nand UO_1061 (O_1061,N_11592,N_10189);
or UO_1062 (O_1062,N_10751,N_13665);
nor UO_1063 (O_1063,N_11861,N_11862);
or UO_1064 (O_1064,N_11746,N_12363);
and UO_1065 (O_1065,N_11868,N_12675);
xor UO_1066 (O_1066,N_14039,N_14294);
or UO_1067 (O_1067,N_11102,N_11565);
nand UO_1068 (O_1068,N_12007,N_13466);
or UO_1069 (O_1069,N_12837,N_14226);
xnor UO_1070 (O_1070,N_12766,N_12284);
or UO_1071 (O_1071,N_14339,N_10836);
or UO_1072 (O_1072,N_12447,N_10920);
nor UO_1073 (O_1073,N_12533,N_13807);
xnor UO_1074 (O_1074,N_10499,N_12402);
and UO_1075 (O_1075,N_14973,N_11418);
xnor UO_1076 (O_1076,N_11852,N_12334);
and UO_1077 (O_1077,N_12548,N_14255);
xor UO_1078 (O_1078,N_10102,N_13313);
xnor UO_1079 (O_1079,N_11042,N_11415);
and UO_1080 (O_1080,N_12270,N_10788);
and UO_1081 (O_1081,N_13857,N_10770);
or UO_1082 (O_1082,N_12070,N_10023);
and UO_1083 (O_1083,N_13663,N_13420);
and UO_1084 (O_1084,N_11576,N_13844);
nor UO_1085 (O_1085,N_10200,N_10454);
or UO_1086 (O_1086,N_12953,N_11556);
or UO_1087 (O_1087,N_12368,N_10064);
and UO_1088 (O_1088,N_13808,N_14746);
nor UO_1089 (O_1089,N_14453,N_11045);
and UO_1090 (O_1090,N_12377,N_12281);
nor UO_1091 (O_1091,N_11393,N_10524);
nand UO_1092 (O_1092,N_12771,N_11847);
nor UO_1093 (O_1093,N_14148,N_10638);
or UO_1094 (O_1094,N_13641,N_11428);
nand UO_1095 (O_1095,N_11249,N_11352);
and UO_1096 (O_1096,N_12469,N_12806);
nand UO_1097 (O_1097,N_14050,N_14174);
or UO_1098 (O_1098,N_11035,N_10183);
and UO_1099 (O_1099,N_14729,N_11619);
nor UO_1100 (O_1100,N_11617,N_12981);
xnor UO_1101 (O_1101,N_11902,N_11120);
nand UO_1102 (O_1102,N_14795,N_14374);
nand UO_1103 (O_1103,N_10362,N_12246);
and UO_1104 (O_1104,N_12492,N_14263);
nand UO_1105 (O_1105,N_11304,N_12117);
or UO_1106 (O_1106,N_13881,N_12910);
or UO_1107 (O_1107,N_14623,N_13371);
or UO_1108 (O_1108,N_10905,N_11007);
xor UO_1109 (O_1109,N_11037,N_14447);
xnor UO_1110 (O_1110,N_14881,N_13131);
or UO_1111 (O_1111,N_12537,N_12950);
and UO_1112 (O_1112,N_10672,N_11496);
xor UO_1113 (O_1113,N_11277,N_11408);
nor UO_1114 (O_1114,N_13403,N_11101);
nor UO_1115 (O_1115,N_10674,N_13195);
nor UO_1116 (O_1116,N_13929,N_10032);
nor UO_1117 (O_1117,N_10899,N_12373);
or UO_1118 (O_1118,N_12332,N_13988);
nand UO_1119 (O_1119,N_10968,N_13959);
and UO_1120 (O_1120,N_10045,N_11348);
xnor UO_1121 (O_1121,N_10365,N_11939);
or UO_1122 (O_1122,N_14601,N_14508);
xor UO_1123 (O_1123,N_11994,N_10973);
and UO_1124 (O_1124,N_11171,N_12593);
nand UO_1125 (O_1125,N_13388,N_11795);
xor UO_1126 (O_1126,N_12415,N_14946);
and UO_1127 (O_1127,N_11507,N_12945);
and UO_1128 (O_1128,N_12558,N_13101);
and UO_1129 (O_1129,N_13103,N_11069);
xor UO_1130 (O_1130,N_12085,N_10271);
or UO_1131 (O_1131,N_11376,N_10134);
and UO_1132 (O_1132,N_10181,N_11086);
or UO_1133 (O_1133,N_11594,N_14495);
xor UO_1134 (O_1134,N_14122,N_12735);
nor UO_1135 (O_1135,N_11768,N_12276);
xor UO_1136 (O_1136,N_13939,N_10029);
xor UO_1137 (O_1137,N_10772,N_11906);
xor UO_1138 (O_1138,N_12023,N_12960);
nand UO_1139 (O_1139,N_13642,N_12125);
nor UO_1140 (O_1140,N_10662,N_13533);
or UO_1141 (O_1141,N_13336,N_11389);
or UO_1142 (O_1142,N_11284,N_11866);
xnor UO_1143 (O_1143,N_13908,N_11072);
nor UO_1144 (O_1144,N_10167,N_10780);
and UO_1145 (O_1145,N_12899,N_14670);
xnor UO_1146 (O_1146,N_14687,N_10555);
nor UO_1147 (O_1147,N_11183,N_13786);
and UO_1148 (O_1148,N_11682,N_11602);
and UO_1149 (O_1149,N_10002,N_12698);
and UO_1150 (O_1150,N_10959,N_11597);
or UO_1151 (O_1151,N_12238,N_11762);
xor UO_1152 (O_1152,N_10390,N_11377);
and UO_1153 (O_1153,N_11536,N_12248);
xnor UO_1154 (O_1154,N_11574,N_11668);
nor UO_1155 (O_1155,N_14742,N_11244);
or UO_1156 (O_1156,N_14157,N_14350);
and UO_1157 (O_1157,N_13237,N_13872);
nand UO_1158 (O_1158,N_13860,N_11801);
nor UO_1159 (O_1159,N_13185,N_13492);
xor UO_1160 (O_1160,N_13526,N_11645);
nand UO_1161 (O_1161,N_11219,N_13778);
nor UO_1162 (O_1162,N_13992,N_14329);
nor UO_1163 (O_1163,N_13767,N_11995);
nor UO_1164 (O_1164,N_14569,N_13050);
nand UO_1165 (O_1165,N_12803,N_12905);
nor UO_1166 (O_1166,N_12530,N_10218);
or UO_1167 (O_1167,N_11053,N_10645);
or UO_1168 (O_1168,N_12684,N_11510);
and UO_1169 (O_1169,N_14469,N_10240);
and UO_1170 (O_1170,N_13811,N_13500);
nor UO_1171 (O_1171,N_13790,N_13031);
nor UO_1172 (O_1172,N_13915,N_10212);
nor UO_1173 (O_1173,N_12001,N_14579);
nand UO_1174 (O_1174,N_13074,N_10509);
xor UO_1175 (O_1175,N_13456,N_12974);
and UO_1176 (O_1176,N_14407,N_10289);
nor UO_1177 (O_1177,N_13515,N_13597);
xnor UO_1178 (O_1178,N_14896,N_11819);
or UO_1179 (O_1179,N_11688,N_11541);
and UO_1180 (O_1180,N_11135,N_13943);
or UO_1181 (O_1181,N_13180,N_12713);
and UO_1182 (O_1182,N_12805,N_10447);
nor UO_1183 (O_1183,N_11162,N_12671);
nor UO_1184 (O_1184,N_13250,N_11250);
and UO_1185 (O_1185,N_10378,N_10026);
or UO_1186 (O_1186,N_11366,N_12217);
nand UO_1187 (O_1187,N_10310,N_14417);
nor UO_1188 (O_1188,N_12236,N_12254);
and UO_1189 (O_1189,N_14904,N_12554);
or UO_1190 (O_1190,N_13883,N_12753);
nor UO_1191 (O_1191,N_13352,N_11877);
xnor UO_1192 (O_1192,N_13121,N_13047);
nand UO_1193 (O_1193,N_11842,N_12182);
nor UO_1194 (O_1194,N_14309,N_13556);
or UO_1195 (O_1195,N_11161,N_10947);
nor UO_1196 (O_1196,N_11761,N_12042);
nor UO_1197 (O_1197,N_10967,N_11087);
xnor UO_1198 (O_1198,N_11061,N_10737);
nor UO_1199 (O_1199,N_10740,N_12473);
xor UO_1200 (O_1200,N_13616,N_10155);
or UO_1201 (O_1201,N_11407,N_12016);
and UO_1202 (O_1202,N_14693,N_14872);
xor UO_1203 (O_1203,N_11494,N_13598);
xnor UO_1204 (O_1204,N_10222,N_12441);
nor UO_1205 (O_1205,N_11587,N_10061);
and UO_1206 (O_1206,N_10072,N_12895);
and UO_1207 (O_1207,N_12250,N_14456);
xnor UO_1208 (O_1208,N_12201,N_14051);
xnor UO_1209 (O_1209,N_10284,N_12754);
or UO_1210 (O_1210,N_14123,N_11350);
and UO_1211 (O_1211,N_14168,N_14643);
nand UO_1212 (O_1212,N_12451,N_12237);
and UO_1213 (O_1213,N_14258,N_12758);
or UO_1214 (O_1214,N_10251,N_11381);
or UO_1215 (O_1215,N_13481,N_12399);
nand UO_1216 (O_1216,N_10368,N_14086);
xor UO_1217 (O_1217,N_13169,N_13884);
nor UO_1218 (O_1218,N_14922,N_12487);
and UO_1219 (O_1219,N_13615,N_14097);
and UO_1220 (O_1220,N_11508,N_12362);
and UO_1221 (O_1221,N_13667,N_10921);
or UO_1222 (O_1222,N_14830,N_14311);
and UO_1223 (O_1223,N_14711,N_14167);
xnor UO_1224 (O_1224,N_10712,N_12172);
and UO_1225 (O_1225,N_11659,N_10991);
nor UO_1226 (O_1226,N_11110,N_11267);
and UO_1227 (O_1227,N_13049,N_13048);
nor UO_1228 (O_1228,N_12425,N_10906);
and UO_1229 (O_1229,N_11165,N_12129);
nand UO_1230 (O_1230,N_11987,N_12132);
or UO_1231 (O_1231,N_12833,N_11650);
nor UO_1232 (O_1232,N_11158,N_14880);
or UO_1233 (O_1233,N_12761,N_12756);
and UO_1234 (O_1234,N_10623,N_14789);
or UO_1235 (O_1235,N_10194,N_10904);
nor UO_1236 (O_1236,N_12784,N_13330);
or UO_1237 (O_1237,N_11406,N_10235);
nand UO_1238 (O_1238,N_14520,N_12343);
nor UO_1239 (O_1239,N_11907,N_13907);
nor UO_1240 (O_1240,N_14913,N_14969);
or UO_1241 (O_1241,N_12470,N_10820);
and UO_1242 (O_1242,N_12029,N_14745);
xor UO_1243 (O_1243,N_10108,N_13562);
nand UO_1244 (O_1244,N_11402,N_10602);
or UO_1245 (O_1245,N_10354,N_14819);
xor UO_1246 (O_1246,N_12460,N_10707);
and UO_1247 (O_1247,N_14012,N_12863);
or UO_1248 (O_1248,N_11932,N_12349);
nand UO_1249 (O_1249,N_12550,N_12153);
nor UO_1250 (O_1250,N_14114,N_11957);
nor UO_1251 (O_1251,N_10534,N_13381);
nand UO_1252 (O_1252,N_13305,N_11005);
xnor UO_1253 (O_1253,N_13299,N_11003);
xnor UO_1254 (O_1254,N_12003,N_14576);
or UO_1255 (O_1255,N_13314,N_10629);
xnor UO_1256 (O_1256,N_11446,N_10901);
nor UO_1257 (O_1257,N_14364,N_10044);
nor UO_1258 (O_1258,N_10160,N_11834);
xor UO_1259 (O_1259,N_10331,N_13068);
and UO_1260 (O_1260,N_11965,N_12106);
or UO_1261 (O_1261,N_13733,N_11412);
and UO_1262 (O_1262,N_11492,N_12832);
nand UO_1263 (O_1263,N_14441,N_10616);
or UO_1264 (O_1264,N_11160,N_11318);
nor UO_1265 (O_1265,N_12992,N_10484);
or UO_1266 (O_1266,N_14217,N_12876);
or UO_1267 (O_1267,N_10714,N_14504);
xor UO_1268 (O_1268,N_14461,N_12497);
xor UO_1269 (O_1269,N_13703,N_14549);
nand UO_1270 (O_1270,N_13674,N_13455);
or UO_1271 (O_1271,N_13233,N_11499);
nand UO_1272 (O_1272,N_10071,N_13817);
and UO_1273 (O_1273,N_13474,N_11306);
and UO_1274 (O_1274,N_13676,N_12567);
nand UO_1275 (O_1275,N_10848,N_13516);
nor UO_1276 (O_1276,N_14408,N_12518);
nor UO_1277 (O_1277,N_14194,N_10758);
nand UO_1278 (O_1278,N_11287,N_12094);
nor UO_1279 (O_1279,N_13006,N_12627);
and UO_1280 (O_1280,N_12378,N_12664);
xnor UO_1281 (O_1281,N_11240,N_13069);
nand UO_1282 (O_1282,N_14272,N_10705);
and UO_1283 (O_1283,N_10556,N_14985);
nand UO_1284 (O_1284,N_10912,N_11890);
or UO_1285 (O_1285,N_10261,N_13661);
and UO_1286 (O_1286,N_13392,N_13027);
nand UO_1287 (O_1287,N_11865,N_14548);
nand UO_1288 (O_1288,N_14924,N_12653);
nand UO_1289 (O_1289,N_14698,N_10138);
and UO_1290 (O_1290,N_13270,N_13871);
or UO_1291 (O_1291,N_14462,N_13558);
and UO_1292 (O_1292,N_11210,N_13935);
nor UO_1293 (O_1293,N_12918,N_14471);
xor UO_1294 (O_1294,N_12092,N_12660);
and UO_1295 (O_1295,N_12494,N_14522);
nor UO_1296 (O_1296,N_10690,N_13470);
or UO_1297 (O_1297,N_11128,N_14616);
nand UO_1298 (O_1298,N_10769,N_13781);
xor UO_1299 (O_1299,N_13090,N_14211);
nand UO_1300 (O_1300,N_10260,N_12708);
or UO_1301 (O_1301,N_10477,N_11334);
or UO_1302 (O_1302,N_11057,N_13014);
or UO_1303 (O_1303,N_10958,N_10798);
nand UO_1304 (O_1304,N_11437,N_11694);
and UO_1305 (O_1305,N_11274,N_10576);
or UO_1306 (O_1306,N_13944,N_14960);
xor UO_1307 (O_1307,N_11949,N_14935);
and UO_1308 (O_1308,N_14929,N_13086);
or UO_1309 (O_1309,N_10689,N_14058);
nand UO_1310 (O_1310,N_12940,N_11708);
xor UO_1311 (O_1311,N_13965,N_14386);
and UO_1312 (O_1312,N_10451,N_13876);
and UO_1313 (O_1313,N_10649,N_13476);
and UO_1314 (O_1314,N_10501,N_14054);
or UO_1315 (O_1315,N_12408,N_14753);
nand UO_1316 (O_1316,N_11454,N_10316);
and UO_1317 (O_1317,N_11567,N_13713);
xor UO_1318 (O_1318,N_10735,N_11502);
nand UO_1319 (O_1319,N_14502,N_13689);
xor UO_1320 (O_1320,N_12065,N_10307);
xnor UO_1321 (O_1321,N_14437,N_10301);
or UO_1322 (O_1322,N_14921,N_12951);
nor UO_1323 (O_1323,N_13142,N_13836);
or UO_1324 (O_1324,N_14891,N_13722);
or UO_1325 (O_1325,N_10618,N_12317);
xnor UO_1326 (O_1326,N_13970,N_13165);
and UO_1327 (O_1327,N_14588,N_11854);
nand UO_1328 (O_1328,N_14518,N_10895);
nand UO_1329 (O_1329,N_13726,N_14378);
nand UO_1330 (O_1330,N_13574,N_13868);
nand UO_1331 (O_1331,N_14225,N_12636);
or UO_1332 (O_1332,N_14382,N_13141);
xnor UO_1333 (O_1333,N_13110,N_12198);
nand UO_1334 (O_1334,N_12521,N_13507);
nor UO_1335 (O_1335,N_13427,N_12439);
nand UO_1336 (O_1336,N_13400,N_13060);
and UO_1337 (O_1337,N_12549,N_14867);
xnor UO_1338 (O_1338,N_12506,N_10280);
nor UO_1339 (O_1339,N_12862,N_13691);
nand UO_1340 (O_1340,N_10481,N_12504);
nor UO_1341 (O_1341,N_14663,N_13033);
or UO_1342 (O_1342,N_10983,N_12626);
xor UO_1343 (O_1343,N_12781,N_14261);
or UO_1344 (O_1344,N_14726,N_10605);
nor UO_1345 (O_1345,N_11531,N_11675);
nor UO_1346 (O_1346,N_12512,N_13053);
xnor UO_1347 (O_1347,N_10809,N_11079);
xor UO_1348 (O_1348,N_11121,N_11884);
nand UO_1349 (O_1349,N_11649,N_14483);
nand UO_1350 (O_1350,N_13845,N_12389);
nand UO_1351 (O_1351,N_12475,N_11364);
nor UO_1352 (O_1352,N_14352,N_12922);
or UO_1353 (O_1353,N_12437,N_10432);
or UO_1354 (O_1354,N_10174,N_14127);
xnor UO_1355 (O_1355,N_14981,N_12275);
nand UO_1356 (O_1356,N_13968,N_11013);
or UO_1357 (O_1357,N_10355,N_12079);
nand UO_1358 (O_1358,N_11396,N_11124);
nor UO_1359 (O_1359,N_14426,N_11815);
and UO_1360 (O_1360,N_10188,N_12167);
nor UO_1361 (O_1361,N_11552,N_11647);
nand UO_1362 (O_1362,N_14047,N_12662);
or UO_1363 (O_1363,N_14916,N_14843);
nor UO_1364 (O_1364,N_10233,N_10214);
xnor UO_1365 (O_1365,N_13711,N_13573);
xor UO_1366 (O_1366,N_13440,N_11620);
nor UO_1367 (O_1367,N_14181,N_14222);
xnor UO_1368 (O_1368,N_12900,N_13213);
and UO_1369 (O_1369,N_11400,N_10118);
nor UO_1370 (O_1370,N_13622,N_14848);
or UO_1371 (O_1371,N_11298,N_13709);
nor UO_1372 (O_1372,N_11094,N_11078);
or UO_1373 (O_1373,N_12958,N_13382);
and UO_1374 (O_1374,N_12136,N_12025);
nor UO_1375 (O_1375,N_12773,N_12261);
nand UO_1376 (O_1376,N_10981,N_12995);
xor UO_1377 (O_1377,N_13290,N_14035);
and UO_1378 (O_1378,N_11478,N_11549);
xnor UO_1379 (O_1379,N_11017,N_14177);
nand UO_1380 (O_1380,N_12809,N_14128);
nand UO_1381 (O_1381,N_12937,N_11450);
and UO_1382 (O_1382,N_12393,N_13548);
nor UO_1383 (O_1383,N_12948,N_13266);
nor UO_1384 (O_1384,N_14393,N_14928);
nand UO_1385 (O_1385,N_11876,N_11753);
nor UO_1386 (O_1386,N_14080,N_14626);
xor UO_1387 (O_1387,N_13405,N_11498);
nand UO_1388 (O_1388,N_13255,N_12076);
nand UO_1389 (O_1389,N_10789,N_14827);
or UO_1390 (O_1390,N_10648,N_14027);
nand UO_1391 (O_1391,N_12534,N_13896);
xor UO_1392 (O_1392,N_13453,N_12139);
nand UO_1393 (O_1393,N_12145,N_14224);
and UO_1394 (O_1394,N_11461,N_11247);
or UO_1395 (O_1395,N_10907,N_12765);
and UO_1396 (O_1396,N_13317,N_10611);
nor UO_1397 (O_1397,N_14335,N_14093);
nand UO_1398 (O_1398,N_14610,N_12556);
nand UO_1399 (O_1399,N_14372,N_11754);
or UO_1400 (O_1400,N_13818,N_11016);
or UO_1401 (O_1401,N_14545,N_13188);
nor UO_1402 (O_1402,N_14499,N_11540);
or UO_1403 (O_1403,N_12736,N_11143);
or UO_1404 (O_1404,N_10898,N_13536);
xor UO_1405 (O_1405,N_13216,N_11797);
nor UO_1406 (O_1406,N_13451,N_12522);
nand UO_1407 (O_1407,N_12637,N_13496);
nor UO_1408 (O_1408,N_14696,N_13699);
or UO_1409 (O_1409,N_14076,N_13798);
or UO_1410 (O_1410,N_14534,N_11775);
nor UO_1411 (O_1411,N_11323,N_13125);
nor UO_1412 (O_1412,N_14883,N_11031);
nor UO_1413 (O_1413,N_11584,N_13039);
xnor UO_1414 (O_1414,N_12096,N_10369);
xnor UO_1415 (O_1415,N_10211,N_10048);
and UO_1416 (O_1416,N_13095,N_10213);
nand UO_1417 (O_1417,N_12651,N_11825);
or UO_1418 (O_1418,N_13508,N_10658);
nand UO_1419 (O_1419,N_10851,N_14129);
nor UO_1420 (O_1420,N_10008,N_10065);
and UO_1421 (O_1421,N_12505,N_12327);
or UO_1422 (O_1422,N_13377,N_13327);
nand UO_1423 (O_1423,N_10074,N_12223);
nand UO_1424 (O_1424,N_11152,N_10563);
or UO_1425 (O_1425,N_11986,N_11342);
xor UO_1426 (O_1426,N_14142,N_10441);
xnor UO_1427 (O_1427,N_14111,N_12949);
nand UO_1428 (O_1428,N_14492,N_13221);
nand UO_1429 (O_1429,N_12608,N_10884);
or UO_1430 (O_1430,N_14065,N_11457);
and UO_1431 (O_1431,N_14590,N_14828);
xnor UO_1432 (O_1432,N_10632,N_10062);
xnor UO_1433 (O_1433,N_14621,N_11976);
xnor UO_1434 (O_1434,N_14715,N_13911);
nand UO_1435 (O_1435,N_14717,N_12693);
and UO_1436 (O_1436,N_13565,N_10496);
or UO_1437 (O_1437,N_14568,N_11080);
or UO_1438 (O_1438,N_14767,N_10553);
or UO_1439 (O_1439,N_13729,N_11613);
xnor UO_1440 (O_1440,N_11044,N_12335);
and UO_1441 (O_1441,N_13159,N_13179);
xor UO_1442 (O_1442,N_13483,N_13802);
and UO_1443 (O_1443,N_14566,N_14552);
or UO_1444 (O_1444,N_14042,N_11060);
and UO_1445 (O_1445,N_12263,N_12392);
nor UO_1446 (O_1446,N_13363,N_14899);
xnor UO_1447 (O_1447,N_13930,N_13529);
nor UO_1448 (O_1448,N_12396,N_14004);
xor UO_1449 (O_1449,N_12618,N_13479);
nor UO_1450 (O_1450,N_12621,N_11073);
and UO_1451 (O_1451,N_13581,N_14278);
xor UO_1452 (O_1452,N_10265,N_10114);
nand UO_1453 (O_1453,N_12776,N_13282);
nor UO_1454 (O_1454,N_10317,N_12925);
nor UO_1455 (O_1455,N_11251,N_10151);
or UO_1456 (O_1456,N_14253,N_14028);
xnor UO_1457 (O_1457,N_12313,N_13319);
nor UO_1458 (O_1458,N_14156,N_11063);
and UO_1459 (O_1459,N_12199,N_10970);
and UO_1460 (O_1460,N_14151,N_10364);
and UO_1461 (O_1461,N_13728,N_10762);
xor UO_1462 (O_1462,N_14216,N_11071);
nand UO_1463 (O_1463,N_13409,N_13325);
and UO_1464 (O_1464,N_11681,N_14497);
and UO_1465 (O_1465,N_12163,N_10230);
or UO_1466 (O_1466,N_12703,N_12152);
nand UO_1467 (O_1467,N_10094,N_14939);
nand UO_1468 (O_1468,N_14106,N_10764);
xor UO_1469 (O_1469,N_14479,N_12871);
and UO_1470 (O_1470,N_13238,N_12727);
nand UO_1471 (O_1471,N_12641,N_12242);
and UO_1472 (O_1472,N_14257,N_12090);
nor UO_1473 (O_1473,N_12486,N_11671);
or UO_1474 (O_1474,N_14608,N_14066);
xnor UO_1475 (O_1475,N_12151,N_12680);
and UO_1476 (O_1476,N_14683,N_14118);
nor UO_1477 (O_1477,N_11011,N_12902);
nor UO_1478 (O_1478,N_11123,N_11760);
and UO_1479 (O_1479,N_12367,N_14266);
and UO_1480 (O_1480,N_10272,N_11084);
and UO_1481 (O_1481,N_10526,N_11558);
xor UO_1482 (O_1482,N_12541,N_11564);
and UO_1483 (O_1483,N_10433,N_12866);
nor UO_1484 (O_1484,N_14221,N_11788);
and UO_1485 (O_1485,N_10075,N_14641);
nand UO_1486 (O_1486,N_13472,N_14586);
and UO_1487 (O_1487,N_14609,N_12307);
and UO_1488 (O_1488,N_11291,N_12032);
nand UO_1489 (O_1489,N_11254,N_11134);
or UO_1490 (O_1490,N_10480,N_13354);
and UO_1491 (O_1491,N_10842,N_12762);
xnor UO_1492 (O_1492,N_10242,N_13633);
nand UO_1493 (O_1493,N_13814,N_11491);
nand UO_1494 (O_1494,N_12687,N_14397);
xor UO_1495 (O_1495,N_14527,N_11319);
or UO_1496 (O_1496,N_10949,N_13746);
nand UO_1497 (O_1497,N_11505,N_12464);
xor UO_1498 (O_1498,N_11264,N_10043);
xnor UO_1499 (O_1499,N_14574,N_14459);
and UO_1500 (O_1500,N_14434,N_10370);
and UO_1501 (O_1501,N_12792,N_10752);
or UO_1502 (O_1502,N_12433,N_10217);
and UO_1503 (O_1503,N_10017,N_12594);
xor UO_1504 (O_1504,N_12817,N_13173);
nor UO_1505 (O_1505,N_14684,N_14914);
and UO_1506 (O_1506,N_11424,N_11848);
xnor UO_1507 (O_1507,N_10677,N_12947);
nor UO_1508 (O_1508,N_13184,N_14957);
xnor UO_1509 (O_1509,N_14689,N_12161);
and UO_1510 (O_1510,N_11719,N_14821);
or UO_1511 (O_1511,N_13957,N_13076);
or UO_1512 (O_1512,N_14885,N_10231);
xor UO_1513 (O_1513,N_10147,N_11723);
or UO_1514 (O_1514,N_14444,N_11635);
nor UO_1515 (O_1515,N_12987,N_10011);
nor UO_1516 (O_1516,N_10173,N_11780);
or UO_1517 (O_1517,N_11946,N_14911);
nand UO_1518 (O_1518,N_13582,N_12459);
and UO_1519 (O_1519,N_13231,N_13096);
nor UO_1520 (O_1520,N_14112,N_10642);
nor UO_1521 (O_1521,N_12531,N_11872);
or UO_1522 (O_1522,N_12150,N_13147);
nor UO_1523 (O_1523,N_11463,N_12663);
xor UO_1524 (O_1524,N_11633,N_13993);
or UO_1525 (O_1525,N_11833,N_10653);
and UO_1526 (O_1526,N_11327,N_14558);
or UO_1527 (O_1527,N_11004,N_13662);
and UO_1528 (O_1528,N_13947,N_10995);
or UO_1529 (O_1529,N_11113,N_12581);
xnor UO_1530 (O_1530,N_14541,N_11956);
nor UO_1531 (O_1531,N_13575,N_14801);
nor UO_1532 (O_1532,N_13856,N_14734);
xor UO_1533 (O_1533,N_13851,N_11435);
or UO_1534 (O_1534,N_14519,N_14964);
or UO_1535 (O_1535,N_13077,N_13682);
or UO_1536 (O_1536,N_12344,N_14203);
and UO_1537 (O_1537,N_10012,N_13418);
nor UO_1538 (O_1538,N_10281,N_11950);
nor UO_1539 (O_1539,N_11871,N_13660);
and UO_1540 (O_1540,N_11637,N_10350);
nor UO_1541 (O_1541,N_14200,N_10080);
and UO_1542 (O_1542,N_14844,N_14805);
or UO_1543 (O_1543,N_10598,N_11724);
xnor UO_1544 (O_1544,N_11578,N_11607);
and UO_1545 (O_1545,N_12502,N_10915);
xor UO_1546 (O_1546,N_14763,N_10931);
and UO_1547 (O_1547,N_12652,N_14030);
and UO_1548 (O_1548,N_14084,N_12811);
nand UO_1549 (O_1549,N_13977,N_14432);
nand UO_1550 (O_1550,N_14597,N_12113);
nand UO_1551 (O_1551,N_13066,N_12936);
xor UO_1552 (O_1552,N_12836,N_12683);
xor UO_1553 (O_1553,N_11225,N_10051);
or UO_1554 (O_1554,N_10145,N_11353);
nor UO_1555 (O_1555,N_13404,N_11166);
and UO_1556 (O_1556,N_14796,N_13365);
and UO_1557 (O_1557,N_12955,N_11090);
nor UO_1558 (O_1558,N_14606,N_13484);
and UO_1559 (O_1559,N_12580,N_11330);
or UO_1560 (O_1560,N_10482,N_14984);
nand UO_1561 (O_1561,N_11859,N_11231);
nand UO_1562 (O_1562,N_11206,N_11807);
nor UO_1563 (O_1563,N_14375,N_14301);
or UO_1564 (O_1564,N_13463,N_14906);
or UO_1565 (O_1565,N_11253,N_11278);
or UO_1566 (O_1566,N_14733,N_12642);
nand UO_1567 (O_1567,N_12498,N_11763);
or UO_1568 (O_1568,N_10667,N_14219);
or UO_1569 (O_1569,N_12689,N_10733);
or UO_1570 (O_1570,N_14107,N_14525);
xnor UO_1571 (O_1571,N_10448,N_14920);
nor UO_1572 (O_1572,N_12183,N_10205);
xor UO_1573 (O_1573,N_11303,N_10241);
and UO_1574 (O_1574,N_13742,N_11422);
nand UO_1575 (O_1575,N_14769,N_12728);
nand UO_1576 (O_1576,N_10357,N_11276);
and UO_1577 (O_1577,N_13602,N_11015);
and UO_1578 (O_1578,N_14832,N_13593);
nor UO_1579 (O_1579,N_10381,N_12084);
or UO_1580 (O_1580,N_10777,N_13546);
and UO_1581 (O_1581,N_10158,N_11333);
xnor UO_1582 (O_1582,N_13643,N_10548);
nand UO_1583 (O_1583,N_12966,N_14494);
xor UO_1584 (O_1584,N_12724,N_10879);
and UO_1585 (O_1585,N_12639,N_10852);
nor UO_1586 (O_1586,N_12400,N_14036);
nand UO_1587 (O_1587,N_13583,N_13333);
and UO_1588 (O_1588,N_12859,N_11026);
nor UO_1589 (O_1589,N_11217,N_13140);
nor UO_1590 (O_1590,N_13132,N_10282);
nor UO_1591 (O_1591,N_11504,N_12115);
xor UO_1592 (O_1592,N_10079,N_10431);
xor UO_1593 (O_1593,N_10550,N_13153);
nand UO_1594 (O_1594,N_14900,N_11769);
xor UO_1595 (O_1595,N_11483,N_10473);
xnor UO_1596 (O_1596,N_14307,N_13843);
or UO_1597 (O_1597,N_13361,N_10069);
nor UO_1598 (O_1598,N_14271,N_12725);
and UO_1599 (O_1599,N_10977,N_13716);
or UO_1600 (O_1600,N_13399,N_10803);
nand UO_1601 (O_1601,N_13655,N_12391);
or UO_1602 (O_1602,N_11545,N_11503);
and UO_1603 (O_1603,N_14943,N_13099);
nor UO_1604 (O_1604,N_10946,N_14241);
xnor UO_1605 (O_1605,N_12071,N_11703);
and UO_1606 (O_1606,N_13397,N_14446);
or UO_1607 (O_1607,N_11542,N_13846);
or UO_1608 (O_1608,N_11538,N_11118);
xnor UO_1609 (O_1609,N_12911,N_10757);
nand UO_1610 (O_1610,N_10107,N_13422);
nand UO_1611 (O_1611,N_10989,N_12889);
or UO_1612 (O_1612,N_10727,N_10198);
and UO_1613 (O_1613,N_13357,N_13083);
nand UO_1614 (O_1614,N_10144,N_14808);
or UO_1615 (O_1615,N_10601,N_14451);
nand UO_1616 (O_1616,N_12287,N_11501);
xnor UO_1617 (O_1617,N_11598,N_13839);
and UO_1618 (O_1618,N_14242,N_10786);
or UO_1619 (O_1619,N_11676,N_14589);
xnor UO_1620 (O_1620,N_14671,N_14033);
and UO_1621 (O_1621,N_14649,N_10651);
and UO_1622 (O_1622,N_13596,N_13619);
and UO_1623 (O_1623,N_11455,N_11476);
nor UO_1624 (O_1624,N_13701,N_13162);
xor UO_1625 (O_1625,N_13419,N_10122);
xnor UO_1626 (O_1626,N_14857,N_11023);
nand UO_1627 (O_1627,N_10542,N_13129);
nand UO_1628 (O_1628,N_14790,N_12782);
and UO_1629 (O_1629,N_13172,N_11924);
nand UO_1630 (O_1630,N_13176,N_14150);
nand UO_1631 (O_1631,N_13302,N_12835);
nor UO_1632 (O_1632,N_11830,N_14467);
nor UO_1633 (O_1633,N_14713,N_14448);
xnor UO_1634 (O_1634,N_13469,N_12184);
or UO_1635 (O_1635,N_13854,N_12213);
nand UO_1636 (O_1636,N_13710,N_10171);
and UO_1637 (O_1637,N_12352,N_13738);
nor UO_1638 (O_1638,N_12933,N_13520);
nor UO_1639 (O_1639,N_11429,N_10082);
or UO_1640 (O_1640,N_14048,N_11758);
nor UO_1641 (O_1641,N_14365,N_13932);
nand UO_1642 (O_1642,N_11809,N_12584);
nor UO_1643 (O_1643,N_12174,N_11419);
or UO_1644 (O_1644,N_10192,N_10461);
and UO_1645 (O_1645,N_12069,N_14571);
nand UO_1646 (O_1646,N_13627,N_14628);
and UO_1647 (O_1647,N_10275,N_11187);
nand UO_1648 (O_1648,N_11922,N_11997);
nand UO_1649 (O_1649,N_11256,N_14591);
nor UO_1650 (O_1650,N_11599,N_14991);
nor UO_1651 (O_1651,N_12609,N_11164);
xor UO_1652 (O_1652,N_13295,N_14787);
xnor UO_1653 (O_1653,N_13088,N_14053);
nand UO_1654 (O_1654,N_12501,N_11216);
xor UO_1655 (O_1655,N_10854,N_13983);
nor UO_1656 (O_1656,N_14965,N_10857);
nor UO_1657 (O_1657,N_12980,N_13137);
nor UO_1658 (O_1658,N_10185,N_12472);
xor UO_1659 (O_1659,N_10016,N_13964);
and UO_1660 (O_1660,N_10093,N_12908);
xor UO_1661 (O_1661,N_13750,N_10633);
or UO_1662 (O_1662,N_12483,N_10243);
or UO_1663 (O_1663,N_10152,N_12105);
nor UO_1664 (O_1664,N_11627,N_14293);
nor UO_1665 (O_1665,N_10825,N_14144);
or UO_1666 (O_1666,N_13489,N_13164);
nand UO_1667 (O_1667,N_14978,N_10400);
nor UO_1668 (O_1668,N_14298,N_13473);
xnor UO_1669 (O_1669,N_12148,N_14101);
nor UO_1670 (O_1670,N_13645,N_13063);
xnor UO_1671 (O_1671,N_12097,N_13106);
nor UO_1672 (O_1672,N_11716,N_10263);
xor UO_1673 (O_1673,N_11258,N_12602);
xnor UO_1674 (O_1674,N_10408,N_13104);
and UO_1675 (O_1675,N_10941,N_10800);
nand UO_1676 (O_1676,N_11632,N_11245);
and UO_1677 (O_1677,N_14008,N_11983);
or UO_1678 (O_1678,N_10443,N_12279);
and UO_1679 (O_1679,N_12337,N_11106);
nand UO_1680 (O_1680,N_12849,N_11641);
or UO_1681 (O_1681,N_14854,N_10630);
xor UO_1682 (O_1682,N_10345,N_14672);
or UO_1683 (O_1683,N_11019,N_10838);
and UO_1684 (O_1684,N_13705,N_10221);
xnor UO_1685 (O_1685,N_11479,N_11099);
or UO_1686 (O_1686,N_14220,N_14542);
and UO_1687 (O_1687,N_14691,N_14115);
or UO_1688 (O_1688,N_13435,N_10224);
or UO_1689 (O_1689,N_11465,N_10244);
or UO_1690 (O_1690,N_11977,N_13281);
and UO_1691 (O_1691,N_14645,N_11595);
nor UO_1692 (O_1692,N_13369,N_11493);
or UO_1693 (O_1693,N_14056,N_11718);
nor UO_1694 (O_1694,N_13519,N_12093);
and UO_1695 (O_1695,N_12984,N_12743);
nand UO_1696 (O_1696,N_13603,N_13996);
and UO_1697 (O_1697,N_13084,N_13273);
nor UO_1698 (O_1698,N_11175,N_11728);
nor UO_1699 (O_1699,N_11521,N_14947);
nand UO_1700 (O_1700,N_11961,N_12173);
nand UO_1701 (O_1701,N_13962,N_12416);
xor UO_1702 (O_1702,N_13398,N_14068);
and UO_1703 (O_1703,N_14458,N_13747);
nand UO_1704 (O_1704,N_13501,N_11609);
or UO_1705 (O_1705,N_10225,N_14959);
nand UO_1706 (O_1706,N_14146,N_13564);
nand UO_1707 (O_1707,N_13787,N_10067);
or UO_1708 (O_1708,N_11782,N_11917);
and UO_1709 (O_1709,N_12994,N_12255);
and UO_1710 (O_1710,N_11982,N_14223);
nor UO_1711 (O_1711,N_13638,N_14651);
and UO_1712 (O_1712,N_12382,N_12049);
or UO_1713 (O_1713,N_13143,N_14284);
nand UO_1714 (O_1714,N_11375,N_13741);
nand UO_1715 (O_1715,N_14580,N_11340);
xnor UO_1716 (O_1716,N_11662,N_12801);
or UO_1717 (O_1717,N_11841,N_11098);
and UO_1718 (O_1718,N_14442,N_13192);
nand UO_1719 (O_1719,N_12286,N_11960);
and UO_1720 (O_1720,N_14481,N_13842);
nand UO_1721 (O_1721,N_13956,N_13599);
or UO_1722 (O_1722,N_13700,N_12570);
nand UO_1723 (O_1723,N_12881,N_13203);
nand UO_1724 (O_1724,N_10323,N_12579);
nor UO_1725 (O_1725,N_14771,N_10805);
nand UO_1726 (O_1726,N_10341,N_13462);
xor UO_1727 (O_1727,N_14820,N_11212);
nand UO_1728 (O_1728,N_11840,N_14598);
and UO_1729 (O_1729,N_11974,N_12536);
xnor UO_1730 (O_1730,N_12696,N_12686);
xor UO_1731 (O_1731,N_12599,N_13278);
nand UO_1732 (O_1732,N_11755,N_13512);
and UO_1733 (O_1733,N_12017,N_13997);
nand UO_1734 (O_1734,N_13262,N_13450);
nand UO_1735 (O_1735,N_10287,N_12365);
and UO_1736 (O_1736,N_14138,N_11184);
or UO_1737 (O_1737,N_11273,N_14774);
and UO_1738 (O_1738,N_14953,N_12251);
nor UO_1739 (O_1739,N_13864,N_14812);
xor UO_1740 (O_1740,N_13010,N_12138);
and UO_1741 (O_1741,N_11808,N_10109);
nand UO_1742 (O_1742,N_14353,N_10366);
xnor UO_1743 (O_1743,N_14280,N_10715);
or UO_1744 (O_1744,N_14889,N_13820);
nor UO_1745 (O_1745,N_10219,N_12508);
nand UO_1746 (O_1746,N_10908,N_10068);
and UO_1747 (O_1747,N_13065,N_12012);
nor UO_1748 (O_1748,N_13827,N_13677);
and UO_1749 (O_1749,N_13446,N_13694);
nor UO_1750 (O_1750,N_12166,N_12654);
nor UO_1751 (O_1751,N_12310,N_13756);
or UO_1752 (O_1752,N_12598,N_10976);
or UO_1753 (O_1753,N_11097,N_12603);
xnor UO_1754 (O_1754,N_14934,N_13963);
and UO_1755 (O_1755,N_13356,N_11539);
and UO_1756 (O_1756,N_13120,N_14533);
nand UO_1757 (O_1757,N_12620,N_11177);
and UO_1758 (O_1758,N_13004,N_12372);
or UO_1759 (O_1759,N_14834,N_10565);
or UO_1760 (O_1760,N_12033,N_13429);
nor UO_1761 (O_1761,N_10283,N_10215);
nand UO_1762 (O_1762,N_11234,N_10471);
and UO_1763 (O_1763,N_14358,N_14305);
nand UO_1764 (O_1764,N_11709,N_10829);
or UO_1765 (O_1765,N_13659,N_14477);
and UO_1766 (O_1766,N_14303,N_10695);
nor UO_1767 (O_1767,N_11747,N_11354);
xnor UO_1768 (O_1768,N_12410,N_13760);
nor UO_1769 (O_1769,N_11711,N_13675);
nor UO_1770 (O_1770,N_12454,N_11497);
nor UO_1771 (O_1771,N_11816,N_10305);
and UO_1772 (O_1772,N_10382,N_10754);
nor UO_1773 (O_1773,N_14793,N_13912);
nor UO_1774 (O_1774,N_14501,N_12818);
or UO_1775 (O_1775,N_14126,N_14273);
xnor UO_1776 (O_1776,N_12440,N_11149);
and UO_1777 (O_1777,N_13240,N_12695);
or UO_1778 (O_1778,N_14809,N_11692);
or UO_1779 (O_1779,N_13704,N_11579);
and UO_1780 (O_1780,N_12140,N_13032);
xnor UO_1781 (O_1781,N_10559,N_14171);
nand UO_1782 (O_1782,N_13551,N_13210);
nand UO_1783 (O_1783,N_11436,N_11908);
xnor UO_1784 (O_1784,N_11525,N_12575);
nand UO_1785 (O_1785,N_13205,N_10730);
or UO_1786 (O_1786,N_13918,N_11142);
nor UO_1787 (O_1787,N_12613,N_11038);
or UO_1788 (O_1788,N_12212,N_10141);
nand UO_1789 (O_1789,N_12043,N_13861);
xor UO_1790 (O_1790,N_10483,N_12356);
nand UO_1791 (O_1791,N_12840,N_13177);
xnor UO_1792 (O_1792,N_13630,N_12882);
or UO_1793 (O_1793,N_14405,N_14951);
nor UO_1794 (O_1794,N_12775,N_14105);
xnor UO_1795 (O_1795,N_10876,N_10514);
xnor UO_1796 (O_1796,N_11093,N_12155);
and UO_1797 (O_1797,N_12878,N_12260);
and UO_1798 (O_1798,N_11308,N_14037);
or UO_1799 (O_1799,N_13771,N_12374);
nor UO_1800 (O_1800,N_13566,N_13920);
nand UO_1801 (O_1801,N_11480,N_12162);
nand UO_1802 (O_1802,N_12030,N_11236);
or UO_1803 (O_1803,N_13485,N_13608);
nor UO_1804 (O_1804,N_14837,N_11196);
or UO_1805 (O_1805,N_12104,N_14500);
and UO_1806 (O_1806,N_10902,N_14762);
xnor UO_1807 (O_1807,N_14846,N_13980);
nor UO_1808 (O_1808,N_14480,N_10722);
nand UO_1809 (O_1809,N_11232,N_11566);
xor UO_1810 (O_1810,N_12318,N_12045);
and UO_1811 (O_1811,N_12705,N_11881);
xor UO_1812 (O_1812,N_14680,N_10353);
xor UO_1813 (O_1813,N_11361,N_10266);
xnor UO_1814 (O_1814,N_10646,N_10207);
or UO_1815 (O_1815,N_10037,N_11968);
xor UO_1816 (O_1816,N_14855,N_10025);
and UO_1817 (O_1817,N_12462,N_12401);
or UO_1818 (O_1818,N_14317,N_12325);
and UO_1819 (O_1819,N_14806,N_12359);
nor UO_1820 (O_1820,N_11846,N_13025);
or UO_1821 (O_1821,N_13437,N_13277);
xnor UO_1822 (O_1822,N_10493,N_10466);
xnor UO_1823 (O_1823,N_14537,N_14354);
nor UO_1824 (O_1824,N_11878,N_12293);
or UO_1825 (O_1825,N_13960,N_12628);
nor UO_1826 (O_1826,N_12977,N_14239);
or UO_1827 (O_1827,N_12222,N_12640);
and UO_1828 (O_1828,N_13668,N_14422);
or UO_1829 (O_1829,N_14605,N_13753);
and UO_1830 (O_1830,N_10389,N_10533);
xor UO_1831 (O_1831,N_13324,N_13612);
nand UO_1832 (O_1832,N_11810,N_12519);
or UO_1833 (O_1833,N_12510,N_11642);
nand UO_1834 (O_1834,N_13015,N_12019);
and UO_1835 (O_1835,N_11943,N_13740);
nand UO_1836 (O_1836,N_13618,N_14059);
nand UO_1837 (O_1837,N_13938,N_12202);
nand UO_1838 (O_1838,N_10641,N_13953);
xor UO_1839 (O_1839,N_14778,N_11315);
nand UO_1840 (O_1840,N_14077,N_12716);
nor UO_1841 (O_1841,N_12412,N_10536);
nand UO_1842 (O_1842,N_13878,N_13686);
xnor UO_1843 (O_1843,N_11773,N_11481);
nand UO_1844 (O_1844,N_14810,N_14704);
and UO_1845 (O_1845,N_11529,N_11915);
or UO_1846 (O_1846,N_10637,N_11136);
xnor UO_1847 (O_1847,N_12171,N_14000);
nand UO_1848 (O_1848,N_14513,N_11307);
and UO_1849 (O_1849,N_11929,N_11105);
nor UO_1850 (O_1850,N_11518,N_12864);
nand UO_1851 (O_1851,N_12560,N_13532);
nor UO_1852 (O_1852,N_11853,N_11188);
nand UO_1853 (O_1853,N_13155,N_14858);
nand UO_1854 (O_1854,N_10041,N_11283);
and UO_1855 (O_1855,N_14075,N_10150);
nand UO_1856 (O_1856,N_14233,N_11686);
or UO_1857 (O_1857,N_14125,N_11112);
and UO_1858 (O_1858,N_14323,N_11616);
nand UO_1859 (O_1859,N_11900,N_10395);
nor UO_1860 (O_1860,N_14905,N_14980);
nor UO_1861 (O_1861,N_10844,N_12623);
nand UO_1862 (O_1862,N_11215,N_12672);
xnor UO_1863 (O_1863,N_12108,N_14267);
or UO_1864 (O_1864,N_14781,N_10543);
and UO_1865 (O_1865,N_10923,N_10148);
or UO_1866 (O_1866,N_14256,N_11033);
or UO_1867 (O_1867,N_14988,N_11174);
and UO_1868 (O_1868,N_10595,N_14506);
xnor UO_1869 (O_1869,N_10897,N_14104);
xor UO_1870 (O_1870,N_10154,N_12149);
nand UO_1871 (O_1871,N_11670,N_11172);
nand UO_1872 (O_1872,N_10612,N_11199);
xnor UO_1873 (O_1873,N_10801,N_12385);
nand UO_1874 (O_1874,N_11367,N_12369);
nor UO_1875 (O_1875,N_13822,N_12796);
and UO_1876 (O_1876,N_11395,N_13994);
and UO_1877 (O_1877,N_10833,N_12884);
and UO_1878 (O_1878,N_10237,N_14240);
nor UO_1879 (O_1879,N_14614,N_10403);
or UO_1880 (O_1880,N_13459,N_10728);
nor UO_1881 (O_1881,N_13345,N_13590);
or UO_1882 (O_1882,N_13149,N_11568);
and UO_1883 (O_1883,N_14530,N_10582);
or UO_1884 (O_1884,N_11472,N_12929);
xor UO_1885 (O_1885,N_10518,N_10692);
nand UO_1886 (O_1886,N_12883,N_13552);
xnor UO_1887 (O_1887,N_11663,N_13788);
nor UO_1888 (O_1888,N_12763,N_13757);
nand UO_1889 (O_1889,N_12707,N_11012);
nand UO_1890 (O_1890,N_13416,N_11634);
and UO_1891 (O_1891,N_12700,N_12221);
and UO_1892 (O_1892,N_10617,N_10311);
xor UO_1893 (O_1893,N_14091,N_12566);
xor UO_1894 (O_1894,N_14772,N_13664);
and UO_1895 (O_1895,N_14038,N_11391);
xnor UO_1896 (O_1896,N_13776,N_10349);
nand UO_1897 (O_1897,N_14315,N_12923);
xnor UO_1898 (O_1898,N_11928,N_11117);
or UO_1899 (O_1899,N_10129,N_12258);
nor UO_1900 (O_1900,N_12193,N_11735);
or UO_1901 (O_1901,N_11103,N_13358);
or UO_1902 (O_1902,N_14823,N_12670);
nand UO_1903 (O_1903,N_10781,N_14320);
xor UO_1904 (O_1904,N_12904,N_11471);
nand UO_1905 (O_1905,N_11357,N_11159);
xor UO_1906 (O_1906,N_11262,N_10202);
and UO_1907 (O_1907,N_11317,N_13222);
nand UO_1908 (O_1908,N_11629,N_14950);
nand UO_1909 (O_1909,N_11104,N_12553);
and UO_1910 (O_1910,N_12511,N_14865);
or UO_1911 (O_1911,N_10834,N_13874);
xor UO_1912 (O_1912,N_11281,N_13236);
xor UO_1913 (O_1913,N_10420,N_11710);
and UO_1914 (O_1914,N_11947,N_12648);
or UO_1915 (O_1915,N_11874,N_12006);
or UO_1916 (O_1916,N_14755,N_14773);
nand UO_1917 (O_1917,N_12734,N_14594);
and UO_1918 (O_1918,N_13311,N_10404);
nor UO_1919 (O_1919,N_12164,N_13840);
xnor UO_1920 (O_1920,N_14833,N_14015);
nand UO_1921 (O_1921,N_12574,N_11040);
and UO_1922 (O_1922,N_10771,N_11644);
or UO_1923 (O_1923,N_12529,N_10169);
and UO_1924 (O_1924,N_14554,N_10101);
nor UO_1925 (O_1925,N_11506,N_12804);
nand UO_1926 (O_1926,N_11850,N_14498);
or UO_1927 (O_1927,N_11482,N_14538);
nor UO_1928 (O_1928,N_12778,N_13190);
xnor UO_1929 (O_1929,N_13653,N_11226);
and UO_1930 (O_1930,N_10092,N_13749);
or UO_1931 (O_1931,N_11148,N_12037);
xor UO_1932 (O_1932,N_14536,N_13012);
and UO_1933 (O_1933,N_12755,N_13852);
and UO_1934 (O_1934,N_11697,N_13035);
or UO_1935 (O_1935,N_10971,N_12427);
xor UO_1936 (O_1936,N_12331,N_10410);
and UO_1937 (O_1937,N_13267,N_10232);
and UO_1938 (O_1938,N_14158,N_12851);
xor UO_1939 (O_1939,N_14496,N_11163);
nand UO_1940 (O_1940,N_10761,N_14901);
nand UO_1941 (O_1941,N_10575,N_13580);
nand UO_1942 (O_1942,N_11942,N_10175);
xor UO_1943 (O_1943,N_10116,N_13146);
nand UO_1944 (O_1944,N_13632,N_13537);
and UO_1945 (O_1945,N_14029,N_12606);
or UO_1946 (O_1946,N_11238,N_14347);
nand UO_1947 (O_1947,N_11190,N_12326);
and UO_1948 (O_1948,N_11467,N_12668);
and UO_1949 (O_1949,N_11324,N_11715);
nor UO_1950 (O_1950,N_13972,N_14143);
and UO_1951 (O_1951,N_11661,N_14436);
nand UO_1952 (O_1952,N_14132,N_11991);
xnor UO_1953 (O_1953,N_10249,N_11669);
nor UO_1954 (O_1954,N_10325,N_14852);
nor UO_1955 (O_1955,N_12256,N_12176);
nand UO_1956 (O_1956,N_10636,N_11603);
or UO_1957 (O_1957,N_12719,N_14788);
nand UO_1958 (O_1958,N_14646,N_13226);
and UO_1959 (O_1959,N_14340,N_13666);
nand UO_1960 (O_1960,N_14544,N_12666);
or UO_1961 (O_1961,N_11512,N_14941);
xnor UO_1962 (O_1962,N_12965,N_10309);
nand UO_1963 (O_1963,N_12973,N_13154);
nand UO_1964 (O_1964,N_13847,N_13239);
xor UO_1965 (O_1965,N_14903,N_13877);
xor UO_1966 (O_1966,N_12297,N_12991);
or UO_1967 (O_1967,N_10296,N_11904);
xnor UO_1968 (O_1968,N_13777,N_11562);
or UO_1969 (O_1969,N_11132,N_10504);
or UO_1970 (O_1970,N_13865,N_12324);
nor UO_1971 (O_1971,N_14676,N_13193);
nand UO_1972 (O_1972,N_14187,N_10100);
or UO_1973 (O_1973,N_13948,N_11299);
nand UO_1974 (O_1974,N_12885,N_12316);
and UO_1975 (O_1975,N_11485,N_14411);
nand UO_1976 (O_1976,N_13477,N_10647);
or UO_1977 (O_1977,N_14719,N_14201);
and UO_1978 (O_1978,N_11717,N_12191);
nor UO_1979 (O_1979,N_13214,N_10285);
xnor UO_1980 (O_1980,N_14707,N_14249);
nand UO_1981 (O_1981,N_12491,N_13340);
and UO_1982 (O_1982,N_13745,N_14351);
nand UO_1983 (O_1983,N_12848,N_11056);
nor UO_1984 (O_1984,N_10322,N_11628);
and UO_1985 (O_1985,N_11039,N_10180);
or UO_1986 (O_1986,N_12845,N_13646);
nor UO_1987 (O_1987,N_10295,N_12390);
xor UO_1988 (O_1988,N_12932,N_12546);
nor UO_1989 (O_1989,N_12585,N_10720);
or UO_1990 (O_1990,N_10303,N_11456);
nand UO_1991 (O_1991,N_12896,N_12692);
and UO_1992 (O_1992,N_10528,N_13505);
nor UO_1993 (O_1993,N_14139,N_14640);
nand UO_1994 (O_1994,N_10562,N_13407);
nor UO_1995 (O_1995,N_13981,N_13123);
nor UO_1996 (O_1996,N_13126,N_12230);
xor UO_1997 (O_1997,N_11698,N_10040);
or UO_1998 (O_1998,N_11870,N_10290);
nor UO_1999 (O_1999,N_13072,N_10870);
endmodule