module basic_750_5000_1000_2_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2507,N_2508,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2553,N_2554,N_2557,N_2558,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2568,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2582,N_2583,N_2585,N_2586,N_2587,N_2588,N_2590,N_2593,N_2595,N_2596,N_2597,N_2598,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2610,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2637,N_2638,N_2640,N_2642,N_2643,N_2644,N_2645,N_2647,N_2648,N_2649,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2658,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2697,N_2698,N_2699,N_2701,N_2702,N_2703,N_2705,N_2706,N_2707,N_2709,N_2710,N_2711,N_2712,N_2713,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2743,N_2744,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2755,N_2756,N_2758,N_2760,N_2761,N_2763,N_2764,N_2765,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2795,N_2796,N_2797,N_2798,N_2799,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2819,N_2820,N_2821,N_2822,N_2823,N_2825,N_2827,N_2828,N_2829,N_2830,N_2831,N_2833,N_2834,N_2835,N_2837,N_2839,N_2842,N_2843,N_2844,N_2845,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2859,N_2860,N_2861,N_2862,N_2864,N_2865,N_2866,N_2867,N_2868,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2880,N_2881,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2913,N_2914,N_2915,N_2916,N_2917,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2936,N_2937,N_2938,N_2940,N_2941,N_2942,N_2943,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2952,N_2953,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3062,N_3063,N_3064,N_3065,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3076,N_3077,N_3078,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3089,N_3090,N_3094,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3113,N_3115,N_3116,N_3118,N_3119,N_3121,N_3122,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3140,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3152,N_3154,N_3155,N_3156,N_3157,N_3158,N_3160,N_3161,N_3162,N_3163,N_3165,N_3166,N_3167,N_3170,N_3171,N_3172,N_3173,N_3175,N_3176,N_3177,N_3178,N_3180,N_3182,N_3183,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3200,N_3201,N_3202,N_3203,N_3205,N_3206,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3226,N_3227,N_3228,N_3229,N_3231,N_3232,N_3233,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3243,N_3244,N_3245,N_3246,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3275,N_3276,N_3277,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3297,N_3298,N_3300,N_3301,N_3302,N_3303,N_3305,N_3306,N_3307,N_3309,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3325,N_3326,N_3327,N_3328,N_3329,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3341,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3355,N_3356,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3365,N_3366,N_3367,N_3369,N_3370,N_3371,N_3373,N_3375,N_3377,N_3378,N_3379,N_3381,N_3382,N_3384,N_3385,N_3387,N_3388,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3399,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3426,N_3427,N_3428,N_3429,N_3430,N_3432,N_3435,N_3436,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3457,N_3458,N_3460,N_3461,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3480,N_3481,N_3482,N_3483,N_3485,N_3486,N_3487,N_3488,N_3489,N_3491,N_3492,N_3493,N_3494,N_3498,N_3499,N_3501,N_3502,N_3503,N_3504,N_3506,N_3507,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3526,N_3527,N_3528,N_3529,N_3530,N_3533,N_3534,N_3535,N_3536,N_3538,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3547,N_3548,N_3549,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3563,N_3564,N_3567,N_3568,N_3569,N_3570,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3587,N_3588,N_3589,N_3590,N_3591,N_3593,N_3594,N_3595,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3609,N_3610,N_3612,N_3614,N_3616,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3637,N_3638,N_3639,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3653,N_3654,N_3656,N_3659,N_3660,N_3661,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3688,N_3689,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3711,N_3712,N_3713,N_3715,N_3716,N_3717,N_3718,N_3719,N_3721,N_3723,N_3724,N_3725,N_3726,N_3727,N_3729,N_3730,N_3731,N_3732,N_3734,N_3735,N_3736,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3746,N_3747,N_3748,N_3749,N_3750,N_3752,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3779,N_3780,N_3783,N_3784,N_3788,N_3789,N_3791,N_3793,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3803,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3813,N_3814,N_3815,N_3817,N_3818,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3841,N_3843,N_3844,N_3845,N_3847,N_3849,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3860,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3881,N_3883,N_3885,N_3886,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3900,N_3901,N_3902,N_3903,N_3905,N_3906,N_3907,N_3909,N_3912,N_3913,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3922,N_3923,N_3924,N_3925,N_3926,N_3928,N_3929,N_3931,N_3932,N_3933,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3943,N_3944,N_3946,N_3947,N_3948,N_3949,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3992,N_3993,N_3997,N_3998,N_3999,N_4000,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4015,N_4017,N_4018,N_4019,N_4020,N_4021,N_4024,N_4025,N_4026,N_4027,N_4028,N_4030,N_4031,N_4032,N_4033,N_4034,N_4036,N_4038,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4050,N_4051,N_4052,N_4053,N_4054,N_4056,N_4059,N_4060,N_4061,N_4062,N_4063,N_4065,N_4067,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4081,N_4083,N_4084,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4093,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4108,N_4110,N_4112,N_4113,N_4115,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4133,N_4134,N_4135,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4147,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4156,N_4157,N_4158,N_4159,N_4161,N_4162,N_4163,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4230,N_4231,N_4233,N_4234,N_4236,N_4237,N_4238,N_4239,N_4240,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4269,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4281,N_4284,N_4285,N_4286,N_4290,N_4294,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4320,N_4322,N_4323,N_4324,N_4325,N_4326,N_4328,N_4329,N_4330,N_4331,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4343,N_4344,N_4346,N_4347,N_4349,N_4350,N_4352,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4370,N_4371,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4380,N_4381,N_4382,N_4383,N_4384,N_4386,N_4388,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4399,N_4401,N_4402,N_4403,N_4404,N_4408,N_4410,N_4411,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4430,N_4431,N_4434,N_4435,N_4436,N_4438,N_4439,N_4440,N_4441,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4475,N_4476,N_4479,N_4480,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4524,N_4525,N_4527,N_4528,N_4529,N_4530,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4565,N_4566,N_4567,N_4568,N_4570,N_4572,N_4573,N_4574,N_4575,N_4578,N_4579,N_4580,N_4581,N_4582,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4602,N_4604,N_4605,N_4606,N_4607,N_4609,N_4611,N_4612,N_4613,N_4615,N_4616,N_4618,N_4619,N_4620,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4632,N_4633,N_4634,N_4635,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4647,N_4649,N_4650,N_4652,N_4653,N_4654,N_4655,N_4656,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4671,N_4672,N_4673,N_4674,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4696,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4708,N_4709,N_4710,N_4711,N_4713,N_4714,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4733,N_4734,N_4736,N_4739,N_4740,N_4742,N_4743,N_4745,N_4746,N_4748,N_4749,N_4750,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4762,N_4763,N_4765,N_4766,N_4767,N_4768,N_4770,N_4772,N_4774,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4804,N_4807,N_4808,N_4810,N_4812,N_4814,N_4815,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4839,N_4844,N_4845,N_4847,N_4848,N_4849,N_4850,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4860,N_4861,N_4862,N_4863,N_4864,N_4866,N_4867,N_4869,N_4870,N_4871,N_4872,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4893,N_4894,N_4896,N_4897,N_4898,N_4900,N_4904,N_4905,N_4906,N_4908,N_4909,N_4910,N_4912,N_4914,N_4916,N_4917,N_4919,N_4920,N_4921,N_4922,N_4925,N_4927,N_4928,N_4931,N_4932,N_4933,N_4936,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4951,N_4952,N_4953,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4966,N_4969,N_4970,N_4972,N_4973,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4988,N_4989,N_4990,N_4992,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xor U0 (N_0,In_534,In_666);
nand U1 (N_1,In_725,In_187);
xnor U2 (N_2,In_548,In_736);
xor U3 (N_3,In_81,In_110);
nand U4 (N_4,In_108,In_562);
nand U5 (N_5,In_721,In_346);
nor U6 (N_6,In_602,In_583);
and U7 (N_7,In_268,In_642);
xor U8 (N_8,In_481,In_317);
xnor U9 (N_9,In_485,In_295);
nand U10 (N_10,In_680,In_115);
and U11 (N_11,In_409,In_80);
nor U12 (N_12,In_297,In_271);
nor U13 (N_13,In_202,In_383);
or U14 (N_14,In_586,In_255);
nand U15 (N_15,In_274,In_307);
xor U16 (N_16,In_28,In_660);
nor U17 (N_17,In_167,In_665);
nand U18 (N_18,In_125,In_510);
or U19 (N_19,In_31,In_209);
or U20 (N_20,In_243,In_121);
xor U21 (N_21,In_474,In_0);
or U22 (N_22,In_264,In_433);
or U23 (N_23,In_476,In_114);
nor U24 (N_24,In_691,In_422);
xnor U25 (N_25,In_22,In_281);
or U26 (N_26,In_570,In_61);
and U27 (N_27,In_643,In_13);
nand U28 (N_28,In_531,In_97);
xnor U29 (N_29,In_457,In_630);
xor U30 (N_30,In_616,In_1);
nand U31 (N_31,In_464,In_161);
xor U32 (N_32,In_75,In_126);
xnor U33 (N_33,In_214,In_77);
xnor U34 (N_34,In_546,In_674);
and U35 (N_35,In_607,In_318);
nor U36 (N_36,In_479,In_564);
xnor U37 (N_37,In_399,In_105);
nor U38 (N_38,In_94,In_312);
nor U39 (N_39,In_449,In_522);
nand U40 (N_40,In_85,In_462);
and U41 (N_41,In_732,In_171);
and U42 (N_42,In_56,In_23);
or U43 (N_43,In_468,In_406);
or U44 (N_44,In_613,In_168);
or U45 (N_45,In_153,In_84);
and U46 (N_46,In_661,In_141);
or U47 (N_47,In_689,In_742);
xnor U48 (N_48,In_194,In_208);
xor U49 (N_49,In_190,In_175);
or U50 (N_50,In_70,In_552);
and U51 (N_51,In_477,In_396);
nand U52 (N_52,In_48,In_402);
xor U53 (N_53,In_335,In_263);
or U54 (N_54,In_192,In_359);
and U55 (N_55,In_235,In_18);
xor U56 (N_56,In_96,In_219);
and U57 (N_57,In_256,In_143);
or U58 (N_58,In_499,In_431);
xnor U59 (N_59,In_709,In_198);
xnor U60 (N_60,In_129,In_500);
nor U61 (N_61,In_63,In_511);
and U62 (N_62,In_461,In_130);
and U63 (N_63,In_700,In_25);
or U64 (N_64,In_65,In_412);
or U65 (N_65,In_526,In_387);
and U66 (N_66,In_726,In_506);
xnor U67 (N_67,In_614,In_322);
nor U68 (N_68,In_539,In_354);
and U69 (N_69,In_581,In_184);
nand U70 (N_70,In_372,In_38);
or U71 (N_71,In_486,In_701);
and U72 (N_72,In_142,In_279);
or U73 (N_73,In_357,In_553);
nor U74 (N_74,In_528,In_43);
xnor U75 (N_75,In_106,In_26);
and U76 (N_76,In_544,In_180);
xnor U77 (N_77,In_748,In_735);
nand U78 (N_78,In_708,In_555);
and U79 (N_79,In_532,In_254);
and U80 (N_80,In_656,In_340);
nor U81 (N_81,In_728,In_269);
nand U82 (N_82,In_344,In_645);
or U83 (N_83,In_266,In_634);
and U84 (N_84,In_440,In_494);
xnor U85 (N_85,In_542,In_111);
xor U86 (N_86,In_195,In_128);
or U87 (N_87,In_53,In_90);
nor U88 (N_88,In_107,In_738);
or U89 (N_89,In_439,In_154);
nor U90 (N_90,In_566,In_603);
nor U91 (N_91,In_186,In_624);
nor U92 (N_92,In_628,In_46);
xor U93 (N_93,In_27,In_580);
nor U94 (N_94,In_390,In_682);
xor U95 (N_95,In_467,In_326);
and U96 (N_96,In_368,In_291);
xnor U97 (N_97,In_151,In_52);
and U98 (N_98,In_147,In_426);
xor U99 (N_99,In_73,In_329);
and U100 (N_100,In_137,In_465);
nor U101 (N_101,In_188,In_491);
nand U102 (N_102,In_641,In_239);
and U103 (N_103,In_724,In_668);
and U104 (N_104,In_410,In_554);
nand U105 (N_105,In_421,In_530);
nand U106 (N_106,In_231,In_218);
nand U107 (N_107,In_658,In_463);
and U108 (N_108,In_571,In_127);
nor U109 (N_109,In_471,In_286);
and U110 (N_110,In_694,In_71);
xnor U111 (N_111,In_631,In_621);
xnor U112 (N_112,In_206,In_159);
nand U113 (N_113,In_398,In_520);
nor U114 (N_114,In_565,In_419);
or U115 (N_115,In_425,In_653);
or U116 (N_116,In_47,In_388);
and U117 (N_117,In_6,In_144);
and U118 (N_118,In_193,In_537);
or U119 (N_119,In_8,In_389);
nand U120 (N_120,In_191,In_623);
nor U121 (N_121,In_210,In_249);
nor U122 (N_122,In_377,In_2);
nor U123 (N_123,In_201,In_514);
and U124 (N_124,In_288,In_617);
xnor U125 (N_125,In_152,In_181);
and U126 (N_126,In_712,In_667);
and U127 (N_127,In_685,In_540);
xor U128 (N_128,In_595,In_415);
and U129 (N_129,In_258,In_743);
nor U130 (N_130,In_89,In_220);
and U131 (N_131,In_610,In_189);
nand U132 (N_132,In_212,In_637);
nand U133 (N_133,In_333,In_484);
nor U134 (N_134,In_584,In_234);
or U135 (N_135,In_604,In_325);
or U136 (N_136,In_640,In_86);
nand U137 (N_137,In_104,In_686);
nand U138 (N_138,In_718,In_132);
nor U139 (N_139,In_698,In_339);
nand U140 (N_140,In_678,In_293);
xor U141 (N_141,In_699,In_238);
nand U142 (N_142,In_558,In_587);
and U143 (N_143,In_556,In_331);
nor U144 (N_144,In_550,In_460);
or U145 (N_145,In_40,In_582);
or U146 (N_146,In_237,In_619);
and U147 (N_147,In_138,In_21);
nor U148 (N_148,In_729,In_480);
and U149 (N_149,In_221,In_58);
xnor U150 (N_150,In_44,In_670);
nor U151 (N_151,In_622,In_29);
xor U152 (N_152,In_252,In_343);
nand U153 (N_153,In_118,In_713);
xnor U154 (N_154,In_299,In_64);
and U155 (N_155,In_224,In_145);
nand U156 (N_156,In_240,In_527);
nand U157 (N_157,In_253,In_478);
nand U158 (N_158,In_273,In_493);
xnor U159 (N_159,In_405,In_606);
xnor U160 (N_160,In_332,In_458);
nand U161 (N_161,In_676,In_639);
xor U162 (N_162,In_599,In_275);
nor U163 (N_163,In_102,In_515);
nor U164 (N_164,In_225,In_717);
or U165 (N_165,In_657,In_386);
and U166 (N_166,In_683,In_644);
nand U167 (N_167,In_232,In_310);
or U168 (N_168,In_401,In_294);
xnor U169 (N_169,In_513,In_597);
nand U170 (N_170,In_543,In_4);
nor U171 (N_171,In_696,In_349);
xnor U172 (N_172,In_677,In_78);
xnor U173 (N_173,In_262,In_336);
and U174 (N_174,In_367,In_523);
or U175 (N_175,In_385,In_632);
or U176 (N_176,In_663,In_598);
nor U177 (N_177,In_216,In_693);
xor U178 (N_178,In_320,In_400);
nand U179 (N_179,In_423,In_39);
or U180 (N_180,In_3,In_747);
nor U181 (N_181,In_98,In_17);
and U182 (N_182,In_139,In_135);
and U183 (N_183,In_611,In_376);
nor U184 (N_184,In_148,In_170);
xnor U185 (N_185,In_734,In_495);
and U186 (N_186,In_469,In_350);
nor U187 (N_187,In_549,In_472);
and U188 (N_188,In_436,In_156);
and U189 (N_189,In_267,In_83);
and U190 (N_190,In_117,In_375);
nor U191 (N_191,In_560,In_716);
or U192 (N_192,In_524,In_92);
xnor U193 (N_193,In_62,In_733);
nor U194 (N_194,In_690,In_384);
nand U195 (N_195,In_577,In_706);
nand U196 (N_196,In_596,In_482);
and U197 (N_197,In_516,In_538);
xnor U198 (N_198,In_35,In_146);
and U199 (N_199,In_711,In_20);
xnor U200 (N_200,In_620,In_638);
or U201 (N_201,In_448,In_217);
nor U202 (N_202,In_172,In_173);
nand U203 (N_203,In_633,In_730);
xnor U204 (N_204,In_629,In_120);
xor U205 (N_205,In_233,In_594);
and U206 (N_206,In_313,In_124);
or U207 (N_207,In_298,In_563);
nand U208 (N_208,In_334,In_704);
or U209 (N_209,In_119,In_205);
or U210 (N_210,In_723,In_392);
xnor U211 (N_211,In_379,In_455);
and U212 (N_212,In_420,In_533);
nor U213 (N_213,In_703,In_551);
nor U214 (N_214,In_408,In_112);
nand U215 (N_215,In_272,In_287);
nor U216 (N_216,In_380,In_369);
or U217 (N_217,In_547,In_162);
and U218 (N_218,In_741,In_183);
nor U219 (N_219,In_705,In_103);
nand U220 (N_220,In_45,In_328);
nor U221 (N_221,In_36,In_15);
nand U222 (N_222,In_358,In_285);
nand U223 (N_223,In_67,In_122);
xor U224 (N_224,In_24,In_197);
or U225 (N_225,In_215,In_150);
and U226 (N_226,In_95,In_306);
nor U227 (N_227,In_608,In_59);
xnor U228 (N_228,In_483,In_567);
nor U229 (N_229,In_438,In_251);
xnor U230 (N_230,In_200,In_497);
nor U231 (N_231,In_155,In_282);
and U232 (N_232,In_158,In_362);
xnor U233 (N_233,In_5,In_348);
xor U234 (N_234,In_174,In_648);
xor U235 (N_235,In_475,In_626);
nor U236 (N_236,In_196,In_270);
xnor U237 (N_237,In_211,In_204);
nand U238 (N_238,In_341,In_671);
nor U239 (N_239,In_227,In_7);
nor U240 (N_240,In_568,In_746);
nand U241 (N_241,In_69,In_116);
nor U242 (N_242,In_12,In_347);
or U243 (N_243,In_11,In_179);
and U244 (N_244,In_600,In_160);
xor U245 (N_245,In_444,In_418);
nand U246 (N_246,In_57,In_34);
nand U247 (N_247,In_625,In_246);
nand U248 (N_248,In_572,In_487);
xor U249 (N_249,In_697,In_403);
or U250 (N_250,In_283,In_207);
nor U251 (N_251,In_9,In_652);
nand U252 (N_252,In_361,In_10);
nand U253 (N_253,In_647,In_672);
and U254 (N_254,In_308,In_618);
xnor U255 (N_255,In_501,In_601);
nor U256 (N_256,In_33,In_302);
and U257 (N_257,In_50,In_374);
xnor U258 (N_258,In_536,In_578);
xnor U259 (N_259,In_437,In_569);
nor U260 (N_260,In_55,In_447);
nand U261 (N_261,In_473,In_178);
or U262 (N_262,In_337,In_427);
and U263 (N_263,In_429,In_589);
and U264 (N_264,In_428,In_397);
nor U265 (N_265,In_378,In_241);
nor U266 (N_266,In_199,In_615);
and U267 (N_267,In_371,In_673);
or U268 (N_268,In_261,In_373);
xor U269 (N_269,In_276,In_679);
nor U270 (N_270,In_250,In_257);
or U271 (N_271,In_731,In_488);
or U272 (N_272,In_545,In_498);
and U273 (N_273,In_627,In_442);
nand U274 (N_274,In_675,In_76);
nor U275 (N_275,In_176,In_324);
xor U276 (N_276,In_445,In_659);
nor U277 (N_277,In_327,In_68);
nor U278 (N_278,In_507,In_123);
nand U279 (N_279,In_684,In_163);
nand U280 (N_280,In_230,In_432);
or U281 (N_281,In_722,In_177);
and U282 (N_282,In_292,In_692);
and U283 (N_283,In_454,In_100);
or U284 (N_284,In_424,In_355);
or U285 (N_285,In_248,In_301);
nand U286 (N_286,In_353,In_280);
xnor U287 (N_287,In_311,In_688);
xor U288 (N_288,In_740,In_707);
and U289 (N_289,In_74,In_635);
or U290 (N_290,In_140,In_32);
nor U291 (N_291,In_451,In_309);
or U292 (N_292,In_702,In_681);
nand U293 (N_293,In_19,In_93);
xnor U294 (N_294,In_591,In_541);
or U295 (N_295,In_650,In_557);
and U296 (N_296,In_588,In_737);
nor U297 (N_297,In_305,In_456);
or U298 (N_298,In_66,In_393);
nand U299 (N_299,In_72,In_435);
and U300 (N_300,In_213,In_521);
and U301 (N_301,In_304,In_654);
and U302 (N_302,In_323,In_593);
or U303 (N_303,In_338,In_87);
or U304 (N_304,In_363,In_508);
nor U305 (N_305,In_365,In_303);
xnor U306 (N_306,In_370,In_290);
xnor U307 (N_307,In_529,In_413);
nand U308 (N_308,In_91,In_79);
nor U309 (N_309,In_41,In_503);
or U310 (N_310,In_394,In_664);
or U311 (N_311,In_446,In_296);
or U312 (N_312,In_164,In_687);
nor U313 (N_313,In_715,In_518);
nand U314 (N_314,In_185,In_719);
nor U315 (N_315,In_749,In_739);
xnor U316 (N_316,In_223,In_284);
nand U317 (N_317,In_609,In_37);
xnor U318 (N_318,In_450,In_592);
nor U319 (N_319,In_242,In_351);
xor U320 (N_320,In_381,In_590);
and U321 (N_321,In_576,In_278);
nor U322 (N_322,In_131,In_136);
nand U323 (N_323,In_517,In_459);
nor U324 (N_324,In_585,In_417);
nor U325 (N_325,In_575,In_165);
and U326 (N_326,In_54,In_99);
xor U327 (N_327,In_649,In_382);
or U328 (N_328,In_655,In_605);
xnor U329 (N_329,In_574,In_236);
xor U330 (N_330,In_42,In_489);
and U331 (N_331,In_51,In_470);
xnor U332 (N_332,In_404,In_134);
and U333 (N_333,In_330,In_504);
nor U334 (N_334,In_166,In_443);
xnor U335 (N_335,In_453,In_714);
and U336 (N_336,In_356,In_289);
nand U337 (N_337,In_492,In_109);
nand U338 (N_338,In_744,In_157);
and U339 (N_339,In_636,In_502);
nand U340 (N_340,In_247,In_222);
and U341 (N_341,In_316,In_260);
and U342 (N_342,In_669,In_720);
nand U343 (N_343,In_366,In_14);
xor U344 (N_344,In_391,In_49);
xnor U345 (N_345,In_505,In_345);
xnor U346 (N_346,In_319,In_244);
and U347 (N_347,In_407,In_441);
or U348 (N_348,In_30,In_646);
or U349 (N_349,In_496,In_228);
nor U350 (N_350,In_452,In_535);
nand U351 (N_351,In_315,In_509);
nor U352 (N_352,In_519,In_662);
nand U353 (N_353,In_612,In_16);
nor U354 (N_354,In_352,In_133);
nand U355 (N_355,In_430,In_169);
xor U356 (N_356,In_342,In_60);
or U357 (N_357,In_395,In_203);
nand U358 (N_358,In_414,In_579);
and U359 (N_359,In_182,In_149);
nor U360 (N_360,In_434,In_561);
nor U361 (N_361,In_559,In_364);
or U362 (N_362,In_300,In_265);
nand U363 (N_363,In_360,In_416);
xnor U364 (N_364,In_411,In_277);
or U365 (N_365,In_101,In_321);
and U366 (N_366,In_727,In_490);
nand U367 (N_367,In_82,In_651);
nor U368 (N_368,In_573,In_525);
or U369 (N_369,In_466,In_229);
and U370 (N_370,In_113,In_512);
nand U371 (N_371,In_245,In_745);
xnor U372 (N_372,In_314,In_710);
xor U373 (N_373,In_259,In_88);
and U374 (N_374,In_226,In_695);
xnor U375 (N_375,In_600,In_174);
nor U376 (N_376,In_363,In_312);
xnor U377 (N_377,In_576,In_1);
nand U378 (N_378,In_711,In_577);
xnor U379 (N_379,In_441,In_408);
and U380 (N_380,In_178,In_580);
and U381 (N_381,In_121,In_501);
xnor U382 (N_382,In_7,In_173);
xor U383 (N_383,In_233,In_100);
nand U384 (N_384,In_13,In_734);
and U385 (N_385,In_232,In_142);
and U386 (N_386,In_385,In_340);
or U387 (N_387,In_441,In_557);
or U388 (N_388,In_209,In_297);
nand U389 (N_389,In_419,In_580);
xnor U390 (N_390,In_169,In_608);
xnor U391 (N_391,In_522,In_519);
and U392 (N_392,In_53,In_455);
xnor U393 (N_393,In_88,In_363);
nand U394 (N_394,In_220,In_283);
nor U395 (N_395,In_470,In_586);
xnor U396 (N_396,In_518,In_537);
nor U397 (N_397,In_28,In_68);
and U398 (N_398,In_60,In_270);
nand U399 (N_399,In_616,In_54);
xnor U400 (N_400,In_616,In_386);
and U401 (N_401,In_737,In_133);
nand U402 (N_402,In_189,In_326);
and U403 (N_403,In_205,In_229);
or U404 (N_404,In_111,In_599);
xnor U405 (N_405,In_478,In_218);
nor U406 (N_406,In_380,In_94);
and U407 (N_407,In_128,In_17);
and U408 (N_408,In_323,In_488);
and U409 (N_409,In_492,In_369);
or U410 (N_410,In_591,In_451);
xor U411 (N_411,In_472,In_494);
nor U412 (N_412,In_511,In_698);
nor U413 (N_413,In_373,In_225);
and U414 (N_414,In_388,In_611);
and U415 (N_415,In_691,In_598);
and U416 (N_416,In_72,In_8);
or U417 (N_417,In_565,In_573);
nor U418 (N_418,In_138,In_2);
xnor U419 (N_419,In_490,In_623);
or U420 (N_420,In_157,In_101);
xor U421 (N_421,In_552,In_566);
xor U422 (N_422,In_719,In_113);
or U423 (N_423,In_354,In_255);
nor U424 (N_424,In_347,In_664);
nor U425 (N_425,In_213,In_684);
nand U426 (N_426,In_315,In_212);
or U427 (N_427,In_424,In_261);
nor U428 (N_428,In_679,In_668);
nor U429 (N_429,In_42,In_540);
and U430 (N_430,In_660,In_349);
nand U431 (N_431,In_502,In_405);
and U432 (N_432,In_36,In_499);
nor U433 (N_433,In_11,In_76);
nor U434 (N_434,In_257,In_353);
or U435 (N_435,In_594,In_330);
nor U436 (N_436,In_260,In_741);
nand U437 (N_437,In_651,In_244);
and U438 (N_438,In_376,In_2);
nand U439 (N_439,In_183,In_656);
nor U440 (N_440,In_581,In_434);
nor U441 (N_441,In_568,In_165);
nand U442 (N_442,In_469,In_472);
xnor U443 (N_443,In_60,In_429);
xor U444 (N_444,In_55,In_432);
and U445 (N_445,In_399,In_343);
or U446 (N_446,In_255,In_643);
or U447 (N_447,In_31,In_70);
or U448 (N_448,In_674,In_483);
nand U449 (N_449,In_70,In_336);
xor U450 (N_450,In_382,In_76);
and U451 (N_451,In_558,In_733);
nand U452 (N_452,In_542,In_166);
and U453 (N_453,In_405,In_168);
or U454 (N_454,In_445,In_240);
xnor U455 (N_455,In_709,In_637);
xnor U456 (N_456,In_311,In_7);
nand U457 (N_457,In_125,In_629);
xor U458 (N_458,In_254,In_650);
xor U459 (N_459,In_483,In_409);
nor U460 (N_460,In_558,In_284);
or U461 (N_461,In_342,In_119);
or U462 (N_462,In_399,In_357);
nor U463 (N_463,In_521,In_313);
nand U464 (N_464,In_747,In_378);
xnor U465 (N_465,In_365,In_125);
nand U466 (N_466,In_243,In_67);
and U467 (N_467,In_167,In_346);
and U468 (N_468,In_74,In_640);
nor U469 (N_469,In_694,In_330);
xor U470 (N_470,In_41,In_323);
xor U471 (N_471,In_596,In_474);
or U472 (N_472,In_121,In_691);
nand U473 (N_473,In_306,In_325);
and U474 (N_474,In_522,In_620);
and U475 (N_475,In_633,In_334);
or U476 (N_476,In_430,In_245);
xnor U477 (N_477,In_294,In_305);
xnor U478 (N_478,In_160,In_571);
xor U479 (N_479,In_510,In_143);
or U480 (N_480,In_43,In_338);
nor U481 (N_481,In_189,In_67);
or U482 (N_482,In_408,In_742);
xnor U483 (N_483,In_116,In_537);
xor U484 (N_484,In_18,In_403);
and U485 (N_485,In_234,In_332);
or U486 (N_486,In_363,In_292);
and U487 (N_487,In_453,In_309);
or U488 (N_488,In_12,In_405);
or U489 (N_489,In_415,In_342);
xor U490 (N_490,In_737,In_117);
or U491 (N_491,In_533,In_137);
nand U492 (N_492,In_514,In_121);
and U493 (N_493,In_515,In_384);
nor U494 (N_494,In_315,In_222);
and U495 (N_495,In_50,In_21);
nor U496 (N_496,In_554,In_308);
xnor U497 (N_497,In_235,In_266);
nor U498 (N_498,In_177,In_25);
xnor U499 (N_499,In_145,In_600);
and U500 (N_500,In_586,In_588);
xnor U501 (N_501,In_52,In_335);
nor U502 (N_502,In_617,In_725);
nor U503 (N_503,In_563,In_339);
and U504 (N_504,In_169,In_653);
nand U505 (N_505,In_685,In_488);
xnor U506 (N_506,In_74,In_701);
and U507 (N_507,In_401,In_316);
xor U508 (N_508,In_233,In_556);
xnor U509 (N_509,In_456,In_201);
nor U510 (N_510,In_625,In_309);
nand U511 (N_511,In_303,In_235);
nand U512 (N_512,In_721,In_385);
and U513 (N_513,In_202,In_638);
nor U514 (N_514,In_639,In_329);
xor U515 (N_515,In_324,In_511);
nor U516 (N_516,In_402,In_700);
nand U517 (N_517,In_574,In_490);
xnor U518 (N_518,In_340,In_354);
or U519 (N_519,In_636,In_651);
or U520 (N_520,In_528,In_84);
nand U521 (N_521,In_120,In_421);
and U522 (N_522,In_730,In_13);
and U523 (N_523,In_261,In_508);
nand U524 (N_524,In_87,In_506);
nand U525 (N_525,In_424,In_716);
nor U526 (N_526,In_683,In_739);
nand U527 (N_527,In_383,In_443);
or U528 (N_528,In_207,In_277);
and U529 (N_529,In_236,In_369);
nand U530 (N_530,In_389,In_564);
and U531 (N_531,In_512,In_281);
nand U532 (N_532,In_241,In_389);
and U533 (N_533,In_692,In_438);
xnor U534 (N_534,In_568,In_113);
or U535 (N_535,In_195,In_62);
nor U536 (N_536,In_98,In_285);
or U537 (N_537,In_654,In_384);
or U538 (N_538,In_100,In_427);
or U539 (N_539,In_666,In_681);
or U540 (N_540,In_177,In_299);
or U541 (N_541,In_345,In_131);
or U542 (N_542,In_687,In_116);
nand U543 (N_543,In_655,In_352);
xor U544 (N_544,In_336,In_539);
and U545 (N_545,In_424,In_658);
xor U546 (N_546,In_439,In_335);
or U547 (N_547,In_724,In_552);
xor U548 (N_548,In_451,In_731);
or U549 (N_549,In_592,In_92);
or U550 (N_550,In_336,In_242);
nor U551 (N_551,In_451,In_419);
nand U552 (N_552,In_22,In_595);
and U553 (N_553,In_630,In_524);
nand U554 (N_554,In_208,In_473);
xor U555 (N_555,In_298,In_24);
nor U556 (N_556,In_104,In_580);
or U557 (N_557,In_516,In_515);
and U558 (N_558,In_387,In_8);
nor U559 (N_559,In_200,In_309);
xnor U560 (N_560,In_592,In_728);
nor U561 (N_561,In_608,In_636);
xnor U562 (N_562,In_327,In_64);
xnor U563 (N_563,In_289,In_160);
nor U564 (N_564,In_551,In_745);
and U565 (N_565,In_533,In_222);
and U566 (N_566,In_511,In_550);
nor U567 (N_567,In_635,In_353);
or U568 (N_568,In_615,In_705);
or U569 (N_569,In_197,In_458);
nor U570 (N_570,In_339,In_593);
or U571 (N_571,In_360,In_699);
xor U572 (N_572,In_206,In_487);
nor U573 (N_573,In_721,In_387);
xnor U574 (N_574,In_592,In_609);
and U575 (N_575,In_337,In_324);
or U576 (N_576,In_413,In_185);
nand U577 (N_577,In_60,In_612);
xor U578 (N_578,In_2,In_438);
xor U579 (N_579,In_83,In_575);
xor U580 (N_580,In_456,In_222);
nor U581 (N_581,In_420,In_3);
or U582 (N_582,In_520,In_515);
xor U583 (N_583,In_741,In_611);
or U584 (N_584,In_71,In_610);
and U585 (N_585,In_353,In_181);
xnor U586 (N_586,In_154,In_610);
nor U587 (N_587,In_142,In_365);
and U588 (N_588,In_182,In_408);
nor U589 (N_589,In_386,In_316);
nand U590 (N_590,In_258,In_68);
and U591 (N_591,In_725,In_717);
or U592 (N_592,In_227,In_164);
or U593 (N_593,In_471,In_291);
nand U594 (N_594,In_314,In_212);
nor U595 (N_595,In_715,In_55);
nor U596 (N_596,In_170,In_461);
and U597 (N_597,In_433,In_279);
xnor U598 (N_598,In_654,In_88);
nand U599 (N_599,In_472,In_322);
or U600 (N_600,In_315,In_258);
and U601 (N_601,In_236,In_193);
nand U602 (N_602,In_695,In_59);
and U603 (N_603,In_175,In_637);
or U604 (N_604,In_16,In_227);
nand U605 (N_605,In_686,In_423);
xor U606 (N_606,In_343,In_731);
xnor U607 (N_607,In_631,In_243);
nor U608 (N_608,In_699,In_496);
nor U609 (N_609,In_15,In_316);
nand U610 (N_610,In_105,In_405);
and U611 (N_611,In_351,In_661);
nand U612 (N_612,In_515,In_288);
or U613 (N_613,In_5,In_657);
nand U614 (N_614,In_460,In_364);
nor U615 (N_615,In_435,In_127);
and U616 (N_616,In_499,In_359);
nand U617 (N_617,In_176,In_82);
nor U618 (N_618,In_351,In_544);
nor U619 (N_619,In_102,In_470);
and U620 (N_620,In_595,In_600);
or U621 (N_621,In_396,In_566);
or U622 (N_622,In_268,In_447);
xor U623 (N_623,In_140,In_265);
xor U624 (N_624,In_699,In_593);
xor U625 (N_625,In_301,In_413);
nor U626 (N_626,In_357,In_187);
or U627 (N_627,In_255,In_358);
or U628 (N_628,In_545,In_166);
nand U629 (N_629,In_676,In_686);
and U630 (N_630,In_491,In_8);
xor U631 (N_631,In_374,In_257);
nand U632 (N_632,In_193,In_569);
and U633 (N_633,In_274,In_389);
or U634 (N_634,In_287,In_394);
xor U635 (N_635,In_168,In_509);
or U636 (N_636,In_618,In_296);
nand U637 (N_637,In_250,In_47);
and U638 (N_638,In_583,In_721);
and U639 (N_639,In_51,In_59);
nor U640 (N_640,In_484,In_62);
nand U641 (N_641,In_323,In_475);
and U642 (N_642,In_642,In_182);
or U643 (N_643,In_400,In_458);
nand U644 (N_644,In_254,In_576);
or U645 (N_645,In_682,In_83);
or U646 (N_646,In_469,In_493);
and U647 (N_647,In_273,In_309);
nand U648 (N_648,In_585,In_246);
xnor U649 (N_649,In_482,In_615);
nand U650 (N_650,In_580,In_106);
or U651 (N_651,In_292,In_707);
or U652 (N_652,In_71,In_679);
and U653 (N_653,In_459,In_401);
nor U654 (N_654,In_152,In_589);
nand U655 (N_655,In_116,In_703);
or U656 (N_656,In_284,In_349);
and U657 (N_657,In_428,In_351);
and U658 (N_658,In_438,In_500);
xnor U659 (N_659,In_23,In_678);
nor U660 (N_660,In_93,In_421);
or U661 (N_661,In_121,In_46);
nand U662 (N_662,In_505,In_74);
and U663 (N_663,In_404,In_583);
xnor U664 (N_664,In_580,In_285);
nand U665 (N_665,In_428,In_189);
and U666 (N_666,In_227,In_521);
nor U667 (N_667,In_15,In_121);
and U668 (N_668,In_633,In_162);
xnor U669 (N_669,In_484,In_356);
nand U670 (N_670,In_81,In_738);
nand U671 (N_671,In_732,In_55);
or U672 (N_672,In_347,In_420);
xor U673 (N_673,In_316,In_457);
or U674 (N_674,In_694,In_661);
and U675 (N_675,In_569,In_318);
xnor U676 (N_676,In_192,In_356);
xnor U677 (N_677,In_748,In_505);
nor U678 (N_678,In_315,In_506);
or U679 (N_679,In_610,In_345);
nand U680 (N_680,In_442,In_194);
or U681 (N_681,In_17,In_312);
and U682 (N_682,In_72,In_693);
or U683 (N_683,In_171,In_631);
or U684 (N_684,In_412,In_333);
nand U685 (N_685,In_192,In_399);
nor U686 (N_686,In_434,In_603);
and U687 (N_687,In_262,In_543);
nor U688 (N_688,In_671,In_746);
or U689 (N_689,In_715,In_21);
nor U690 (N_690,In_524,In_97);
nand U691 (N_691,In_33,In_733);
xor U692 (N_692,In_720,In_202);
or U693 (N_693,In_287,In_406);
nand U694 (N_694,In_310,In_387);
nand U695 (N_695,In_126,In_21);
or U696 (N_696,In_211,In_695);
nor U697 (N_697,In_573,In_342);
xnor U698 (N_698,In_133,In_172);
or U699 (N_699,In_521,In_73);
and U700 (N_700,In_583,In_498);
and U701 (N_701,In_698,In_357);
xor U702 (N_702,In_735,In_210);
xor U703 (N_703,In_680,In_10);
nand U704 (N_704,In_85,In_198);
nand U705 (N_705,In_749,In_237);
xnor U706 (N_706,In_345,In_568);
xnor U707 (N_707,In_434,In_736);
nand U708 (N_708,In_424,In_45);
nand U709 (N_709,In_16,In_425);
nor U710 (N_710,In_264,In_131);
nand U711 (N_711,In_628,In_12);
xor U712 (N_712,In_240,In_577);
nor U713 (N_713,In_610,In_728);
or U714 (N_714,In_697,In_679);
and U715 (N_715,In_36,In_91);
nor U716 (N_716,In_38,In_596);
nand U717 (N_717,In_274,In_688);
xor U718 (N_718,In_158,In_284);
and U719 (N_719,In_592,In_608);
nor U720 (N_720,In_662,In_3);
nor U721 (N_721,In_265,In_383);
nand U722 (N_722,In_426,In_247);
nand U723 (N_723,In_63,In_726);
nand U724 (N_724,In_603,In_671);
or U725 (N_725,In_132,In_223);
xnor U726 (N_726,In_296,In_652);
and U727 (N_727,In_360,In_248);
nand U728 (N_728,In_288,In_127);
nor U729 (N_729,In_119,In_95);
nand U730 (N_730,In_192,In_62);
nor U731 (N_731,In_364,In_446);
nor U732 (N_732,In_462,In_273);
nor U733 (N_733,In_182,In_334);
xor U734 (N_734,In_289,In_428);
nor U735 (N_735,In_50,In_687);
nand U736 (N_736,In_625,In_519);
or U737 (N_737,In_602,In_620);
xnor U738 (N_738,In_637,In_743);
or U739 (N_739,In_324,In_581);
or U740 (N_740,In_501,In_389);
and U741 (N_741,In_712,In_286);
nor U742 (N_742,In_299,In_339);
xnor U743 (N_743,In_311,In_259);
and U744 (N_744,In_28,In_498);
or U745 (N_745,In_380,In_726);
and U746 (N_746,In_284,In_566);
or U747 (N_747,In_607,In_369);
and U748 (N_748,In_273,In_221);
nand U749 (N_749,In_544,In_35);
xnor U750 (N_750,In_643,In_735);
or U751 (N_751,In_206,In_208);
and U752 (N_752,In_95,In_608);
nor U753 (N_753,In_414,In_173);
xnor U754 (N_754,In_13,In_473);
xor U755 (N_755,In_640,In_371);
or U756 (N_756,In_534,In_207);
xnor U757 (N_757,In_474,In_637);
xnor U758 (N_758,In_161,In_405);
nand U759 (N_759,In_320,In_345);
nand U760 (N_760,In_542,In_291);
nand U761 (N_761,In_498,In_505);
nand U762 (N_762,In_545,In_359);
or U763 (N_763,In_551,In_179);
and U764 (N_764,In_349,In_550);
xnor U765 (N_765,In_683,In_347);
or U766 (N_766,In_491,In_427);
nand U767 (N_767,In_26,In_580);
nor U768 (N_768,In_609,In_506);
nand U769 (N_769,In_428,In_358);
and U770 (N_770,In_673,In_52);
and U771 (N_771,In_355,In_651);
and U772 (N_772,In_297,In_717);
nor U773 (N_773,In_157,In_695);
and U774 (N_774,In_168,In_42);
xnor U775 (N_775,In_7,In_619);
nand U776 (N_776,In_533,In_650);
nand U777 (N_777,In_55,In_35);
or U778 (N_778,In_433,In_593);
or U779 (N_779,In_450,In_442);
xor U780 (N_780,In_423,In_87);
nand U781 (N_781,In_196,In_560);
nand U782 (N_782,In_327,In_175);
nand U783 (N_783,In_486,In_184);
and U784 (N_784,In_19,In_95);
nand U785 (N_785,In_643,In_636);
nand U786 (N_786,In_554,In_458);
nor U787 (N_787,In_365,In_91);
and U788 (N_788,In_631,In_184);
nand U789 (N_789,In_484,In_239);
nand U790 (N_790,In_726,In_722);
and U791 (N_791,In_419,In_508);
xnor U792 (N_792,In_19,In_83);
nand U793 (N_793,In_263,In_271);
xor U794 (N_794,In_743,In_620);
xnor U795 (N_795,In_559,In_738);
nor U796 (N_796,In_699,In_510);
nand U797 (N_797,In_534,In_374);
or U798 (N_798,In_123,In_591);
and U799 (N_799,In_719,In_95);
nand U800 (N_800,In_489,In_95);
and U801 (N_801,In_194,In_722);
xor U802 (N_802,In_704,In_259);
and U803 (N_803,In_493,In_629);
nor U804 (N_804,In_528,In_687);
or U805 (N_805,In_179,In_125);
and U806 (N_806,In_192,In_45);
xnor U807 (N_807,In_299,In_544);
or U808 (N_808,In_662,In_6);
nand U809 (N_809,In_525,In_454);
nand U810 (N_810,In_734,In_173);
and U811 (N_811,In_76,In_116);
and U812 (N_812,In_639,In_159);
and U813 (N_813,In_544,In_230);
or U814 (N_814,In_371,In_641);
xor U815 (N_815,In_468,In_102);
nand U816 (N_816,In_111,In_530);
nand U817 (N_817,In_38,In_615);
xnor U818 (N_818,In_342,In_427);
nand U819 (N_819,In_537,In_695);
nor U820 (N_820,In_414,In_361);
nand U821 (N_821,In_248,In_638);
xor U822 (N_822,In_354,In_562);
nor U823 (N_823,In_307,In_409);
xor U824 (N_824,In_85,In_202);
nor U825 (N_825,In_52,In_541);
and U826 (N_826,In_457,In_488);
xor U827 (N_827,In_574,In_388);
nor U828 (N_828,In_736,In_653);
nor U829 (N_829,In_685,In_283);
and U830 (N_830,In_431,In_118);
or U831 (N_831,In_391,In_575);
and U832 (N_832,In_293,In_439);
or U833 (N_833,In_735,In_290);
and U834 (N_834,In_562,In_362);
or U835 (N_835,In_49,In_565);
nand U836 (N_836,In_54,In_574);
or U837 (N_837,In_497,In_382);
nor U838 (N_838,In_76,In_674);
nor U839 (N_839,In_192,In_214);
and U840 (N_840,In_636,In_151);
nor U841 (N_841,In_81,In_714);
or U842 (N_842,In_612,In_524);
nor U843 (N_843,In_388,In_115);
nor U844 (N_844,In_368,In_109);
or U845 (N_845,In_45,In_744);
and U846 (N_846,In_65,In_526);
nor U847 (N_847,In_133,In_435);
xnor U848 (N_848,In_82,In_670);
nor U849 (N_849,In_356,In_507);
xor U850 (N_850,In_90,In_260);
nand U851 (N_851,In_559,In_365);
nor U852 (N_852,In_580,In_701);
nand U853 (N_853,In_484,In_197);
and U854 (N_854,In_511,In_237);
and U855 (N_855,In_590,In_644);
xnor U856 (N_856,In_95,In_470);
and U857 (N_857,In_570,In_363);
or U858 (N_858,In_322,In_202);
and U859 (N_859,In_562,In_79);
or U860 (N_860,In_87,In_239);
xnor U861 (N_861,In_590,In_650);
nand U862 (N_862,In_499,In_461);
nand U863 (N_863,In_13,In_296);
xnor U864 (N_864,In_145,In_98);
xor U865 (N_865,In_615,In_30);
and U866 (N_866,In_157,In_450);
xor U867 (N_867,In_364,In_101);
and U868 (N_868,In_670,In_714);
nor U869 (N_869,In_476,In_81);
nor U870 (N_870,In_167,In_507);
xor U871 (N_871,In_651,In_204);
xor U872 (N_872,In_702,In_37);
or U873 (N_873,In_188,In_124);
nand U874 (N_874,In_470,In_195);
or U875 (N_875,In_599,In_304);
xor U876 (N_876,In_350,In_433);
nor U877 (N_877,In_671,In_38);
or U878 (N_878,In_416,In_140);
xnor U879 (N_879,In_180,In_167);
or U880 (N_880,In_261,In_157);
nand U881 (N_881,In_45,In_63);
nand U882 (N_882,In_370,In_147);
xor U883 (N_883,In_507,In_60);
or U884 (N_884,In_244,In_693);
and U885 (N_885,In_711,In_316);
nor U886 (N_886,In_235,In_87);
nand U887 (N_887,In_75,In_187);
and U888 (N_888,In_260,In_711);
xnor U889 (N_889,In_250,In_653);
or U890 (N_890,In_596,In_570);
nor U891 (N_891,In_407,In_163);
or U892 (N_892,In_569,In_132);
or U893 (N_893,In_536,In_644);
and U894 (N_894,In_585,In_693);
nor U895 (N_895,In_644,In_179);
and U896 (N_896,In_174,In_461);
nand U897 (N_897,In_378,In_9);
nor U898 (N_898,In_70,In_520);
or U899 (N_899,In_701,In_610);
and U900 (N_900,In_379,In_578);
and U901 (N_901,In_12,In_354);
or U902 (N_902,In_97,In_659);
and U903 (N_903,In_667,In_331);
nor U904 (N_904,In_254,In_374);
or U905 (N_905,In_525,In_536);
or U906 (N_906,In_635,In_316);
or U907 (N_907,In_218,In_703);
nand U908 (N_908,In_276,In_744);
xnor U909 (N_909,In_732,In_683);
or U910 (N_910,In_363,In_253);
and U911 (N_911,In_399,In_220);
and U912 (N_912,In_516,In_323);
and U913 (N_913,In_671,In_403);
and U914 (N_914,In_386,In_97);
xnor U915 (N_915,In_174,In_641);
nor U916 (N_916,In_408,In_278);
xor U917 (N_917,In_211,In_171);
and U918 (N_918,In_436,In_116);
and U919 (N_919,In_14,In_612);
or U920 (N_920,In_405,In_176);
nor U921 (N_921,In_108,In_543);
nor U922 (N_922,In_38,In_73);
nor U923 (N_923,In_86,In_677);
nor U924 (N_924,In_638,In_121);
or U925 (N_925,In_728,In_125);
nor U926 (N_926,In_0,In_716);
and U927 (N_927,In_737,In_708);
nand U928 (N_928,In_317,In_590);
and U929 (N_929,In_243,In_655);
and U930 (N_930,In_439,In_176);
or U931 (N_931,In_741,In_729);
or U932 (N_932,In_341,In_668);
or U933 (N_933,In_140,In_743);
nor U934 (N_934,In_132,In_708);
xor U935 (N_935,In_652,In_687);
and U936 (N_936,In_534,In_301);
or U937 (N_937,In_385,In_591);
nand U938 (N_938,In_747,In_416);
xor U939 (N_939,In_151,In_452);
or U940 (N_940,In_293,In_490);
nor U941 (N_941,In_545,In_122);
nor U942 (N_942,In_318,In_606);
nor U943 (N_943,In_600,In_657);
and U944 (N_944,In_205,In_76);
or U945 (N_945,In_475,In_104);
xnor U946 (N_946,In_743,In_672);
nand U947 (N_947,In_400,In_121);
xor U948 (N_948,In_170,In_112);
nand U949 (N_949,In_105,In_464);
xor U950 (N_950,In_30,In_207);
nand U951 (N_951,In_573,In_696);
nor U952 (N_952,In_221,In_379);
nand U953 (N_953,In_500,In_651);
or U954 (N_954,In_165,In_4);
nor U955 (N_955,In_260,In_495);
or U956 (N_956,In_31,In_599);
nand U957 (N_957,In_350,In_361);
and U958 (N_958,In_660,In_684);
and U959 (N_959,In_356,In_132);
nor U960 (N_960,In_13,In_701);
xor U961 (N_961,In_655,In_583);
nor U962 (N_962,In_588,In_297);
or U963 (N_963,In_597,In_72);
nand U964 (N_964,In_568,In_212);
xor U965 (N_965,In_566,In_189);
and U966 (N_966,In_31,In_501);
or U967 (N_967,In_75,In_324);
xnor U968 (N_968,In_508,In_124);
xnor U969 (N_969,In_110,In_577);
nor U970 (N_970,In_448,In_246);
or U971 (N_971,In_0,In_34);
xnor U972 (N_972,In_217,In_301);
xor U973 (N_973,In_10,In_491);
and U974 (N_974,In_132,In_319);
nor U975 (N_975,In_325,In_572);
and U976 (N_976,In_712,In_496);
xnor U977 (N_977,In_520,In_287);
nand U978 (N_978,In_609,In_407);
nor U979 (N_979,In_642,In_493);
xor U980 (N_980,In_572,In_588);
nor U981 (N_981,In_165,In_447);
nor U982 (N_982,In_691,In_725);
nor U983 (N_983,In_147,In_310);
xor U984 (N_984,In_682,In_376);
nor U985 (N_985,In_455,In_554);
or U986 (N_986,In_493,In_242);
nand U987 (N_987,In_80,In_699);
xor U988 (N_988,In_746,In_90);
or U989 (N_989,In_234,In_657);
xor U990 (N_990,In_229,In_388);
xor U991 (N_991,In_34,In_303);
nand U992 (N_992,In_610,In_343);
or U993 (N_993,In_125,In_234);
nand U994 (N_994,In_327,In_513);
nand U995 (N_995,In_564,In_609);
nor U996 (N_996,In_381,In_591);
xor U997 (N_997,In_267,In_575);
or U998 (N_998,In_138,In_711);
nand U999 (N_999,In_688,In_421);
nand U1000 (N_1000,In_229,In_734);
nor U1001 (N_1001,In_548,In_152);
and U1002 (N_1002,In_496,In_442);
nor U1003 (N_1003,In_636,In_4);
or U1004 (N_1004,In_164,In_180);
or U1005 (N_1005,In_191,In_254);
nor U1006 (N_1006,In_348,In_251);
or U1007 (N_1007,In_261,In_473);
or U1008 (N_1008,In_84,In_653);
or U1009 (N_1009,In_441,In_708);
or U1010 (N_1010,In_465,In_744);
or U1011 (N_1011,In_122,In_17);
nor U1012 (N_1012,In_600,In_610);
and U1013 (N_1013,In_439,In_307);
nor U1014 (N_1014,In_206,In_142);
nor U1015 (N_1015,In_196,In_237);
xnor U1016 (N_1016,In_1,In_678);
or U1017 (N_1017,In_115,In_518);
nand U1018 (N_1018,In_435,In_398);
nand U1019 (N_1019,In_591,In_631);
nor U1020 (N_1020,In_42,In_581);
nor U1021 (N_1021,In_243,In_607);
or U1022 (N_1022,In_100,In_83);
and U1023 (N_1023,In_452,In_641);
nand U1024 (N_1024,In_738,In_313);
nand U1025 (N_1025,In_198,In_535);
nor U1026 (N_1026,In_531,In_207);
nor U1027 (N_1027,In_617,In_172);
or U1028 (N_1028,In_439,In_340);
or U1029 (N_1029,In_182,In_467);
nand U1030 (N_1030,In_139,In_9);
nand U1031 (N_1031,In_350,In_64);
xnor U1032 (N_1032,In_388,In_324);
xor U1033 (N_1033,In_239,In_500);
nor U1034 (N_1034,In_136,In_604);
or U1035 (N_1035,In_8,In_626);
xnor U1036 (N_1036,In_250,In_715);
xnor U1037 (N_1037,In_340,In_339);
and U1038 (N_1038,In_660,In_587);
or U1039 (N_1039,In_721,In_392);
nor U1040 (N_1040,In_328,In_532);
nand U1041 (N_1041,In_61,In_528);
and U1042 (N_1042,In_476,In_710);
and U1043 (N_1043,In_116,In_30);
nor U1044 (N_1044,In_701,In_123);
or U1045 (N_1045,In_107,In_472);
or U1046 (N_1046,In_251,In_7);
nor U1047 (N_1047,In_486,In_244);
nand U1048 (N_1048,In_312,In_554);
xor U1049 (N_1049,In_142,In_421);
xnor U1050 (N_1050,In_295,In_61);
xnor U1051 (N_1051,In_35,In_674);
or U1052 (N_1052,In_622,In_230);
or U1053 (N_1053,In_428,In_524);
or U1054 (N_1054,In_139,In_363);
nor U1055 (N_1055,In_65,In_6);
and U1056 (N_1056,In_392,In_706);
or U1057 (N_1057,In_717,In_100);
or U1058 (N_1058,In_69,In_585);
and U1059 (N_1059,In_744,In_487);
nand U1060 (N_1060,In_743,In_296);
nand U1061 (N_1061,In_354,In_611);
xnor U1062 (N_1062,In_332,In_126);
nor U1063 (N_1063,In_200,In_73);
nor U1064 (N_1064,In_433,In_581);
nand U1065 (N_1065,In_182,In_418);
nand U1066 (N_1066,In_715,In_325);
or U1067 (N_1067,In_203,In_470);
nor U1068 (N_1068,In_220,In_443);
and U1069 (N_1069,In_140,In_718);
nor U1070 (N_1070,In_307,In_99);
xor U1071 (N_1071,In_253,In_617);
or U1072 (N_1072,In_19,In_157);
and U1073 (N_1073,In_489,In_422);
or U1074 (N_1074,In_595,In_692);
nand U1075 (N_1075,In_462,In_111);
xnor U1076 (N_1076,In_480,In_225);
xor U1077 (N_1077,In_80,In_185);
xor U1078 (N_1078,In_191,In_60);
nor U1079 (N_1079,In_665,In_115);
or U1080 (N_1080,In_497,In_21);
nor U1081 (N_1081,In_11,In_475);
or U1082 (N_1082,In_83,In_270);
and U1083 (N_1083,In_463,In_653);
and U1084 (N_1084,In_378,In_645);
or U1085 (N_1085,In_355,In_700);
or U1086 (N_1086,In_593,In_169);
xor U1087 (N_1087,In_236,In_536);
nor U1088 (N_1088,In_652,In_336);
nor U1089 (N_1089,In_66,In_717);
and U1090 (N_1090,In_78,In_518);
xnor U1091 (N_1091,In_88,In_329);
nand U1092 (N_1092,In_555,In_192);
nand U1093 (N_1093,In_198,In_602);
nand U1094 (N_1094,In_682,In_19);
nand U1095 (N_1095,In_535,In_479);
and U1096 (N_1096,In_286,In_19);
nor U1097 (N_1097,In_517,In_257);
nand U1098 (N_1098,In_441,In_235);
nand U1099 (N_1099,In_721,In_647);
and U1100 (N_1100,In_332,In_43);
or U1101 (N_1101,In_276,In_691);
and U1102 (N_1102,In_64,In_550);
nor U1103 (N_1103,In_704,In_355);
xnor U1104 (N_1104,In_15,In_740);
nand U1105 (N_1105,In_13,In_38);
nand U1106 (N_1106,In_265,In_640);
xnor U1107 (N_1107,In_724,In_416);
or U1108 (N_1108,In_732,In_133);
nor U1109 (N_1109,In_603,In_139);
and U1110 (N_1110,In_185,In_208);
nor U1111 (N_1111,In_27,In_170);
or U1112 (N_1112,In_359,In_522);
and U1113 (N_1113,In_171,In_686);
nand U1114 (N_1114,In_554,In_510);
or U1115 (N_1115,In_661,In_573);
and U1116 (N_1116,In_654,In_22);
nand U1117 (N_1117,In_321,In_260);
or U1118 (N_1118,In_596,In_320);
nand U1119 (N_1119,In_465,In_65);
and U1120 (N_1120,In_26,In_573);
nor U1121 (N_1121,In_425,In_162);
nor U1122 (N_1122,In_537,In_17);
or U1123 (N_1123,In_678,In_430);
and U1124 (N_1124,In_13,In_302);
or U1125 (N_1125,In_514,In_219);
nor U1126 (N_1126,In_160,In_13);
or U1127 (N_1127,In_136,In_621);
nand U1128 (N_1128,In_211,In_727);
nor U1129 (N_1129,In_96,In_490);
and U1130 (N_1130,In_573,In_112);
or U1131 (N_1131,In_293,In_368);
nor U1132 (N_1132,In_360,In_278);
xnor U1133 (N_1133,In_515,In_328);
or U1134 (N_1134,In_229,In_394);
nor U1135 (N_1135,In_328,In_143);
xnor U1136 (N_1136,In_233,In_419);
and U1137 (N_1137,In_623,In_298);
and U1138 (N_1138,In_704,In_710);
xor U1139 (N_1139,In_50,In_89);
nand U1140 (N_1140,In_561,In_270);
and U1141 (N_1141,In_328,In_610);
or U1142 (N_1142,In_186,In_162);
nand U1143 (N_1143,In_637,In_550);
or U1144 (N_1144,In_467,In_654);
nor U1145 (N_1145,In_454,In_68);
nor U1146 (N_1146,In_171,In_691);
xnor U1147 (N_1147,In_451,In_148);
nor U1148 (N_1148,In_689,In_335);
xnor U1149 (N_1149,In_112,In_66);
nor U1150 (N_1150,In_106,In_551);
or U1151 (N_1151,In_634,In_12);
xnor U1152 (N_1152,In_325,In_589);
and U1153 (N_1153,In_545,In_375);
xnor U1154 (N_1154,In_23,In_165);
nand U1155 (N_1155,In_40,In_708);
nand U1156 (N_1156,In_721,In_371);
and U1157 (N_1157,In_324,In_273);
or U1158 (N_1158,In_389,In_32);
or U1159 (N_1159,In_730,In_532);
or U1160 (N_1160,In_421,In_733);
nand U1161 (N_1161,In_551,In_502);
and U1162 (N_1162,In_524,In_111);
and U1163 (N_1163,In_203,In_411);
xor U1164 (N_1164,In_208,In_313);
nand U1165 (N_1165,In_210,In_13);
or U1166 (N_1166,In_505,In_86);
nor U1167 (N_1167,In_302,In_246);
and U1168 (N_1168,In_627,In_543);
xor U1169 (N_1169,In_475,In_93);
and U1170 (N_1170,In_219,In_215);
nor U1171 (N_1171,In_31,In_626);
nand U1172 (N_1172,In_723,In_551);
and U1173 (N_1173,In_141,In_257);
nand U1174 (N_1174,In_445,In_709);
xnor U1175 (N_1175,In_304,In_694);
and U1176 (N_1176,In_237,In_340);
xnor U1177 (N_1177,In_127,In_84);
nor U1178 (N_1178,In_546,In_586);
xor U1179 (N_1179,In_384,In_671);
and U1180 (N_1180,In_375,In_187);
and U1181 (N_1181,In_377,In_689);
and U1182 (N_1182,In_552,In_57);
nand U1183 (N_1183,In_93,In_259);
nor U1184 (N_1184,In_717,In_452);
nor U1185 (N_1185,In_329,In_118);
or U1186 (N_1186,In_212,In_428);
and U1187 (N_1187,In_565,In_692);
and U1188 (N_1188,In_99,In_6);
nand U1189 (N_1189,In_493,In_618);
and U1190 (N_1190,In_33,In_203);
or U1191 (N_1191,In_79,In_614);
nand U1192 (N_1192,In_38,In_30);
nand U1193 (N_1193,In_7,In_428);
nand U1194 (N_1194,In_60,In_571);
or U1195 (N_1195,In_414,In_619);
nor U1196 (N_1196,In_470,In_353);
nor U1197 (N_1197,In_468,In_651);
and U1198 (N_1198,In_134,In_312);
nand U1199 (N_1199,In_149,In_186);
nand U1200 (N_1200,In_591,In_3);
nand U1201 (N_1201,In_427,In_478);
nor U1202 (N_1202,In_146,In_718);
or U1203 (N_1203,In_574,In_343);
nand U1204 (N_1204,In_139,In_164);
nand U1205 (N_1205,In_439,In_712);
nor U1206 (N_1206,In_569,In_80);
and U1207 (N_1207,In_17,In_591);
or U1208 (N_1208,In_725,In_600);
nand U1209 (N_1209,In_541,In_291);
xor U1210 (N_1210,In_468,In_163);
and U1211 (N_1211,In_86,In_666);
and U1212 (N_1212,In_524,In_143);
xnor U1213 (N_1213,In_147,In_686);
xor U1214 (N_1214,In_606,In_207);
or U1215 (N_1215,In_352,In_586);
nand U1216 (N_1216,In_518,In_284);
nand U1217 (N_1217,In_309,In_540);
nand U1218 (N_1218,In_90,In_602);
nand U1219 (N_1219,In_271,In_286);
nor U1220 (N_1220,In_7,In_113);
or U1221 (N_1221,In_175,In_529);
or U1222 (N_1222,In_222,In_697);
and U1223 (N_1223,In_140,In_81);
nand U1224 (N_1224,In_661,In_605);
or U1225 (N_1225,In_108,In_427);
nor U1226 (N_1226,In_132,In_627);
or U1227 (N_1227,In_315,In_225);
nor U1228 (N_1228,In_538,In_1);
nor U1229 (N_1229,In_611,In_401);
or U1230 (N_1230,In_233,In_133);
nor U1231 (N_1231,In_376,In_540);
or U1232 (N_1232,In_63,In_551);
nand U1233 (N_1233,In_145,In_2);
or U1234 (N_1234,In_470,In_381);
nand U1235 (N_1235,In_51,In_308);
nor U1236 (N_1236,In_234,In_606);
and U1237 (N_1237,In_546,In_393);
xnor U1238 (N_1238,In_179,In_637);
and U1239 (N_1239,In_407,In_555);
nor U1240 (N_1240,In_702,In_385);
xor U1241 (N_1241,In_351,In_602);
xnor U1242 (N_1242,In_513,In_292);
and U1243 (N_1243,In_121,In_398);
nor U1244 (N_1244,In_175,In_492);
nor U1245 (N_1245,In_76,In_505);
and U1246 (N_1246,In_477,In_512);
xnor U1247 (N_1247,In_19,In_57);
and U1248 (N_1248,In_22,In_354);
nor U1249 (N_1249,In_14,In_456);
xor U1250 (N_1250,In_421,In_368);
nand U1251 (N_1251,In_102,In_672);
nand U1252 (N_1252,In_450,In_570);
nor U1253 (N_1253,In_691,In_650);
nor U1254 (N_1254,In_54,In_716);
and U1255 (N_1255,In_749,In_48);
or U1256 (N_1256,In_601,In_711);
nor U1257 (N_1257,In_100,In_266);
nor U1258 (N_1258,In_68,In_420);
nor U1259 (N_1259,In_82,In_169);
or U1260 (N_1260,In_519,In_145);
and U1261 (N_1261,In_380,In_320);
nor U1262 (N_1262,In_569,In_109);
or U1263 (N_1263,In_654,In_179);
xor U1264 (N_1264,In_473,In_563);
nor U1265 (N_1265,In_294,In_415);
nand U1266 (N_1266,In_633,In_112);
nand U1267 (N_1267,In_620,In_228);
or U1268 (N_1268,In_447,In_318);
nand U1269 (N_1269,In_337,In_509);
nor U1270 (N_1270,In_82,In_482);
or U1271 (N_1271,In_580,In_468);
xor U1272 (N_1272,In_232,In_375);
or U1273 (N_1273,In_529,In_696);
xnor U1274 (N_1274,In_341,In_503);
nand U1275 (N_1275,In_161,In_189);
or U1276 (N_1276,In_135,In_381);
nor U1277 (N_1277,In_231,In_68);
nor U1278 (N_1278,In_626,In_244);
nor U1279 (N_1279,In_649,In_731);
nand U1280 (N_1280,In_428,In_622);
nor U1281 (N_1281,In_14,In_507);
nand U1282 (N_1282,In_383,In_15);
nor U1283 (N_1283,In_687,In_454);
or U1284 (N_1284,In_523,In_219);
and U1285 (N_1285,In_579,In_415);
nand U1286 (N_1286,In_139,In_744);
nor U1287 (N_1287,In_368,In_332);
xor U1288 (N_1288,In_407,In_304);
nor U1289 (N_1289,In_30,In_91);
and U1290 (N_1290,In_637,In_282);
nor U1291 (N_1291,In_420,In_49);
xor U1292 (N_1292,In_704,In_420);
or U1293 (N_1293,In_169,In_168);
xnor U1294 (N_1294,In_346,In_130);
xor U1295 (N_1295,In_140,In_111);
or U1296 (N_1296,In_236,In_1);
xnor U1297 (N_1297,In_657,In_207);
xnor U1298 (N_1298,In_341,In_356);
or U1299 (N_1299,In_450,In_282);
xnor U1300 (N_1300,In_517,In_364);
and U1301 (N_1301,In_342,In_534);
or U1302 (N_1302,In_703,In_139);
and U1303 (N_1303,In_293,In_364);
and U1304 (N_1304,In_79,In_452);
nor U1305 (N_1305,In_144,In_669);
and U1306 (N_1306,In_118,In_55);
and U1307 (N_1307,In_548,In_499);
nand U1308 (N_1308,In_580,In_700);
and U1309 (N_1309,In_617,In_622);
nor U1310 (N_1310,In_518,In_226);
and U1311 (N_1311,In_712,In_82);
xor U1312 (N_1312,In_94,In_4);
and U1313 (N_1313,In_357,In_707);
or U1314 (N_1314,In_625,In_568);
nand U1315 (N_1315,In_624,In_294);
nand U1316 (N_1316,In_673,In_188);
xnor U1317 (N_1317,In_729,In_710);
nor U1318 (N_1318,In_246,In_370);
or U1319 (N_1319,In_350,In_121);
or U1320 (N_1320,In_41,In_705);
xor U1321 (N_1321,In_182,In_696);
nor U1322 (N_1322,In_340,In_94);
and U1323 (N_1323,In_47,In_631);
or U1324 (N_1324,In_529,In_20);
nand U1325 (N_1325,In_616,In_246);
nor U1326 (N_1326,In_159,In_262);
xnor U1327 (N_1327,In_12,In_392);
or U1328 (N_1328,In_45,In_141);
nor U1329 (N_1329,In_241,In_119);
xnor U1330 (N_1330,In_310,In_705);
xor U1331 (N_1331,In_221,In_567);
xor U1332 (N_1332,In_19,In_715);
nor U1333 (N_1333,In_534,In_359);
nand U1334 (N_1334,In_267,In_739);
or U1335 (N_1335,In_613,In_503);
or U1336 (N_1336,In_228,In_33);
nor U1337 (N_1337,In_3,In_339);
xor U1338 (N_1338,In_458,In_647);
nand U1339 (N_1339,In_129,In_343);
or U1340 (N_1340,In_157,In_285);
nand U1341 (N_1341,In_133,In_298);
xor U1342 (N_1342,In_48,In_660);
or U1343 (N_1343,In_92,In_404);
nand U1344 (N_1344,In_291,In_268);
nand U1345 (N_1345,In_163,In_47);
and U1346 (N_1346,In_291,In_99);
nand U1347 (N_1347,In_55,In_277);
xor U1348 (N_1348,In_331,In_356);
or U1349 (N_1349,In_261,In_624);
and U1350 (N_1350,In_497,In_125);
nand U1351 (N_1351,In_56,In_263);
and U1352 (N_1352,In_441,In_313);
or U1353 (N_1353,In_295,In_470);
nor U1354 (N_1354,In_694,In_73);
or U1355 (N_1355,In_729,In_358);
and U1356 (N_1356,In_504,In_17);
and U1357 (N_1357,In_304,In_573);
xnor U1358 (N_1358,In_20,In_344);
xor U1359 (N_1359,In_679,In_196);
nand U1360 (N_1360,In_53,In_328);
nor U1361 (N_1361,In_692,In_334);
xnor U1362 (N_1362,In_34,In_411);
nor U1363 (N_1363,In_231,In_428);
xnor U1364 (N_1364,In_95,In_735);
nor U1365 (N_1365,In_472,In_234);
or U1366 (N_1366,In_584,In_380);
or U1367 (N_1367,In_475,In_166);
or U1368 (N_1368,In_321,In_580);
nor U1369 (N_1369,In_263,In_31);
nor U1370 (N_1370,In_243,In_72);
and U1371 (N_1371,In_35,In_114);
or U1372 (N_1372,In_376,In_723);
or U1373 (N_1373,In_396,In_470);
nand U1374 (N_1374,In_52,In_182);
nand U1375 (N_1375,In_3,In_107);
nor U1376 (N_1376,In_252,In_292);
nand U1377 (N_1377,In_50,In_166);
and U1378 (N_1378,In_169,In_446);
nand U1379 (N_1379,In_429,In_591);
or U1380 (N_1380,In_132,In_576);
nor U1381 (N_1381,In_442,In_207);
nor U1382 (N_1382,In_275,In_257);
nand U1383 (N_1383,In_522,In_176);
and U1384 (N_1384,In_327,In_690);
nand U1385 (N_1385,In_459,In_86);
or U1386 (N_1386,In_581,In_352);
or U1387 (N_1387,In_13,In_350);
or U1388 (N_1388,In_298,In_745);
or U1389 (N_1389,In_462,In_39);
nor U1390 (N_1390,In_346,In_728);
or U1391 (N_1391,In_443,In_38);
or U1392 (N_1392,In_289,In_117);
and U1393 (N_1393,In_461,In_704);
xnor U1394 (N_1394,In_71,In_267);
nor U1395 (N_1395,In_452,In_443);
nand U1396 (N_1396,In_299,In_294);
nand U1397 (N_1397,In_367,In_199);
or U1398 (N_1398,In_529,In_619);
nor U1399 (N_1399,In_224,In_287);
and U1400 (N_1400,In_523,In_651);
nand U1401 (N_1401,In_691,In_123);
and U1402 (N_1402,In_9,In_145);
or U1403 (N_1403,In_5,In_621);
nand U1404 (N_1404,In_689,In_460);
and U1405 (N_1405,In_713,In_87);
and U1406 (N_1406,In_191,In_396);
and U1407 (N_1407,In_517,In_493);
and U1408 (N_1408,In_543,In_166);
nor U1409 (N_1409,In_302,In_144);
xor U1410 (N_1410,In_508,In_420);
or U1411 (N_1411,In_607,In_537);
xnor U1412 (N_1412,In_576,In_604);
nand U1413 (N_1413,In_631,In_703);
nor U1414 (N_1414,In_550,In_514);
and U1415 (N_1415,In_411,In_280);
xor U1416 (N_1416,In_69,In_621);
xnor U1417 (N_1417,In_402,In_221);
nand U1418 (N_1418,In_446,In_206);
nor U1419 (N_1419,In_31,In_329);
or U1420 (N_1420,In_748,In_606);
nor U1421 (N_1421,In_299,In_34);
xnor U1422 (N_1422,In_108,In_698);
or U1423 (N_1423,In_455,In_439);
xor U1424 (N_1424,In_450,In_538);
nor U1425 (N_1425,In_276,In_318);
xnor U1426 (N_1426,In_512,In_544);
nand U1427 (N_1427,In_573,In_446);
nor U1428 (N_1428,In_646,In_66);
or U1429 (N_1429,In_80,In_35);
or U1430 (N_1430,In_511,In_280);
nor U1431 (N_1431,In_525,In_331);
or U1432 (N_1432,In_292,In_75);
nor U1433 (N_1433,In_333,In_449);
nor U1434 (N_1434,In_717,In_101);
nor U1435 (N_1435,In_644,In_144);
and U1436 (N_1436,In_117,In_357);
nand U1437 (N_1437,In_519,In_537);
nand U1438 (N_1438,In_617,In_322);
xnor U1439 (N_1439,In_190,In_671);
nand U1440 (N_1440,In_532,In_157);
nand U1441 (N_1441,In_634,In_135);
and U1442 (N_1442,In_48,In_400);
nor U1443 (N_1443,In_280,In_410);
or U1444 (N_1444,In_412,In_560);
and U1445 (N_1445,In_36,In_575);
nand U1446 (N_1446,In_556,In_175);
xor U1447 (N_1447,In_352,In_323);
and U1448 (N_1448,In_704,In_264);
and U1449 (N_1449,In_628,In_715);
nor U1450 (N_1450,In_172,In_698);
nand U1451 (N_1451,In_671,In_57);
and U1452 (N_1452,In_154,In_260);
nor U1453 (N_1453,In_60,In_615);
xnor U1454 (N_1454,In_560,In_606);
nand U1455 (N_1455,In_475,In_318);
nor U1456 (N_1456,In_724,In_697);
or U1457 (N_1457,In_61,In_175);
or U1458 (N_1458,In_543,In_672);
or U1459 (N_1459,In_352,In_331);
and U1460 (N_1460,In_561,In_25);
nor U1461 (N_1461,In_698,In_743);
and U1462 (N_1462,In_441,In_569);
or U1463 (N_1463,In_30,In_362);
and U1464 (N_1464,In_666,In_106);
xor U1465 (N_1465,In_287,In_703);
xor U1466 (N_1466,In_568,In_687);
or U1467 (N_1467,In_256,In_363);
nor U1468 (N_1468,In_76,In_501);
nor U1469 (N_1469,In_341,In_509);
or U1470 (N_1470,In_462,In_232);
xor U1471 (N_1471,In_661,In_469);
nor U1472 (N_1472,In_579,In_225);
xnor U1473 (N_1473,In_429,In_684);
nor U1474 (N_1474,In_525,In_290);
nor U1475 (N_1475,In_432,In_541);
or U1476 (N_1476,In_474,In_739);
nor U1477 (N_1477,In_728,In_534);
or U1478 (N_1478,In_443,In_136);
xor U1479 (N_1479,In_670,In_482);
xnor U1480 (N_1480,In_393,In_221);
and U1481 (N_1481,In_42,In_234);
nor U1482 (N_1482,In_479,In_88);
or U1483 (N_1483,In_414,In_440);
nor U1484 (N_1484,In_449,In_461);
xor U1485 (N_1485,In_397,In_662);
or U1486 (N_1486,In_622,In_359);
or U1487 (N_1487,In_169,In_552);
xor U1488 (N_1488,In_512,In_325);
xor U1489 (N_1489,In_722,In_331);
nand U1490 (N_1490,In_297,In_93);
nor U1491 (N_1491,In_118,In_481);
xor U1492 (N_1492,In_572,In_707);
and U1493 (N_1493,In_124,In_598);
nand U1494 (N_1494,In_61,In_368);
and U1495 (N_1495,In_212,In_192);
and U1496 (N_1496,In_710,In_648);
xor U1497 (N_1497,In_612,In_36);
nor U1498 (N_1498,In_133,In_291);
nor U1499 (N_1499,In_6,In_461);
and U1500 (N_1500,In_563,In_722);
and U1501 (N_1501,In_279,In_334);
nor U1502 (N_1502,In_379,In_685);
or U1503 (N_1503,In_257,In_453);
or U1504 (N_1504,In_487,In_403);
or U1505 (N_1505,In_80,In_348);
and U1506 (N_1506,In_341,In_290);
nor U1507 (N_1507,In_404,In_22);
nand U1508 (N_1508,In_408,In_319);
and U1509 (N_1509,In_224,In_352);
nand U1510 (N_1510,In_119,In_400);
xnor U1511 (N_1511,In_278,In_97);
and U1512 (N_1512,In_296,In_445);
nand U1513 (N_1513,In_38,In_442);
nand U1514 (N_1514,In_516,In_552);
xor U1515 (N_1515,In_53,In_18);
nor U1516 (N_1516,In_258,In_242);
and U1517 (N_1517,In_524,In_736);
nand U1518 (N_1518,In_289,In_0);
or U1519 (N_1519,In_341,In_101);
nand U1520 (N_1520,In_91,In_620);
and U1521 (N_1521,In_102,In_79);
xor U1522 (N_1522,In_453,In_588);
nand U1523 (N_1523,In_330,In_494);
or U1524 (N_1524,In_714,In_341);
nor U1525 (N_1525,In_329,In_307);
or U1526 (N_1526,In_83,In_300);
nor U1527 (N_1527,In_360,In_109);
nor U1528 (N_1528,In_609,In_65);
nand U1529 (N_1529,In_159,In_94);
nand U1530 (N_1530,In_22,In_460);
nand U1531 (N_1531,In_133,In_590);
nor U1532 (N_1532,In_387,In_430);
nand U1533 (N_1533,In_666,In_321);
nand U1534 (N_1534,In_595,In_425);
and U1535 (N_1535,In_524,In_527);
nor U1536 (N_1536,In_208,In_213);
and U1537 (N_1537,In_4,In_713);
or U1538 (N_1538,In_460,In_596);
xor U1539 (N_1539,In_544,In_82);
nand U1540 (N_1540,In_284,In_570);
xnor U1541 (N_1541,In_31,In_722);
xnor U1542 (N_1542,In_144,In_404);
and U1543 (N_1543,In_397,In_39);
xnor U1544 (N_1544,In_310,In_503);
xnor U1545 (N_1545,In_129,In_414);
xnor U1546 (N_1546,In_483,In_171);
nor U1547 (N_1547,In_201,In_276);
or U1548 (N_1548,In_325,In_692);
or U1549 (N_1549,In_451,In_425);
nand U1550 (N_1550,In_286,In_696);
xnor U1551 (N_1551,In_26,In_611);
and U1552 (N_1552,In_456,In_349);
and U1553 (N_1553,In_614,In_626);
or U1554 (N_1554,In_241,In_251);
xor U1555 (N_1555,In_241,In_32);
and U1556 (N_1556,In_20,In_186);
and U1557 (N_1557,In_735,In_283);
and U1558 (N_1558,In_515,In_459);
or U1559 (N_1559,In_663,In_442);
xor U1560 (N_1560,In_681,In_96);
xor U1561 (N_1561,In_43,In_623);
or U1562 (N_1562,In_150,In_533);
nor U1563 (N_1563,In_301,In_95);
xor U1564 (N_1564,In_374,In_194);
xnor U1565 (N_1565,In_319,In_531);
or U1566 (N_1566,In_287,In_713);
or U1567 (N_1567,In_424,In_151);
and U1568 (N_1568,In_699,In_733);
nand U1569 (N_1569,In_737,In_689);
nor U1570 (N_1570,In_184,In_612);
nand U1571 (N_1571,In_522,In_15);
nor U1572 (N_1572,In_729,In_150);
or U1573 (N_1573,In_392,In_717);
or U1574 (N_1574,In_728,In_470);
or U1575 (N_1575,In_595,In_126);
nor U1576 (N_1576,In_550,In_539);
nor U1577 (N_1577,In_272,In_192);
xor U1578 (N_1578,In_281,In_147);
nand U1579 (N_1579,In_675,In_16);
and U1580 (N_1580,In_45,In_491);
xnor U1581 (N_1581,In_379,In_207);
nand U1582 (N_1582,In_287,In_6);
nand U1583 (N_1583,In_678,In_69);
nor U1584 (N_1584,In_639,In_121);
nand U1585 (N_1585,In_244,In_717);
or U1586 (N_1586,In_590,In_524);
nand U1587 (N_1587,In_534,In_678);
or U1588 (N_1588,In_372,In_357);
and U1589 (N_1589,In_514,In_161);
or U1590 (N_1590,In_53,In_22);
xnor U1591 (N_1591,In_379,In_412);
or U1592 (N_1592,In_149,In_120);
or U1593 (N_1593,In_226,In_378);
nand U1594 (N_1594,In_554,In_13);
nor U1595 (N_1595,In_568,In_490);
nor U1596 (N_1596,In_614,In_74);
nand U1597 (N_1597,In_494,In_293);
or U1598 (N_1598,In_466,In_732);
xnor U1599 (N_1599,In_748,In_541);
or U1600 (N_1600,In_614,In_628);
and U1601 (N_1601,In_82,In_704);
nor U1602 (N_1602,In_689,In_431);
and U1603 (N_1603,In_3,In_259);
and U1604 (N_1604,In_689,In_79);
nor U1605 (N_1605,In_298,In_455);
and U1606 (N_1606,In_691,In_91);
xnor U1607 (N_1607,In_260,In_652);
nand U1608 (N_1608,In_107,In_462);
nor U1609 (N_1609,In_193,In_41);
and U1610 (N_1610,In_142,In_520);
and U1611 (N_1611,In_549,In_716);
nand U1612 (N_1612,In_183,In_688);
or U1613 (N_1613,In_501,In_210);
or U1614 (N_1614,In_292,In_147);
nand U1615 (N_1615,In_502,In_734);
nor U1616 (N_1616,In_505,In_663);
xnor U1617 (N_1617,In_215,In_698);
xor U1618 (N_1618,In_130,In_308);
or U1619 (N_1619,In_283,In_29);
or U1620 (N_1620,In_559,In_91);
or U1621 (N_1621,In_511,In_94);
xnor U1622 (N_1622,In_66,In_379);
or U1623 (N_1623,In_383,In_43);
nor U1624 (N_1624,In_128,In_120);
or U1625 (N_1625,In_14,In_135);
nor U1626 (N_1626,In_271,In_725);
nor U1627 (N_1627,In_427,In_392);
or U1628 (N_1628,In_497,In_710);
or U1629 (N_1629,In_86,In_144);
xnor U1630 (N_1630,In_360,In_735);
nor U1631 (N_1631,In_269,In_573);
xor U1632 (N_1632,In_391,In_610);
or U1633 (N_1633,In_646,In_460);
xnor U1634 (N_1634,In_565,In_467);
xnor U1635 (N_1635,In_457,In_527);
or U1636 (N_1636,In_454,In_127);
nand U1637 (N_1637,In_735,In_746);
or U1638 (N_1638,In_528,In_317);
nand U1639 (N_1639,In_448,In_279);
or U1640 (N_1640,In_525,In_363);
and U1641 (N_1641,In_68,In_673);
nor U1642 (N_1642,In_343,In_628);
nor U1643 (N_1643,In_75,In_42);
nor U1644 (N_1644,In_82,In_283);
or U1645 (N_1645,In_91,In_140);
nor U1646 (N_1646,In_34,In_168);
nor U1647 (N_1647,In_415,In_644);
or U1648 (N_1648,In_6,In_538);
xnor U1649 (N_1649,In_167,In_571);
and U1650 (N_1650,In_145,In_633);
or U1651 (N_1651,In_166,In_307);
nand U1652 (N_1652,In_130,In_618);
xor U1653 (N_1653,In_268,In_383);
xnor U1654 (N_1654,In_123,In_164);
and U1655 (N_1655,In_411,In_459);
nand U1656 (N_1656,In_400,In_99);
nand U1657 (N_1657,In_485,In_198);
or U1658 (N_1658,In_591,In_620);
xor U1659 (N_1659,In_265,In_332);
or U1660 (N_1660,In_458,In_224);
nand U1661 (N_1661,In_313,In_187);
nor U1662 (N_1662,In_22,In_411);
and U1663 (N_1663,In_30,In_716);
and U1664 (N_1664,In_135,In_306);
xnor U1665 (N_1665,In_39,In_14);
or U1666 (N_1666,In_625,In_480);
nor U1667 (N_1667,In_400,In_283);
and U1668 (N_1668,In_601,In_619);
nor U1669 (N_1669,In_599,In_505);
nand U1670 (N_1670,In_235,In_348);
xnor U1671 (N_1671,In_496,In_331);
or U1672 (N_1672,In_129,In_166);
or U1673 (N_1673,In_620,In_662);
nand U1674 (N_1674,In_197,In_598);
nor U1675 (N_1675,In_177,In_307);
nand U1676 (N_1676,In_367,In_368);
and U1677 (N_1677,In_488,In_539);
and U1678 (N_1678,In_205,In_610);
xor U1679 (N_1679,In_371,In_134);
nor U1680 (N_1680,In_108,In_281);
or U1681 (N_1681,In_333,In_175);
nor U1682 (N_1682,In_332,In_52);
or U1683 (N_1683,In_334,In_138);
xnor U1684 (N_1684,In_403,In_144);
xnor U1685 (N_1685,In_298,In_732);
xnor U1686 (N_1686,In_387,In_254);
nor U1687 (N_1687,In_123,In_114);
xor U1688 (N_1688,In_211,In_284);
and U1689 (N_1689,In_470,In_443);
or U1690 (N_1690,In_691,In_225);
xnor U1691 (N_1691,In_161,In_253);
and U1692 (N_1692,In_477,In_429);
nand U1693 (N_1693,In_193,In_513);
nand U1694 (N_1694,In_238,In_407);
xnor U1695 (N_1695,In_205,In_425);
or U1696 (N_1696,In_514,In_698);
nor U1697 (N_1697,In_316,In_570);
xor U1698 (N_1698,In_66,In_209);
nand U1699 (N_1699,In_592,In_102);
xor U1700 (N_1700,In_522,In_581);
nor U1701 (N_1701,In_675,In_499);
nand U1702 (N_1702,In_310,In_69);
and U1703 (N_1703,In_86,In_2);
or U1704 (N_1704,In_61,In_519);
and U1705 (N_1705,In_641,In_736);
or U1706 (N_1706,In_95,In_71);
nor U1707 (N_1707,In_438,In_141);
nor U1708 (N_1708,In_195,In_359);
nor U1709 (N_1709,In_470,In_645);
xor U1710 (N_1710,In_376,In_359);
xnor U1711 (N_1711,In_289,In_155);
or U1712 (N_1712,In_377,In_289);
or U1713 (N_1713,In_548,In_404);
and U1714 (N_1714,In_133,In_61);
or U1715 (N_1715,In_563,In_644);
nand U1716 (N_1716,In_678,In_652);
or U1717 (N_1717,In_695,In_119);
nand U1718 (N_1718,In_749,In_9);
nor U1719 (N_1719,In_250,In_44);
nand U1720 (N_1720,In_432,In_390);
nand U1721 (N_1721,In_161,In_382);
or U1722 (N_1722,In_314,In_243);
and U1723 (N_1723,In_79,In_166);
xnor U1724 (N_1724,In_396,In_252);
nand U1725 (N_1725,In_195,In_79);
nor U1726 (N_1726,In_696,In_502);
or U1727 (N_1727,In_156,In_277);
nand U1728 (N_1728,In_382,In_373);
xor U1729 (N_1729,In_733,In_134);
and U1730 (N_1730,In_38,In_617);
nor U1731 (N_1731,In_0,In_1);
or U1732 (N_1732,In_483,In_465);
and U1733 (N_1733,In_353,In_423);
xnor U1734 (N_1734,In_454,In_222);
nand U1735 (N_1735,In_152,In_465);
nand U1736 (N_1736,In_617,In_140);
xor U1737 (N_1737,In_385,In_654);
nand U1738 (N_1738,In_582,In_348);
nand U1739 (N_1739,In_309,In_272);
and U1740 (N_1740,In_50,In_168);
and U1741 (N_1741,In_102,In_443);
nand U1742 (N_1742,In_501,In_192);
nand U1743 (N_1743,In_116,In_240);
or U1744 (N_1744,In_544,In_730);
nand U1745 (N_1745,In_395,In_656);
nand U1746 (N_1746,In_278,In_635);
nor U1747 (N_1747,In_47,In_545);
or U1748 (N_1748,In_607,In_11);
xor U1749 (N_1749,In_31,In_528);
or U1750 (N_1750,In_489,In_485);
and U1751 (N_1751,In_504,In_344);
xnor U1752 (N_1752,In_221,In_56);
nand U1753 (N_1753,In_615,In_559);
and U1754 (N_1754,In_285,In_384);
nor U1755 (N_1755,In_694,In_70);
xor U1756 (N_1756,In_506,In_134);
xnor U1757 (N_1757,In_218,In_708);
or U1758 (N_1758,In_17,In_712);
nor U1759 (N_1759,In_169,In_347);
xnor U1760 (N_1760,In_511,In_105);
nand U1761 (N_1761,In_247,In_176);
or U1762 (N_1762,In_464,In_260);
xor U1763 (N_1763,In_443,In_103);
nor U1764 (N_1764,In_429,In_471);
or U1765 (N_1765,In_149,In_98);
xnor U1766 (N_1766,In_227,In_339);
xor U1767 (N_1767,In_531,In_404);
nor U1768 (N_1768,In_245,In_592);
nor U1769 (N_1769,In_345,In_400);
or U1770 (N_1770,In_204,In_235);
xor U1771 (N_1771,In_423,In_581);
and U1772 (N_1772,In_621,In_23);
or U1773 (N_1773,In_235,In_462);
nand U1774 (N_1774,In_576,In_562);
nor U1775 (N_1775,In_313,In_711);
and U1776 (N_1776,In_237,In_542);
nand U1777 (N_1777,In_312,In_406);
nand U1778 (N_1778,In_264,In_356);
nor U1779 (N_1779,In_696,In_454);
and U1780 (N_1780,In_441,In_541);
nor U1781 (N_1781,In_446,In_562);
nand U1782 (N_1782,In_622,In_597);
and U1783 (N_1783,In_587,In_112);
nand U1784 (N_1784,In_175,In_724);
and U1785 (N_1785,In_200,In_278);
and U1786 (N_1786,In_497,In_298);
nor U1787 (N_1787,In_130,In_89);
nor U1788 (N_1788,In_154,In_366);
xor U1789 (N_1789,In_293,In_538);
xor U1790 (N_1790,In_744,In_101);
or U1791 (N_1791,In_455,In_341);
or U1792 (N_1792,In_384,In_322);
nor U1793 (N_1793,In_641,In_26);
xnor U1794 (N_1794,In_117,In_196);
nand U1795 (N_1795,In_683,In_530);
and U1796 (N_1796,In_35,In_583);
nor U1797 (N_1797,In_276,In_424);
and U1798 (N_1798,In_717,In_197);
xor U1799 (N_1799,In_94,In_531);
or U1800 (N_1800,In_480,In_680);
xnor U1801 (N_1801,In_349,In_178);
and U1802 (N_1802,In_453,In_716);
nor U1803 (N_1803,In_189,In_388);
nor U1804 (N_1804,In_335,In_560);
nand U1805 (N_1805,In_432,In_44);
nand U1806 (N_1806,In_105,In_741);
nor U1807 (N_1807,In_304,In_385);
and U1808 (N_1808,In_246,In_231);
nand U1809 (N_1809,In_746,In_537);
or U1810 (N_1810,In_51,In_689);
nand U1811 (N_1811,In_564,In_126);
or U1812 (N_1812,In_499,In_412);
or U1813 (N_1813,In_481,In_261);
nor U1814 (N_1814,In_499,In_167);
nand U1815 (N_1815,In_543,In_299);
nand U1816 (N_1816,In_653,In_249);
and U1817 (N_1817,In_746,In_376);
xor U1818 (N_1818,In_226,In_28);
nor U1819 (N_1819,In_470,In_606);
xnor U1820 (N_1820,In_339,In_356);
and U1821 (N_1821,In_155,In_687);
nor U1822 (N_1822,In_424,In_650);
and U1823 (N_1823,In_166,In_397);
or U1824 (N_1824,In_301,In_512);
and U1825 (N_1825,In_244,In_180);
or U1826 (N_1826,In_599,In_669);
and U1827 (N_1827,In_72,In_177);
and U1828 (N_1828,In_311,In_97);
and U1829 (N_1829,In_499,In_617);
and U1830 (N_1830,In_245,In_397);
or U1831 (N_1831,In_421,In_369);
xor U1832 (N_1832,In_191,In_170);
and U1833 (N_1833,In_227,In_186);
nor U1834 (N_1834,In_641,In_678);
or U1835 (N_1835,In_117,In_592);
nand U1836 (N_1836,In_97,In_166);
or U1837 (N_1837,In_595,In_290);
xnor U1838 (N_1838,In_426,In_360);
nor U1839 (N_1839,In_412,In_524);
nor U1840 (N_1840,In_41,In_633);
nor U1841 (N_1841,In_505,In_164);
nand U1842 (N_1842,In_221,In_452);
xnor U1843 (N_1843,In_600,In_169);
or U1844 (N_1844,In_701,In_288);
or U1845 (N_1845,In_48,In_172);
or U1846 (N_1846,In_273,In_202);
and U1847 (N_1847,In_529,In_694);
nand U1848 (N_1848,In_418,In_133);
xnor U1849 (N_1849,In_496,In_155);
or U1850 (N_1850,In_276,In_520);
or U1851 (N_1851,In_195,In_482);
or U1852 (N_1852,In_125,In_719);
xor U1853 (N_1853,In_156,In_609);
or U1854 (N_1854,In_648,In_76);
nor U1855 (N_1855,In_43,In_122);
xnor U1856 (N_1856,In_735,In_522);
xnor U1857 (N_1857,In_563,In_667);
nand U1858 (N_1858,In_184,In_243);
nand U1859 (N_1859,In_241,In_447);
xor U1860 (N_1860,In_85,In_475);
nand U1861 (N_1861,In_666,In_301);
nand U1862 (N_1862,In_572,In_14);
or U1863 (N_1863,In_144,In_121);
or U1864 (N_1864,In_67,In_600);
nand U1865 (N_1865,In_652,In_610);
xnor U1866 (N_1866,In_628,In_61);
xor U1867 (N_1867,In_18,In_421);
nor U1868 (N_1868,In_30,In_579);
and U1869 (N_1869,In_138,In_748);
and U1870 (N_1870,In_74,In_109);
nor U1871 (N_1871,In_723,In_65);
xor U1872 (N_1872,In_186,In_207);
nor U1873 (N_1873,In_404,In_660);
nand U1874 (N_1874,In_744,In_689);
and U1875 (N_1875,In_155,In_364);
nand U1876 (N_1876,In_425,In_506);
nor U1877 (N_1877,In_582,In_45);
nor U1878 (N_1878,In_392,In_48);
or U1879 (N_1879,In_192,In_594);
and U1880 (N_1880,In_60,In_296);
and U1881 (N_1881,In_491,In_311);
xor U1882 (N_1882,In_667,In_721);
or U1883 (N_1883,In_636,In_363);
and U1884 (N_1884,In_343,In_183);
or U1885 (N_1885,In_469,In_500);
nor U1886 (N_1886,In_106,In_516);
xnor U1887 (N_1887,In_230,In_46);
nor U1888 (N_1888,In_321,In_149);
and U1889 (N_1889,In_707,In_311);
nand U1890 (N_1890,In_18,In_239);
and U1891 (N_1891,In_146,In_703);
nand U1892 (N_1892,In_191,In_102);
nor U1893 (N_1893,In_285,In_693);
nand U1894 (N_1894,In_665,In_28);
xnor U1895 (N_1895,In_284,In_364);
xor U1896 (N_1896,In_431,In_75);
nand U1897 (N_1897,In_664,In_633);
xor U1898 (N_1898,In_576,In_602);
xor U1899 (N_1899,In_744,In_706);
nor U1900 (N_1900,In_40,In_346);
xnor U1901 (N_1901,In_746,In_379);
or U1902 (N_1902,In_163,In_691);
nand U1903 (N_1903,In_391,In_361);
nor U1904 (N_1904,In_138,In_628);
xnor U1905 (N_1905,In_733,In_476);
nand U1906 (N_1906,In_231,In_516);
nor U1907 (N_1907,In_333,In_174);
or U1908 (N_1908,In_229,In_515);
or U1909 (N_1909,In_14,In_597);
nor U1910 (N_1910,In_687,In_336);
and U1911 (N_1911,In_302,In_151);
or U1912 (N_1912,In_396,In_100);
or U1913 (N_1913,In_595,In_324);
nand U1914 (N_1914,In_264,In_608);
nor U1915 (N_1915,In_582,In_505);
nor U1916 (N_1916,In_281,In_393);
nor U1917 (N_1917,In_542,In_218);
and U1918 (N_1918,In_653,In_31);
xnor U1919 (N_1919,In_708,In_655);
nor U1920 (N_1920,In_585,In_334);
xnor U1921 (N_1921,In_617,In_731);
nor U1922 (N_1922,In_306,In_669);
and U1923 (N_1923,In_483,In_639);
nor U1924 (N_1924,In_81,In_711);
nor U1925 (N_1925,In_79,In_174);
nor U1926 (N_1926,In_544,In_123);
or U1927 (N_1927,In_389,In_653);
nor U1928 (N_1928,In_413,In_710);
or U1929 (N_1929,In_713,In_269);
xnor U1930 (N_1930,In_747,In_136);
and U1931 (N_1931,In_517,In_304);
and U1932 (N_1932,In_145,In_324);
or U1933 (N_1933,In_725,In_687);
nor U1934 (N_1934,In_333,In_111);
and U1935 (N_1935,In_212,In_649);
xor U1936 (N_1936,In_504,In_429);
nor U1937 (N_1937,In_123,In_553);
xor U1938 (N_1938,In_365,In_2);
nor U1939 (N_1939,In_261,In_426);
xor U1940 (N_1940,In_137,In_207);
nand U1941 (N_1941,In_194,In_592);
or U1942 (N_1942,In_689,In_213);
or U1943 (N_1943,In_462,In_95);
and U1944 (N_1944,In_361,In_471);
nand U1945 (N_1945,In_589,In_351);
xnor U1946 (N_1946,In_265,In_160);
nand U1947 (N_1947,In_28,In_467);
nor U1948 (N_1948,In_191,In_316);
and U1949 (N_1949,In_718,In_599);
or U1950 (N_1950,In_329,In_53);
nand U1951 (N_1951,In_230,In_49);
nand U1952 (N_1952,In_449,In_249);
xnor U1953 (N_1953,In_603,In_690);
xnor U1954 (N_1954,In_385,In_484);
and U1955 (N_1955,In_15,In_607);
xor U1956 (N_1956,In_465,In_457);
xnor U1957 (N_1957,In_451,In_440);
nor U1958 (N_1958,In_261,In_590);
nand U1959 (N_1959,In_166,In_64);
nand U1960 (N_1960,In_346,In_250);
nand U1961 (N_1961,In_41,In_124);
or U1962 (N_1962,In_696,In_419);
nor U1963 (N_1963,In_186,In_194);
and U1964 (N_1964,In_668,In_592);
xnor U1965 (N_1965,In_369,In_540);
or U1966 (N_1966,In_377,In_310);
and U1967 (N_1967,In_487,In_171);
xnor U1968 (N_1968,In_72,In_709);
and U1969 (N_1969,In_341,In_429);
xor U1970 (N_1970,In_453,In_194);
nand U1971 (N_1971,In_344,In_140);
or U1972 (N_1972,In_293,In_177);
or U1973 (N_1973,In_150,In_175);
xor U1974 (N_1974,In_267,In_718);
nor U1975 (N_1975,In_141,In_67);
nand U1976 (N_1976,In_719,In_214);
nor U1977 (N_1977,In_385,In_231);
xnor U1978 (N_1978,In_461,In_605);
xnor U1979 (N_1979,In_177,In_536);
and U1980 (N_1980,In_207,In_68);
nor U1981 (N_1981,In_29,In_328);
or U1982 (N_1982,In_570,In_185);
or U1983 (N_1983,In_628,In_55);
and U1984 (N_1984,In_713,In_442);
or U1985 (N_1985,In_242,In_286);
nand U1986 (N_1986,In_98,In_301);
nand U1987 (N_1987,In_501,In_177);
xnor U1988 (N_1988,In_653,In_646);
nor U1989 (N_1989,In_600,In_562);
or U1990 (N_1990,In_73,In_590);
nand U1991 (N_1991,In_337,In_516);
xor U1992 (N_1992,In_177,In_49);
nand U1993 (N_1993,In_519,In_517);
or U1994 (N_1994,In_155,In_94);
nor U1995 (N_1995,In_416,In_88);
xor U1996 (N_1996,In_98,In_104);
xnor U1997 (N_1997,In_172,In_703);
and U1998 (N_1998,In_230,In_379);
or U1999 (N_1999,In_380,In_479);
nor U2000 (N_2000,In_3,In_292);
nor U2001 (N_2001,In_457,In_526);
and U2002 (N_2002,In_19,In_397);
nor U2003 (N_2003,In_154,In_594);
nand U2004 (N_2004,In_716,In_268);
xor U2005 (N_2005,In_700,In_514);
and U2006 (N_2006,In_62,In_288);
or U2007 (N_2007,In_673,In_719);
and U2008 (N_2008,In_390,In_191);
xor U2009 (N_2009,In_557,In_135);
xor U2010 (N_2010,In_34,In_180);
and U2011 (N_2011,In_678,In_671);
and U2012 (N_2012,In_563,In_735);
nand U2013 (N_2013,In_630,In_26);
xor U2014 (N_2014,In_250,In_538);
xor U2015 (N_2015,In_121,In_364);
or U2016 (N_2016,In_515,In_541);
nor U2017 (N_2017,In_692,In_736);
and U2018 (N_2018,In_316,In_146);
xnor U2019 (N_2019,In_28,In_90);
nor U2020 (N_2020,In_306,In_185);
and U2021 (N_2021,In_257,In_526);
nand U2022 (N_2022,In_542,In_235);
or U2023 (N_2023,In_374,In_22);
nor U2024 (N_2024,In_82,In_38);
and U2025 (N_2025,In_154,In_727);
nor U2026 (N_2026,In_92,In_157);
nor U2027 (N_2027,In_449,In_725);
or U2028 (N_2028,In_87,In_311);
nor U2029 (N_2029,In_630,In_4);
or U2030 (N_2030,In_624,In_13);
or U2031 (N_2031,In_106,In_319);
nand U2032 (N_2032,In_112,In_49);
nor U2033 (N_2033,In_731,In_4);
nor U2034 (N_2034,In_537,In_254);
or U2035 (N_2035,In_238,In_244);
xor U2036 (N_2036,In_485,In_229);
nand U2037 (N_2037,In_495,In_335);
and U2038 (N_2038,In_98,In_502);
or U2039 (N_2039,In_572,In_431);
or U2040 (N_2040,In_339,In_455);
xor U2041 (N_2041,In_218,In_445);
nor U2042 (N_2042,In_420,In_425);
xnor U2043 (N_2043,In_74,In_355);
and U2044 (N_2044,In_222,In_106);
xor U2045 (N_2045,In_468,In_682);
xor U2046 (N_2046,In_159,In_150);
xnor U2047 (N_2047,In_24,In_209);
nor U2048 (N_2048,In_422,In_215);
xor U2049 (N_2049,In_616,In_504);
and U2050 (N_2050,In_28,In_336);
nand U2051 (N_2051,In_191,In_743);
nor U2052 (N_2052,In_176,In_371);
and U2053 (N_2053,In_241,In_155);
and U2054 (N_2054,In_575,In_640);
or U2055 (N_2055,In_173,In_478);
and U2056 (N_2056,In_589,In_326);
xnor U2057 (N_2057,In_360,In_666);
nand U2058 (N_2058,In_273,In_540);
xnor U2059 (N_2059,In_633,In_564);
nor U2060 (N_2060,In_741,In_115);
or U2061 (N_2061,In_539,In_311);
or U2062 (N_2062,In_446,In_671);
nand U2063 (N_2063,In_506,In_309);
nor U2064 (N_2064,In_353,In_672);
nor U2065 (N_2065,In_490,In_312);
nor U2066 (N_2066,In_724,In_226);
nand U2067 (N_2067,In_608,In_649);
or U2068 (N_2068,In_378,In_420);
or U2069 (N_2069,In_518,In_292);
or U2070 (N_2070,In_219,In_571);
nand U2071 (N_2071,In_379,In_665);
and U2072 (N_2072,In_130,In_498);
nor U2073 (N_2073,In_397,In_474);
nor U2074 (N_2074,In_389,In_353);
or U2075 (N_2075,In_265,In_654);
nor U2076 (N_2076,In_116,In_92);
or U2077 (N_2077,In_570,In_128);
and U2078 (N_2078,In_134,In_741);
and U2079 (N_2079,In_679,In_695);
nor U2080 (N_2080,In_297,In_154);
nand U2081 (N_2081,In_683,In_38);
and U2082 (N_2082,In_722,In_323);
or U2083 (N_2083,In_711,In_597);
nand U2084 (N_2084,In_210,In_425);
nand U2085 (N_2085,In_542,In_372);
xor U2086 (N_2086,In_671,In_98);
nand U2087 (N_2087,In_298,In_312);
xor U2088 (N_2088,In_477,In_425);
xor U2089 (N_2089,In_481,In_228);
or U2090 (N_2090,In_599,In_497);
xor U2091 (N_2091,In_389,In_548);
nand U2092 (N_2092,In_243,In_635);
and U2093 (N_2093,In_410,In_370);
nand U2094 (N_2094,In_85,In_177);
or U2095 (N_2095,In_303,In_400);
nand U2096 (N_2096,In_469,In_735);
or U2097 (N_2097,In_58,In_621);
and U2098 (N_2098,In_352,In_299);
or U2099 (N_2099,In_440,In_306);
and U2100 (N_2100,In_91,In_557);
and U2101 (N_2101,In_704,In_696);
and U2102 (N_2102,In_704,In_189);
nand U2103 (N_2103,In_136,In_607);
or U2104 (N_2104,In_69,In_453);
or U2105 (N_2105,In_474,In_168);
nand U2106 (N_2106,In_704,In_645);
and U2107 (N_2107,In_377,In_679);
nor U2108 (N_2108,In_66,In_10);
nor U2109 (N_2109,In_519,In_360);
and U2110 (N_2110,In_735,In_729);
nor U2111 (N_2111,In_418,In_689);
xor U2112 (N_2112,In_409,In_283);
or U2113 (N_2113,In_144,In_90);
xnor U2114 (N_2114,In_402,In_21);
nand U2115 (N_2115,In_569,In_472);
nor U2116 (N_2116,In_174,In_304);
and U2117 (N_2117,In_597,In_427);
xnor U2118 (N_2118,In_420,In_231);
xor U2119 (N_2119,In_361,In_100);
nand U2120 (N_2120,In_635,In_708);
or U2121 (N_2121,In_424,In_273);
and U2122 (N_2122,In_593,In_464);
and U2123 (N_2123,In_155,In_315);
nor U2124 (N_2124,In_106,In_199);
nand U2125 (N_2125,In_345,In_117);
nor U2126 (N_2126,In_558,In_27);
nor U2127 (N_2127,In_558,In_572);
or U2128 (N_2128,In_34,In_130);
and U2129 (N_2129,In_524,In_629);
nor U2130 (N_2130,In_748,In_707);
and U2131 (N_2131,In_377,In_283);
nand U2132 (N_2132,In_20,In_434);
xnor U2133 (N_2133,In_610,In_580);
nand U2134 (N_2134,In_722,In_511);
nand U2135 (N_2135,In_525,In_100);
nand U2136 (N_2136,In_573,In_416);
or U2137 (N_2137,In_359,In_600);
nand U2138 (N_2138,In_649,In_467);
xnor U2139 (N_2139,In_577,In_549);
or U2140 (N_2140,In_181,In_464);
nor U2141 (N_2141,In_112,In_480);
nand U2142 (N_2142,In_539,In_588);
and U2143 (N_2143,In_143,In_298);
nor U2144 (N_2144,In_268,In_159);
or U2145 (N_2145,In_647,In_444);
nand U2146 (N_2146,In_174,In_226);
xnor U2147 (N_2147,In_135,In_349);
and U2148 (N_2148,In_652,In_700);
and U2149 (N_2149,In_84,In_707);
nand U2150 (N_2150,In_617,In_427);
nand U2151 (N_2151,In_106,In_340);
nor U2152 (N_2152,In_709,In_674);
or U2153 (N_2153,In_148,In_498);
xnor U2154 (N_2154,In_699,In_670);
or U2155 (N_2155,In_425,In_56);
nand U2156 (N_2156,In_108,In_346);
nand U2157 (N_2157,In_187,In_654);
or U2158 (N_2158,In_509,In_686);
xnor U2159 (N_2159,In_194,In_39);
and U2160 (N_2160,In_121,In_478);
xnor U2161 (N_2161,In_152,In_354);
xor U2162 (N_2162,In_349,In_652);
or U2163 (N_2163,In_93,In_108);
nand U2164 (N_2164,In_359,In_575);
or U2165 (N_2165,In_118,In_379);
or U2166 (N_2166,In_546,In_706);
nor U2167 (N_2167,In_295,In_46);
and U2168 (N_2168,In_204,In_692);
and U2169 (N_2169,In_177,In_655);
nor U2170 (N_2170,In_63,In_289);
nor U2171 (N_2171,In_285,In_483);
and U2172 (N_2172,In_82,In_33);
nand U2173 (N_2173,In_431,In_671);
or U2174 (N_2174,In_618,In_66);
or U2175 (N_2175,In_480,In_213);
and U2176 (N_2176,In_54,In_627);
xor U2177 (N_2177,In_66,In_437);
xnor U2178 (N_2178,In_331,In_391);
nor U2179 (N_2179,In_293,In_134);
nor U2180 (N_2180,In_214,In_288);
or U2181 (N_2181,In_307,In_35);
and U2182 (N_2182,In_174,In_9);
nor U2183 (N_2183,In_247,In_616);
or U2184 (N_2184,In_596,In_738);
nor U2185 (N_2185,In_152,In_73);
nor U2186 (N_2186,In_117,In_607);
nand U2187 (N_2187,In_364,In_521);
xnor U2188 (N_2188,In_465,In_598);
xor U2189 (N_2189,In_50,In_86);
nor U2190 (N_2190,In_733,In_680);
and U2191 (N_2191,In_176,In_305);
or U2192 (N_2192,In_741,In_314);
nand U2193 (N_2193,In_556,In_532);
or U2194 (N_2194,In_164,In_206);
or U2195 (N_2195,In_201,In_125);
nor U2196 (N_2196,In_47,In_742);
and U2197 (N_2197,In_288,In_145);
xor U2198 (N_2198,In_326,In_574);
and U2199 (N_2199,In_424,In_419);
nand U2200 (N_2200,In_557,In_642);
nor U2201 (N_2201,In_303,In_520);
nand U2202 (N_2202,In_112,In_118);
xnor U2203 (N_2203,In_443,In_723);
and U2204 (N_2204,In_253,In_335);
and U2205 (N_2205,In_281,In_23);
nand U2206 (N_2206,In_546,In_196);
nor U2207 (N_2207,In_691,In_255);
or U2208 (N_2208,In_21,In_293);
nand U2209 (N_2209,In_179,In_254);
nor U2210 (N_2210,In_555,In_501);
nor U2211 (N_2211,In_568,In_168);
xnor U2212 (N_2212,In_561,In_6);
nand U2213 (N_2213,In_378,In_11);
nor U2214 (N_2214,In_544,In_616);
or U2215 (N_2215,In_192,In_140);
xnor U2216 (N_2216,In_702,In_112);
and U2217 (N_2217,In_35,In_30);
and U2218 (N_2218,In_547,In_297);
nor U2219 (N_2219,In_32,In_448);
or U2220 (N_2220,In_327,In_691);
and U2221 (N_2221,In_644,In_320);
and U2222 (N_2222,In_687,In_618);
nand U2223 (N_2223,In_589,In_297);
and U2224 (N_2224,In_565,In_164);
nand U2225 (N_2225,In_713,In_53);
or U2226 (N_2226,In_197,In_736);
nand U2227 (N_2227,In_254,In_446);
or U2228 (N_2228,In_398,In_530);
or U2229 (N_2229,In_68,In_615);
xor U2230 (N_2230,In_341,In_49);
xor U2231 (N_2231,In_662,In_491);
xor U2232 (N_2232,In_656,In_217);
or U2233 (N_2233,In_449,In_566);
nand U2234 (N_2234,In_673,In_609);
nand U2235 (N_2235,In_694,In_262);
or U2236 (N_2236,In_723,In_737);
and U2237 (N_2237,In_621,In_47);
or U2238 (N_2238,In_248,In_550);
and U2239 (N_2239,In_334,In_433);
xnor U2240 (N_2240,In_496,In_168);
nor U2241 (N_2241,In_695,In_195);
and U2242 (N_2242,In_392,In_221);
nor U2243 (N_2243,In_562,In_111);
nor U2244 (N_2244,In_481,In_476);
xnor U2245 (N_2245,In_530,In_112);
nor U2246 (N_2246,In_69,In_251);
nor U2247 (N_2247,In_637,In_568);
nor U2248 (N_2248,In_501,In_462);
xor U2249 (N_2249,In_732,In_302);
xor U2250 (N_2250,In_339,In_128);
xor U2251 (N_2251,In_71,In_193);
or U2252 (N_2252,In_533,In_506);
and U2253 (N_2253,In_540,In_456);
and U2254 (N_2254,In_347,In_684);
nor U2255 (N_2255,In_660,In_399);
or U2256 (N_2256,In_331,In_681);
or U2257 (N_2257,In_661,In_689);
nor U2258 (N_2258,In_558,In_36);
nand U2259 (N_2259,In_411,In_233);
nor U2260 (N_2260,In_92,In_742);
nand U2261 (N_2261,In_256,In_457);
nand U2262 (N_2262,In_724,In_257);
nand U2263 (N_2263,In_241,In_233);
or U2264 (N_2264,In_617,In_570);
xor U2265 (N_2265,In_473,In_259);
nor U2266 (N_2266,In_642,In_604);
nor U2267 (N_2267,In_70,In_0);
xor U2268 (N_2268,In_194,In_708);
nor U2269 (N_2269,In_541,In_183);
xnor U2270 (N_2270,In_45,In_156);
nand U2271 (N_2271,In_727,In_52);
or U2272 (N_2272,In_178,In_176);
and U2273 (N_2273,In_721,In_358);
and U2274 (N_2274,In_485,In_14);
nor U2275 (N_2275,In_615,In_728);
nor U2276 (N_2276,In_41,In_599);
nor U2277 (N_2277,In_164,In_2);
and U2278 (N_2278,In_683,In_171);
or U2279 (N_2279,In_314,In_66);
xor U2280 (N_2280,In_677,In_470);
nor U2281 (N_2281,In_676,In_582);
or U2282 (N_2282,In_747,In_538);
nand U2283 (N_2283,In_437,In_349);
nand U2284 (N_2284,In_474,In_429);
or U2285 (N_2285,In_675,In_75);
nand U2286 (N_2286,In_304,In_659);
and U2287 (N_2287,In_57,In_209);
nor U2288 (N_2288,In_464,In_259);
and U2289 (N_2289,In_462,In_115);
nor U2290 (N_2290,In_176,In_186);
nand U2291 (N_2291,In_472,In_664);
and U2292 (N_2292,In_129,In_75);
nand U2293 (N_2293,In_460,In_741);
or U2294 (N_2294,In_58,In_494);
and U2295 (N_2295,In_231,In_296);
or U2296 (N_2296,In_508,In_187);
xnor U2297 (N_2297,In_699,In_370);
and U2298 (N_2298,In_490,In_324);
nand U2299 (N_2299,In_197,In_32);
nor U2300 (N_2300,In_191,In_422);
nand U2301 (N_2301,In_362,In_228);
and U2302 (N_2302,In_277,In_310);
xnor U2303 (N_2303,In_607,In_169);
xor U2304 (N_2304,In_465,In_398);
and U2305 (N_2305,In_329,In_338);
nor U2306 (N_2306,In_379,In_132);
xor U2307 (N_2307,In_466,In_273);
and U2308 (N_2308,In_398,In_676);
xor U2309 (N_2309,In_280,In_109);
nand U2310 (N_2310,In_242,In_245);
xor U2311 (N_2311,In_38,In_461);
xnor U2312 (N_2312,In_453,In_176);
nor U2313 (N_2313,In_525,In_714);
and U2314 (N_2314,In_557,In_583);
or U2315 (N_2315,In_192,In_622);
nand U2316 (N_2316,In_628,In_464);
nor U2317 (N_2317,In_656,In_723);
nor U2318 (N_2318,In_545,In_121);
xnor U2319 (N_2319,In_708,In_175);
or U2320 (N_2320,In_55,In_200);
or U2321 (N_2321,In_682,In_294);
and U2322 (N_2322,In_480,In_666);
nand U2323 (N_2323,In_104,In_188);
nand U2324 (N_2324,In_207,In_524);
nand U2325 (N_2325,In_721,In_711);
nand U2326 (N_2326,In_710,In_681);
nor U2327 (N_2327,In_658,In_434);
xnor U2328 (N_2328,In_745,In_391);
or U2329 (N_2329,In_610,In_0);
and U2330 (N_2330,In_241,In_503);
or U2331 (N_2331,In_325,In_189);
nand U2332 (N_2332,In_732,In_603);
nand U2333 (N_2333,In_608,In_459);
or U2334 (N_2334,In_309,In_370);
or U2335 (N_2335,In_523,In_581);
or U2336 (N_2336,In_601,In_51);
or U2337 (N_2337,In_491,In_560);
and U2338 (N_2338,In_343,In_134);
or U2339 (N_2339,In_459,In_501);
and U2340 (N_2340,In_690,In_676);
and U2341 (N_2341,In_105,In_397);
xor U2342 (N_2342,In_463,In_453);
xor U2343 (N_2343,In_83,In_431);
and U2344 (N_2344,In_301,In_444);
xnor U2345 (N_2345,In_518,In_256);
nor U2346 (N_2346,In_462,In_154);
and U2347 (N_2347,In_489,In_578);
and U2348 (N_2348,In_366,In_3);
and U2349 (N_2349,In_266,In_446);
xnor U2350 (N_2350,In_416,In_683);
and U2351 (N_2351,In_122,In_583);
xnor U2352 (N_2352,In_361,In_105);
and U2353 (N_2353,In_227,In_393);
or U2354 (N_2354,In_137,In_576);
or U2355 (N_2355,In_734,In_642);
xor U2356 (N_2356,In_100,In_688);
or U2357 (N_2357,In_79,In_101);
or U2358 (N_2358,In_134,In_179);
nor U2359 (N_2359,In_616,In_696);
xnor U2360 (N_2360,In_621,In_330);
nor U2361 (N_2361,In_292,In_717);
xor U2362 (N_2362,In_736,In_526);
nand U2363 (N_2363,In_273,In_251);
nor U2364 (N_2364,In_89,In_746);
and U2365 (N_2365,In_380,In_246);
or U2366 (N_2366,In_155,In_623);
xnor U2367 (N_2367,In_263,In_310);
xor U2368 (N_2368,In_498,In_549);
nand U2369 (N_2369,In_367,In_80);
and U2370 (N_2370,In_689,In_297);
and U2371 (N_2371,In_390,In_195);
and U2372 (N_2372,In_149,In_527);
xnor U2373 (N_2373,In_185,In_658);
and U2374 (N_2374,In_391,In_121);
nand U2375 (N_2375,In_425,In_35);
nor U2376 (N_2376,In_387,In_693);
and U2377 (N_2377,In_680,In_124);
and U2378 (N_2378,In_419,In_71);
nor U2379 (N_2379,In_336,In_272);
nand U2380 (N_2380,In_77,In_164);
or U2381 (N_2381,In_692,In_598);
nand U2382 (N_2382,In_415,In_494);
or U2383 (N_2383,In_200,In_443);
and U2384 (N_2384,In_545,In_109);
or U2385 (N_2385,In_467,In_18);
and U2386 (N_2386,In_739,In_504);
nand U2387 (N_2387,In_432,In_367);
nand U2388 (N_2388,In_264,In_649);
xor U2389 (N_2389,In_178,In_378);
nand U2390 (N_2390,In_107,In_518);
and U2391 (N_2391,In_746,In_14);
nor U2392 (N_2392,In_32,In_494);
and U2393 (N_2393,In_702,In_447);
and U2394 (N_2394,In_463,In_111);
nand U2395 (N_2395,In_688,In_130);
nor U2396 (N_2396,In_482,In_652);
or U2397 (N_2397,In_380,In_319);
and U2398 (N_2398,In_278,In_335);
xnor U2399 (N_2399,In_747,In_692);
nand U2400 (N_2400,In_550,In_565);
or U2401 (N_2401,In_385,In_363);
and U2402 (N_2402,In_409,In_102);
or U2403 (N_2403,In_238,In_418);
or U2404 (N_2404,In_43,In_542);
xor U2405 (N_2405,In_63,In_181);
xor U2406 (N_2406,In_735,In_378);
nand U2407 (N_2407,In_177,In_650);
or U2408 (N_2408,In_708,In_613);
nor U2409 (N_2409,In_681,In_371);
or U2410 (N_2410,In_749,In_524);
nand U2411 (N_2411,In_383,In_282);
or U2412 (N_2412,In_9,In_327);
and U2413 (N_2413,In_242,In_687);
nand U2414 (N_2414,In_485,In_618);
and U2415 (N_2415,In_434,In_668);
xor U2416 (N_2416,In_490,In_542);
nor U2417 (N_2417,In_580,In_481);
and U2418 (N_2418,In_272,In_333);
nor U2419 (N_2419,In_579,In_134);
xnor U2420 (N_2420,In_348,In_387);
and U2421 (N_2421,In_214,In_413);
nand U2422 (N_2422,In_520,In_358);
and U2423 (N_2423,In_499,In_284);
and U2424 (N_2424,In_172,In_493);
xnor U2425 (N_2425,In_365,In_113);
nor U2426 (N_2426,In_241,In_318);
xnor U2427 (N_2427,In_627,In_225);
xnor U2428 (N_2428,In_155,In_716);
nand U2429 (N_2429,In_68,In_688);
and U2430 (N_2430,In_486,In_384);
nand U2431 (N_2431,In_217,In_672);
nor U2432 (N_2432,In_66,In_459);
or U2433 (N_2433,In_741,In_716);
xnor U2434 (N_2434,In_563,In_597);
or U2435 (N_2435,In_493,In_672);
or U2436 (N_2436,In_10,In_110);
or U2437 (N_2437,In_307,In_424);
xor U2438 (N_2438,In_35,In_296);
nor U2439 (N_2439,In_460,In_287);
or U2440 (N_2440,In_624,In_627);
nand U2441 (N_2441,In_309,In_535);
nor U2442 (N_2442,In_466,In_460);
nor U2443 (N_2443,In_264,In_403);
xnor U2444 (N_2444,In_734,In_40);
nand U2445 (N_2445,In_741,In_707);
xor U2446 (N_2446,In_276,In_604);
or U2447 (N_2447,In_384,In_635);
and U2448 (N_2448,In_397,In_529);
nor U2449 (N_2449,In_479,In_87);
and U2450 (N_2450,In_674,In_184);
or U2451 (N_2451,In_346,In_105);
and U2452 (N_2452,In_192,In_508);
or U2453 (N_2453,In_408,In_410);
nor U2454 (N_2454,In_162,In_586);
and U2455 (N_2455,In_474,In_457);
nand U2456 (N_2456,In_481,In_578);
nand U2457 (N_2457,In_461,In_527);
or U2458 (N_2458,In_708,In_712);
nor U2459 (N_2459,In_89,In_254);
nor U2460 (N_2460,In_309,In_445);
nand U2461 (N_2461,In_54,In_264);
or U2462 (N_2462,In_301,In_297);
and U2463 (N_2463,In_363,In_120);
xnor U2464 (N_2464,In_373,In_455);
nor U2465 (N_2465,In_490,In_82);
xor U2466 (N_2466,In_418,In_688);
or U2467 (N_2467,In_364,In_316);
nor U2468 (N_2468,In_327,In_377);
nand U2469 (N_2469,In_629,In_681);
nor U2470 (N_2470,In_287,In_318);
nand U2471 (N_2471,In_536,In_158);
nor U2472 (N_2472,In_659,In_417);
nor U2473 (N_2473,In_73,In_540);
or U2474 (N_2474,In_144,In_426);
xor U2475 (N_2475,In_59,In_263);
xor U2476 (N_2476,In_364,In_280);
nand U2477 (N_2477,In_285,In_691);
and U2478 (N_2478,In_35,In_246);
and U2479 (N_2479,In_50,In_266);
and U2480 (N_2480,In_535,In_114);
and U2481 (N_2481,In_41,In_432);
and U2482 (N_2482,In_724,In_285);
nor U2483 (N_2483,In_721,In_502);
nor U2484 (N_2484,In_148,In_394);
and U2485 (N_2485,In_447,In_743);
xnor U2486 (N_2486,In_390,In_49);
xnor U2487 (N_2487,In_681,In_124);
xnor U2488 (N_2488,In_280,In_600);
or U2489 (N_2489,In_113,In_112);
xor U2490 (N_2490,In_572,In_557);
xnor U2491 (N_2491,In_66,In_165);
nand U2492 (N_2492,In_24,In_425);
xnor U2493 (N_2493,In_692,In_253);
and U2494 (N_2494,In_591,In_554);
and U2495 (N_2495,In_368,In_749);
or U2496 (N_2496,In_460,In_325);
nand U2497 (N_2497,In_540,In_1);
nand U2498 (N_2498,In_112,In_294);
and U2499 (N_2499,In_421,In_194);
and U2500 (N_2500,N_776,N_480);
nor U2501 (N_2501,N_1910,N_546);
nand U2502 (N_2502,N_1631,N_453);
nor U2503 (N_2503,N_1502,N_726);
xor U2504 (N_2504,N_1990,N_1758);
or U2505 (N_2505,N_331,N_1794);
xor U2506 (N_2506,N_1720,N_937);
nor U2507 (N_2507,N_2395,N_323);
nand U2508 (N_2508,N_243,N_1243);
and U2509 (N_2509,N_2013,N_255);
and U2510 (N_2510,N_1163,N_1275);
xor U2511 (N_2511,N_466,N_2198);
nand U2512 (N_2512,N_2300,N_1467);
or U2513 (N_2513,N_2233,N_229);
and U2514 (N_2514,N_2025,N_2019);
xor U2515 (N_2515,N_1276,N_858);
or U2516 (N_2516,N_1301,N_2235);
and U2517 (N_2517,N_1581,N_2325);
nand U2518 (N_2518,N_1180,N_215);
nand U2519 (N_2519,N_586,N_1297);
and U2520 (N_2520,N_1368,N_345);
nand U2521 (N_2521,N_905,N_2211);
or U2522 (N_2522,N_2255,N_147);
or U2523 (N_2523,N_1436,N_1088);
or U2524 (N_2524,N_1189,N_1204);
or U2525 (N_2525,N_1733,N_1448);
xnor U2526 (N_2526,N_661,N_2127);
xnor U2527 (N_2527,N_1353,N_1024);
or U2528 (N_2528,N_1125,N_1688);
and U2529 (N_2529,N_2212,N_1772);
nand U2530 (N_2530,N_240,N_923);
nor U2531 (N_2531,N_188,N_2075);
and U2532 (N_2532,N_512,N_1615);
xor U2533 (N_2533,N_575,N_556);
nor U2534 (N_2534,N_1273,N_1317);
or U2535 (N_2535,N_1337,N_1768);
xor U2536 (N_2536,N_1068,N_1672);
xnor U2537 (N_2537,N_1922,N_48);
and U2538 (N_2538,N_1637,N_1251);
and U2539 (N_2539,N_543,N_1349);
and U2540 (N_2540,N_2204,N_72);
nor U2541 (N_2541,N_414,N_2236);
nor U2542 (N_2542,N_2432,N_2320);
nand U2543 (N_2543,N_1008,N_872);
and U2544 (N_2544,N_561,N_1139);
or U2545 (N_2545,N_675,N_1712);
nand U2546 (N_2546,N_1030,N_1583);
and U2547 (N_2547,N_1623,N_141);
nor U2548 (N_2548,N_416,N_1962);
and U2549 (N_2549,N_2216,N_452);
nor U2550 (N_2550,N_1646,N_1263);
and U2551 (N_2551,N_226,N_807);
nor U2552 (N_2552,N_230,N_84);
xnor U2553 (N_2553,N_1878,N_975);
nor U2554 (N_2554,N_442,N_2433);
or U2555 (N_2555,N_588,N_2452);
nor U2556 (N_2556,N_1966,N_2413);
nand U2557 (N_2557,N_1240,N_327);
and U2558 (N_2558,N_601,N_438);
and U2559 (N_2559,N_131,N_1464);
and U2560 (N_2560,N_813,N_2172);
nor U2561 (N_2561,N_2188,N_2499);
or U2562 (N_2562,N_2478,N_1557);
nor U2563 (N_2563,N_1985,N_821);
nor U2564 (N_2564,N_1744,N_689);
or U2565 (N_2565,N_105,N_2047);
nand U2566 (N_2566,N_1134,N_739);
nand U2567 (N_2567,N_790,N_885);
xnor U2568 (N_2568,N_894,N_307);
nor U2569 (N_2569,N_1509,N_1282);
and U2570 (N_2570,N_1094,N_1763);
xor U2571 (N_2571,N_705,N_1736);
nand U2572 (N_2572,N_1657,N_338);
nor U2573 (N_2573,N_1304,N_2438);
or U2574 (N_2574,N_1359,N_1288);
or U2575 (N_2575,N_1913,N_985);
nor U2576 (N_2576,N_2455,N_391);
and U2577 (N_2577,N_190,N_2283);
or U2578 (N_2578,N_2383,N_1049);
nand U2579 (N_2579,N_1724,N_98);
nor U2580 (N_2580,N_1812,N_1063);
nor U2581 (N_2581,N_679,N_1735);
nor U2582 (N_2582,N_922,N_1746);
and U2583 (N_2583,N_1221,N_195);
nor U2584 (N_2584,N_1328,N_745);
or U2585 (N_2585,N_36,N_2372);
xnor U2586 (N_2586,N_403,N_2250);
and U2587 (N_2587,N_1466,N_201);
xnor U2588 (N_2588,N_101,N_1549);
or U2589 (N_2589,N_2289,N_92);
xnor U2590 (N_2590,N_429,N_236);
nand U2591 (N_2591,N_55,N_1460);
xnor U2592 (N_2592,N_1222,N_664);
and U2593 (N_2593,N_2482,N_1983);
nor U2594 (N_2594,N_1331,N_1479);
or U2595 (N_2595,N_1806,N_6);
xor U2596 (N_2596,N_369,N_2051);
nand U2597 (N_2597,N_669,N_2392);
nand U2598 (N_2598,N_1148,N_748);
nor U2599 (N_2599,N_1504,N_305);
nor U2600 (N_2600,N_2215,N_781);
or U2601 (N_2601,N_1601,N_2001);
nand U2602 (N_2602,N_1056,N_2314);
and U2603 (N_2603,N_1072,N_390);
or U2604 (N_2604,N_2374,N_751);
nor U2605 (N_2605,N_854,N_2268);
xor U2606 (N_2606,N_1086,N_2224);
nor U2607 (N_2607,N_1099,N_275);
xnor U2608 (N_2608,N_491,N_1930);
nor U2609 (N_2609,N_370,N_701);
and U2610 (N_2610,N_1028,N_1032);
nor U2611 (N_2611,N_1462,N_1151);
xnor U2612 (N_2612,N_421,N_1386);
nor U2613 (N_2613,N_1062,N_163);
nor U2614 (N_2614,N_1608,N_1058);
nor U2615 (N_2615,N_1394,N_1627);
xor U2616 (N_2616,N_633,N_1868);
nor U2617 (N_2617,N_335,N_2107);
nor U2618 (N_2618,N_1731,N_2201);
and U2619 (N_2619,N_826,N_1803);
and U2620 (N_2620,N_1843,N_1571);
or U2621 (N_2621,N_511,N_649);
xor U2622 (N_2622,N_2386,N_548);
nor U2623 (N_2623,N_613,N_2185);
or U2624 (N_2624,N_1400,N_2114);
and U2625 (N_2625,N_1122,N_2409);
and U2626 (N_2626,N_60,N_1891);
nand U2627 (N_2627,N_2281,N_2072);
and U2628 (N_2628,N_1461,N_804);
xor U2629 (N_2629,N_1272,N_1184);
and U2630 (N_2630,N_1604,N_259);
nor U2631 (N_2631,N_1059,N_866);
nand U2632 (N_2632,N_1664,N_1997);
nand U2633 (N_2633,N_2387,N_1654);
or U2634 (N_2634,N_474,N_2396);
or U2635 (N_2635,N_2479,N_1773);
and U2636 (N_2636,N_2108,N_1612);
xor U2637 (N_2637,N_541,N_2113);
nor U2638 (N_2638,N_1360,N_1920);
and U2639 (N_2639,N_2117,N_2184);
xor U2640 (N_2640,N_612,N_1991);
nor U2641 (N_2641,N_2306,N_949);
or U2642 (N_2642,N_2166,N_747);
xor U2643 (N_2643,N_1884,N_1454);
and U2644 (N_2644,N_1551,N_520);
xnor U2645 (N_2645,N_1012,N_944);
xor U2646 (N_2646,N_1090,N_470);
nor U2647 (N_2647,N_607,N_926);
nand U2648 (N_2648,N_1591,N_2103);
xnor U2649 (N_2649,N_2470,N_320);
nand U2650 (N_2650,N_1231,N_684);
and U2651 (N_2651,N_992,N_1338);
and U2652 (N_2652,N_531,N_547);
or U2653 (N_2653,N_214,N_2243);
nand U2654 (N_2654,N_1484,N_674);
or U2655 (N_2655,N_1396,N_456);
nand U2656 (N_2656,N_969,N_2456);
or U2657 (N_2657,N_931,N_447);
nor U2658 (N_2658,N_2459,N_1630);
nor U2659 (N_2659,N_908,N_1605);
xnor U2660 (N_2660,N_899,N_329);
or U2661 (N_2661,N_1468,N_843);
and U2662 (N_2662,N_1432,N_979);
xnor U2663 (N_2663,N_2170,N_2408);
xnor U2664 (N_2664,N_1948,N_1410);
and U2665 (N_2665,N_344,N_2178);
nor U2666 (N_2666,N_1677,N_2488);
nor U2667 (N_2667,N_404,N_1770);
nor U2668 (N_2668,N_1314,N_1934);
nor U2669 (N_2669,N_2335,N_2089);
or U2670 (N_2670,N_410,N_904);
and U2671 (N_2671,N_1413,N_1707);
and U2672 (N_2672,N_1723,N_964);
xnor U2673 (N_2673,N_1682,N_2315);
and U2674 (N_2674,N_2393,N_623);
or U2675 (N_2675,N_1442,N_206);
or U2676 (N_2676,N_93,N_1170);
or U2677 (N_2677,N_1738,N_1405);
and U2678 (N_2678,N_755,N_1636);
xnor U2679 (N_2679,N_2385,N_2147);
nor U2680 (N_2680,N_341,N_642);
and U2681 (N_2681,N_870,N_95);
and U2682 (N_2682,N_280,N_2071);
nand U2683 (N_2683,N_1004,N_337);
or U2684 (N_2684,N_1530,N_203);
nor U2685 (N_2685,N_662,N_1164);
nor U2686 (N_2686,N_768,N_1117);
or U2687 (N_2687,N_100,N_2168);
and U2688 (N_2688,N_510,N_2077);
xnor U2689 (N_2689,N_1310,N_994);
and U2690 (N_2690,N_673,N_657);
or U2691 (N_2691,N_1401,N_2378);
nor U2692 (N_2692,N_875,N_2181);
nor U2693 (N_2693,N_2132,N_1217);
nand U2694 (N_2694,N_890,N_2274);
xnor U2695 (N_2695,N_2021,N_2157);
nand U2696 (N_2696,N_1833,N_782);
or U2697 (N_2697,N_914,N_1190);
xor U2698 (N_2698,N_539,N_1980);
xnor U2699 (N_2699,N_1575,N_1266);
or U2700 (N_2700,N_1269,N_1777);
or U2701 (N_2701,N_2015,N_1346);
xnor U2702 (N_2702,N_1989,N_2231);
nand U2703 (N_2703,N_974,N_1416);
nor U2704 (N_2704,N_1584,N_2337);
xor U2705 (N_2705,N_606,N_1617);
or U2706 (N_2706,N_2050,N_2263);
nor U2707 (N_2707,N_250,N_1907);
nor U2708 (N_2708,N_1898,N_2126);
nand U2709 (N_2709,N_1610,N_256);
xnor U2710 (N_2710,N_1241,N_2327);
xor U2711 (N_2711,N_2405,N_1185);
nor U2712 (N_2712,N_650,N_1728);
nand U2713 (N_2713,N_721,N_1261);
nand U2714 (N_2714,N_1455,N_655);
or U2715 (N_2715,N_1207,N_1371);
xor U2716 (N_2716,N_2056,N_326);
xnor U2717 (N_2717,N_151,N_115);
nand U2718 (N_2718,N_433,N_574);
nor U2719 (N_2719,N_682,N_1671);
nand U2720 (N_2720,N_296,N_698);
nor U2721 (N_2721,N_621,N_257);
or U2722 (N_2722,N_2331,N_486);
xnor U2723 (N_2723,N_498,N_232);
xor U2724 (N_2724,N_1205,N_902);
and U2725 (N_2725,N_1113,N_1043);
nand U2726 (N_2726,N_1474,N_882);
xor U2727 (N_2727,N_2343,N_1246);
or U2728 (N_2728,N_2276,N_17);
and U2729 (N_2729,N_1296,N_2298);
or U2730 (N_2730,N_774,N_114);
or U2731 (N_2731,N_1018,N_597);
xnor U2732 (N_2732,N_819,N_1312);
xor U2733 (N_2733,N_1558,N_1813);
xnor U2734 (N_2734,N_1285,N_1831);
nor U2735 (N_2735,N_2318,N_2038);
nand U2736 (N_2736,N_224,N_1109);
xnor U2737 (N_2737,N_604,N_306);
or U2738 (N_2738,N_1755,N_1093);
and U2739 (N_2739,N_2205,N_1574);
xnor U2740 (N_2740,N_783,N_1235);
and U2741 (N_2741,N_1822,N_1882);
xnor U2742 (N_2742,N_1078,N_1006);
or U2743 (N_2743,N_2146,N_1650);
nor U2744 (N_2744,N_1259,N_437);
xor U2745 (N_2745,N_2173,N_2034);
and U2746 (N_2746,N_756,N_1387);
nand U2747 (N_2747,N_572,N_1080);
xor U2748 (N_2748,N_715,N_1749);
nand U2749 (N_2749,N_176,N_876);
xor U2750 (N_2750,N_1459,N_353);
nand U2751 (N_2751,N_1219,N_360);
and U2752 (N_2752,N_262,N_681);
nand U2753 (N_2753,N_1695,N_1960);
nor U2754 (N_2754,N_900,N_2422);
and U2755 (N_2755,N_420,N_1804);
nor U2756 (N_2756,N_428,N_177);
or U2757 (N_2757,N_2042,N_2164);
or U2758 (N_2758,N_1716,N_1002);
nor U2759 (N_2759,N_2118,N_142);
and U2760 (N_2760,N_1667,N_986);
or U2761 (N_2761,N_1007,N_2024);
xor U2762 (N_2762,N_2085,N_300);
or U2763 (N_2763,N_1722,N_473);
nor U2764 (N_2764,N_281,N_2099);
nand U2765 (N_2765,N_1258,N_1105);
xor U2766 (N_2766,N_785,N_963);
nand U2767 (N_2767,N_1091,N_1641);
xor U2768 (N_2768,N_1489,N_1510);
or U2769 (N_2769,N_1175,N_2293);
nor U2770 (N_2770,N_4,N_637);
and U2771 (N_2771,N_202,N_1174);
nand U2772 (N_2772,N_1977,N_1865);
nand U2773 (N_2773,N_1188,N_643);
nand U2774 (N_2774,N_129,N_2119);
xor U2775 (N_2775,N_47,N_2302);
nor U2776 (N_2776,N_1748,N_94);
and U2777 (N_2777,N_753,N_127);
xnor U2778 (N_2778,N_96,N_608);
or U2779 (N_2779,N_1743,N_559);
or U2780 (N_2780,N_487,N_1412);
xnor U2781 (N_2781,N_2154,N_1986);
or U2782 (N_2782,N_181,N_1225);
and U2783 (N_2783,N_958,N_75);
xor U2784 (N_2784,N_2330,N_2415);
nand U2785 (N_2785,N_1710,N_2149);
xor U2786 (N_2786,N_1963,N_2088);
and U2787 (N_2787,N_394,N_599);
xor U2788 (N_2788,N_628,N_685);
nand U2789 (N_2789,N_1052,N_557);
nor U2790 (N_2790,N_617,N_1936);
or U2791 (N_2791,N_1766,N_1661);
nand U2792 (N_2792,N_156,N_310);
and U2793 (N_2793,N_1384,N_2260);
or U2794 (N_2794,N_1673,N_793);
nor U2795 (N_2795,N_1197,N_704);
nand U2796 (N_2796,N_1166,N_1996);
nor U2797 (N_2797,N_2246,N_806);
nor U2798 (N_2798,N_1481,N_2017);
xnor U2799 (N_2799,N_1172,N_1932);
and U2800 (N_2800,N_1662,N_971);
and U2801 (N_2801,N_610,N_1611);
or U2802 (N_2802,N_401,N_213);
nor U2803 (N_2803,N_524,N_2037);
nor U2804 (N_2804,N_2262,N_1177);
and U2805 (N_2805,N_1536,N_1051);
nor U2806 (N_2806,N_378,N_1832);
or U2807 (N_2807,N_1789,N_1929);
and U2808 (N_2808,N_1161,N_1694);
or U2809 (N_2809,N_1194,N_2495);
and U2810 (N_2810,N_24,N_150);
xor U2811 (N_2811,N_2312,N_283);
and U2812 (N_2812,N_58,N_1638);
or U2813 (N_2813,N_122,N_878);
or U2814 (N_2814,N_375,N_173);
and U2815 (N_2815,N_1862,N_1887);
and U2816 (N_2816,N_2238,N_1995);
and U2817 (N_2817,N_2139,N_1552);
nand U2818 (N_2818,N_696,N_99);
nor U2819 (N_2819,N_334,N_1529);
nor U2820 (N_2820,N_919,N_454);
nor U2821 (N_2821,N_171,N_1588);
xnor U2822 (N_2822,N_1419,N_102);
or U2823 (N_2823,N_737,N_89);
xor U2824 (N_2824,N_1152,N_2102);
or U2825 (N_2825,N_1528,N_57);
xnor U2826 (N_2826,N_1928,N_2186);
nand U2827 (N_2827,N_2443,N_2497);
and U2828 (N_2828,N_1840,N_2041);
nand U2829 (N_2829,N_66,N_49);
xor U2830 (N_2830,N_761,N_2053);
nand U2831 (N_2831,N_2403,N_569);
and U2832 (N_2832,N_2493,N_1038);
or U2833 (N_2833,N_1594,N_1362);
and U2834 (N_2834,N_2048,N_1801);
xor U2835 (N_2835,N_915,N_809);
xor U2836 (N_2836,N_1771,N_2059);
nand U2837 (N_2837,N_2296,N_1345);
and U2838 (N_2838,N_1234,N_2060);
or U2839 (N_2839,N_377,N_2434);
or U2840 (N_2840,N_205,N_663);
nor U2841 (N_2841,N_443,N_431);
and U2842 (N_2842,N_2279,N_1104);
nor U2843 (N_2843,N_2096,N_591);
or U2844 (N_2844,N_2189,N_1944);
or U2845 (N_2845,N_1923,N_81);
or U2846 (N_2846,N_1182,N_566);
and U2847 (N_2847,N_7,N_1909);
nor U2848 (N_2848,N_494,N_1856);
nor U2849 (N_2849,N_2498,N_45);
or U2850 (N_2850,N_1517,N_249);
nor U2851 (N_2851,N_2428,N_1788);
nand U2852 (N_2852,N_1752,N_677);
or U2853 (N_2853,N_2237,N_1550);
and U2854 (N_2854,N_1848,N_2208);
or U2855 (N_2855,N_1674,N_2301);
nand U2856 (N_2856,N_1477,N_1702);
nor U2857 (N_2857,N_193,N_1508);
nor U2858 (N_2858,N_234,N_2120);
nor U2859 (N_2859,N_1914,N_1855);
and U2860 (N_2860,N_311,N_2319);
and U2861 (N_2861,N_140,N_1064);
nor U2862 (N_2862,N_1844,N_2133);
nor U2863 (N_2863,N_1042,N_697);
or U2864 (N_2864,N_1787,N_125);
or U2865 (N_2865,N_2464,N_1469);
and U2866 (N_2866,N_1970,N_1001);
or U2867 (N_2867,N_2079,N_1227);
nor U2868 (N_2868,N_506,N_426);
nor U2869 (N_2869,N_977,N_1513);
xnor U2870 (N_2870,N_62,N_869);
nor U2871 (N_2871,N_1663,N_840);
and U2872 (N_2872,N_1377,N_1237);
nor U2873 (N_2873,N_2339,N_1146);
and U2874 (N_2874,N_2039,N_165);
and U2875 (N_2875,N_1711,N_2);
nor U2876 (N_2876,N_1976,N_39);
or U2877 (N_2877,N_411,N_1306);
nand U2878 (N_2878,N_1993,N_2258);
or U2879 (N_2879,N_644,N_1277);
and U2880 (N_2880,N_1429,N_1793);
or U2881 (N_2881,N_935,N_848);
or U2882 (N_2882,N_137,N_1713);
nand U2883 (N_2883,N_219,N_818);
or U2884 (N_2884,N_1539,N_1280);
nor U2885 (N_2885,N_74,N_1961);
or U2886 (N_2886,N_2480,N_1298);
nor U2887 (N_2887,N_170,N_2259);
nor U2888 (N_2888,N_2109,N_152);
nand U2889 (N_2889,N_1992,N_117);
nor U2890 (N_2890,N_738,N_168);
xnor U2891 (N_2891,N_162,N_1435);
or U2892 (N_2892,N_717,N_290);
nor U2893 (N_2893,N_2098,N_1208);
and U2894 (N_2894,N_1559,N_2031);
nor U2895 (N_2895,N_656,N_820);
or U2896 (N_2896,N_2449,N_2003);
nor U2897 (N_2897,N_2288,N_856);
nor U2898 (N_2898,N_917,N_1547);
or U2899 (N_2899,N_196,N_2492);
and U2900 (N_2900,N_497,N_1344);
nand U2901 (N_2901,N_504,N_1257);
nand U2902 (N_2902,N_1013,N_2286);
or U2903 (N_2903,N_273,N_78);
nand U2904 (N_2904,N_1655,N_235);
or U2905 (N_2905,N_357,N_1382);
or U2906 (N_2906,N_1077,N_880);
nand U2907 (N_2907,N_1411,N_1561);
and U2908 (N_2908,N_1973,N_2419);
and U2909 (N_2909,N_1998,N_2049);
or U2910 (N_2910,N_2196,N_2329);
nor U2911 (N_2911,N_740,N_1560);
xnor U2912 (N_2912,N_319,N_1329);
xor U2913 (N_2913,N_1507,N_1691);
nor U2914 (N_2914,N_1406,N_406);
xnor U2915 (N_2915,N_1252,N_1703);
nand U2916 (N_2916,N_1096,N_2371);
and U2917 (N_2917,N_1589,N_1181);
or U2918 (N_2918,N_618,N_169);
or U2919 (N_2919,N_2087,N_1421);
nor U2920 (N_2920,N_130,N_2266);
nand U2921 (N_2921,N_1135,N_20);
xor U2922 (N_2922,N_1355,N_476);
nand U2923 (N_2923,N_1132,N_1356);
xor U2924 (N_2924,N_581,N_712);
and U2925 (N_2925,N_1430,N_787);
nand U2926 (N_2926,N_2180,N_2360);
nor U2927 (N_2927,N_1186,N_830);
nor U2928 (N_2928,N_2394,N_1145);
xnor U2929 (N_2929,N_1570,N_1089);
or U2930 (N_2930,N_1879,N_2440);
nor U2931 (N_2931,N_2167,N_1248);
nor U2932 (N_2932,N_1532,N_1780);
and U2933 (N_2933,N_1942,N_709);
and U2934 (N_2934,N_2202,N_2161);
xor U2935 (N_2935,N_553,N_28);
xnor U2936 (N_2936,N_356,N_2481);
nand U2937 (N_2937,N_1965,N_788);
or U2938 (N_2938,N_1541,N_2082);
nor U2939 (N_2939,N_1238,N_1103);
xnor U2940 (N_2940,N_970,N_1343);
nand U2941 (N_2941,N_1745,N_1364);
or U2942 (N_2942,N_741,N_446);
nor U2943 (N_2943,N_711,N_441);
xnor U2944 (N_2944,N_1506,N_814);
xor U2945 (N_2945,N_2439,N_727);
and U2946 (N_2946,N_2155,N_913);
xor U2947 (N_2947,N_1587,N_112);
or U2948 (N_2948,N_324,N_772);
or U2949 (N_2949,N_760,N_688);
nor U2950 (N_2950,N_1439,N_651);
and U2951 (N_2951,N_605,N_1573);
xnor U2952 (N_2952,N_2278,N_630);
nor U2953 (N_2953,N_1034,N_1863);
or U2954 (N_2954,N_359,N_1171);
xor U2955 (N_2955,N_308,N_1392);
nor U2956 (N_2956,N_2036,N_530);
or U2957 (N_2957,N_1625,N_1434);
nand U2958 (N_2958,N_457,N_231);
nand U2959 (N_2959,N_1579,N_1624);
xnor U2960 (N_2960,N_780,N_2285);
nand U2961 (N_2961,N_2010,N_947);
nand U2962 (N_2962,N_1830,N_488);
nand U2963 (N_2963,N_1516,N_528);
and U2964 (N_2964,N_1471,N_1690);
xnor U2965 (N_2965,N_522,N_1810);
and U2966 (N_2966,N_1108,N_798);
or U2967 (N_2967,N_2183,N_413);
xnor U2968 (N_2968,N_309,N_0);
nor U2969 (N_2969,N_1046,N_1653);
nand U2970 (N_2970,N_27,N_945);
xor U2971 (N_2971,N_1366,N_632);
and U2972 (N_2972,N_1418,N_1719);
nand U2973 (N_2973,N_1417,N_1737);
nor U2974 (N_2974,N_1150,N_1926);
xnor U2975 (N_2975,N_1873,N_1683);
nand U2976 (N_2976,N_620,N_2425);
and U2977 (N_2977,N_545,N_301);
xor U2978 (N_2978,N_1950,N_1534);
or U2979 (N_2979,N_1302,N_1451);
and U2980 (N_2980,N_2134,N_109);
nand U2981 (N_2981,N_1358,N_533);
xnor U2982 (N_2982,N_2303,N_1747);
or U2983 (N_2983,N_405,N_1332);
nand U2984 (N_2984,N_133,N_1142);
nor U2985 (N_2985,N_2290,N_2277);
or U2986 (N_2986,N_1676,N_1488);
nand U2987 (N_2987,N_434,N_23);
nand U2988 (N_2988,N_1952,N_2052);
or U2989 (N_2989,N_2177,N_540);
xnor U2990 (N_2990,N_149,N_1374);
nor U2991 (N_2991,N_1894,N_1857);
nand U2992 (N_2992,N_998,N_354);
nor U2993 (N_2993,N_641,N_1003);
or U2994 (N_2994,N_2441,N_1498);
and U2995 (N_2995,N_1326,N_5);
nor U2996 (N_2996,N_2412,N_631);
xnor U2997 (N_2997,N_322,N_965);
and U2998 (N_2998,N_1255,N_412);
nor U2999 (N_2999,N_1022,N_2160);
nor U3000 (N_3000,N_1981,N_2299);
or U3001 (N_3001,N_824,N_1635);
xor U3002 (N_3002,N_455,N_576);
and U3003 (N_3003,N_962,N_1778);
xor U3004 (N_3004,N_2225,N_710);
nor U3005 (N_3005,N_449,N_427);
and U3006 (N_3006,N_379,N_2450);
xnor U3007 (N_3007,N_1520,N_1178);
nand U3008 (N_3008,N_1260,N_728);
nand U3009 (N_3009,N_953,N_2226);
or U3010 (N_3010,N_1757,N_2080);
xor U3011 (N_3011,N_289,N_1389);
or U3012 (N_3012,N_26,N_383);
and U3013 (N_3013,N_1082,N_138);
xor U3014 (N_3014,N_1011,N_2399);
or U3015 (N_3015,N_279,N_676);
nand U3016 (N_3016,N_1390,N_263);
nand U3017 (N_3017,N_1687,N_2365);
nand U3018 (N_3018,N_693,N_853);
nor U3019 (N_3019,N_1054,N_1501);
or U3020 (N_3020,N_2199,N_587);
and U3021 (N_3021,N_1896,N_816);
nand U3022 (N_3022,N_1972,N_1851);
or U3023 (N_3023,N_552,N_502);
nor U3024 (N_3024,N_248,N_1734);
nor U3025 (N_3025,N_1141,N_912);
xnor U3026 (N_3026,N_1750,N_2364);
nand U3027 (N_3027,N_616,N_185);
nor U3028 (N_3028,N_1503,N_2227);
or U3029 (N_3029,N_1889,N_1372);
and U3030 (N_3030,N_1020,N_2472);
nor U3031 (N_3031,N_1223,N_2151);
nand U3032 (N_3032,N_1074,N_1629);
xor U3033 (N_3033,N_1697,N_948);
xnor U3034 (N_3034,N_2163,N_479);
xor U3035 (N_3035,N_2035,N_2484);
or U3036 (N_3036,N_1162,N_204);
and U3037 (N_3037,N_2192,N_2138);
nand U3038 (N_3038,N_2256,N_1839);
and U3039 (N_3039,N_1721,N_2054);
or U3040 (N_3040,N_2328,N_1198);
or U3041 (N_3041,N_1675,N_887);
nor U3042 (N_3042,N_2485,N_223);
nor U3043 (N_3043,N_2029,N_2011);
nand U3044 (N_3044,N_625,N_797);
nor U3045 (N_3045,N_2055,N_86);
nand U3046 (N_3046,N_1933,N_626);
nor U3047 (N_3047,N_2027,N_1872);
xnor U3048 (N_3048,N_477,N_1290);
xnor U3049 (N_3049,N_2125,N_1576);
and U3050 (N_3050,N_865,N_1299);
nor U3051 (N_3051,N_784,N_1265);
xnor U3052 (N_3052,N_718,N_966);
or U3053 (N_3053,N_1823,N_1835);
nand U3054 (N_3054,N_1480,N_730);
nor U3055 (N_3055,N_1206,N_680);
nor U3056 (N_3056,N_734,N_1956);
or U3057 (N_3057,N_1505,N_367);
xnor U3058 (N_3058,N_2148,N_1315);
nor U3059 (N_3059,N_1200,N_261);
nor U3060 (N_3060,N_277,N_1380);
xor U3061 (N_3061,N_1341,N_1656);
and U3062 (N_3062,N_1069,N_1585);
xnor U3063 (N_3063,N_729,N_2214);
xnor U3064 (N_3064,N_1979,N_1478);
xnor U3065 (N_3065,N_382,N_603);
or U3066 (N_3066,N_2321,N_2018);
nor U3067 (N_3067,N_35,N_1495);
xor U3068 (N_3068,N_1279,N_1669);
or U3069 (N_3069,N_1048,N_1569);
nor U3070 (N_3070,N_2326,N_513);
xnor U3071 (N_3071,N_145,N_469);
or U3072 (N_3072,N_116,N_881);
or U3073 (N_3073,N_767,N_1453);
or U3074 (N_3074,N_600,N_1945);
or U3075 (N_3075,N_1875,N_2095);
nand U3076 (N_3076,N_1765,N_1363);
and U3077 (N_3077,N_1639,N_519);
or U3078 (N_3078,N_278,N_1634);
nand U3079 (N_3079,N_799,N_1836);
xor U3080 (N_3080,N_1869,N_2142);
nor U3081 (N_3081,N_2352,N_860);
nand U3082 (N_3082,N_2219,N_918);
or U3083 (N_3083,N_276,N_838);
and U3084 (N_3084,N_51,N_515);
or U3085 (N_3085,N_1271,N_526);
and U3086 (N_3086,N_1754,N_179);
and U3087 (N_3087,N_2115,N_287);
xnor U3088 (N_3088,N_1562,N_580);
nor U3089 (N_3089,N_2270,N_1596);
or U3090 (N_3090,N_1250,N_754);
or U3091 (N_3091,N_2213,N_371);
nand U3092 (N_3092,N_1876,N_1781);
nand U3093 (N_3093,N_1566,N_366);
and U3094 (N_3094,N_217,N_1106);
nand U3095 (N_3095,N_828,N_463);
nor U3096 (N_3096,N_645,N_811);
or U3097 (N_3097,N_2310,N_573);
xor U3098 (N_3098,N_1500,N_2152);
nand U3099 (N_3099,N_419,N_1397);
xor U3100 (N_3100,N_1075,N_313);
nand U3101 (N_3101,N_925,N_1751);
xor U3102 (N_3102,N_535,N_25);
or U3103 (N_3103,N_355,N_1640);
nor U3104 (N_3104,N_1626,N_1519);
xor U3105 (N_3105,N_1892,N_2333);
nor U3106 (N_3106,N_636,N_1701);
nand U3107 (N_3107,N_1537,N_934);
xor U3108 (N_3108,N_514,N_417);
or U3109 (N_3109,N_509,N_1906);
nand U3110 (N_3110,N_1883,N_1785);
and U3111 (N_3111,N_609,N_2282);
xor U3112 (N_3112,N_267,N_1809);
and U3113 (N_3113,N_11,N_1262);
and U3114 (N_3114,N_2334,N_2458);
and U3115 (N_3115,N_1514,N_2389);
nand U3116 (N_3116,N_1652,N_2411);
and U3117 (N_3117,N_796,N_1555);
or U3118 (N_3118,N_672,N_2287);
xor U3119 (N_3119,N_624,N_831);
nand U3120 (N_3120,N_2407,N_1978);
and U3121 (N_3121,N_916,N_2101);
xnor U3122 (N_3122,N_22,N_2073);
xnor U3123 (N_3123,N_328,N_2012);
nor U3124 (N_3124,N_2254,N_627);
nand U3125 (N_3125,N_1643,N_1939);
nand U3126 (N_3126,N_1158,N_1404);
nand U3127 (N_3127,N_863,N_54);
xor U3128 (N_3128,N_126,N_461);
nor U3129 (N_3129,N_2404,N_8);
and U3130 (N_3130,N_1292,N_83);
and U3131 (N_3131,N_2234,N_490);
xnor U3132 (N_3132,N_29,N_2332);
and U3133 (N_3133,N_1616,N_1483);
and U3134 (N_3134,N_1764,N_846);
and U3135 (N_3135,N_1119,N_1704);
nand U3136 (N_3136,N_1324,N_1919);
nand U3137 (N_3137,N_1233,N_1228);
and U3138 (N_3138,N_892,N_71);
nor U3139 (N_3139,N_1515,N_2217);
or U3140 (N_3140,N_3,N_629);
nand U3141 (N_3141,N_2240,N_2065);
xor U3142 (N_3142,N_2083,N_1287);
and U3143 (N_3143,N_161,N_1016);
or U3144 (N_3144,N_233,N_184);
or U3145 (N_3145,N_1511,N_1070);
xnor U3146 (N_3146,N_987,N_1473);
and U3147 (N_3147,N_1212,N_79);
or U3148 (N_3148,N_2379,N_1437);
nand U3149 (N_3149,N_749,N_1431);
xnor U3150 (N_3150,N_1947,N_2223);
or U3151 (N_3151,N_1847,N_2361);
nor U3152 (N_3152,N_167,N_815);
and U3153 (N_3153,N_40,N_445);
and U3154 (N_3154,N_1244,N_1917);
nand U3155 (N_3155,N_2005,N_759);
or U3156 (N_3156,N_186,N_1370);
nor U3157 (N_3157,N_1821,N_725);
or U3158 (N_3158,N_2261,N_1239);
nor U3159 (N_3159,N_658,N_1375);
and U3160 (N_3160,N_595,N_53);
nand U3161 (N_3161,N_1648,N_33);
or U3162 (N_3162,N_302,N_239);
xnor U3163 (N_3163,N_2135,N_9);
and U3164 (N_3164,N_1157,N_1458);
and U3165 (N_3165,N_2473,N_121);
and U3166 (N_3166,N_2308,N_376);
and U3167 (N_3167,N_568,N_2150);
nand U3168 (N_3168,N_1696,N_647);
nor U3169 (N_3169,N_346,N_1632);
and U3170 (N_3170,N_2032,N_695);
nand U3171 (N_3171,N_1791,N_2093);
nor U3172 (N_3172,N_1774,N_1678);
or U3173 (N_3173,N_1620,N_735);
nor U3174 (N_3174,N_2451,N_1854);
nand U3175 (N_3175,N_2462,N_2496);
and U3176 (N_3176,N_1138,N_1179);
and U3177 (N_3177,N_2137,N_888);
nand U3178 (N_3178,N_1121,N_555);
or U3179 (N_3179,N_959,N_330);
or U3180 (N_3180,N_1420,N_1447);
nand U3181 (N_3181,N_159,N_1321);
or U3182 (N_3182,N_2220,N_2206);
nand U3183 (N_3183,N_1247,N_343);
nor U3184 (N_3184,N_15,N_2435);
or U3185 (N_3185,N_157,N_1548);
or U3186 (N_3186,N_2209,N_1095);
xnor U3187 (N_3187,N_52,N_1457);
or U3188 (N_3188,N_44,N_284);
xnor U3189 (N_3189,N_2207,N_1742);
or U3190 (N_3190,N_423,N_687);
or U3191 (N_3191,N_1381,N_318);
or U3192 (N_3192,N_2002,N_238);
and U3193 (N_3193,N_2086,N_736);
and U3194 (N_3194,N_2368,N_425);
nand U3195 (N_3195,N_2307,N_1567);
and U3196 (N_3196,N_1167,N_1027);
nor U3197 (N_3197,N_1320,N_333);
or U3198 (N_3198,N_1092,N_478);
and U3199 (N_3199,N_2347,N_907);
xnor U3200 (N_3200,N_2230,N_1902);
or U3201 (N_3201,N_594,N_1367);
and U3202 (N_3202,N_583,N_1126);
or U3203 (N_3203,N_1305,N_1137);
xnor U3204 (N_3204,N_2193,N_1);
and U3205 (N_3205,N_1874,N_825);
xnor U3206 (N_3206,N_653,N_791);
or U3207 (N_3207,N_1005,N_667);
xor U3208 (N_3208,N_1039,N_2381);
xnor U3209 (N_3209,N_1201,N_1545);
nor U3210 (N_3210,N_1149,N_1021);
xor U3211 (N_3211,N_1921,N_743);
nor U3212 (N_3212,N_200,N_2295);
xnor U3213 (N_3213,N_1168,N_2291);
xnor U3214 (N_3214,N_1911,N_1073);
xnor U3215 (N_3215,N_1522,N_2363);
nand U3216 (N_3216,N_365,N_436);
or U3217 (N_3217,N_2474,N_1409);
nor U3218 (N_3218,N_565,N_304);
nand U3219 (N_3219,N_1597,N_460);
xnor U3220 (N_3220,N_1365,N_1901);
nand U3221 (N_3221,N_1805,N_1313);
nor U3222 (N_3222,N_352,N_237);
and U3223 (N_3223,N_2158,N_1815);
xnor U3224 (N_3224,N_210,N_1937);
xor U3225 (N_3225,N_495,N_1057);
and U3226 (N_3226,N_1123,N_332);
xor U3227 (N_3227,N_1586,N_1642);
and U3228 (N_3228,N_1666,N_1693);
or U3229 (N_3229,N_1443,N_1533);
and U3230 (N_3230,N_90,N_485);
nand U3231 (N_3231,N_2247,N_532);
nor U3232 (N_3232,N_362,N_1971);
xor U3233 (N_3233,N_812,N_482);
and U3234 (N_3234,N_132,N_1322);
or U3235 (N_3235,N_1700,N_2203);
xnor U3236 (N_3236,N_794,N_554);
xnor U3237 (N_3237,N_1689,N_212);
or U3238 (N_3238,N_1543,N_402);
and U3239 (N_3239,N_2391,N_134);
xor U3240 (N_3240,N_2143,N_1957);
and U3241 (N_3241,N_1025,N_12);
nand U3242 (N_3242,N_1415,N_291);
nor U3243 (N_3243,N_646,N_2322);
or U3244 (N_3244,N_508,N_2468);
nor U3245 (N_3245,N_1023,N_395);
and U3246 (N_3246,N_2402,N_192);
or U3247 (N_3247,N_832,N_562);
or U3248 (N_3248,N_1987,N_1881);
or U3249 (N_3249,N_946,N_1120);
xnor U3250 (N_3250,N_1598,N_1325);
or U3251 (N_3251,N_686,N_227);
xnor U3252 (N_3252,N_1609,N_2367);
and U3253 (N_3253,N_1352,N_252);
and U3254 (N_3254,N_1592,N_468);
and U3255 (N_3255,N_1097,N_2067);
nand U3256 (N_3256,N_73,N_1154);
and U3257 (N_3257,N_692,N_1779);
nand U3258 (N_3258,N_2429,N_2317);
xor U3259 (N_3259,N_1490,N_2008);
nand U3260 (N_3260,N_2272,N_1422);
nor U3261 (N_3261,N_2190,N_1647);
xnor U3262 (N_3262,N_340,N_91);
xnor U3263 (N_3263,N_2465,N_400);
and U3264 (N_3264,N_871,N_241);
xor U3265 (N_3265,N_898,N_1215);
nor U3266 (N_3266,N_1739,N_1224);
or U3267 (N_3267,N_2323,N_2195);
or U3268 (N_3268,N_1614,N_744);
xnor U3269 (N_3269,N_1159,N_2370);
or U3270 (N_3270,N_1336,N_368);
or U3271 (N_3271,N_1268,N_387);
xor U3272 (N_3272,N_1143,N_1931);
nor U3273 (N_3273,N_2251,N_164);
nand U3274 (N_3274,N_218,N_2074);
and U3275 (N_3275,N_317,N_285);
and U3276 (N_3276,N_269,N_766);
xnor U3277 (N_3277,N_1850,N_1156);
xor U3278 (N_3278,N_635,N_1846);
xnor U3279 (N_3279,N_1173,N_1014);
nand U3280 (N_3280,N_1951,N_652);
nand U3281 (N_3281,N_2269,N_757);
xor U3282 (N_3282,N_381,N_2090);
and U3283 (N_3283,N_1802,N_570);
and U3284 (N_3284,N_778,N_1491);
nor U3285 (N_3285,N_1084,N_1784);
xnor U3286 (N_3286,N_2271,N_911);
xnor U3287 (N_3287,N_392,N_297);
and U3288 (N_3288,N_991,N_1209);
and U3289 (N_3289,N_1334,N_1193);
nand U3290 (N_3290,N_2171,N_1767);
or U3291 (N_3291,N_251,N_1544);
nor U3292 (N_3292,N_1727,N_2249);
or U3293 (N_3293,N_325,N_2338);
or U3294 (N_3294,N_993,N_148);
nor U3295 (N_3295,N_1799,N_801);
nor U3296 (N_3296,N_63,N_665);
and U3297 (N_3297,N_1087,N_678);
nor U3298 (N_3298,N_982,N_1114);
xnor U3299 (N_3299,N_808,N_1590);
xnor U3300 (N_3300,N_68,N_2446);
or U3301 (N_3301,N_1291,N_1408);
xnor U3302 (N_3302,N_957,N_700);
nor U3303 (N_3303,N_2275,N_2410);
nand U3304 (N_3304,N_802,N_614);
nor U3305 (N_3305,N_350,N_660);
xor U3306 (N_3306,N_2200,N_222);
nand U3307 (N_3307,N_955,N_385);
and U3308 (N_3308,N_927,N_1388);
nor U3309 (N_3309,N_1210,N_1741);
and U3310 (N_3310,N_1714,N_1818);
nand U3311 (N_3311,N_1493,N_59);
and U3312 (N_3312,N_2356,N_1808);
nor U3313 (N_3313,N_2194,N_1607);
or U3314 (N_3314,N_1230,N_1354);
or U3315 (N_3315,N_450,N_2179);
and U3316 (N_3316,N_260,N_2084);
nand U3317 (N_3317,N_144,N_2130);
xnor U3318 (N_3318,N_2156,N_874);
and U3319 (N_3319,N_194,N_542);
or U3320 (N_3320,N_1619,N_1441);
xnor U3321 (N_3321,N_996,N_841);
or U3322 (N_3322,N_1242,N_2111);
xnor U3323 (N_3323,N_1465,N_2414);
and U3324 (N_3324,N_2044,N_430);
or U3325 (N_3325,N_1797,N_124);
or U3326 (N_3326,N_1031,N_1044);
nand U3327 (N_3327,N_207,N_551);
nand U3328 (N_3328,N_2416,N_1118);
xor U3329 (N_3329,N_2354,N_1786);
xnor U3330 (N_3330,N_2366,N_1554);
nor U3331 (N_3331,N_590,N_910);
nand U3332 (N_3332,N_1893,N_1568);
or U3333 (N_3333,N_1867,N_1213);
xor U3334 (N_3334,N_842,N_1649);
and U3335 (N_3335,N_496,N_713);
or U3336 (N_3336,N_1155,N_2026);
or U3337 (N_3337,N_16,N_1216);
or U3338 (N_3338,N_107,N_1128);
or U3339 (N_3339,N_2028,N_493);
xnor U3340 (N_3340,N_316,N_1281);
and U3341 (N_3341,N_1740,N_771);
and U3342 (N_3342,N_1029,N_2218);
nand U3343 (N_3343,N_1187,N_2357);
or U3344 (N_3344,N_1318,N_2182);
or U3345 (N_3345,N_1129,N_111);
and U3346 (N_3346,N_61,N_1563);
nand U3347 (N_3347,N_1946,N_2466);
or U3348 (N_3348,N_1407,N_1895);
or U3349 (N_3349,N_2313,N_972);
xor U3350 (N_3350,N_980,N_1398);
and U3351 (N_3351,N_1726,N_1817);
and U3352 (N_3352,N_1732,N_348);
or U3353 (N_3353,N_777,N_1414);
nand U3354 (N_3354,N_732,N_2377);
nor U3355 (N_3355,N_1053,N_191);
and U3356 (N_3356,N_1169,N_719);
nand U3357 (N_3357,N_2489,N_2123);
xor U3358 (N_3358,N_1866,N_1795);
and U3359 (N_3359,N_2121,N_46);
or U3360 (N_3360,N_775,N_1327);
and U3361 (N_3361,N_465,N_1602);
xor U3362 (N_3362,N_119,N_852);
and U3363 (N_3363,N_1294,N_1841);
or U3364 (N_3364,N_2063,N_2424);
nand U3365 (N_3365,N_2460,N_139);
and U3366 (N_3366,N_41,N_374);
nand U3367 (N_3367,N_393,N_2304);
nor U3368 (N_3368,N_1834,N_1903);
nor U3369 (N_3369,N_2162,N_699);
xnor U3370 (N_3370,N_1482,N_363);
and U3371 (N_3371,N_244,N_1692);
nand U3372 (N_3372,N_593,N_503);
nand U3373 (N_3373,N_896,N_2445);
and U3374 (N_3374,N_2140,N_770);
nor U3375 (N_3375,N_622,N_2483);
and U3376 (N_3376,N_128,N_1445);
nor U3377 (N_3377,N_1393,N_2461);
nand U3378 (N_3378,N_1603,N_891);
and U3379 (N_3379,N_2316,N_868);
nor U3380 (N_3380,N_242,N_1659);
xnor U3381 (N_3381,N_2153,N_1838);
nor U3382 (N_3382,N_2486,N_1428);
xor U3383 (N_3383,N_1880,N_1858);
nor U3384 (N_3384,N_1426,N_1111);
xnor U3385 (N_3385,N_823,N_1924);
and U3386 (N_3386,N_2197,N_2131);
and U3387 (N_3387,N_1908,N_1645);
nor U3388 (N_3388,N_2248,N_2078);
or U3389 (N_3389,N_1982,N_1680);
or U3390 (N_3390,N_2376,N_2221);
nand U3391 (N_3391,N_1218,N_517);
and U3392 (N_3392,N_1323,N_1307);
xor U3393 (N_3393,N_1101,N_845);
xor U3394 (N_3394,N_1079,N_1102);
xnor U3395 (N_3395,N_1402,N_1842);
or U3396 (N_3396,N_21,N_1176);
and U3397 (N_3397,N_564,N_984);
nand U3398 (N_3398,N_50,N_70);
nor U3399 (N_3399,N_2418,N_750);
and U3400 (N_3400,N_2229,N_1497);
and U3401 (N_3401,N_1308,N_1796);
and U3402 (N_3402,N_1035,N_1994);
or U3403 (N_3403,N_722,N_187);
nand U3404 (N_3404,N_1829,N_1725);
and U3405 (N_3405,N_1775,N_2058);
and U3406 (N_3406,N_1191,N_1311);
nand U3407 (N_3407,N_534,N_1679);
and U3408 (N_3408,N_1523,N_989);
nand U3409 (N_3409,N_2490,N_523);
nor U3410 (N_3410,N_292,N_2004);
nor U3411 (N_3411,N_2292,N_166);
and U3412 (N_3412,N_76,N_800);
or U3413 (N_3413,N_859,N_861);
nand U3414 (N_3414,N_2241,N_596);
or U3415 (N_3415,N_567,N_1379);
xor U3416 (N_3416,N_2475,N_104);
nor U3417 (N_3417,N_995,N_1580);
nand U3418 (N_3418,N_2165,N_764);
xor U3419 (N_3419,N_2380,N_2159);
and U3420 (N_3420,N_847,N_936);
xnor U3421 (N_3421,N_1730,N_2104);
and U3422 (N_3422,N_2176,N_2349);
and U3423 (N_3423,N_1512,N_1904);
or U3424 (N_3424,N_1165,N_619);
and U3425 (N_3425,N_1026,N_1350);
or U3426 (N_3426,N_245,N_929);
xnor U3427 (N_3427,N_2061,N_2491);
nand U3428 (N_3428,N_1214,N_103);
and U3429 (N_3429,N_2145,N_851);
nand U3430 (N_3430,N_1706,N_2420);
nand U3431 (N_3431,N_1153,N_1760);
nand U3432 (N_3432,N_435,N_1927);
nand U3433 (N_3433,N_1621,N_2253);
or U3434 (N_3434,N_1644,N_1853);
and U3435 (N_3435,N_2477,N_1811);
or U3436 (N_3436,N_1256,N_82);
and U3437 (N_3437,N_670,N_123);
and U3438 (N_3438,N_2469,N_1319);
nor U3439 (N_3439,N_769,N_444);
or U3440 (N_3440,N_1783,N_960);
nor U3441 (N_3441,N_763,N_1759);
nor U3442 (N_3442,N_2297,N_87);
and U3443 (N_3443,N_1373,N_1264);
and U3444 (N_3444,N_1685,N_1475);
xor U3445 (N_3445,N_143,N_2487);
nand U3446 (N_3446,N_1890,N_303);
nand U3447 (N_3447,N_2057,N_180);
or U3448 (N_3448,N_786,N_440);
and U3449 (N_3449,N_1476,N_1236);
and U3450 (N_3450,N_2373,N_462);
or U3451 (N_3451,N_2066,N_1715);
nand U3452 (N_3452,N_1226,N_2311);
nor U3453 (N_3453,N_1229,N_183);
and U3454 (N_3454,N_877,N_294);
nand U3455 (N_3455,N_1283,N_2309);
nand U3456 (N_3456,N_1958,N_1253);
xnor U3457 (N_3457,N_1470,N_978);
or U3458 (N_3458,N_708,N_2340);
xor U3459 (N_3459,N_810,N_397);
nor U3460 (N_3460,N_714,N_2430);
nand U3461 (N_3461,N_1144,N_1357);
xnor U3462 (N_3462,N_415,N_1140);
or U3463 (N_3463,N_1595,N_439);
nand U3464 (N_3464,N_889,N_1660);
nand U3465 (N_3465,N_1015,N_1107);
and U3466 (N_3466,N_855,N_2294);
nor U3467 (N_3467,N_723,N_1037);
nor U3468 (N_3468,N_1347,N_1953);
or U3469 (N_3469,N_1565,N_1403);
or U3470 (N_3470,N_2210,N_839);
nand U3471 (N_3471,N_199,N_146);
nor U3472 (N_3472,N_1100,N_13);
and U3473 (N_3473,N_2257,N_1009);
nand U3474 (N_3474,N_389,N_247);
or U3475 (N_3475,N_2069,N_951);
or U3476 (N_3476,N_2342,N_64);
or U3477 (N_3477,N_1232,N_1284);
nand U3478 (N_3478,N_857,N_266);
nor U3479 (N_3479,N_1399,N_529);
and U3480 (N_3480,N_579,N_1861);
or U3481 (N_3481,N_1270,N_833);
and U3482 (N_3482,N_1494,N_475);
or U3483 (N_3483,N_34,N_611);
nor U3484 (N_3484,N_1613,N_1599);
nand U3485 (N_3485,N_408,N_286);
nand U3486 (N_3486,N_32,N_19);
xor U3487 (N_3487,N_1606,N_1199);
and U3488 (N_3488,N_1527,N_837);
nand U3489 (N_3489,N_1081,N_836);
and U3490 (N_3490,N_1130,N_1538);
or U3491 (N_3491,N_2348,N_1814);
xnor U3492 (N_3492,N_2040,N_2265);
nor U3493 (N_3493,N_1061,N_1472);
nand U3494 (N_3494,N_582,N_106);
nor U3495 (N_3495,N_500,N_1340);
nand U3496 (N_3496,N_954,N_1938);
nor U3497 (N_3497,N_879,N_1160);
and U3498 (N_3498,N_1133,N_2350);
nand U3499 (N_3499,N_516,N_1826);
nand U3500 (N_3500,N_1935,N_999);
nor U3501 (N_3501,N_2222,N_1967);
or U3502 (N_3502,N_56,N_1968);
nor U3503 (N_3503,N_762,N_1351);
nand U3504 (N_3504,N_1449,N_1019);
or U3505 (N_3505,N_549,N_2033);
nor U3506 (N_3506,N_483,N_779);
and U3507 (N_3507,N_2426,N_2000);
or U3508 (N_3508,N_282,N_2239);
or U3509 (N_3509,N_867,N_873);
or U3510 (N_3510,N_1220,N_351);
or U3511 (N_3511,N_211,N_264);
nand U3512 (N_3512,N_2068,N_358);
nand U3513 (N_3513,N_720,N_598);
or U3514 (N_3514,N_1578,N_459);
xor U3515 (N_3515,N_1274,N_518);
xnor U3516 (N_3516,N_1800,N_174);
nor U3517 (N_3517,N_2436,N_2030);
nand U3518 (N_3518,N_347,N_198);
or U3519 (N_3519,N_1886,N_943);
nor U3520 (N_3520,N_2401,N_2341);
nand U3521 (N_3521,N_571,N_2324);
nand U3522 (N_3522,N_602,N_2423);
nor U3523 (N_3523,N_2007,N_932);
or U3524 (N_3524,N_2105,N_407);
nor U3525 (N_3525,N_585,N_208);
nand U3526 (N_3526,N_1542,N_1556);
xor U3527 (N_3527,N_1050,N_2454);
or U3528 (N_3528,N_2174,N_2397);
nor U3529 (N_3529,N_424,N_1487);
xor U3530 (N_3530,N_1828,N_1267);
or U3531 (N_3531,N_2023,N_2245);
nand U3532 (N_3532,N_288,N_822);
and U3533 (N_3533,N_589,N_14);
or U3534 (N_3534,N_422,N_458);
nand U3535 (N_3535,N_2081,N_2228);
or U3536 (N_3536,N_1192,N_924);
and U3537 (N_3537,N_1708,N_1705);
xor U3538 (N_3538,N_1665,N_80);
or U3539 (N_3539,N_2094,N_2267);
nor U3540 (N_3540,N_2169,N_1698);
xor U3541 (N_3541,N_396,N_2020);
xnor U3542 (N_3542,N_2467,N_1790);
nand U3543 (N_3543,N_1540,N_1798);
nand U3544 (N_3544,N_988,N_1776);
xor U3545 (N_3545,N_906,N_221);
or U3546 (N_3546,N_1816,N_1289);
nor U3547 (N_3547,N_18,N_2124);
or U3548 (N_3548,N_158,N_850);
or U3549 (N_3549,N_903,N_1618);
and U3550 (N_3550,N_691,N_1974);
nand U3551 (N_3551,N_930,N_2175);
nor U3552 (N_3552,N_1333,N_472);
nor U3553 (N_3553,N_1916,N_2421);
nor U3554 (N_3554,N_1955,N_1112);
nor U3555 (N_3555,N_638,N_2191);
and U3556 (N_3556,N_893,N_2112);
nor U3557 (N_3557,N_265,N_254);
and U3558 (N_3558,N_2444,N_862);
nor U3559 (N_3559,N_1792,N_2406);
and U3560 (N_3560,N_1718,N_1316);
or U3561 (N_3561,N_2400,N_77);
nor U3562 (N_3562,N_817,N_216);
nand U3563 (N_3563,N_1753,N_2273);
and U3564 (N_3564,N_1651,N_448);
nor U3565 (N_3565,N_968,N_1083);
and U3566 (N_3566,N_2110,N_1147);
and U3567 (N_3567,N_1915,N_1984);
nor U3568 (N_3568,N_640,N_703);
nor U3569 (N_3569,N_342,N_451);
nor U3570 (N_3570,N_537,N_1827);
nand U3571 (N_3571,N_1553,N_1195);
and U3572 (N_3572,N_1593,N_1423);
and U3573 (N_3573,N_2006,N_1017);
nand U3574 (N_3574,N_558,N_1300);
nand U3575 (N_3575,N_1203,N_1076);
and U3576 (N_3576,N_1249,N_2398);
or U3577 (N_3577,N_1668,N_1954);
nand U3578 (N_3578,N_1463,N_1684);
and U3579 (N_3579,N_792,N_1633);
xor U3580 (N_3580,N_983,N_1859);
nand U3581 (N_3581,N_2046,N_349);
nor U3582 (N_3582,N_1060,N_2116);
nand U3583 (N_3583,N_42,N_384);
xnor U3584 (N_3584,N_1361,N_1433);
xnor U3585 (N_3585,N_961,N_258);
and U3586 (N_3586,N_1067,N_1999);
xor U3587 (N_3587,N_1709,N_1033);
nand U3588 (N_3588,N_1782,N_1040);
xor U3589 (N_3589,N_298,N_2494);
and U3590 (N_3590,N_499,N_928);
nand U3591 (N_3591,N_2457,N_268);
nor U3592 (N_3592,N_1825,N_1871);
nand U3593 (N_3593,N_2141,N_175);
xor U3594 (N_3594,N_136,N_364);
xnor U3595 (N_3595,N_2382,N_2043);
nor U3596 (N_3596,N_789,N_507);
xor U3597 (N_3597,N_246,N_666);
xor U3598 (N_3598,N_380,N_1348);
nor U3599 (N_3599,N_154,N_432);
nand U3600 (N_3600,N_118,N_706);
nand U3601 (N_3601,N_648,N_1837);
nand U3602 (N_3602,N_742,N_69);
nor U3603 (N_3603,N_1524,N_2106);
and U3604 (N_3604,N_271,N_189);
nor U3605 (N_3605,N_501,N_694);
or U3606 (N_3606,N_1900,N_253);
nor U3607 (N_3607,N_2476,N_1885);
or U3608 (N_3608,N_886,N_2453);
and U3609 (N_3609,N_2388,N_38);
or U3610 (N_3610,N_1531,N_1925);
nand U3611 (N_3611,N_312,N_2345);
nand U3612 (N_3612,N_1756,N_1116);
xnor U3613 (N_3613,N_1124,N_1385);
xnor U3614 (N_3614,N_120,N_178);
nand U3615 (N_3615,N_758,N_1988);
or U3616 (N_3616,N_690,N_1085);
or U3617 (N_3617,N_716,N_1047);
and U3618 (N_3618,N_197,N_950);
nand U3619 (N_3619,N_65,N_1196);
xnor U3620 (N_3620,N_2359,N_1492);
and U3621 (N_3621,N_1824,N_1335);
or U3622 (N_3622,N_1518,N_10);
nand U3623 (N_3623,N_1127,N_1245);
and U3624 (N_3624,N_1761,N_2353);
nor U3625 (N_3625,N_1582,N_1860);
and U3626 (N_3626,N_659,N_2128);
and U3627 (N_3627,N_1969,N_639);
or U3628 (N_3628,N_1572,N_1717);
xnor U3629 (N_3629,N_2252,N_1852);
xor U3630 (N_3630,N_270,N_577);
or U3631 (N_3631,N_521,N_1376);
nor U3632 (N_3632,N_2355,N_933);
or U3633 (N_3633,N_2417,N_43);
nand U3634 (N_3634,N_2144,N_1045);
nor U3635 (N_3635,N_1959,N_1521);
nand U3636 (N_3636,N_1888,N_1202);
and U3637 (N_3637,N_895,N_1964);
and U3638 (N_3638,N_1295,N_295);
nor U3639 (N_3639,N_293,N_2122);
and U3640 (N_3640,N_1845,N_1136);
and U3641 (N_3641,N_2427,N_2100);
or U3642 (N_3642,N_399,N_901);
and U3643 (N_3643,N_1450,N_339);
or U3644 (N_3644,N_1622,N_1066);
nor U3645 (N_3645,N_578,N_920);
nor U3646 (N_3646,N_2437,N_1293);
xor U3647 (N_3647,N_1877,N_2062);
nand U3648 (N_3648,N_1369,N_373);
and U3649 (N_3649,N_1342,N_155);
or U3650 (N_3650,N_2448,N_1211);
and U3651 (N_3651,N_1425,N_864);
nor U3652 (N_3652,N_2305,N_2097);
nor U3653 (N_3653,N_2022,N_897);
xor U3654 (N_3654,N_110,N_941);
nand U3655 (N_3655,N_805,N_683);
or U3656 (N_3656,N_1485,N_550);
nand U3657 (N_3657,N_505,N_884);
or U3658 (N_3658,N_765,N_2280);
nand U3659 (N_3659,N_1339,N_997);
and U3660 (N_3660,N_844,N_1098);
or U3661 (N_3661,N_37,N_834);
xor U3662 (N_3662,N_2070,N_1670);
or U3663 (N_3663,N_2431,N_615);
nor U3664 (N_3664,N_724,N_938);
nor U3665 (N_3665,N_592,N_1941);
or U3666 (N_3666,N_1943,N_1041);
or U3667 (N_3667,N_1286,N_733);
and U3668 (N_3668,N_2129,N_2375);
nor U3669 (N_3669,N_2232,N_2242);
or U3670 (N_3670,N_2362,N_1729);
or U3671 (N_3671,N_1036,N_1330);
nor U3672 (N_3672,N_1303,N_1278);
nor U3673 (N_3673,N_484,N_220);
nand U3674 (N_3674,N_321,N_97);
xor U3675 (N_3675,N_1183,N_921);
xnor U3676 (N_3676,N_153,N_1899);
xnor U3677 (N_3677,N_707,N_1600);
and U3678 (N_3678,N_952,N_1115);
nand U3679 (N_3679,N_1000,N_634);
xor U3680 (N_3680,N_1686,N_1071);
nand U3681 (N_3681,N_85,N_939);
nor U3682 (N_3682,N_671,N_967);
nor U3683 (N_3683,N_827,N_702);
nand U3684 (N_3684,N_1383,N_1010);
or U3685 (N_3685,N_67,N_1819);
nor U3686 (N_3686,N_2447,N_563);
nor U3687 (N_3687,N_2284,N_1864);
and U3688 (N_3688,N_1486,N_1065);
or U3689 (N_3689,N_209,N_976);
xnor U3690 (N_3690,N_1762,N_1897);
and U3691 (N_3691,N_1849,N_849);
xor U3692 (N_3692,N_544,N_1395);
xnor U3693 (N_3693,N_2016,N_829);
xor U3694 (N_3694,N_1564,N_752);
or U3695 (N_3695,N_746,N_274);
nand U3696 (N_3696,N_1254,N_361);
nor U3697 (N_3697,N_2358,N_1681);
xnor U3698 (N_3698,N_315,N_388);
and U3699 (N_3699,N_1496,N_1870);
xor U3700 (N_3700,N_2344,N_942);
xnor U3701 (N_3701,N_527,N_990);
and U3702 (N_3702,N_731,N_795);
or U3703 (N_3703,N_981,N_2384);
nand U3704 (N_3704,N_1820,N_1769);
xor U3705 (N_3705,N_88,N_1807);
nand U3706 (N_3706,N_2351,N_909);
and U3707 (N_3707,N_2369,N_1309);
nand U3708 (N_3708,N_2442,N_398);
or U3709 (N_3709,N_1446,N_2064);
nand U3710 (N_3710,N_481,N_1391);
nand U3711 (N_3711,N_2346,N_1975);
nand U3712 (N_3712,N_1628,N_113);
or U3713 (N_3713,N_803,N_2076);
nand U3714 (N_3714,N_1378,N_1546);
nor U3715 (N_3715,N_2187,N_1110);
or U3716 (N_3716,N_1444,N_1940);
nand U3717 (N_3717,N_1658,N_1905);
xnor U3718 (N_3718,N_2463,N_973);
or U3719 (N_3719,N_471,N_1577);
or U3720 (N_3720,N_883,N_956);
nand U3721 (N_3721,N_386,N_668);
and U3722 (N_3722,N_2471,N_492);
nand U3723 (N_3723,N_464,N_2045);
xor U3724 (N_3724,N_1424,N_2244);
nand U3725 (N_3725,N_135,N_1699);
or U3726 (N_3726,N_228,N_1055);
xor U3727 (N_3727,N_182,N_2091);
nor U3728 (N_3728,N_1456,N_1525);
xnor U3729 (N_3729,N_489,N_835);
nor U3730 (N_3730,N_160,N_225);
nand U3731 (N_3731,N_525,N_418);
nand U3732 (N_3732,N_1438,N_314);
or U3733 (N_3733,N_1427,N_1535);
or U3734 (N_3734,N_31,N_30);
or U3735 (N_3735,N_108,N_2264);
xnor U3736 (N_3736,N_409,N_1949);
nor U3737 (N_3737,N_299,N_654);
and U3738 (N_3738,N_1918,N_2009);
nand U3739 (N_3739,N_2092,N_336);
and U3740 (N_3740,N_172,N_773);
nand U3741 (N_3741,N_2390,N_2014);
xor U3742 (N_3742,N_538,N_272);
nand U3743 (N_3743,N_467,N_1131);
nand U3744 (N_3744,N_1912,N_2136);
nand U3745 (N_3745,N_940,N_1452);
or U3746 (N_3746,N_2336,N_584);
and U3747 (N_3747,N_1526,N_1499);
nor U3748 (N_3748,N_560,N_536);
nor U3749 (N_3749,N_372,N_1440);
nand U3750 (N_3750,N_1019,N_1492);
and U3751 (N_3751,N_2043,N_278);
nand U3752 (N_3752,N_572,N_2134);
nor U3753 (N_3753,N_2241,N_2045);
nand U3754 (N_3754,N_966,N_2279);
xor U3755 (N_3755,N_847,N_1831);
nand U3756 (N_3756,N_957,N_568);
nand U3757 (N_3757,N_936,N_814);
xnor U3758 (N_3758,N_580,N_1639);
nor U3759 (N_3759,N_2209,N_1286);
or U3760 (N_3760,N_2405,N_1861);
xnor U3761 (N_3761,N_1446,N_222);
and U3762 (N_3762,N_678,N_1878);
xnor U3763 (N_3763,N_874,N_637);
xnor U3764 (N_3764,N_2361,N_618);
nor U3765 (N_3765,N_52,N_1409);
xnor U3766 (N_3766,N_1766,N_2284);
and U3767 (N_3767,N_208,N_1938);
and U3768 (N_3768,N_2129,N_1486);
xnor U3769 (N_3769,N_244,N_792);
and U3770 (N_3770,N_1018,N_142);
and U3771 (N_3771,N_1456,N_2318);
nand U3772 (N_3772,N_704,N_23);
xnor U3773 (N_3773,N_378,N_2409);
or U3774 (N_3774,N_1606,N_1109);
nand U3775 (N_3775,N_1646,N_1122);
nand U3776 (N_3776,N_2043,N_1920);
nand U3777 (N_3777,N_1781,N_2252);
nor U3778 (N_3778,N_2195,N_1062);
and U3779 (N_3779,N_1649,N_153);
or U3780 (N_3780,N_1566,N_406);
nand U3781 (N_3781,N_1525,N_1506);
xor U3782 (N_3782,N_320,N_1974);
and U3783 (N_3783,N_1144,N_473);
nor U3784 (N_3784,N_542,N_1808);
xor U3785 (N_3785,N_1154,N_2341);
nor U3786 (N_3786,N_2233,N_1557);
and U3787 (N_3787,N_1747,N_2092);
or U3788 (N_3788,N_1350,N_907);
or U3789 (N_3789,N_1677,N_819);
and U3790 (N_3790,N_1638,N_1436);
nand U3791 (N_3791,N_1234,N_55);
nor U3792 (N_3792,N_2134,N_477);
nor U3793 (N_3793,N_660,N_1599);
or U3794 (N_3794,N_1603,N_1323);
xnor U3795 (N_3795,N_2044,N_743);
nand U3796 (N_3796,N_2391,N_1247);
nor U3797 (N_3797,N_435,N_188);
or U3798 (N_3798,N_1082,N_1134);
nand U3799 (N_3799,N_2177,N_1594);
nand U3800 (N_3800,N_941,N_1596);
nand U3801 (N_3801,N_1740,N_1019);
xnor U3802 (N_3802,N_1328,N_1451);
nor U3803 (N_3803,N_517,N_2474);
or U3804 (N_3804,N_2262,N_1973);
and U3805 (N_3805,N_825,N_381);
nand U3806 (N_3806,N_1959,N_2398);
or U3807 (N_3807,N_316,N_48);
or U3808 (N_3808,N_277,N_871);
nand U3809 (N_3809,N_1213,N_1289);
and U3810 (N_3810,N_2243,N_285);
nand U3811 (N_3811,N_672,N_2213);
nand U3812 (N_3812,N_1181,N_1042);
nand U3813 (N_3813,N_878,N_641);
nor U3814 (N_3814,N_2175,N_1880);
or U3815 (N_3815,N_2425,N_2131);
nand U3816 (N_3816,N_1713,N_973);
xor U3817 (N_3817,N_912,N_957);
or U3818 (N_3818,N_98,N_1420);
and U3819 (N_3819,N_2213,N_2054);
nand U3820 (N_3820,N_343,N_2317);
and U3821 (N_3821,N_1273,N_1358);
xor U3822 (N_3822,N_1404,N_805);
and U3823 (N_3823,N_1455,N_1473);
xor U3824 (N_3824,N_1640,N_2406);
nor U3825 (N_3825,N_1705,N_602);
or U3826 (N_3826,N_1453,N_410);
nand U3827 (N_3827,N_2168,N_2408);
nor U3828 (N_3828,N_1415,N_1844);
nand U3829 (N_3829,N_441,N_2423);
nand U3830 (N_3830,N_193,N_1843);
xnor U3831 (N_3831,N_1943,N_441);
or U3832 (N_3832,N_2253,N_1698);
and U3833 (N_3833,N_2167,N_1039);
nor U3834 (N_3834,N_2109,N_1656);
nand U3835 (N_3835,N_276,N_667);
or U3836 (N_3836,N_1395,N_2014);
nor U3837 (N_3837,N_1364,N_761);
and U3838 (N_3838,N_225,N_1958);
nor U3839 (N_3839,N_1236,N_853);
xnor U3840 (N_3840,N_1699,N_1861);
nor U3841 (N_3841,N_9,N_424);
nor U3842 (N_3842,N_2465,N_2093);
and U3843 (N_3843,N_1676,N_64);
or U3844 (N_3844,N_1732,N_1316);
nor U3845 (N_3845,N_901,N_2248);
and U3846 (N_3846,N_709,N_1947);
or U3847 (N_3847,N_255,N_773);
xor U3848 (N_3848,N_39,N_1589);
nor U3849 (N_3849,N_463,N_1981);
nor U3850 (N_3850,N_2114,N_2229);
nor U3851 (N_3851,N_530,N_2037);
nand U3852 (N_3852,N_1812,N_2355);
xnor U3853 (N_3853,N_1666,N_31);
xor U3854 (N_3854,N_326,N_100);
nor U3855 (N_3855,N_959,N_223);
and U3856 (N_3856,N_1936,N_389);
nand U3857 (N_3857,N_1020,N_20);
or U3858 (N_3858,N_1125,N_337);
or U3859 (N_3859,N_1232,N_373);
nand U3860 (N_3860,N_657,N_716);
or U3861 (N_3861,N_1518,N_2007);
and U3862 (N_3862,N_2113,N_1928);
nor U3863 (N_3863,N_511,N_170);
xor U3864 (N_3864,N_2447,N_1517);
xor U3865 (N_3865,N_2060,N_172);
xnor U3866 (N_3866,N_2353,N_354);
or U3867 (N_3867,N_1648,N_570);
or U3868 (N_3868,N_1827,N_1561);
nand U3869 (N_3869,N_673,N_477);
or U3870 (N_3870,N_2140,N_696);
nand U3871 (N_3871,N_1280,N_2473);
nand U3872 (N_3872,N_268,N_1698);
nor U3873 (N_3873,N_1783,N_1712);
or U3874 (N_3874,N_1518,N_1273);
or U3875 (N_3875,N_2291,N_1861);
and U3876 (N_3876,N_133,N_1378);
or U3877 (N_3877,N_757,N_1300);
or U3878 (N_3878,N_966,N_2472);
nand U3879 (N_3879,N_523,N_484);
or U3880 (N_3880,N_620,N_2323);
nor U3881 (N_3881,N_692,N_1125);
xnor U3882 (N_3882,N_2040,N_1718);
and U3883 (N_3883,N_1406,N_1630);
xor U3884 (N_3884,N_72,N_2245);
nor U3885 (N_3885,N_701,N_735);
nor U3886 (N_3886,N_493,N_1520);
nand U3887 (N_3887,N_1877,N_1058);
xor U3888 (N_3888,N_1127,N_624);
xor U3889 (N_3889,N_1569,N_1037);
and U3890 (N_3890,N_996,N_1700);
xor U3891 (N_3891,N_1700,N_1359);
and U3892 (N_3892,N_2364,N_2363);
nand U3893 (N_3893,N_2307,N_35);
xor U3894 (N_3894,N_2307,N_1266);
xor U3895 (N_3895,N_577,N_1088);
and U3896 (N_3896,N_1103,N_1021);
or U3897 (N_3897,N_2272,N_2073);
or U3898 (N_3898,N_555,N_212);
xnor U3899 (N_3899,N_1989,N_1691);
nor U3900 (N_3900,N_213,N_335);
xnor U3901 (N_3901,N_1775,N_1288);
or U3902 (N_3902,N_5,N_1598);
nand U3903 (N_3903,N_701,N_960);
xor U3904 (N_3904,N_702,N_2397);
and U3905 (N_3905,N_2165,N_392);
and U3906 (N_3906,N_60,N_2283);
or U3907 (N_3907,N_1369,N_2271);
xnor U3908 (N_3908,N_680,N_857);
or U3909 (N_3909,N_1424,N_1146);
nand U3910 (N_3910,N_2373,N_846);
xnor U3911 (N_3911,N_1160,N_1043);
nand U3912 (N_3912,N_959,N_1685);
nor U3913 (N_3913,N_2388,N_1964);
xor U3914 (N_3914,N_1576,N_1114);
or U3915 (N_3915,N_1430,N_1440);
or U3916 (N_3916,N_2411,N_1736);
nor U3917 (N_3917,N_1996,N_1700);
or U3918 (N_3918,N_919,N_72);
xor U3919 (N_3919,N_173,N_1059);
nor U3920 (N_3920,N_1525,N_863);
xor U3921 (N_3921,N_1115,N_115);
nor U3922 (N_3922,N_2136,N_432);
nand U3923 (N_3923,N_1526,N_640);
or U3924 (N_3924,N_1293,N_622);
or U3925 (N_3925,N_1825,N_1184);
xor U3926 (N_3926,N_2309,N_2297);
xor U3927 (N_3927,N_1027,N_925);
or U3928 (N_3928,N_1022,N_279);
and U3929 (N_3929,N_116,N_713);
nand U3930 (N_3930,N_1970,N_2419);
nor U3931 (N_3931,N_1086,N_1004);
nand U3932 (N_3932,N_656,N_238);
nand U3933 (N_3933,N_1043,N_2258);
or U3934 (N_3934,N_677,N_640);
xnor U3935 (N_3935,N_176,N_731);
nand U3936 (N_3936,N_926,N_2242);
nand U3937 (N_3937,N_311,N_2078);
xnor U3938 (N_3938,N_2308,N_511);
nor U3939 (N_3939,N_2061,N_1352);
and U3940 (N_3940,N_2121,N_1850);
nor U3941 (N_3941,N_195,N_1672);
nand U3942 (N_3942,N_1152,N_704);
nor U3943 (N_3943,N_289,N_2264);
and U3944 (N_3944,N_1006,N_1348);
and U3945 (N_3945,N_2083,N_2274);
nor U3946 (N_3946,N_1549,N_1876);
nor U3947 (N_3947,N_1413,N_741);
nand U3948 (N_3948,N_1563,N_1652);
or U3949 (N_3949,N_1472,N_1735);
nor U3950 (N_3950,N_471,N_30);
or U3951 (N_3951,N_1252,N_594);
xor U3952 (N_3952,N_2127,N_1954);
nor U3953 (N_3953,N_488,N_1573);
xnor U3954 (N_3954,N_2393,N_2021);
nand U3955 (N_3955,N_153,N_1258);
xnor U3956 (N_3956,N_2213,N_2381);
and U3957 (N_3957,N_1576,N_1266);
nand U3958 (N_3958,N_2076,N_1416);
xnor U3959 (N_3959,N_207,N_763);
xor U3960 (N_3960,N_781,N_787);
xnor U3961 (N_3961,N_447,N_1205);
xor U3962 (N_3962,N_1877,N_2250);
and U3963 (N_3963,N_422,N_798);
nand U3964 (N_3964,N_2318,N_1022);
nand U3965 (N_3965,N_763,N_1149);
nand U3966 (N_3966,N_2453,N_688);
and U3967 (N_3967,N_198,N_1090);
nor U3968 (N_3968,N_281,N_1486);
and U3969 (N_3969,N_2125,N_1059);
nand U3970 (N_3970,N_1370,N_1196);
xnor U3971 (N_3971,N_201,N_64);
nand U3972 (N_3972,N_1992,N_48);
nor U3973 (N_3973,N_1567,N_567);
nor U3974 (N_3974,N_1744,N_2245);
nand U3975 (N_3975,N_261,N_2000);
nor U3976 (N_3976,N_1696,N_2124);
nor U3977 (N_3977,N_1935,N_1481);
nor U3978 (N_3978,N_219,N_130);
or U3979 (N_3979,N_1535,N_644);
xnor U3980 (N_3980,N_240,N_309);
and U3981 (N_3981,N_2485,N_1676);
xnor U3982 (N_3982,N_1038,N_977);
or U3983 (N_3983,N_1904,N_551);
nand U3984 (N_3984,N_350,N_592);
or U3985 (N_3985,N_1559,N_1335);
xor U3986 (N_3986,N_57,N_1359);
xnor U3987 (N_3987,N_231,N_73);
nor U3988 (N_3988,N_2392,N_1224);
nor U3989 (N_3989,N_2028,N_832);
and U3990 (N_3990,N_1218,N_1581);
xnor U3991 (N_3991,N_2167,N_1262);
or U3992 (N_3992,N_2171,N_20);
xnor U3993 (N_3993,N_22,N_1308);
xor U3994 (N_3994,N_1337,N_661);
or U3995 (N_3995,N_788,N_1089);
nor U3996 (N_3996,N_482,N_238);
or U3997 (N_3997,N_968,N_2211);
and U3998 (N_3998,N_650,N_997);
and U3999 (N_3999,N_172,N_643);
nor U4000 (N_4000,N_273,N_146);
xnor U4001 (N_4001,N_744,N_181);
nand U4002 (N_4002,N_480,N_53);
nor U4003 (N_4003,N_2151,N_1349);
or U4004 (N_4004,N_1735,N_28);
xor U4005 (N_4005,N_625,N_1562);
nand U4006 (N_4006,N_1752,N_183);
or U4007 (N_4007,N_437,N_1060);
nor U4008 (N_4008,N_938,N_1436);
xnor U4009 (N_4009,N_581,N_1807);
and U4010 (N_4010,N_2268,N_2108);
nor U4011 (N_4011,N_1009,N_1104);
xnor U4012 (N_4012,N_1378,N_330);
and U4013 (N_4013,N_1840,N_2457);
nor U4014 (N_4014,N_688,N_1480);
xor U4015 (N_4015,N_333,N_1327);
or U4016 (N_4016,N_909,N_1039);
or U4017 (N_4017,N_1109,N_2409);
or U4018 (N_4018,N_2448,N_1549);
xnor U4019 (N_4019,N_2146,N_1149);
nor U4020 (N_4020,N_1304,N_1338);
nor U4021 (N_4021,N_1287,N_1695);
nor U4022 (N_4022,N_1337,N_607);
nand U4023 (N_4023,N_832,N_2238);
nor U4024 (N_4024,N_1139,N_147);
nor U4025 (N_4025,N_1994,N_1180);
xnor U4026 (N_4026,N_372,N_2118);
and U4027 (N_4027,N_743,N_1619);
and U4028 (N_4028,N_641,N_2234);
xor U4029 (N_4029,N_2495,N_914);
or U4030 (N_4030,N_1819,N_732);
xor U4031 (N_4031,N_543,N_2115);
xor U4032 (N_4032,N_12,N_1104);
and U4033 (N_4033,N_181,N_290);
or U4034 (N_4034,N_1454,N_2175);
nor U4035 (N_4035,N_1519,N_804);
xnor U4036 (N_4036,N_1257,N_103);
or U4037 (N_4037,N_277,N_928);
nor U4038 (N_4038,N_1819,N_1757);
xor U4039 (N_4039,N_536,N_993);
nor U4040 (N_4040,N_2299,N_1851);
nor U4041 (N_4041,N_1641,N_1935);
xor U4042 (N_4042,N_1289,N_2035);
nand U4043 (N_4043,N_1593,N_209);
nor U4044 (N_4044,N_671,N_1214);
nor U4045 (N_4045,N_540,N_1637);
nand U4046 (N_4046,N_2123,N_99);
or U4047 (N_4047,N_2254,N_1454);
nand U4048 (N_4048,N_89,N_1038);
nand U4049 (N_4049,N_1105,N_1995);
nand U4050 (N_4050,N_2397,N_2047);
nand U4051 (N_4051,N_870,N_1074);
and U4052 (N_4052,N_2469,N_993);
or U4053 (N_4053,N_1990,N_354);
nand U4054 (N_4054,N_2209,N_1038);
or U4055 (N_4055,N_1202,N_412);
nand U4056 (N_4056,N_802,N_2345);
nor U4057 (N_4057,N_1009,N_556);
and U4058 (N_4058,N_2280,N_2198);
nand U4059 (N_4059,N_2100,N_932);
or U4060 (N_4060,N_1057,N_1428);
nor U4061 (N_4061,N_263,N_2293);
and U4062 (N_4062,N_1465,N_2115);
xnor U4063 (N_4063,N_1305,N_725);
and U4064 (N_4064,N_519,N_693);
and U4065 (N_4065,N_213,N_1205);
and U4066 (N_4066,N_2307,N_1551);
xor U4067 (N_4067,N_817,N_1672);
and U4068 (N_4068,N_561,N_1490);
nor U4069 (N_4069,N_400,N_892);
and U4070 (N_4070,N_370,N_1829);
nand U4071 (N_4071,N_2468,N_1537);
nand U4072 (N_4072,N_1286,N_1200);
or U4073 (N_4073,N_412,N_1948);
xor U4074 (N_4074,N_181,N_1828);
xor U4075 (N_4075,N_1796,N_2412);
nor U4076 (N_4076,N_1473,N_2119);
nor U4077 (N_4077,N_955,N_2088);
or U4078 (N_4078,N_2030,N_1123);
or U4079 (N_4079,N_1280,N_1811);
nand U4080 (N_4080,N_1189,N_466);
or U4081 (N_4081,N_1947,N_685);
nand U4082 (N_4082,N_627,N_1708);
or U4083 (N_4083,N_1600,N_991);
nor U4084 (N_4084,N_663,N_1971);
nand U4085 (N_4085,N_2222,N_2346);
or U4086 (N_4086,N_1503,N_940);
nor U4087 (N_4087,N_2490,N_436);
xor U4088 (N_4088,N_1626,N_1231);
xnor U4089 (N_4089,N_654,N_1462);
nand U4090 (N_4090,N_1663,N_1612);
nor U4091 (N_4091,N_2151,N_774);
nor U4092 (N_4092,N_1602,N_290);
and U4093 (N_4093,N_1203,N_1337);
and U4094 (N_4094,N_543,N_1184);
or U4095 (N_4095,N_2102,N_1063);
and U4096 (N_4096,N_325,N_1221);
xnor U4097 (N_4097,N_1876,N_2257);
and U4098 (N_4098,N_1516,N_1266);
xnor U4099 (N_4099,N_2170,N_498);
and U4100 (N_4100,N_1054,N_1435);
and U4101 (N_4101,N_2177,N_968);
xor U4102 (N_4102,N_908,N_1163);
and U4103 (N_4103,N_824,N_1056);
and U4104 (N_4104,N_2368,N_1376);
nor U4105 (N_4105,N_218,N_2072);
xor U4106 (N_4106,N_5,N_2009);
and U4107 (N_4107,N_516,N_685);
xor U4108 (N_4108,N_1984,N_687);
or U4109 (N_4109,N_530,N_1439);
or U4110 (N_4110,N_2404,N_1343);
xnor U4111 (N_4111,N_607,N_2053);
or U4112 (N_4112,N_1244,N_1035);
and U4113 (N_4113,N_1189,N_100);
and U4114 (N_4114,N_1378,N_1458);
and U4115 (N_4115,N_1069,N_510);
nand U4116 (N_4116,N_602,N_1140);
and U4117 (N_4117,N_2194,N_669);
nor U4118 (N_4118,N_2263,N_477);
xnor U4119 (N_4119,N_2202,N_1615);
and U4120 (N_4120,N_710,N_1750);
xor U4121 (N_4121,N_2214,N_861);
or U4122 (N_4122,N_1713,N_1536);
xor U4123 (N_4123,N_810,N_2417);
nand U4124 (N_4124,N_1508,N_1504);
nand U4125 (N_4125,N_427,N_63);
nor U4126 (N_4126,N_307,N_827);
xnor U4127 (N_4127,N_1478,N_428);
or U4128 (N_4128,N_2361,N_1117);
nand U4129 (N_4129,N_563,N_390);
nand U4130 (N_4130,N_196,N_331);
nor U4131 (N_4131,N_668,N_1918);
nand U4132 (N_4132,N_144,N_1133);
nor U4133 (N_4133,N_2256,N_1522);
xnor U4134 (N_4134,N_1868,N_527);
and U4135 (N_4135,N_2003,N_270);
xor U4136 (N_4136,N_695,N_237);
and U4137 (N_4137,N_309,N_1342);
xor U4138 (N_4138,N_2387,N_1989);
nand U4139 (N_4139,N_637,N_745);
nand U4140 (N_4140,N_2208,N_263);
and U4141 (N_4141,N_280,N_948);
xnor U4142 (N_4142,N_1451,N_161);
nand U4143 (N_4143,N_757,N_1616);
nor U4144 (N_4144,N_120,N_147);
xor U4145 (N_4145,N_1890,N_810);
and U4146 (N_4146,N_2174,N_1991);
xnor U4147 (N_4147,N_2063,N_42);
nand U4148 (N_4148,N_1261,N_2055);
nand U4149 (N_4149,N_979,N_1228);
nand U4150 (N_4150,N_84,N_1365);
nand U4151 (N_4151,N_26,N_2024);
nor U4152 (N_4152,N_617,N_1088);
and U4153 (N_4153,N_222,N_12);
or U4154 (N_4154,N_614,N_959);
nand U4155 (N_4155,N_1767,N_2298);
or U4156 (N_4156,N_1464,N_498);
and U4157 (N_4157,N_550,N_1906);
nor U4158 (N_4158,N_884,N_1585);
nor U4159 (N_4159,N_1337,N_663);
or U4160 (N_4160,N_548,N_282);
nor U4161 (N_4161,N_366,N_530);
nor U4162 (N_4162,N_1143,N_1038);
xor U4163 (N_4163,N_694,N_2040);
nand U4164 (N_4164,N_578,N_1647);
nor U4165 (N_4165,N_396,N_631);
or U4166 (N_4166,N_2413,N_666);
or U4167 (N_4167,N_844,N_184);
or U4168 (N_4168,N_375,N_2196);
or U4169 (N_4169,N_1157,N_1595);
and U4170 (N_4170,N_1161,N_643);
or U4171 (N_4171,N_2330,N_592);
nand U4172 (N_4172,N_951,N_1054);
nor U4173 (N_4173,N_2370,N_1715);
nor U4174 (N_4174,N_854,N_690);
and U4175 (N_4175,N_2235,N_857);
or U4176 (N_4176,N_1833,N_1526);
or U4177 (N_4177,N_522,N_1791);
xnor U4178 (N_4178,N_190,N_87);
nor U4179 (N_4179,N_1762,N_270);
or U4180 (N_4180,N_1343,N_915);
nor U4181 (N_4181,N_1456,N_1524);
xor U4182 (N_4182,N_574,N_373);
or U4183 (N_4183,N_66,N_1042);
and U4184 (N_4184,N_2001,N_2457);
and U4185 (N_4185,N_1414,N_1652);
nor U4186 (N_4186,N_2116,N_963);
and U4187 (N_4187,N_443,N_1533);
and U4188 (N_4188,N_924,N_2024);
xor U4189 (N_4189,N_1179,N_1002);
nand U4190 (N_4190,N_2445,N_1215);
and U4191 (N_4191,N_2288,N_616);
nor U4192 (N_4192,N_123,N_430);
xnor U4193 (N_4193,N_233,N_561);
xor U4194 (N_4194,N_2452,N_451);
or U4195 (N_4195,N_1399,N_263);
nand U4196 (N_4196,N_506,N_2107);
xnor U4197 (N_4197,N_1295,N_2466);
xor U4198 (N_4198,N_1002,N_124);
xnor U4199 (N_4199,N_2397,N_1093);
nor U4200 (N_4200,N_742,N_1033);
nor U4201 (N_4201,N_1826,N_1751);
nor U4202 (N_4202,N_2092,N_1788);
and U4203 (N_4203,N_214,N_1423);
nor U4204 (N_4204,N_2289,N_593);
or U4205 (N_4205,N_1807,N_2427);
nand U4206 (N_4206,N_1343,N_2191);
and U4207 (N_4207,N_1311,N_1082);
nand U4208 (N_4208,N_1031,N_1447);
nand U4209 (N_4209,N_1025,N_456);
and U4210 (N_4210,N_1682,N_502);
and U4211 (N_4211,N_326,N_1480);
or U4212 (N_4212,N_1301,N_931);
or U4213 (N_4213,N_2304,N_1127);
xnor U4214 (N_4214,N_488,N_1887);
xor U4215 (N_4215,N_1409,N_1716);
and U4216 (N_4216,N_1956,N_783);
or U4217 (N_4217,N_1613,N_1856);
nor U4218 (N_4218,N_960,N_349);
or U4219 (N_4219,N_1886,N_137);
nand U4220 (N_4220,N_2194,N_492);
nor U4221 (N_4221,N_430,N_1305);
nor U4222 (N_4222,N_2440,N_905);
or U4223 (N_4223,N_2318,N_415);
and U4224 (N_4224,N_2033,N_1904);
or U4225 (N_4225,N_1281,N_311);
or U4226 (N_4226,N_1723,N_840);
xor U4227 (N_4227,N_666,N_550);
nand U4228 (N_4228,N_2432,N_856);
nand U4229 (N_4229,N_310,N_79);
xnor U4230 (N_4230,N_1385,N_2269);
nor U4231 (N_4231,N_2190,N_1542);
and U4232 (N_4232,N_2295,N_185);
nand U4233 (N_4233,N_77,N_714);
xnor U4234 (N_4234,N_1297,N_135);
or U4235 (N_4235,N_844,N_1333);
xor U4236 (N_4236,N_218,N_2324);
xnor U4237 (N_4237,N_2134,N_1058);
xnor U4238 (N_4238,N_2427,N_459);
or U4239 (N_4239,N_112,N_2210);
or U4240 (N_4240,N_1269,N_1239);
or U4241 (N_4241,N_980,N_2479);
nor U4242 (N_4242,N_2058,N_1372);
xnor U4243 (N_4243,N_2000,N_2058);
or U4244 (N_4244,N_256,N_2222);
nor U4245 (N_4245,N_885,N_2369);
and U4246 (N_4246,N_2156,N_1656);
nor U4247 (N_4247,N_597,N_1665);
nand U4248 (N_4248,N_2238,N_300);
nor U4249 (N_4249,N_1451,N_1947);
nand U4250 (N_4250,N_1955,N_1206);
and U4251 (N_4251,N_817,N_2142);
and U4252 (N_4252,N_1590,N_568);
xor U4253 (N_4253,N_252,N_613);
nor U4254 (N_4254,N_380,N_2050);
or U4255 (N_4255,N_1511,N_1661);
and U4256 (N_4256,N_359,N_934);
nand U4257 (N_4257,N_1966,N_1913);
nor U4258 (N_4258,N_1151,N_612);
nor U4259 (N_4259,N_787,N_81);
nand U4260 (N_4260,N_437,N_796);
or U4261 (N_4261,N_2013,N_1544);
xor U4262 (N_4262,N_1229,N_274);
nand U4263 (N_4263,N_623,N_73);
xor U4264 (N_4264,N_2343,N_2016);
or U4265 (N_4265,N_742,N_540);
xor U4266 (N_4266,N_1794,N_643);
nor U4267 (N_4267,N_2318,N_797);
and U4268 (N_4268,N_112,N_670);
or U4269 (N_4269,N_1258,N_2179);
and U4270 (N_4270,N_2110,N_915);
nor U4271 (N_4271,N_2243,N_974);
nand U4272 (N_4272,N_945,N_871);
or U4273 (N_4273,N_1129,N_932);
or U4274 (N_4274,N_534,N_91);
nor U4275 (N_4275,N_2143,N_1854);
and U4276 (N_4276,N_1374,N_512);
or U4277 (N_4277,N_1438,N_616);
nand U4278 (N_4278,N_338,N_1157);
and U4279 (N_4279,N_1899,N_60);
or U4280 (N_4280,N_1098,N_1628);
xnor U4281 (N_4281,N_1122,N_30);
nand U4282 (N_4282,N_1431,N_2314);
nor U4283 (N_4283,N_343,N_1512);
nand U4284 (N_4284,N_73,N_1717);
nand U4285 (N_4285,N_2272,N_802);
nor U4286 (N_4286,N_536,N_1180);
xnor U4287 (N_4287,N_1666,N_2218);
nor U4288 (N_4288,N_1723,N_160);
nor U4289 (N_4289,N_1608,N_1808);
xnor U4290 (N_4290,N_810,N_1706);
nor U4291 (N_4291,N_1736,N_1094);
and U4292 (N_4292,N_965,N_2247);
nand U4293 (N_4293,N_716,N_520);
or U4294 (N_4294,N_1231,N_1340);
nor U4295 (N_4295,N_1085,N_603);
xor U4296 (N_4296,N_1001,N_1442);
or U4297 (N_4297,N_649,N_1119);
nand U4298 (N_4298,N_1139,N_225);
nand U4299 (N_4299,N_463,N_1153);
nand U4300 (N_4300,N_1046,N_724);
nand U4301 (N_4301,N_1328,N_2020);
nor U4302 (N_4302,N_1812,N_258);
xnor U4303 (N_4303,N_428,N_1004);
or U4304 (N_4304,N_1744,N_826);
xor U4305 (N_4305,N_2288,N_1462);
and U4306 (N_4306,N_966,N_1748);
and U4307 (N_4307,N_2392,N_1629);
nor U4308 (N_4308,N_871,N_2329);
and U4309 (N_4309,N_940,N_1318);
xor U4310 (N_4310,N_1186,N_1021);
nand U4311 (N_4311,N_1105,N_1814);
nand U4312 (N_4312,N_1999,N_454);
nand U4313 (N_4313,N_374,N_2151);
and U4314 (N_4314,N_1728,N_2467);
xor U4315 (N_4315,N_922,N_1121);
or U4316 (N_4316,N_989,N_1415);
or U4317 (N_4317,N_1388,N_1619);
and U4318 (N_4318,N_2262,N_2243);
xor U4319 (N_4319,N_231,N_383);
and U4320 (N_4320,N_1682,N_1336);
xnor U4321 (N_4321,N_1633,N_2385);
or U4322 (N_4322,N_1841,N_1439);
nor U4323 (N_4323,N_155,N_2315);
or U4324 (N_4324,N_2292,N_1897);
and U4325 (N_4325,N_2138,N_1550);
xor U4326 (N_4326,N_332,N_831);
and U4327 (N_4327,N_390,N_1438);
or U4328 (N_4328,N_1260,N_512);
and U4329 (N_4329,N_1236,N_1696);
nand U4330 (N_4330,N_758,N_1996);
xor U4331 (N_4331,N_414,N_2097);
and U4332 (N_4332,N_2187,N_432);
xnor U4333 (N_4333,N_131,N_870);
nand U4334 (N_4334,N_1609,N_737);
nand U4335 (N_4335,N_1042,N_1383);
or U4336 (N_4336,N_2173,N_1298);
nand U4337 (N_4337,N_2007,N_2160);
or U4338 (N_4338,N_1128,N_2049);
nor U4339 (N_4339,N_1020,N_746);
nor U4340 (N_4340,N_395,N_2144);
nor U4341 (N_4341,N_1885,N_1189);
xnor U4342 (N_4342,N_1772,N_1795);
nand U4343 (N_4343,N_2440,N_768);
xor U4344 (N_4344,N_1508,N_720);
nor U4345 (N_4345,N_649,N_1954);
xor U4346 (N_4346,N_1556,N_1424);
or U4347 (N_4347,N_540,N_756);
nand U4348 (N_4348,N_1867,N_2298);
or U4349 (N_4349,N_680,N_1290);
nor U4350 (N_4350,N_2497,N_263);
and U4351 (N_4351,N_2083,N_1835);
and U4352 (N_4352,N_2325,N_2094);
xnor U4353 (N_4353,N_625,N_1785);
and U4354 (N_4354,N_2271,N_1317);
nor U4355 (N_4355,N_2499,N_1399);
nor U4356 (N_4356,N_1489,N_278);
nand U4357 (N_4357,N_1863,N_1073);
nand U4358 (N_4358,N_276,N_705);
nor U4359 (N_4359,N_921,N_1446);
xnor U4360 (N_4360,N_2323,N_437);
or U4361 (N_4361,N_234,N_357);
nand U4362 (N_4362,N_329,N_1156);
xor U4363 (N_4363,N_1428,N_2227);
or U4364 (N_4364,N_1451,N_986);
xor U4365 (N_4365,N_425,N_1881);
or U4366 (N_4366,N_636,N_1223);
and U4367 (N_4367,N_1538,N_1363);
nor U4368 (N_4368,N_2041,N_1149);
and U4369 (N_4369,N_2384,N_2475);
xnor U4370 (N_4370,N_2085,N_2);
or U4371 (N_4371,N_1927,N_1239);
nor U4372 (N_4372,N_1577,N_2270);
xor U4373 (N_4373,N_99,N_1501);
nand U4374 (N_4374,N_2294,N_1261);
xnor U4375 (N_4375,N_32,N_600);
or U4376 (N_4376,N_2367,N_2273);
nor U4377 (N_4377,N_1910,N_2266);
nand U4378 (N_4378,N_934,N_1739);
nor U4379 (N_4379,N_996,N_726);
nand U4380 (N_4380,N_45,N_2248);
xor U4381 (N_4381,N_166,N_641);
nand U4382 (N_4382,N_1691,N_1659);
xor U4383 (N_4383,N_1259,N_1555);
nand U4384 (N_4384,N_1092,N_2462);
and U4385 (N_4385,N_495,N_1182);
or U4386 (N_4386,N_2212,N_1984);
and U4387 (N_4387,N_171,N_478);
xnor U4388 (N_4388,N_92,N_888);
nand U4389 (N_4389,N_1165,N_1154);
and U4390 (N_4390,N_2268,N_224);
or U4391 (N_4391,N_1644,N_2283);
nor U4392 (N_4392,N_1074,N_971);
nor U4393 (N_4393,N_2269,N_1021);
nand U4394 (N_4394,N_1918,N_224);
nor U4395 (N_4395,N_1488,N_309);
nand U4396 (N_4396,N_456,N_2478);
nand U4397 (N_4397,N_1521,N_1505);
nand U4398 (N_4398,N_2497,N_1489);
nor U4399 (N_4399,N_102,N_1474);
nor U4400 (N_4400,N_257,N_1499);
nand U4401 (N_4401,N_2073,N_883);
xnor U4402 (N_4402,N_890,N_1066);
nand U4403 (N_4403,N_2085,N_486);
and U4404 (N_4404,N_1557,N_1142);
xor U4405 (N_4405,N_800,N_2478);
nor U4406 (N_4406,N_2362,N_1000);
nor U4407 (N_4407,N_368,N_507);
nand U4408 (N_4408,N_555,N_575);
nor U4409 (N_4409,N_2471,N_1523);
nor U4410 (N_4410,N_1291,N_2080);
nand U4411 (N_4411,N_944,N_2362);
xor U4412 (N_4412,N_524,N_69);
nor U4413 (N_4413,N_670,N_755);
xor U4414 (N_4414,N_1203,N_103);
nand U4415 (N_4415,N_1267,N_931);
and U4416 (N_4416,N_200,N_1747);
and U4417 (N_4417,N_2091,N_432);
nand U4418 (N_4418,N_1342,N_1042);
or U4419 (N_4419,N_207,N_31);
nor U4420 (N_4420,N_336,N_633);
nor U4421 (N_4421,N_604,N_2229);
nor U4422 (N_4422,N_1092,N_1809);
nor U4423 (N_4423,N_931,N_244);
nand U4424 (N_4424,N_917,N_2015);
or U4425 (N_4425,N_1440,N_442);
nand U4426 (N_4426,N_1822,N_816);
or U4427 (N_4427,N_2025,N_1507);
and U4428 (N_4428,N_2047,N_563);
or U4429 (N_4429,N_1533,N_2141);
and U4430 (N_4430,N_1110,N_1109);
nand U4431 (N_4431,N_1797,N_1422);
nor U4432 (N_4432,N_37,N_1656);
or U4433 (N_4433,N_458,N_541);
or U4434 (N_4434,N_1470,N_185);
or U4435 (N_4435,N_1085,N_438);
nor U4436 (N_4436,N_2013,N_2278);
nor U4437 (N_4437,N_1773,N_448);
nor U4438 (N_4438,N_1271,N_1370);
xor U4439 (N_4439,N_2491,N_1986);
or U4440 (N_4440,N_1864,N_592);
nand U4441 (N_4441,N_571,N_293);
xor U4442 (N_4442,N_769,N_936);
nand U4443 (N_4443,N_1340,N_109);
and U4444 (N_4444,N_1213,N_1488);
xor U4445 (N_4445,N_1951,N_601);
nor U4446 (N_4446,N_892,N_2459);
and U4447 (N_4447,N_746,N_76);
nor U4448 (N_4448,N_1639,N_1287);
xnor U4449 (N_4449,N_1197,N_1333);
and U4450 (N_4450,N_105,N_369);
nand U4451 (N_4451,N_2432,N_143);
nand U4452 (N_4452,N_2242,N_498);
nand U4453 (N_4453,N_741,N_560);
nor U4454 (N_4454,N_395,N_1171);
xnor U4455 (N_4455,N_1310,N_155);
nand U4456 (N_4456,N_2311,N_2313);
nor U4457 (N_4457,N_354,N_525);
nor U4458 (N_4458,N_727,N_2318);
nor U4459 (N_4459,N_1007,N_864);
nand U4460 (N_4460,N_1469,N_1831);
or U4461 (N_4461,N_1138,N_1904);
nor U4462 (N_4462,N_1500,N_976);
nor U4463 (N_4463,N_1415,N_1866);
nor U4464 (N_4464,N_2027,N_1918);
or U4465 (N_4465,N_1032,N_2099);
xnor U4466 (N_4466,N_795,N_2427);
xnor U4467 (N_4467,N_1397,N_2261);
nand U4468 (N_4468,N_574,N_2459);
nor U4469 (N_4469,N_1016,N_1529);
or U4470 (N_4470,N_2292,N_139);
nor U4471 (N_4471,N_355,N_36);
nor U4472 (N_4472,N_1556,N_889);
xnor U4473 (N_4473,N_383,N_792);
nand U4474 (N_4474,N_1661,N_1208);
xor U4475 (N_4475,N_1395,N_621);
nand U4476 (N_4476,N_867,N_36);
xnor U4477 (N_4477,N_365,N_571);
nor U4478 (N_4478,N_1649,N_2457);
xor U4479 (N_4479,N_735,N_817);
nor U4480 (N_4480,N_2421,N_1311);
xor U4481 (N_4481,N_536,N_345);
nand U4482 (N_4482,N_1809,N_1169);
nand U4483 (N_4483,N_1774,N_2200);
and U4484 (N_4484,N_58,N_1701);
xnor U4485 (N_4485,N_416,N_1353);
and U4486 (N_4486,N_616,N_1119);
nor U4487 (N_4487,N_172,N_1463);
nand U4488 (N_4488,N_1202,N_1892);
or U4489 (N_4489,N_1296,N_657);
nor U4490 (N_4490,N_2139,N_1897);
and U4491 (N_4491,N_2162,N_1296);
xnor U4492 (N_4492,N_879,N_2089);
or U4493 (N_4493,N_2370,N_458);
nand U4494 (N_4494,N_2343,N_584);
or U4495 (N_4495,N_2310,N_1650);
nand U4496 (N_4496,N_2235,N_1466);
nor U4497 (N_4497,N_1667,N_2245);
and U4498 (N_4498,N_1073,N_2337);
nand U4499 (N_4499,N_2092,N_665);
nor U4500 (N_4500,N_2408,N_230);
nand U4501 (N_4501,N_1718,N_154);
nand U4502 (N_4502,N_1433,N_446);
or U4503 (N_4503,N_230,N_309);
nand U4504 (N_4504,N_486,N_37);
nor U4505 (N_4505,N_2114,N_827);
xnor U4506 (N_4506,N_1116,N_555);
nor U4507 (N_4507,N_27,N_229);
xor U4508 (N_4508,N_1834,N_1918);
nand U4509 (N_4509,N_1412,N_1373);
or U4510 (N_4510,N_882,N_1232);
xor U4511 (N_4511,N_2231,N_1770);
xnor U4512 (N_4512,N_2240,N_2484);
or U4513 (N_4513,N_176,N_1393);
nor U4514 (N_4514,N_1336,N_1362);
nor U4515 (N_4515,N_2367,N_2198);
or U4516 (N_4516,N_1746,N_1991);
nand U4517 (N_4517,N_1556,N_1490);
xor U4518 (N_4518,N_1767,N_591);
or U4519 (N_4519,N_2170,N_1661);
nor U4520 (N_4520,N_338,N_61);
and U4521 (N_4521,N_1761,N_1113);
nor U4522 (N_4522,N_1812,N_1204);
nand U4523 (N_4523,N_1219,N_684);
or U4524 (N_4524,N_2284,N_895);
and U4525 (N_4525,N_1372,N_77);
and U4526 (N_4526,N_1337,N_1190);
nand U4527 (N_4527,N_358,N_1631);
nor U4528 (N_4528,N_1936,N_115);
or U4529 (N_4529,N_594,N_779);
and U4530 (N_4530,N_205,N_951);
nand U4531 (N_4531,N_2266,N_108);
nor U4532 (N_4532,N_2164,N_1083);
nand U4533 (N_4533,N_2169,N_1989);
or U4534 (N_4534,N_2306,N_844);
xor U4535 (N_4535,N_2144,N_1869);
nor U4536 (N_4536,N_685,N_1880);
nand U4537 (N_4537,N_1588,N_2124);
nor U4538 (N_4538,N_1705,N_2252);
nand U4539 (N_4539,N_876,N_1860);
or U4540 (N_4540,N_2138,N_870);
and U4541 (N_4541,N_966,N_667);
xnor U4542 (N_4542,N_2229,N_1355);
nand U4543 (N_4543,N_1625,N_1694);
and U4544 (N_4544,N_1189,N_2216);
and U4545 (N_4545,N_2379,N_81);
or U4546 (N_4546,N_1637,N_1314);
nand U4547 (N_4547,N_437,N_667);
and U4548 (N_4548,N_199,N_20);
or U4549 (N_4549,N_2359,N_346);
and U4550 (N_4550,N_300,N_703);
or U4551 (N_4551,N_2007,N_1011);
nand U4552 (N_4552,N_2345,N_1279);
nor U4553 (N_4553,N_1254,N_996);
and U4554 (N_4554,N_2262,N_1757);
or U4555 (N_4555,N_146,N_1116);
nor U4556 (N_4556,N_294,N_1226);
xor U4557 (N_4557,N_2142,N_806);
or U4558 (N_4558,N_2165,N_332);
nand U4559 (N_4559,N_2330,N_1477);
and U4560 (N_4560,N_2343,N_1498);
xor U4561 (N_4561,N_665,N_1918);
xnor U4562 (N_4562,N_1097,N_382);
xnor U4563 (N_4563,N_1791,N_1447);
or U4564 (N_4564,N_1222,N_87);
or U4565 (N_4565,N_858,N_2098);
and U4566 (N_4566,N_1047,N_228);
nand U4567 (N_4567,N_354,N_1992);
or U4568 (N_4568,N_187,N_1548);
xor U4569 (N_4569,N_1189,N_2095);
nor U4570 (N_4570,N_192,N_1876);
xnor U4571 (N_4571,N_1891,N_1254);
nor U4572 (N_4572,N_639,N_1531);
xnor U4573 (N_4573,N_2355,N_1735);
xnor U4574 (N_4574,N_843,N_44);
or U4575 (N_4575,N_820,N_621);
xnor U4576 (N_4576,N_1960,N_482);
and U4577 (N_4577,N_814,N_1715);
and U4578 (N_4578,N_588,N_469);
and U4579 (N_4579,N_1181,N_2211);
and U4580 (N_4580,N_1333,N_1626);
xnor U4581 (N_4581,N_2211,N_262);
and U4582 (N_4582,N_1890,N_431);
and U4583 (N_4583,N_694,N_2476);
and U4584 (N_4584,N_1459,N_1787);
nand U4585 (N_4585,N_1642,N_2479);
xor U4586 (N_4586,N_505,N_598);
nand U4587 (N_4587,N_17,N_267);
nand U4588 (N_4588,N_2020,N_898);
xor U4589 (N_4589,N_1626,N_2106);
nand U4590 (N_4590,N_2072,N_1034);
nand U4591 (N_4591,N_996,N_421);
nand U4592 (N_4592,N_1279,N_2460);
nor U4593 (N_4593,N_1576,N_2218);
xnor U4594 (N_4594,N_2,N_558);
or U4595 (N_4595,N_314,N_134);
nor U4596 (N_4596,N_1474,N_970);
nand U4597 (N_4597,N_2242,N_1278);
and U4598 (N_4598,N_1279,N_76);
nand U4599 (N_4599,N_237,N_1602);
nand U4600 (N_4600,N_274,N_871);
nor U4601 (N_4601,N_431,N_1702);
xor U4602 (N_4602,N_1726,N_187);
and U4603 (N_4603,N_2216,N_2150);
and U4604 (N_4604,N_979,N_2296);
nor U4605 (N_4605,N_1808,N_11);
and U4606 (N_4606,N_804,N_253);
or U4607 (N_4607,N_1208,N_2356);
or U4608 (N_4608,N_2254,N_2434);
nand U4609 (N_4609,N_453,N_2223);
nand U4610 (N_4610,N_323,N_204);
nor U4611 (N_4611,N_818,N_1177);
and U4612 (N_4612,N_1847,N_1326);
nand U4613 (N_4613,N_2330,N_114);
or U4614 (N_4614,N_1504,N_329);
and U4615 (N_4615,N_1728,N_168);
nand U4616 (N_4616,N_464,N_506);
nand U4617 (N_4617,N_674,N_1918);
or U4618 (N_4618,N_38,N_43);
nor U4619 (N_4619,N_1067,N_901);
or U4620 (N_4620,N_1560,N_1182);
nor U4621 (N_4621,N_766,N_2248);
nor U4622 (N_4622,N_1012,N_1828);
xor U4623 (N_4623,N_2083,N_114);
nor U4624 (N_4624,N_1504,N_1782);
nor U4625 (N_4625,N_1388,N_2291);
xor U4626 (N_4626,N_1940,N_1261);
nor U4627 (N_4627,N_775,N_1264);
and U4628 (N_4628,N_580,N_23);
nor U4629 (N_4629,N_1605,N_1563);
xor U4630 (N_4630,N_692,N_1308);
xnor U4631 (N_4631,N_1201,N_1596);
xnor U4632 (N_4632,N_768,N_248);
nand U4633 (N_4633,N_320,N_600);
nand U4634 (N_4634,N_2374,N_596);
nor U4635 (N_4635,N_2033,N_1680);
nand U4636 (N_4636,N_714,N_106);
and U4637 (N_4637,N_982,N_1939);
and U4638 (N_4638,N_650,N_1041);
or U4639 (N_4639,N_323,N_2165);
nand U4640 (N_4640,N_255,N_2368);
nand U4641 (N_4641,N_157,N_244);
nand U4642 (N_4642,N_901,N_2138);
or U4643 (N_4643,N_2182,N_2115);
or U4644 (N_4644,N_894,N_140);
xnor U4645 (N_4645,N_941,N_1427);
xor U4646 (N_4646,N_1833,N_1218);
or U4647 (N_4647,N_1512,N_1711);
or U4648 (N_4648,N_768,N_1209);
nor U4649 (N_4649,N_1797,N_34);
or U4650 (N_4650,N_719,N_870);
and U4651 (N_4651,N_363,N_139);
nand U4652 (N_4652,N_2208,N_1863);
xnor U4653 (N_4653,N_1124,N_2128);
nand U4654 (N_4654,N_725,N_862);
or U4655 (N_4655,N_2294,N_1036);
and U4656 (N_4656,N_1537,N_1024);
and U4657 (N_4657,N_1413,N_319);
and U4658 (N_4658,N_1352,N_374);
and U4659 (N_4659,N_1885,N_1542);
nand U4660 (N_4660,N_2099,N_1981);
nor U4661 (N_4661,N_1572,N_155);
nand U4662 (N_4662,N_941,N_1);
nor U4663 (N_4663,N_1731,N_634);
nor U4664 (N_4664,N_449,N_1915);
nor U4665 (N_4665,N_567,N_593);
or U4666 (N_4666,N_538,N_1409);
and U4667 (N_4667,N_1996,N_663);
nand U4668 (N_4668,N_985,N_1441);
nand U4669 (N_4669,N_2084,N_1262);
nand U4670 (N_4670,N_2449,N_1986);
nor U4671 (N_4671,N_395,N_612);
or U4672 (N_4672,N_1883,N_135);
and U4673 (N_4673,N_801,N_1695);
and U4674 (N_4674,N_926,N_284);
or U4675 (N_4675,N_1019,N_1054);
or U4676 (N_4676,N_980,N_2322);
nor U4677 (N_4677,N_282,N_2284);
nor U4678 (N_4678,N_48,N_1350);
nor U4679 (N_4679,N_1925,N_2323);
nand U4680 (N_4680,N_37,N_474);
xnor U4681 (N_4681,N_769,N_1395);
nand U4682 (N_4682,N_1704,N_1385);
and U4683 (N_4683,N_1653,N_2134);
nor U4684 (N_4684,N_1333,N_1134);
or U4685 (N_4685,N_755,N_2428);
or U4686 (N_4686,N_1660,N_2298);
or U4687 (N_4687,N_1368,N_1167);
or U4688 (N_4688,N_2159,N_543);
xor U4689 (N_4689,N_91,N_1827);
and U4690 (N_4690,N_698,N_362);
xor U4691 (N_4691,N_998,N_1213);
nor U4692 (N_4692,N_139,N_70);
xor U4693 (N_4693,N_1636,N_38);
nand U4694 (N_4694,N_27,N_1054);
xnor U4695 (N_4695,N_25,N_2222);
or U4696 (N_4696,N_1959,N_1095);
nand U4697 (N_4697,N_2194,N_1497);
nand U4698 (N_4698,N_730,N_1966);
and U4699 (N_4699,N_937,N_543);
nor U4700 (N_4700,N_2028,N_1174);
and U4701 (N_4701,N_132,N_1823);
xor U4702 (N_4702,N_288,N_1878);
nand U4703 (N_4703,N_2409,N_566);
nand U4704 (N_4704,N_346,N_940);
nor U4705 (N_4705,N_691,N_1487);
nor U4706 (N_4706,N_1312,N_1824);
and U4707 (N_4707,N_2113,N_2155);
nor U4708 (N_4708,N_919,N_1193);
nor U4709 (N_4709,N_55,N_842);
or U4710 (N_4710,N_980,N_946);
nor U4711 (N_4711,N_245,N_1888);
or U4712 (N_4712,N_551,N_1412);
xor U4713 (N_4713,N_1977,N_1707);
and U4714 (N_4714,N_1300,N_928);
xor U4715 (N_4715,N_1297,N_1424);
nor U4716 (N_4716,N_1352,N_1070);
and U4717 (N_4717,N_1733,N_1573);
or U4718 (N_4718,N_1618,N_1537);
xor U4719 (N_4719,N_935,N_1132);
nor U4720 (N_4720,N_1962,N_1457);
xor U4721 (N_4721,N_771,N_1712);
nor U4722 (N_4722,N_2208,N_842);
xnor U4723 (N_4723,N_1856,N_661);
xor U4724 (N_4724,N_242,N_2032);
and U4725 (N_4725,N_1441,N_850);
and U4726 (N_4726,N_1949,N_536);
nor U4727 (N_4727,N_2017,N_362);
nand U4728 (N_4728,N_2351,N_62);
and U4729 (N_4729,N_2153,N_626);
or U4730 (N_4730,N_1341,N_1401);
xor U4731 (N_4731,N_71,N_517);
nand U4732 (N_4732,N_1675,N_225);
nand U4733 (N_4733,N_1071,N_1531);
nor U4734 (N_4734,N_1920,N_617);
or U4735 (N_4735,N_1399,N_2362);
nand U4736 (N_4736,N_2265,N_483);
and U4737 (N_4737,N_696,N_333);
nand U4738 (N_4738,N_1864,N_1126);
xnor U4739 (N_4739,N_608,N_1216);
xnor U4740 (N_4740,N_1728,N_225);
nand U4741 (N_4741,N_522,N_1264);
or U4742 (N_4742,N_649,N_189);
xnor U4743 (N_4743,N_547,N_1939);
and U4744 (N_4744,N_948,N_2431);
and U4745 (N_4745,N_2497,N_1058);
nand U4746 (N_4746,N_840,N_1544);
nor U4747 (N_4747,N_429,N_796);
and U4748 (N_4748,N_1121,N_322);
or U4749 (N_4749,N_686,N_2056);
or U4750 (N_4750,N_1645,N_1175);
nor U4751 (N_4751,N_1386,N_2438);
nor U4752 (N_4752,N_2462,N_1008);
nor U4753 (N_4753,N_1778,N_85);
xnor U4754 (N_4754,N_1738,N_1427);
and U4755 (N_4755,N_263,N_1806);
and U4756 (N_4756,N_1305,N_2262);
nor U4757 (N_4757,N_1051,N_426);
nand U4758 (N_4758,N_385,N_1032);
or U4759 (N_4759,N_372,N_1942);
nor U4760 (N_4760,N_486,N_2067);
nor U4761 (N_4761,N_973,N_767);
nand U4762 (N_4762,N_804,N_1307);
or U4763 (N_4763,N_2005,N_1205);
or U4764 (N_4764,N_652,N_1238);
nor U4765 (N_4765,N_941,N_462);
or U4766 (N_4766,N_2177,N_1916);
nand U4767 (N_4767,N_60,N_517);
xor U4768 (N_4768,N_1421,N_340);
xor U4769 (N_4769,N_506,N_497);
and U4770 (N_4770,N_1658,N_2037);
xor U4771 (N_4771,N_1212,N_2295);
xnor U4772 (N_4772,N_644,N_2226);
nand U4773 (N_4773,N_1400,N_1142);
or U4774 (N_4774,N_1461,N_1919);
or U4775 (N_4775,N_962,N_216);
or U4776 (N_4776,N_818,N_956);
or U4777 (N_4777,N_1183,N_2144);
nor U4778 (N_4778,N_282,N_200);
or U4779 (N_4779,N_1964,N_2499);
xor U4780 (N_4780,N_2357,N_1782);
and U4781 (N_4781,N_537,N_1423);
and U4782 (N_4782,N_2113,N_2460);
nor U4783 (N_4783,N_1341,N_2137);
nor U4784 (N_4784,N_1697,N_286);
xor U4785 (N_4785,N_1663,N_515);
xnor U4786 (N_4786,N_233,N_529);
or U4787 (N_4787,N_387,N_2088);
nand U4788 (N_4788,N_120,N_998);
xor U4789 (N_4789,N_2491,N_1020);
and U4790 (N_4790,N_2045,N_85);
nand U4791 (N_4791,N_2253,N_1616);
nand U4792 (N_4792,N_1363,N_1603);
nor U4793 (N_4793,N_2302,N_558);
or U4794 (N_4794,N_2401,N_650);
nor U4795 (N_4795,N_1017,N_349);
and U4796 (N_4796,N_699,N_105);
and U4797 (N_4797,N_702,N_1299);
and U4798 (N_4798,N_2274,N_385);
nand U4799 (N_4799,N_1262,N_2119);
nand U4800 (N_4800,N_1011,N_1224);
xnor U4801 (N_4801,N_1631,N_851);
nor U4802 (N_4802,N_439,N_1898);
or U4803 (N_4803,N_1071,N_847);
xnor U4804 (N_4804,N_2328,N_2093);
and U4805 (N_4805,N_2444,N_2386);
or U4806 (N_4806,N_2396,N_339);
and U4807 (N_4807,N_1250,N_545);
nor U4808 (N_4808,N_1208,N_1388);
nor U4809 (N_4809,N_2163,N_16);
or U4810 (N_4810,N_941,N_111);
and U4811 (N_4811,N_92,N_502);
nor U4812 (N_4812,N_1441,N_665);
or U4813 (N_4813,N_19,N_355);
nand U4814 (N_4814,N_1395,N_755);
xor U4815 (N_4815,N_2465,N_1491);
xor U4816 (N_4816,N_424,N_1235);
xnor U4817 (N_4817,N_2385,N_259);
nand U4818 (N_4818,N_1601,N_1608);
and U4819 (N_4819,N_2273,N_2371);
or U4820 (N_4820,N_1119,N_931);
xnor U4821 (N_4821,N_1869,N_824);
nor U4822 (N_4822,N_130,N_1852);
nor U4823 (N_4823,N_1895,N_798);
or U4824 (N_4824,N_2078,N_2369);
or U4825 (N_4825,N_517,N_962);
and U4826 (N_4826,N_1740,N_1489);
xnor U4827 (N_4827,N_1872,N_1254);
nor U4828 (N_4828,N_1887,N_410);
and U4829 (N_4829,N_1198,N_76);
nand U4830 (N_4830,N_791,N_364);
xnor U4831 (N_4831,N_1793,N_163);
nor U4832 (N_4832,N_443,N_1623);
or U4833 (N_4833,N_2236,N_944);
xnor U4834 (N_4834,N_164,N_1970);
nor U4835 (N_4835,N_52,N_2416);
or U4836 (N_4836,N_1015,N_1300);
xor U4837 (N_4837,N_112,N_2172);
or U4838 (N_4838,N_1742,N_1733);
xor U4839 (N_4839,N_2005,N_647);
nor U4840 (N_4840,N_1713,N_2156);
or U4841 (N_4841,N_1920,N_1664);
and U4842 (N_4842,N_290,N_2139);
xor U4843 (N_4843,N_1741,N_1694);
or U4844 (N_4844,N_948,N_359);
nor U4845 (N_4845,N_1402,N_1958);
or U4846 (N_4846,N_1104,N_488);
nand U4847 (N_4847,N_1543,N_2219);
nand U4848 (N_4848,N_176,N_2031);
or U4849 (N_4849,N_99,N_1824);
nor U4850 (N_4850,N_105,N_2257);
nor U4851 (N_4851,N_929,N_1280);
nor U4852 (N_4852,N_917,N_2343);
nor U4853 (N_4853,N_1338,N_529);
nand U4854 (N_4854,N_2190,N_2038);
or U4855 (N_4855,N_1159,N_1934);
nor U4856 (N_4856,N_1558,N_461);
nand U4857 (N_4857,N_2238,N_438);
and U4858 (N_4858,N_603,N_1391);
and U4859 (N_4859,N_154,N_801);
and U4860 (N_4860,N_1400,N_2107);
or U4861 (N_4861,N_150,N_1482);
or U4862 (N_4862,N_862,N_2102);
and U4863 (N_4863,N_636,N_1818);
and U4864 (N_4864,N_1264,N_1628);
nor U4865 (N_4865,N_1751,N_1934);
xor U4866 (N_4866,N_2276,N_1738);
or U4867 (N_4867,N_2426,N_628);
nor U4868 (N_4868,N_1269,N_747);
nand U4869 (N_4869,N_1942,N_1895);
and U4870 (N_4870,N_2221,N_1744);
nand U4871 (N_4871,N_585,N_1905);
nand U4872 (N_4872,N_1841,N_802);
nand U4873 (N_4873,N_962,N_1594);
nor U4874 (N_4874,N_391,N_1241);
nor U4875 (N_4875,N_44,N_1768);
xor U4876 (N_4876,N_2008,N_1980);
and U4877 (N_4877,N_803,N_2082);
xnor U4878 (N_4878,N_215,N_1769);
xnor U4879 (N_4879,N_2214,N_990);
nand U4880 (N_4880,N_1207,N_1850);
or U4881 (N_4881,N_370,N_606);
and U4882 (N_4882,N_566,N_1861);
nand U4883 (N_4883,N_1742,N_1662);
nand U4884 (N_4884,N_1128,N_1735);
nand U4885 (N_4885,N_1258,N_1870);
or U4886 (N_4886,N_307,N_1666);
nor U4887 (N_4887,N_1158,N_1871);
and U4888 (N_4888,N_2333,N_1035);
xnor U4889 (N_4889,N_1172,N_2112);
xnor U4890 (N_4890,N_1061,N_332);
and U4891 (N_4891,N_1504,N_1262);
xnor U4892 (N_4892,N_713,N_1973);
nor U4893 (N_4893,N_1740,N_1345);
xor U4894 (N_4894,N_650,N_2444);
nor U4895 (N_4895,N_2467,N_513);
nand U4896 (N_4896,N_272,N_913);
nand U4897 (N_4897,N_1732,N_656);
xor U4898 (N_4898,N_1054,N_1127);
and U4899 (N_4899,N_2238,N_288);
nand U4900 (N_4900,N_1841,N_334);
nand U4901 (N_4901,N_1191,N_1984);
nand U4902 (N_4902,N_615,N_1700);
nor U4903 (N_4903,N_1809,N_1730);
nor U4904 (N_4904,N_1876,N_1031);
or U4905 (N_4905,N_7,N_1898);
nand U4906 (N_4906,N_960,N_844);
and U4907 (N_4907,N_1093,N_88);
nand U4908 (N_4908,N_2116,N_1574);
or U4909 (N_4909,N_1150,N_1165);
and U4910 (N_4910,N_1205,N_2000);
and U4911 (N_4911,N_1342,N_1327);
nand U4912 (N_4912,N_2385,N_62);
or U4913 (N_4913,N_200,N_1919);
nand U4914 (N_4914,N_1985,N_698);
nand U4915 (N_4915,N_1598,N_2458);
and U4916 (N_4916,N_59,N_124);
or U4917 (N_4917,N_511,N_1211);
nor U4918 (N_4918,N_2223,N_1096);
xnor U4919 (N_4919,N_462,N_2135);
or U4920 (N_4920,N_1160,N_1982);
and U4921 (N_4921,N_1841,N_247);
xor U4922 (N_4922,N_2228,N_464);
or U4923 (N_4923,N_180,N_2126);
and U4924 (N_4924,N_778,N_894);
or U4925 (N_4925,N_706,N_1896);
nand U4926 (N_4926,N_1599,N_645);
nor U4927 (N_4927,N_1402,N_750);
nand U4928 (N_4928,N_381,N_974);
or U4929 (N_4929,N_2357,N_1529);
and U4930 (N_4930,N_2441,N_1700);
and U4931 (N_4931,N_1135,N_393);
xor U4932 (N_4932,N_1747,N_2209);
and U4933 (N_4933,N_1735,N_429);
nand U4934 (N_4934,N_100,N_673);
and U4935 (N_4935,N_1726,N_1216);
nand U4936 (N_4936,N_1985,N_140);
xor U4937 (N_4937,N_1692,N_2076);
xor U4938 (N_4938,N_2227,N_704);
or U4939 (N_4939,N_3,N_2415);
and U4940 (N_4940,N_2286,N_2326);
nand U4941 (N_4941,N_1444,N_12);
and U4942 (N_4942,N_391,N_522);
xnor U4943 (N_4943,N_420,N_486);
xnor U4944 (N_4944,N_427,N_1639);
xnor U4945 (N_4945,N_150,N_1446);
nand U4946 (N_4946,N_2050,N_1046);
nand U4947 (N_4947,N_547,N_1595);
nor U4948 (N_4948,N_786,N_2075);
nand U4949 (N_4949,N_661,N_296);
nand U4950 (N_4950,N_2172,N_1361);
xnor U4951 (N_4951,N_706,N_943);
nor U4952 (N_4952,N_508,N_1198);
nand U4953 (N_4953,N_962,N_2385);
and U4954 (N_4954,N_1505,N_426);
or U4955 (N_4955,N_1087,N_1796);
nand U4956 (N_4956,N_299,N_2171);
nor U4957 (N_4957,N_1372,N_1223);
nor U4958 (N_4958,N_1168,N_1403);
nand U4959 (N_4959,N_269,N_1009);
or U4960 (N_4960,N_992,N_2106);
nor U4961 (N_4961,N_1030,N_1334);
and U4962 (N_4962,N_2414,N_829);
xnor U4963 (N_4963,N_639,N_2392);
and U4964 (N_4964,N_1643,N_2287);
and U4965 (N_4965,N_2185,N_1656);
nor U4966 (N_4966,N_923,N_1975);
or U4967 (N_4967,N_1891,N_144);
nand U4968 (N_4968,N_1263,N_1765);
xnor U4969 (N_4969,N_854,N_2140);
nor U4970 (N_4970,N_902,N_7);
xnor U4971 (N_4971,N_140,N_1730);
and U4972 (N_4972,N_1055,N_185);
and U4973 (N_4973,N_1559,N_1044);
or U4974 (N_4974,N_302,N_2347);
nand U4975 (N_4975,N_905,N_95);
or U4976 (N_4976,N_497,N_1466);
or U4977 (N_4977,N_804,N_1047);
nor U4978 (N_4978,N_2275,N_1775);
nand U4979 (N_4979,N_2005,N_1172);
or U4980 (N_4980,N_1336,N_1489);
and U4981 (N_4981,N_1685,N_390);
nor U4982 (N_4982,N_552,N_1430);
nand U4983 (N_4983,N_97,N_855);
xor U4984 (N_4984,N_9,N_1559);
xnor U4985 (N_4985,N_1907,N_1122);
or U4986 (N_4986,N_1456,N_320);
or U4987 (N_4987,N_2407,N_554);
xnor U4988 (N_4988,N_1606,N_1454);
and U4989 (N_4989,N_2208,N_1230);
nor U4990 (N_4990,N_813,N_2327);
nor U4991 (N_4991,N_2244,N_2387);
nor U4992 (N_4992,N_1056,N_1031);
xor U4993 (N_4993,N_1981,N_207);
xor U4994 (N_4994,N_1900,N_1632);
or U4995 (N_4995,N_2185,N_1335);
nor U4996 (N_4996,N_1151,N_1103);
nor U4997 (N_4997,N_1125,N_1684);
and U4998 (N_4998,N_65,N_1652);
xnor U4999 (N_4999,N_2058,N_172);
and UO_0 (O_0,N_2613,N_3393);
or UO_1 (O_1,N_4570,N_4197);
nand UO_2 (O_2,N_2664,N_4983);
and UO_3 (O_3,N_4509,N_2923);
xnor UO_4 (O_4,N_3176,N_3985);
or UO_5 (O_5,N_3660,N_2813);
nor UO_6 (O_6,N_2733,N_3757);
and UO_7 (O_7,N_3998,N_3542);
or UO_8 (O_8,N_4871,N_4798);
nor UO_9 (O_9,N_4172,N_2703);
or UO_10 (O_10,N_3827,N_3579);
and UO_11 (O_11,N_4362,N_3852);
and UO_12 (O_12,N_3999,N_3519);
or UO_13 (O_13,N_4361,N_3018);
nor UO_14 (O_14,N_4451,N_3430);
nand UO_15 (O_15,N_2953,N_3984);
xor UO_16 (O_16,N_3167,N_3692);
or UO_17 (O_17,N_4228,N_4248);
and UO_18 (O_18,N_4124,N_2964);
nand UO_19 (O_19,N_3131,N_3074);
xor UO_20 (O_20,N_3055,N_2598);
or UO_21 (O_21,N_2695,N_4122);
xnor UO_22 (O_22,N_3236,N_3416);
nor UO_23 (O_23,N_4236,N_3489);
xnor UO_24 (O_24,N_2624,N_4673);
nor UO_25 (O_25,N_4438,N_3793);
nand UO_26 (O_26,N_4812,N_4457);
xnor UO_27 (O_27,N_3569,N_4684);
xor UO_28 (O_28,N_3736,N_4605);
or UO_29 (O_29,N_3989,N_3319);
nor UO_30 (O_30,N_4959,N_2868);
xnor UO_31 (O_31,N_2604,N_3492);
and UO_32 (O_32,N_2600,N_4883);
and UO_33 (O_33,N_2913,N_2992);
xnor UO_34 (O_34,N_3628,N_2878);
xnor UO_35 (O_35,N_4877,N_4691);
nor UO_36 (O_36,N_2693,N_3633);
nand UO_37 (O_37,N_3249,N_3465);
nor UO_38 (O_38,N_2615,N_3216);
nor UO_39 (O_39,N_3100,N_4978);
and UO_40 (O_40,N_4909,N_4458);
nand UO_41 (O_41,N_4359,N_3873);
and UO_42 (O_42,N_3877,N_2980);
xnor UO_43 (O_43,N_2730,N_4875);
xor UO_44 (O_44,N_4853,N_2656);
xor UO_45 (O_45,N_4337,N_3717);
xor UO_46 (O_46,N_4018,N_3674);
nor UO_47 (O_47,N_3923,N_4650);
xor UO_48 (O_48,N_2871,N_4994);
or UO_49 (O_49,N_3039,N_3370);
or UO_50 (O_50,N_2883,N_2528);
xnor UO_51 (O_51,N_3607,N_4863);
nand UO_52 (O_52,N_3867,N_3598);
nor UO_53 (O_53,N_2525,N_2920);
nand UO_54 (O_54,N_3602,N_4250);
xor UO_55 (O_55,N_2820,N_4521);
or UO_56 (O_56,N_3853,N_4797);
and UO_57 (O_57,N_4062,N_3748);
nor UO_58 (O_58,N_4370,N_4003);
nor UO_59 (O_59,N_4920,N_2501);
xor UO_60 (O_60,N_3501,N_4126);
xor UO_61 (O_61,N_3314,N_2792);
xor UO_62 (O_62,N_4653,N_4760);
and UO_63 (O_63,N_2709,N_4693);
nand UO_64 (O_64,N_4061,N_4940);
xor UO_65 (O_65,N_4543,N_4638);
or UO_66 (O_66,N_3481,N_4135);
xor UO_67 (O_67,N_3208,N_2747);
xor UO_68 (O_68,N_4331,N_3253);
and UO_69 (O_69,N_2614,N_3750);
nand UO_70 (O_70,N_3864,N_4093);
nand UO_71 (O_71,N_4555,N_3218);
and UO_72 (O_72,N_4502,N_2797);
nand UO_73 (O_73,N_3032,N_3452);
xnor UO_74 (O_74,N_4556,N_4517);
or UO_75 (O_75,N_2821,N_4544);
nand UO_76 (O_76,N_3145,N_3766);
nand UO_77 (O_77,N_4349,N_2706);
nor UO_78 (O_78,N_2539,N_3549);
xor UO_79 (O_79,N_3548,N_3629);
xor UO_80 (O_80,N_4017,N_2523);
or UO_81 (O_81,N_3547,N_2961);
nor UO_82 (O_82,N_4204,N_4390);
nor UO_83 (O_83,N_3693,N_2689);
or UO_84 (O_84,N_4498,N_3106);
nand UO_85 (O_85,N_3747,N_2808);
nand UO_86 (O_86,N_3391,N_2680);
xor UO_87 (O_87,N_2972,N_4874);
and UO_88 (O_88,N_4888,N_3132);
and UO_89 (O_89,N_4632,N_3605);
nand UO_90 (O_90,N_2690,N_4944);
and UO_91 (O_91,N_4401,N_4431);
nand UO_92 (O_92,N_4417,N_3022);
or UO_93 (O_93,N_3844,N_4525);
or UO_94 (O_94,N_3740,N_3280);
and UO_95 (O_95,N_4154,N_4393);
or UO_96 (O_96,N_4765,N_3924);
xor UO_97 (O_97,N_3392,N_3591);
nor UO_98 (O_98,N_4835,N_4226);
nand UO_99 (O_99,N_3233,N_2927);
or UO_100 (O_100,N_2666,N_4947);
xnor UO_101 (O_101,N_2653,N_2874);
or UO_102 (O_102,N_3973,N_4101);
or UO_103 (O_103,N_3206,N_4219);
and UO_104 (O_104,N_4002,N_3926);
xor UO_105 (O_105,N_4515,N_2901);
nor UO_106 (O_106,N_3780,N_2860);
xnor UO_107 (O_107,N_4821,N_3774);
and UO_108 (O_108,N_3498,N_4088);
nor UO_109 (O_109,N_3034,N_2867);
or UO_110 (O_110,N_4127,N_3972);
and UO_111 (O_111,N_2776,N_4052);
and UO_112 (O_112,N_4995,N_3735);
or UO_113 (O_113,N_2917,N_2778);
nand UO_114 (O_114,N_4579,N_4034);
nand UO_115 (O_115,N_3186,N_3876);
xor UO_116 (O_116,N_3190,N_2982);
nor UO_117 (O_117,N_3551,N_4470);
or UO_118 (O_118,N_4339,N_3302);
nor UO_119 (O_119,N_4425,N_3860);
xor UO_120 (O_120,N_3679,N_3080);
nor UO_121 (O_121,N_4346,N_3352);
xnor UO_122 (O_122,N_3557,N_3010);
and UO_123 (O_123,N_3920,N_3954);
xnor UO_124 (O_124,N_2833,N_3312);
or UO_125 (O_125,N_4568,N_4831);
nor UO_126 (O_126,N_4882,N_3480);
or UO_127 (O_127,N_2942,N_4820);
xor UO_128 (O_128,N_3311,N_4157);
nor UO_129 (O_129,N_3321,N_2862);
nor UO_130 (O_130,N_3337,N_3711);
and UO_131 (O_131,N_4257,N_3180);
and UO_132 (O_132,N_3110,N_4276);
nand UO_133 (O_133,N_3938,N_4218);
and UO_134 (O_134,N_4958,N_2661);
and UO_135 (O_135,N_4468,N_2897);
and UO_136 (O_136,N_4782,N_2755);
nand UO_137 (O_137,N_2603,N_3062);
or UO_138 (O_138,N_3346,N_3009);
and UO_139 (O_139,N_4652,N_4830);
and UO_140 (O_140,N_2711,N_2831);
nor UO_141 (O_141,N_3901,N_4004);
and UO_142 (O_142,N_4330,N_2617);
or UO_143 (O_143,N_3315,N_4260);
nor UO_144 (O_144,N_4721,N_4495);
or UO_145 (O_145,N_4266,N_4435);
and UO_146 (O_146,N_4787,N_4656);
and UO_147 (O_147,N_2790,N_3033);
or UO_148 (O_148,N_4324,N_2907);
xnor UO_149 (O_149,N_3940,N_4766);
nand UO_150 (O_150,N_2549,N_4700);
or UO_151 (O_151,N_2771,N_4828);
or UO_152 (O_152,N_4343,N_3486);
and UO_153 (O_153,N_3813,N_3036);
nand UO_154 (O_154,N_3192,N_3068);
and UO_155 (O_155,N_4099,N_4180);
or UO_156 (O_156,N_2803,N_4530);
or UO_157 (O_157,N_3245,N_3800);
or UO_158 (O_158,N_3214,N_4674);
xnor UO_159 (O_159,N_4979,N_4780);
and UO_160 (O_160,N_3215,N_2950);
or UO_161 (O_161,N_4886,N_4245);
and UO_162 (O_162,N_4560,N_2859);
or UO_163 (O_163,N_2938,N_3515);
or UO_164 (O_164,N_3196,N_3325);
xnor UO_165 (O_165,N_4561,N_4005);
or UO_166 (O_166,N_3541,N_4480);
xnor UO_167 (O_167,N_4982,N_3158);
nor UO_168 (O_168,N_2537,N_4255);
nor UO_169 (O_169,N_4763,N_2947);
and UO_170 (O_170,N_3659,N_2798);
xnor UO_171 (O_171,N_3344,N_3798);
xnor UO_172 (O_172,N_2572,N_3138);
or UO_173 (O_173,N_3732,N_2532);
or UO_174 (O_174,N_3558,N_2726);
nor UO_175 (O_175,N_2943,N_4665);
or UO_176 (O_176,N_3610,N_3440);
or UO_177 (O_177,N_3854,N_3779);
nand UO_178 (O_178,N_4128,N_4938);
xnor UO_179 (O_179,N_3684,N_2756);
and UO_180 (O_180,N_3444,N_4790);
and UO_181 (O_181,N_2941,N_4628);
and UO_182 (O_182,N_2773,N_4666);
xor UO_183 (O_183,N_4079,N_3408);
nor UO_184 (O_184,N_3203,N_4647);
nand UO_185 (O_185,N_4239,N_3776);
or UO_186 (O_186,N_4258,N_4692);
and UO_187 (O_187,N_4709,N_3081);
nor UO_188 (O_188,N_4312,N_3403);
xor UO_189 (O_189,N_2899,N_3228);
nor UO_190 (O_190,N_3576,N_3683);
or UO_191 (O_191,N_2933,N_3157);
nand UO_192 (O_192,N_4357,N_2580);
or UO_193 (O_193,N_4566,N_3371);
nand UO_194 (O_194,N_2975,N_3504);
nand UO_195 (O_195,N_4981,N_3955);
xnor UO_196 (O_196,N_3815,N_4844);
nand UO_197 (O_197,N_3414,N_3256);
nor UO_198 (O_198,N_2724,N_3499);
nand UO_199 (O_199,N_4044,N_2902);
and UO_200 (O_200,N_3868,N_2959);
nand UO_201 (O_201,N_2535,N_3834);
xor UO_202 (O_202,N_3952,N_3529);
nand UO_203 (O_203,N_2582,N_2981);
xor UO_204 (O_204,N_3246,N_3367);
or UO_205 (O_205,N_3472,N_2585);
or UO_206 (O_206,N_3755,N_4178);
nor UO_207 (O_207,N_4006,N_2885);
or UO_208 (O_208,N_3648,N_3544);
and UO_209 (O_209,N_3202,N_4203);
nor UO_210 (O_210,N_4919,N_3654);
and UO_211 (O_211,N_4338,N_4308);
and UO_212 (O_212,N_3428,N_3518);
or UO_213 (O_213,N_3008,N_3259);
or UO_214 (O_214,N_4589,N_2835);
or UO_215 (O_215,N_3828,N_2767);
nor UO_216 (O_216,N_4256,N_3318);
xnor UO_217 (O_217,N_4997,N_3059);
nand UO_218 (O_218,N_2744,N_4325);
xor UO_219 (O_219,N_3744,N_3359);
xor UO_220 (O_220,N_3507,N_3248);
and UO_221 (O_221,N_3718,N_4520);
and UO_222 (O_222,N_2504,N_2725);
nand UO_223 (O_223,N_3642,N_3052);
xnor UO_224 (O_224,N_4261,N_4939);
or UO_225 (O_225,N_3172,N_2512);
or UO_226 (O_226,N_3661,N_2687);
nand UO_227 (O_227,N_2578,N_3305);
and UO_228 (O_228,N_4942,N_4233);
or UO_229 (O_229,N_3289,N_3412);
or UO_230 (O_230,N_2822,N_3791);
nor UO_231 (O_231,N_2577,N_2631);
nor UO_232 (O_232,N_2527,N_4202);
and UO_233 (O_233,N_3656,N_2634);
nor UO_234 (O_234,N_4162,N_3205);
or UO_235 (O_235,N_4848,N_3178);
xnor UO_236 (O_236,N_3258,N_4591);
nand UO_237 (O_237,N_2705,N_3121);
xnor UO_238 (O_238,N_4649,N_4757);
nor UO_239 (O_239,N_4113,N_4169);
and UO_240 (O_240,N_2852,N_4041);
nor UO_241 (O_241,N_4676,N_3913);
and UO_242 (O_242,N_4810,N_3045);
and UO_243 (O_243,N_2839,N_3060);
nor UO_244 (O_244,N_4242,N_4224);
and UO_245 (O_245,N_4430,N_4225);
xor UO_246 (O_246,N_3822,N_3724);
nand UO_247 (O_247,N_4010,N_3191);
or UO_248 (O_248,N_4476,N_3820);
nand UO_249 (O_249,N_4885,N_4633);
xnor UO_250 (O_250,N_4992,N_3974);
nand UO_251 (O_251,N_4668,N_3016);
or UO_252 (O_252,N_3355,N_3410);
and UO_253 (O_253,N_2999,N_3129);
nand UO_254 (O_254,N_4027,N_3301);
nand UO_255 (O_255,N_4711,N_3026);
nor UO_256 (O_256,N_4972,N_4552);
nand UO_257 (O_257,N_2625,N_4694);
and UO_258 (O_258,N_4269,N_3209);
and UO_259 (O_259,N_4850,N_4252);
and UO_260 (O_260,N_2606,N_3266);
xor UO_261 (O_261,N_2956,N_4645);
or UO_262 (O_262,N_2679,N_3287);
or UO_263 (O_263,N_4300,N_2530);
nor UO_264 (O_264,N_2673,N_3070);
and UO_265 (O_265,N_3013,N_3810);
nand UO_266 (O_266,N_4487,N_4669);
xor UO_267 (O_267,N_3381,N_4328);
and UO_268 (O_268,N_4314,N_2837);
nor UO_269 (O_269,N_3083,N_4922);
nor UO_270 (O_270,N_3028,N_2715);
or UO_271 (O_271,N_3041,N_3935);
and UO_272 (O_272,N_2855,N_4206);
xor UO_273 (O_273,N_3338,N_3446);
nor UO_274 (O_274,N_3270,N_3156);
or UO_275 (O_275,N_4244,N_3360);
nor UO_276 (O_276,N_3906,N_4403);
nor UO_277 (O_277,N_4500,N_2781);
nand UO_278 (O_278,N_3523,N_4415);
and UO_279 (O_279,N_2542,N_2896);
and UO_280 (O_280,N_4089,N_4527);
xor UO_281 (O_281,N_3115,N_2654);
nor UO_282 (O_282,N_4183,N_2783);
and UO_283 (O_283,N_4758,N_2853);
nor UO_284 (O_284,N_2672,N_4081);
and UO_285 (O_285,N_2529,N_4977);
nand UO_286 (O_286,N_4953,N_4402);
or UO_287 (O_287,N_4137,N_4391);
or UO_288 (O_288,N_4825,N_2632);
and UO_289 (O_289,N_3503,N_3421);
and UO_290 (O_290,N_4910,N_3758);
and UO_291 (O_291,N_2669,N_3339);
xor UO_292 (O_292,N_4756,N_3993);
xnor UO_293 (O_293,N_4639,N_2968);
and UO_294 (O_294,N_3616,N_4304);
nand UO_295 (O_295,N_3630,N_4007);
nor UO_296 (O_296,N_4672,N_4683);
nor UO_297 (O_297,N_3291,N_3491);
nor UO_298 (O_298,N_2658,N_4053);
nand UO_299 (O_299,N_2588,N_4047);
or UO_300 (O_300,N_2856,N_4627);
nand UO_301 (O_301,N_2815,N_3650);
or UO_302 (O_302,N_2921,N_3589);
nand UO_303 (O_303,N_3559,N_2983);
nor UO_304 (O_304,N_4818,N_3435);
nand UO_305 (O_305,N_3020,N_4465);
or UO_306 (O_306,N_4833,N_2799);
xor UO_307 (O_307,N_4434,N_4518);
xnor UO_308 (O_308,N_4951,N_3567);
or UO_309 (O_309,N_3925,N_3928);
nand UO_310 (O_310,N_3789,N_3971);
or UO_311 (O_311,N_4999,N_3098);
nor UO_312 (O_312,N_3866,N_3201);
xor UO_313 (O_313,N_4194,N_3454);
nand UO_314 (O_314,N_4395,N_3712);
xor UO_315 (O_315,N_2962,N_3136);
or UO_316 (O_316,N_4708,N_3119);
and UO_317 (O_317,N_4383,N_4916);
or UO_318 (O_318,N_2675,N_4703);
and UO_319 (O_319,N_3603,N_4563);
nand UO_320 (O_320,N_3664,N_4374);
or UO_321 (O_321,N_3941,N_4453);
xnor UO_322 (O_322,N_3963,N_2963);
nand UO_323 (O_323,N_4774,N_3817);
or UO_324 (O_324,N_4344,N_4220);
or UO_325 (O_325,N_4936,N_3273);
nand UO_326 (O_326,N_4772,N_3162);
xnor UO_327 (O_327,N_2932,N_4184);
xor UO_328 (O_328,N_3824,N_4032);
nand UO_329 (O_329,N_4422,N_2678);
nor UO_330 (O_330,N_3574,N_2676);
nand UO_331 (O_331,N_4466,N_2740);
and UO_332 (O_332,N_3478,N_2629);
nor UO_333 (O_333,N_2898,N_4768);
nor UO_334 (O_334,N_3647,N_2795);
and UO_335 (O_335,N_3244,N_4966);
xor UO_336 (O_336,N_4196,N_3983);
nand UO_337 (O_337,N_4011,N_3874);
and UO_338 (O_338,N_4791,N_4964);
or UO_339 (O_339,N_4494,N_3379);
xor UO_340 (O_340,N_2811,N_3885);
xor UO_341 (O_341,N_4644,N_4701);
or UO_342 (O_342,N_2729,N_3232);
or UO_343 (O_343,N_3212,N_3632);
nand UO_344 (O_344,N_4847,N_4870);
xor UO_345 (O_345,N_4723,N_3405);
xnor UO_346 (O_346,N_3439,N_4497);
nand UO_347 (O_347,N_2564,N_4115);
xnor UO_348 (O_348,N_3534,N_3966);
xnor UO_349 (O_349,N_3536,N_3584);
xor UO_350 (O_350,N_4596,N_3290);
and UO_351 (O_351,N_3332,N_4216);
nor UO_352 (O_352,N_3524,N_3965);
or UO_353 (O_353,N_4906,N_4955);
or UO_354 (O_354,N_3897,N_3698);
xor UO_355 (O_355,N_2503,N_3051);
and UO_356 (O_356,N_2994,N_4121);
or UO_357 (O_357,N_4516,N_4504);
and UO_358 (O_358,N_2630,N_3448);
nor UO_359 (O_359,N_3419,N_4026);
and UO_360 (O_360,N_4479,N_4110);
or UO_361 (O_361,N_3105,N_4399);
and UO_362 (O_362,N_3731,N_3575);
nand UO_363 (O_363,N_3823,N_2716);
nand UO_364 (O_364,N_2692,N_2649);
and UO_365 (O_365,N_4364,N_3449);
and UO_366 (O_366,N_3902,N_3577);
nand UO_367 (O_367,N_2545,N_4108);
and UO_368 (O_368,N_3078,N_3967);
xor UO_369 (O_369,N_4444,N_3561);
nor UO_370 (O_370,N_3089,N_2801);
nand UO_371 (O_371,N_3863,N_3847);
and UO_372 (O_372,N_4559,N_3788);
xor UO_373 (O_373,N_4642,N_3471);
xor UO_374 (O_374,N_2924,N_3267);
xnor UO_375 (O_375,N_3021,N_3085);
and UO_376 (O_376,N_4925,N_4176);
nor UO_377 (O_377,N_3533,N_4071);
or UO_378 (O_378,N_2586,N_3933);
or UO_379 (O_379,N_3432,N_3896);
and UO_380 (O_380,N_3189,N_2974);
nand UO_381 (O_381,N_3981,N_4469);
and UO_382 (O_382,N_2522,N_4141);
or UO_383 (O_383,N_2579,N_2566);
and UO_384 (O_384,N_3573,N_3570);
and UO_385 (O_385,N_4414,N_4808);
nor UO_386 (O_386,N_2511,N_4733);
nor UO_387 (O_387,N_3197,N_4251);
xor UO_388 (O_388,N_4789,N_3624);
xor UO_389 (O_389,N_2728,N_3922);
xor UO_390 (O_390,N_4836,N_3126);
xnor UO_391 (O_391,N_3582,N_3856);
or UO_392 (O_392,N_2940,N_4309);
nand UO_393 (O_393,N_2670,N_2660);
or UO_394 (O_394,N_3090,N_4015);
or UO_395 (O_395,N_3704,N_2804);
xor UO_396 (O_396,N_2903,N_4807);
nand UO_397 (O_397,N_3211,N_3317);
nor UO_398 (O_398,N_2727,N_3413);
xnor UO_399 (O_399,N_2575,N_3595);
nor UO_400 (O_400,N_2720,N_3671);
and UO_401 (O_401,N_3721,N_4604);
xnor UO_402 (O_402,N_4253,N_4294);
nor UO_403 (O_403,N_3025,N_2643);
nand UO_404 (O_404,N_3177,N_3445);
and UO_405 (O_405,N_4424,N_4598);
nor UO_406 (O_406,N_3474,N_3451);
and UO_407 (O_407,N_3634,N_2612);
nand UO_408 (O_408,N_3670,N_4637);
or UO_409 (O_409,N_4862,N_2828);
and UO_410 (O_410,N_4501,N_2889);
and UO_411 (O_411,N_3699,N_4686);
xnor UO_412 (O_412,N_2743,N_3356);
or UO_413 (O_413,N_3175,N_4166);
nor UO_414 (O_414,N_3463,N_2990);
nor UO_415 (O_415,N_2683,N_3681);
xor UO_416 (O_416,N_4990,N_3252);
nor UO_417 (O_417,N_3239,N_3705);
nand UO_418 (O_418,N_2909,N_4263);
nor UO_419 (O_419,N_2971,N_4208);
nand UO_420 (O_420,N_4221,N_3843);
nand UO_421 (O_421,N_3895,N_3015);
nor UO_422 (O_422,N_4471,N_4727);
nand UO_423 (O_423,N_4333,N_2684);
nor UO_424 (O_424,N_4031,N_4602);
nand UO_425 (O_425,N_3803,N_4144);
and UO_426 (O_426,N_3394,N_2531);
or UO_427 (O_427,N_3939,N_4839);
nand UO_428 (O_428,N_2685,N_2872);
or UO_429 (O_429,N_4613,N_4750);
nand UO_430 (O_430,N_3685,N_4119);
and UO_431 (O_431,N_4793,N_4679);
nand UO_432 (O_432,N_3422,N_3030);
or UO_433 (O_433,N_4170,N_4599);
xor UO_434 (O_434,N_4822,N_4352);
and UO_435 (O_435,N_4313,N_2554);
xnor UO_436 (O_436,N_3450,N_4008);
and UO_437 (O_437,N_3730,N_3483);
xnor UO_438 (O_438,N_4335,N_3221);
xnor UO_439 (O_439,N_3453,N_2735);
or UO_440 (O_440,N_2946,N_2746);
nor UO_441 (O_441,N_3667,N_3135);
xor UO_442 (O_442,N_2721,N_4590);
and UO_443 (O_443,N_4388,N_3676);
xor UO_444 (O_444,N_4382,N_3771);
nor UO_445 (O_445,N_3522,N_2900);
xor UO_446 (O_446,N_4259,N_4492);
nand UO_447 (O_447,N_2842,N_3932);
or UO_448 (O_448,N_4182,N_2996);
nor UO_449 (O_449,N_3839,N_2645);
xnor UO_450 (O_450,N_3691,N_4040);
nand UO_451 (O_451,N_2583,N_2919);
and UO_452 (O_452,N_3251,N_4445);
nand UO_453 (O_453,N_4240,N_4394);
nand UO_454 (O_454,N_3284,N_3865);
or UO_455 (O_455,N_2602,N_3604);
xnor UO_456 (O_456,N_2779,N_4139);
xor UO_457 (O_457,N_2561,N_3912);
nor UO_458 (O_458,N_2825,N_3978);
xnor UO_459 (O_459,N_4380,N_2601);
nor UO_460 (O_460,N_4404,N_2514);
xor UO_461 (O_461,N_4860,N_2952);
nor UO_462 (O_462,N_3424,N_2915);
nand UO_463 (O_463,N_3614,N_3127);
and UO_464 (O_464,N_4212,N_3269);
nor UO_465 (O_465,N_2969,N_2642);
or UO_466 (O_466,N_3390,N_3326);
or UO_467 (O_467,N_3623,N_4158);
nor UO_468 (O_468,N_4887,N_4819);
or UO_469 (O_469,N_3014,N_4528);
nand UO_470 (O_470,N_3892,N_2780);
xnor UO_471 (O_471,N_3729,N_4984);
nand UO_472 (O_472,N_4746,N_4038);
or UO_473 (O_473,N_4745,N_3709);
and UO_474 (O_474,N_3443,N_4278);
or UO_475 (O_475,N_4145,N_3160);
or UO_476 (O_476,N_2697,N_4496);
or UO_477 (O_477,N_3436,N_4529);
or UO_478 (O_478,N_2809,N_4181);
or UO_479 (O_479,N_3775,N_4375);
nand UO_480 (O_480,N_4754,N_3673);
nor UO_481 (O_481,N_4296,N_2558);
nor UO_482 (O_482,N_3193,N_4320);
nor UO_483 (O_483,N_3903,N_3760);
or UO_484 (O_484,N_3109,N_3680);
xor UO_485 (O_485,N_3053,N_2770);
and UO_486 (O_486,N_4956,N_2540);
xnor UO_487 (O_487,N_4302,N_3149);
xnor UO_488 (O_488,N_2652,N_4696);
nand UO_489 (O_489,N_2691,N_4864);
or UO_490 (O_490,N_4546,N_2626);
and UO_491 (O_491,N_3125,N_4749);
xnor UO_492 (O_492,N_3637,N_3772);
xor UO_493 (O_493,N_4904,N_4281);
or UO_494 (O_494,N_3555,N_4046);
and UO_495 (O_495,N_3696,N_2843);
nor UO_496 (O_496,N_4045,N_3953);
xor UO_497 (O_497,N_2590,N_4508);
nand UO_498 (O_498,N_4043,N_4726);
xor UO_499 (O_499,N_3857,N_2993);
nor UO_500 (O_500,N_4960,N_4748);
and UO_501 (O_501,N_2712,N_2550);
and UO_502 (O_502,N_4609,N_4386);
nor UO_503 (O_503,N_4730,N_4896);
or UO_504 (O_504,N_2516,N_4381);
or UO_505 (O_505,N_3553,N_4606);
nand UO_506 (O_506,N_2880,N_3072);
or UO_507 (O_507,N_3297,N_4586);
nor UO_508 (O_508,N_4168,N_4096);
xnor UO_509 (O_509,N_4371,N_2802);
and UO_510 (O_510,N_2731,N_2787);
nor UO_511 (O_511,N_3005,N_2620);
nor UO_512 (O_512,N_2876,N_4084);
or UO_513 (O_513,N_4699,N_4358);
or UO_514 (O_514,N_3140,N_4187);
xnor UO_515 (O_515,N_4365,N_4230);
nand UO_516 (O_516,N_4625,N_4996);
nand UO_517 (O_517,N_3677,N_2616);
nor UO_518 (O_518,N_4188,N_2719);
nand UO_519 (O_519,N_3946,N_2945);
xor UO_520 (O_520,N_2713,N_3806);
and UO_521 (O_521,N_4592,N_3869);
nand UO_522 (O_522,N_4156,N_4687);
nand UO_523 (O_523,N_2768,N_3734);
xnor UO_524 (O_524,N_3187,N_3276);
and UO_525 (O_525,N_4488,N_4804);
xnor UO_526 (O_526,N_2605,N_3195);
xor UO_527 (O_527,N_2752,N_3378);
or UO_528 (O_528,N_4736,N_4285);
and UO_529 (O_529,N_2978,N_3004);
or UO_530 (O_530,N_4507,N_4073);
or UO_531 (O_531,N_3170,N_4077);
or UO_532 (O_532,N_3765,N_4581);
or UO_533 (O_533,N_2508,N_2510);
nor UO_534 (O_534,N_3007,N_3958);
nor UO_535 (O_535,N_4542,N_3343);
xor UO_536 (O_536,N_3333,N_4076);
nor UO_537 (O_537,N_3476,N_3288);
and UO_538 (O_538,N_4558,N_2595);
or UO_539 (O_539,N_4078,N_4894);
nand UO_540 (O_540,N_3361,N_3801);
xor UO_541 (O_541,N_4410,N_4767);
xor UO_542 (O_542,N_2760,N_3363);
xnor UO_543 (O_543,N_3830,N_3826);
nand UO_544 (O_544,N_4054,N_3011);
and UO_545 (O_545,N_2957,N_3653);
nor UO_546 (O_546,N_3037,N_3303);
xnor UO_547 (O_547,N_3268,N_3675);
nand UO_548 (O_548,N_4659,N_4889);
xnor UO_549 (O_549,N_3883,N_3382);
and UO_550 (O_550,N_4340,N_2737);
xnor UO_551 (O_551,N_4770,N_4519);
or UO_552 (O_552,N_3585,N_2906);
nand UO_553 (O_553,N_2623,N_4941);
or UO_554 (O_554,N_3231,N_2627);
and UO_555 (O_555,N_4456,N_3494);
nand UO_556 (O_556,N_4042,N_2557);
nand UO_557 (O_557,N_3619,N_4588);
and UO_558 (O_558,N_2587,N_3006);
or UO_559 (O_559,N_4446,N_3821);
nand UO_560 (O_560,N_4511,N_4070);
and UO_561 (O_561,N_4512,N_4215);
xor UO_562 (O_562,N_2751,N_4439);
or UO_563 (O_563,N_3841,N_2791);
and UO_564 (O_564,N_2576,N_4355);
and UO_565 (O_565,N_4814,N_3761);
and UO_566 (O_566,N_3351,N_4074);
and UO_567 (O_567,N_2845,N_3102);
or UO_568 (O_568,N_4440,N_2750);
nor UO_569 (O_569,N_3907,N_3407);
and UO_570 (O_570,N_3366,N_3155);
and UO_571 (O_571,N_2987,N_3773);
or UO_572 (O_572,N_4199,N_2807);
or UO_573 (O_573,N_4103,N_2763);
or UO_574 (O_574,N_4083,N_4426);
or UO_575 (O_575,N_2526,N_4829);
nand UO_576 (O_576,N_4275,N_2847);
nand UO_577 (O_577,N_4785,N_4725);
xnor UO_578 (O_578,N_2930,N_3298);
xnor UO_579 (O_579,N_3855,N_3057);
xnor UO_580 (O_580,N_3349,N_4105);
nand UO_581 (O_581,N_4989,N_4729);
nand UO_582 (O_582,N_4616,N_3560);
nor UO_583 (O_583,N_4532,N_2934);
xnor UO_584 (O_584,N_2674,N_2936);
xor UO_585 (O_585,N_3047,N_4150);
and UO_586 (O_586,N_3510,N_3665);
nand UO_587 (O_587,N_4210,N_2565);
xor UO_588 (O_588,N_3612,N_4795);
or UO_589 (O_589,N_3397,N_4493);
nand UO_590 (O_590,N_2543,N_4533);
nand UO_591 (O_591,N_4279,N_4800);
xnor UO_592 (O_592,N_3639,N_4975);
nand UO_593 (O_593,N_2861,N_3134);
or UO_594 (O_594,N_4418,N_2738);
xnor UO_595 (O_595,N_4914,N_2884);
nor UO_596 (O_596,N_4413,N_4858);
nor UO_597 (O_597,N_3171,N_4100);
or UO_598 (O_598,N_4238,N_4483);
or UO_599 (O_599,N_4824,N_4884);
and UO_600 (O_600,N_2834,N_3461);
nand UO_601 (O_601,N_3836,N_4223);
nor UO_602 (O_602,N_3307,N_2638);
nand UO_603 (O_603,N_3909,N_4305);
xnor UO_604 (O_604,N_4969,N_2534);
nor UO_605 (O_605,N_2739,N_2806);
or UO_606 (O_606,N_3423,N_2650);
xor UO_607 (O_607,N_3473,N_3976);
xnor UO_608 (O_608,N_3644,N_4663);
nand UO_609 (O_609,N_4151,N_4306);
and UO_610 (O_610,N_3038,N_3154);
nor UO_611 (O_611,N_4142,N_4783);
or UO_612 (O_612,N_4449,N_4152);
and UO_613 (O_613,N_3521,N_4786);
and UO_614 (O_614,N_4286,N_2988);
and UO_615 (O_615,N_3049,N_4193);
or UO_616 (O_616,N_3282,N_4538);
nor UO_617 (O_617,N_2647,N_2865);
nand UO_618 (O_618,N_4778,N_4277);
nor UO_619 (O_619,N_4378,N_4593);
xnor UO_620 (O_620,N_4067,N_3746);
xnor UO_621 (O_621,N_2628,N_2640);
and UO_622 (O_622,N_4973,N_3845);
nand UO_623 (O_623,N_2893,N_3255);
xor UO_624 (O_624,N_3695,N_4028);
or UO_625 (O_625,N_3427,N_4265);
or UO_626 (O_626,N_3837,N_4460);
nand UO_627 (O_627,N_3460,N_3588);
and UO_628 (O_628,N_4878,N_2849);
and UO_629 (O_629,N_3441,N_3918);
or UO_630 (O_630,N_3292,N_3137);
nand UO_631 (O_631,N_4849,N_2914);
xor UO_632 (O_632,N_3050,N_3982);
xor UO_633 (O_633,N_3743,N_3161);
nand UO_634 (O_634,N_4872,N_3173);
nand UO_635 (O_635,N_4792,N_3464);
or UO_636 (O_636,N_4957,N_4667);
or UO_637 (O_637,N_4867,N_2916);
or UO_638 (O_638,N_4777,N_3277);
or UO_639 (O_639,N_2593,N_3916);
nor UO_640 (O_640,N_4323,N_2644);
nand UO_641 (O_641,N_3905,N_4485);
and UO_642 (O_642,N_4731,N_2753);
xor UO_643 (O_643,N_4097,N_2698);
nand UO_644 (O_644,N_2749,N_3128);
or UO_645 (O_645,N_4329,N_3043);
xor UO_646 (O_646,N_4722,N_3094);
or UO_647 (O_647,N_3829,N_3944);
xnor UO_648 (O_648,N_3986,N_4290);
or UO_649 (O_649,N_3929,N_3341);
nand UO_650 (O_650,N_3024,N_4796);
nor UO_651 (O_651,N_4138,N_4970);
nor UO_652 (O_652,N_4419,N_3593);
and UO_653 (O_653,N_4360,N_3646);
nor UO_654 (O_654,N_3223,N_3420);
and UO_655 (O_655,N_2976,N_4547);
xor UO_656 (O_656,N_2718,N_3900);
nand UO_657 (O_657,N_2597,N_3447);
nand UO_658 (O_658,N_3113,N_4467);
nand UO_659 (O_659,N_3818,N_4447);
and UO_660 (O_660,N_3316,N_4629);
and UO_661 (O_661,N_4091,N_3888);
and UO_662 (O_662,N_2844,N_4854);
nor UO_663 (O_663,N_3556,N_4377);
nor UO_664 (O_664,N_3849,N_3487);
xnor UO_665 (O_665,N_2663,N_4574);
or UO_666 (O_666,N_3152,N_3224);
nand UO_667 (O_667,N_4643,N_4612);
nand UO_668 (O_668,N_4050,N_3502);
xnor UO_669 (O_669,N_3294,N_3992);
nand UO_670 (O_670,N_3350,N_4933);
nand UO_671 (O_671,N_3572,N_3643);
xnor UO_672 (O_672,N_3881,N_4033);
or UO_673 (O_673,N_3262,N_3689);
or UO_674 (O_674,N_4713,N_4689);
nor UO_675 (O_675,N_3200,N_2710);
nor UO_676 (O_676,N_2524,N_3509);
xor UO_677 (O_677,N_3227,N_2857);
and UO_678 (O_678,N_2665,N_3713);
or UO_679 (O_679,N_4505,N_4165);
or UO_680 (O_680,N_3723,N_2734);
and UO_681 (O_681,N_4759,N_2973);
nor UO_682 (O_682,N_4551,N_4211);
and UO_683 (O_683,N_3107,N_3210);
nor UO_684 (O_684,N_4506,N_3649);
xnor UO_685 (O_685,N_2991,N_3552);
or UO_686 (O_686,N_2926,N_4755);
nand UO_687 (O_687,N_4998,N_4350);
xnor UO_688 (O_688,N_3948,N_3358);
nand UO_689 (O_689,N_2895,N_3027);
and UO_690 (O_690,N_2686,N_2769);
xor UO_691 (O_691,N_2507,N_3527);
or UO_692 (O_692,N_4900,N_4861);
nand UO_693 (O_693,N_3369,N_4384);
and UO_694 (O_694,N_2929,N_4462);
xor UO_695 (O_695,N_2892,N_2877);
xor UO_696 (O_696,N_3520,N_4299);
and UO_697 (O_697,N_3606,N_2533);
nand UO_698 (O_698,N_2908,N_3678);
xnor UO_699 (O_699,N_2823,N_4441);
nor UO_700 (O_700,N_4174,N_4660);
and UO_701 (O_701,N_3706,N_3715);
nand UO_702 (O_702,N_4623,N_4567);
nor UO_703 (O_703,N_3651,N_2548);
and UO_704 (O_704,N_3250,N_3807);
xnor UO_705 (O_705,N_3752,N_4661);
nand UO_706 (O_706,N_4143,N_3101);
or UO_707 (O_707,N_3279,N_4163);
or UO_708 (O_708,N_3375,N_3477);
xnor UO_709 (O_709,N_4075,N_4021);
nor UO_710 (O_710,N_2819,N_3493);
xnor UO_711 (O_711,N_2761,N_2911);
xnor UO_712 (O_712,N_2866,N_4264);
nand UO_713 (O_713,N_3596,N_4147);
xnor UO_714 (O_714,N_3962,N_4334);
and UO_715 (O_715,N_3348,N_3042);
and UO_716 (O_716,N_3587,N_2568);
nor UO_717 (O_717,N_4303,N_3563);
and UO_718 (O_718,N_3749,N_2538);
nand UO_719 (O_719,N_4025,N_4195);
nor UO_720 (O_720,N_4020,N_4336);
or UO_721 (O_721,N_3468,N_4262);
and UO_722 (O_722,N_4131,N_2553);
nor UO_723 (O_723,N_2677,N_4565);
and UO_724 (O_724,N_3082,N_4247);
and UO_725 (O_725,N_4718,N_4484);
xnor UO_726 (O_726,N_4680,N_3809);
nor UO_727 (O_727,N_4762,N_4879);
xnor UO_728 (O_728,N_4209,N_4976);
xnor UO_729 (O_729,N_3599,N_2544);
nand UO_730 (O_730,N_3415,N_4740);
and UO_731 (O_731,N_4557,N_2633);
xnor UO_732 (O_732,N_3756,N_4597);
xnor UO_733 (O_733,N_4857,N_3188);
and UO_734 (O_734,N_4192,N_4416);
nand UO_735 (O_735,N_4626,N_3238);
nand UO_736 (O_736,N_2722,N_3347);
nor UO_737 (O_737,N_3281,N_4311);
and UO_738 (O_738,N_3377,N_3458);
or UO_739 (O_739,N_4856,N_4159);
and UO_740 (O_740,N_3029,N_3402);
or UO_741 (O_741,N_4030,N_4681);
nor UO_742 (O_742,N_4310,N_3663);
or UO_743 (O_743,N_4635,N_3528);
or UO_744 (O_744,N_4009,N_4554);
and UO_745 (O_745,N_4534,N_2619);
and UO_746 (O_746,N_4461,N_3467);
and UO_747 (O_747,N_2937,N_4179);
nand UO_748 (O_748,N_4464,N_4249);
and UO_749 (O_749,N_3988,N_3739);
nor UO_750 (O_750,N_4595,N_3144);
and UO_751 (O_751,N_4012,N_4753);
nor UO_752 (O_752,N_3076,N_4580);
and UO_753 (O_753,N_4834,N_2562);
xnor UO_754 (O_754,N_4855,N_3067);
nor UO_755 (O_755,N_3959,N_3387);
or UO_756 (O_756,N_2621,N_3968);
or UO_757 (O_757,N_4123,N_3122);
and UO_758 (O_758,N_4537,N_4832);
xor UO_759 (O_759,N_4690,N_4619);
nand UO_760 (O_760,N_4802,N_3618);
or UO_761 (O_761,N_4539,N_4784);
or UO_762 (O_762,N_2520,N_3668);
nor UO_763 (O_763,N_4363,N_4186);
xor UO_764 (O_764,N_4917,N_2881);
nand UO_765 (O_765,N_2699,N_4912);
xnor UO_766 (O_766,N_3087,N_4963);
xor UO_767 (O_767,N_2655,N_2967);
xor UO_768 (O_768,N_3987,N_4578);
nand UO_769 (O_769,N_4540,N_2989);
and UO_770 (O_770,N_4095,N_3272);
nor UO_771 (O_771,N_4535,N_4274);
and UO_772 (O_772,N_3071,N_3716);
nor UO_773 (O_773,N_3626,N_3568);
xor UO_774 (O_774,N_3226,N_4945);
nor UO_775 (O_775,N_2574,N_4072);
or UO_776 (O_776,N_3385,N_2502);
xor UO_777 (O_777,N_3048,N_4705);
and UO_778 (O_778,N_3631,N_4237);
xor UO_779 (O_779,N_3194,N_3404);
nor UO_780 (O_780,N_4728,N_3645);
and UO_781 (O_781,N_3936,N_2772);
nand UO_782 (O_782,N_2707,N_4273);
nor UO_783 (O_783,N_4943,N_4573);
or UO_784 (O_784,N_3545,N_3742);
and UO_785 (O_785,N_4655,N_4000);
nand UO_786 (O_786,N_4932,N_3069);
nor UO_787 (O_787,N_2736,N_3229);
or UO_788 (O_788,N_4890,N_2732);
nand UO_789 (O_789,N_3012,N_4205);
or UO_790 (O_790,N_4620,N_2970);
or UO_791 (O_791,N_4373,N_4503);
or UO_792 (O_792,N_3956,N_2681);
or UO_793 (O_793,N_3949,N_3951);
xor UO_794 (O_794,N_4090,N_4587);
nor UO_795 (O_795,N_3261,N_3627);
and UO_796 (O_796,N_3871,N_3762);
xnor UO_797 (O_797,N_4234,N_3590);
xnor UO_798 (O_798,N_3764,N_3641);
nor UO_799 (O_799,N_3886,N_4600);
or UO_800 (O_800,N_4553,N_2671);
xnor UO_801 (O_801,N_4217,N_3329);
or UO_802 (O_802,N_3388,N_3741);
nor UO_803 (O_803,N_4246,N_2505);
or UO_804 (O_804,N_2854,N_4171);
xnor UO_805 (O_805,N_3957,N_3000);
xor UO_806 (O_806,N_3725,N_3001);
nand UO_807 (O_807,N_4582,N_2997);
nand UO_808 (O_808,N_4931,N_4817);
and UO_809 (O_809,N_3512,N_2573);
and UO_810 (O_810,N_3890,N_3046);
nand UO_811 (O_811,N_4177,N_3365);
xnor UO_812 (O_812,N_3073,N_3727);
nor UO_813 (O_813,N_4448,N_4607);
xnor UO_814 (O_814,N_4952,N_3784);
or UO_815 (O_815,N_3777,N_3805);
and UO_816 (O_816,N_4455,N_3511);
nor UO_817 (O_817,N_3335,N_2701);
or UO_818 (O_818,N_4214,N_2788);
or UO_819 (O_819,N_3783,N_4298);
xnor UO_820 (O_820,N_4640,N_4490);
or UO_821 (O_821,N_4086,N_4060);
nor UO_822 (O_822,N_2873,N_2541);
nor UO_823 (O_823,N_3457,N_3103);
or UO_824 (O_824,N_3237,N_3894);
nor UO_825 (O_825,N_4059,N_3220);
and UO_826 (O_826,N_3891,N_3063);
nor UO_827 (O_827,N_3254,N_3799);
nand UO_828 (O_828,N_4714,N_4788);
nand UO_829 (O_829,N_4427,N_3019);
or UO_830 (O_830,N_2922,N_4801);
nor UO_831 (O_831,N_4921,N_4189);
and UO_832 (O_832,N_2610,N_2764);
nor UO_833 (O_833,N_4615,N_3814);
and UO_834 (O_834,N_2949,N_3147);
nor UO_835 (O_835,N_2966,N_3373);
and UO_836 (O_836,N_3260,N_3688);
or UO_837 (O_837,N_2905,N_4322);
xor UO_838 (O_838,N_4411,N_2848);
and UO_839 (O_839,N_3832,N_4087);
or UO_840 (O_840,N_3506,N_4284);
nor UO_841 (O_841,N_3286,N_3219);
nor UO_842 (O_842,N_3554,N_2513);
nand UO_843 (O_843,N_2758,N_4962);
nand UO_844 (O_844,N_2827,N_3580);
or UO_845 (O_845,N_3309,N_4618);
and UO_846 (O_846,N_4815,N_3708);
nand UO_847 (O_847,N_3334,N_3384);
nor UO_848 (O_848,N_4366,N_3243);
or UO_849 (O_849,N_2784,N_3031);
or UO_850 (O_850,N_4876,N_4678);
nor UO_851 (O_851,N_4961,N_3399);
nand UO_852 (O_852,N_3666,N_2960);
and UO_853 (O_853,N_2517,N_3065);
nand UO_854 (O_854,N_4482,N_2635);
nor UO_855 (O_855,N_4776,N_3851);
or UO_856 (O_856,N_4779,N_4869);
or UO_857 (O_857,N_2668,N_4118);
nand UO_858 (O_858,N_4065,N_4611);
or UO_859 (O_859,N_4063,N_4454);
nand UO_860 (O_860,N_2816,N_3395);
and UO_861 (O_861,N_4724,N_2851);
xnor UO_862 (O_862,N_2789,N_4098);
and UO_863 (O_863,N_3754,N_4130);
nor UO_864 (O_864,N_3564,N_3535);
and UO_865 (O_865,N_4491,N_3035);
nor UO_866 (O_866,N_3795,N_3833);
or UO_867 (O_867,N_3475,N_4799);
xor UO_868 (O_868,N_3086,N_3044);
xor UO_869 (O_869,N_4685,N_3835);
nand UO_870 (O_870,N_4013,N_3990);
xor UO_871 (O_871,N_3442,N_4463);
xnor UO_872 (O_872,N_3672,N_4140);
xor UO_873 (O_873,N_3838,N_3328);
xnor UO_874 (O_874,N_4396,N_3621);
xnor UO_875 (O_875,N_3058,N_4704);
xor UO_876 (O_876,N_3077,N_3796);
or UO_877 (O_877,N_4624,N_3417);
xnor UO_878 (O_878,N_2864,N_4104);
and UO_879 (O_879,N_3488,N_4198);
nand UO_880 (O_880,N_3336,N_3429);
xnor UO_881 (O_881,N_3185,N_3002);
nand UO_882 (O_882,N_3977,N_4315);
and UO_883 (O_883,N_4051,N_4129);
and UO_884 (O_884,N_2928,N_3331);
and UO_885 (O_885,N_3148,N_3482);
nand UO_886 (O_886,N_3701,N_4898);
nand UO_887 (O_887,N_3694,N_3770);
or UO_888 (O_888,N_4845,N_4019);
xnor UO_889 (O_889,N_4908,N_2886);
nor UO_890 (O_890,N_3872,N_3313);
and UO_891 (O_891,N_3166,N_2931);
or UO_892 (O_892,N_4826,N_4513);
and UO_893 (O_893,N_2748,N_3426);
nor UO_894 (O_894,N_3133,N_4231);
nand UO_895 (O_895,N_4213,N_4781);
xnor UO_896 (O_896,N_2765,N_2887);
and UO_897 (O_897,N_3023,N_2596);
nand UO_898 (O_898,N_3320,N_3538);
nand UO_899 (O_899,N_4562,N_3825);
nand UO_900 (O_900,N_2979,N_4134);
nand UO_901 (O_901,N_4946,N_2547);
and UO_902 (O_902,N_3931,N_3707);
nand UO_903 (O_903,N_3726,N_3401);
nor UO_904 (O_904,N_4545,N_4227);
nand UO_905 (O_905,N_2688,N_2782);
xor UO_906 (O_906,N_3163,N_2958);
or UO_907 (O_907,N_4823,N_3682);
nand UO_908 (O_908,N_2521,N_2723);
and UO_909 (O_909,N_2850,N_4326);
xor UO_910 (O_910,N_2607,N_3300);
xnor UO_911 (O_911,N_4354,N_3213);
or UO_912 (O_912,N_4486,N_3222);
nor UO_913 (O_913,N_3975,N_2986);
and UO_914 (O_914,N_4301,N_3543);
nor UO_915 (O_915,N_3583,N_2812);
nand UO_916 (O_916,N_4167,N_4161);
nor UO_917 (O_917,N_4927,N_4341);
nand UO_918 (O_918,N_3283,N_3235);
and UO_919 (O_919,N_3513,N_3638);
nand UO_920 (O_920,N_2796,N_3943);
or UO_921 (O_921,N_4347,N_4376);
nor UO_922 (O_922,N_4112,N_3600);
nor UO_923 (O_923,N_3327,N_3526);
and UO_924 (O_924,N_4133,N_4897);
and UO_925 (O_925,N_4149,N_4173);
nand UO_926 (O_926,N_3937,N_3104);
nand UO_927 (O_927,N_2662,N_3759);
and UO_928 (O_928,N_3960,N_4117);
nand UO_929 (O_929,N_3514,N_4036);
nor UO_930 (O_930,N_4742,N_3919);
xnor UO_931 (O_931,N_4436,N_4536);
or UO_932 (O_932,N_3275,N_4710);
xor UO_933 (O_933,N_2995,N_2774);
nor UO_934 (O_934,N_4734,N_3362);
nor UO_935 (O_935,N_3609,N_2830);
or UO_936 (O_936,N_3581,N_2637);
and UO_937 (O_937,N_3108,N_3763);
and UO_938 (O_938,N_3466,N_4392);
and UO_939 (O_939,N_3797,N_3893);
nor UO_940 (O_940,N_4572,N_3084);
or UO_941 (O_941,N_3980,N_3150);
and UO_942 (O_942,N_2985,N_4743);
nand UO_943 (O_943,N_2702,N_4120);
nand UO_944 (O_944,N_3064,N_2910);
or UO_945 (O_945,N_3594,N_3517);
and UO_946 (O_946,N_4153,N_3396);
xor UO_947 (O_947,N_3997,N_3697);
and UO_948 (O_948,N_2717,N_3808);
nor UO_949 (O_949,N_3271,N_2694);
or UO_950 (O_950,N_3263,N_2563);
xnor UO_951 (O_951,N_3831,N_3620);
nand UO_952 (O_952,N_2515,N_4423);
or UO_953 (O_953,N_3240,N_2648);
nand UO_954 (O_954,N_4201,N_2618);
xnor UO_955 (O_955,N_2829,N_3970);
nor UO_956 (O_956,N_4837,N_4988);
nor UO_957 (O_957,N_2817,N_3622);
or UO_958 (O_958,N_4662,N_4297);
nor UO_959 (O_959,N_4739,N_3116);
and UO_960 (O_960,N_4664,N_3470);
nand UO_961 (O_961,N_3183,N_2622);
and UO_962 (O_962,N_2608,N_3165);
xnor UO_963 (O_963,N_3345,N_4316);
nand UO_964 (O_964,N_4185,N_3099);
xnor UO_965 (O_965,N_3719,N_2777);
and UO_966 (O_966,N_4905,N_3124);
xor UO_967 (O_967,N_3530,N_4720);
and UO_968 (O_968,N_3146,N_3702);
xnor UO_969 (O_969,N_4472,N_3964);
or UO_970 (O_970,N_4514,N_3700);
nor UO_971 (O_971,N_4641,N_3889);
nor UO_972 (O_972,N_4866,N_2948);
xnor UO_973 (O_973,N_3130,N_2888);
nand UO_974 (O_974,N_3306,N_3406);
and UO_975 (O_975,N_4243,N_4654);
nand UO_976 (O_976,N_4682,N_4421);
and UO_977 (O_977,N_4443,N_3118);
and UO_978 (O_978,N_4980,N_4719);
xor UO_979 (O_979,N_4191,N_4702);
and UO_980 (O_980,N_2814,N_2955);
or UO_981 (O_981,N_4102,N_3601);
xnor UO_982 (O_982,N_3917,N_4125);
or UO_983 (O_983,N_2965,N_4489);
nand UO_984 (O_984,N_2805,N_4893);
xnor UO_985 (O_985,N_3947,N_2500);
or UO_986 (O_986,N_4408,N_3485);
or UO_987 (O_987,N_4928,N_3409);
xor UO_988 (O_988,N_3875,N_3056);
nor UO_989 (O_989,N_3003,N_3182);
or UO_990 (O_990,N_4452,N_3017);
and UO_991 (O_991,N_4671,N_4634);
and UO_992 (O_992,N_3915,N_4677);
nand UO_993 (O_993,N_4475,N_4024);
nand UO_994 (O_994,N_4272,N_3293);
or UO_995 (O_995,N_4356,N_3703);
or UO_996 (O_996,N_2894,N_4575);
nand UO_997 (O_997,N_2875,N_3540);
or UO_998 (O_998,N_4056,N_2546);
nand UO_999 (O_999,N_4524,N_3111);
endmodule