module basic_500_3000_500_40_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_182,In_472);
nor U1 (N_1,In_69,In_240);
nor U2 (N_2,In_63,In_344);
nand U3 (N_3,In_254,In_198);
xor U4 (N_4,In_231,In_28);
xor U5 (N_5,In_295,In_61);
xnor U6 (N_6,In_272,In_477);
or U7 (N_7,In_380,In_283);
and U8 (N_8,In_307,In_335);
nor U9 (N_9,In_441,In_378);
nor U10 (N_10,In_245,In_392);
nor U11 (N_11,In_127,In_442);
nor U12 (N_12,In_81,In_376);
or U13 (N_13,In_457,In_166);
nor U14 (N_14,In_150,In_184);
and U15 (N_15,In_149,In_249);
or U16 (N_16,In_188,In_32);
nand U17 (N_17,In_1,In_93);
nor U18 (N_18,In_315,In_320);
xnor U19 (N_19,In_204,In_257);
and U20 (N_20,In_41,In_387);
or U21 (N_21,In_160,In_403);
nand U22 (N_22,In_480,In_148);
nand U23 (N_23,In_416,In_87);
and U24 (N_24,In_465,In_0);
xnor U25 (N_25,In_132,In_317);
xor U26 (N_26,In_43,In_489);
or U27 (N_27,In_205,In_481);
nor U28 (N_28,In_492,In_45);
or U29 (N_29,In_121,In_279);
nand U30 (N_30,In_299,In_202);
and U31 (N_31,In_330,In_95);
or U32 (N_32,In_301,In_277);
nand U33 (N_33,In_448,In_39);
or U34 (N_34,In_106,In_181);
and U35 (N_35,In_8,In_417);
nor U36 (N_36,In_208,In_109);
nand U37 (N_37,In_209,In_14);
and U38 (N_38,In_398,In_3);
or U39 (N_39,In_185,In_348);
or U40 (N_40,In_289,In_101);
and U41 (N_41,In_88,In_247);
nor U42 (N_42,In_33,In_196);
nand U43 (N_43,In_62,In_18);
or U44 (N_44,In_321,In_189);
nand U45 (N_45,In_130,In_175);
and U46 (N_46,In_486,In_42);
nor U47 (N_47,In_158,In_303);
or U48 (N_48,In_490,In_375);
nor U49 (N_49,In_54,In_355);
and U50 (N_50,In_397,In_74);
xor U51 (N_51,In_329,In_225);
xnor U52 (N_52,In_268,In_361);
nand U53 (N_53,In_30,In_219);
nand U54 (N_54,In_169,In_459);
nor U55 (N_55,In_298,In_126);
nor U56 (N_56,In_168,In_341);
or U57 (N_57,In_151,In_222);
nand U58 (N_58,In_186,In_293);
and U59 (N_59,In_82,In_5);
or U60 (N_60,In_412,In_428);
nor U61 (N_61,In_36,In_438);
nor U62 (N_62,In_450,In_493);
nor U63 (N_63,In_286,In_164);
and U64 (N_64,In_461,In_242);
xor U65 (N_65,In_20,In_251);
nand U66 (N_66,In_64,In_367);
nand U67 (N_67,In_328,In_83);
xnor U68 (N_68,In_302,In_396);
nor U69 (N_69,In_129,In_227);
nand U70 (N_70,In_345,In_498);
or U71 (N_71,In_437,In_371);
nand U72 (N_72,In_294,In_75);
and U73 (N_73,In_53,In_468);
and U74 (N_74,In_147,In_260);
and U75 (N_75,In_218,In_115);
or U76 (N_76,In_449,In_309);
nor U77 (N_77,N_55,N_29);
nand U78 (N_78,In_57,In_215);
nand U79 (N_79,In_281,In_259);
xnor U80 (N_80,In_216,In_278);
and U81 (N_81,In_60,N_17);
or U82 (N_82,In_306,In_84);
and U83 (N_83,In_58,In_25);
nand U84 (N_84,In_10,In_167);
nor U85 (N_85,In_273,In_452);
and U86 (N_86,N_11,In_340);
nor U87 (N_87,N_3,N_2);
nand U88 (N_88,In_332,In_23);
nand U89 (N_89,N_22,In_390);
nand U90 (N_90,In_389,In_161);
or U91 (N_91,In_374,In_79);
nor U92 (N_92,In_19,N_50);
or U93 (N_93,In_322,N_32);
nor U94 (N_94,In_333,In_27);
nor U95 (N_95,In_234,In_427);
nor U96 (N_96,In_409,In_400);
or U97 (N_97,In_9,In_451);
xnor U98 (N_98,In_379,In_102);
xnor U99 (N_99,In_110,In_131);
and U100 (N_100,In_86,In_287);
xnor U101 (N_101,In_76,In_238);
nor U102 (N_102,In_71,N_43);
and U103 (N_103,In_433,In_313);
nand U104 (N_104,In_474,In_165);
xor U105 (N_105,In_246,In_214);
or U106 (N_106,In_37,In_112);
and U107 (N_107,In_352,In_159);
or U108 (N_108,In_310,In_155);
or U109 (N_109,In_235,In_192);
nor U110 (N_110,In_100,N_46);
nor U111 (N_111,In_407,In_264);
or U112 (N_112,In_404,In_377);
or U113 (N_113,In_173,In_402);
and U114 (N_114,N_70,In_228);
nand U115 (N_115,In_354,N_16);
and U116 (N_116,In_72,In_241);
or U117 (N_117,In_12,In_350);
or U118 (N_118,N_42,In_356);
or U119 (N_119,In_410,In_163);
and U120 (N_120,N_49,N_62);
nand U121 (N_121,In_316,In_68);
xnor U122 (N_122,In_203,In_141);
xnor U123 (N_123,In_323,In_291);
nand U124 (N_124,In_117,In_38);
or U125 (N_125,In_373,In_447);
nand U126 (N_126,In_445,In_276);
and U127 (N_127,In_491,In_48);
and U128 (N_128,In_466,In_221);
or U129 (N_129,N_24,In_462);
and U130 (N_130,In_52,In_419);
and U131 (N_131,In_467,In_207);
nor U132 (N_132,In_269,N_45);
nor U133 (N_133,In_334,In_363);
and U134 (N_134,N_31,In_156);
nor U135 (N_135,N_56,In_114);
nand U136 (N_136,In_134,N_1);
nand U137 (N_137,In_425,In_96);
nand U138 (N_138,In_103,In_7);
nand U139 (N_139,In_366,In_499);
and U140 (N_140,In_211,In_290);
or U141 (N_141,In_248,In_413);
and U142 (N_142,In_357,N_44);
nand U143 (N_143,In_411,In_267);
nor U144 (N_144,In_394,In_422);
and U145 (N_145,In_297,In_424);
nand U146 (N_146,In_194,In_78);
nor U147 (N_147,In_319,In_116);
nand U148 (N_148,In_40,In_51);
nand U149 (N_149,In_137,In_111);
or U150 (N_150,In_296,N_126);
and U151 (N_151,In_311,In_460);
nand U152 (N_152,N_112,In_59);
and U153 (N_153,In_31,N_100);
or U154 (N_154,N_147,In_342);
and U155 (N_155,In_372,N_4);
nor U156 (N_156,In_353,In_463);
xnor U157 (N_157,N_54,In_282);
nand U158 (N_158,N_60,In_262);
and U159 (N_159,N_79,N_130);
or U160 (N_160,In_142,N_129);
or U161 (N_161,N_34,In_244);
nand U162 (N_162,N_12,N_73);
or U163 (N_163,In_312,N_92);
or U164 (N_164,In_280,N_9);
nor U165 (N_165,In_469,N_83);
and U166 (N_166,In_258,In_50);
and U167 (N_167,N_82,N_104);
or U168 (N_168,In_201,In_210);
or U169 (N_169,In_261,In_152);
or U170 (N_170,In_29,In_21);
or U171 (N_171,In_243,N_128);
nor U172 (N_172,N_91,In_436);
nand U173 (N_173,N_48,In_16);
nand U174 (N_174,In_415,In_206);
and U175 (N_175,N_89,N_122);
or U176 (N_176,N_37,In_13);
or U177 (N_177,In_143,N_124);
or U178 (N_178,In_140,In_46);
nand U179 (N_179,In_300,In_343);
xnor U180 (N_180,N_117,In_232);
and U181 (N_181,In_431,In_420);
or U182 (N_182,N_40,N_97);
or U183 (N_183,In_146,In_446);
or U184 (N_184,In_133,In_395);
or U185 (N_185,In_108,In_80);
and U186 (N_186,In_144,N_144);
nor U187 (N_187,In_236,In_453);
or U188 (N_188,In_183,N_108);
xnor U189 (N_189,In_456,In_439);
and U190 (N_190,In_128,N_5);
and U191 (N_191,In_47,In_237);
and U192 (N_192,N_28,In_73);
and U193 (N_193,In_200,In_97);
nand U194 (N_194,N_138,In_94);
xnor U195 (N_195,N_137,N_65);
nor U196 (N_196,In_124,In_429);
nand U197 (N_197,N_57,N_98);
and U198 (N_198,In_263,In_275);
nor U199 (N_199,N_0,In_107);
or U200 (N_200,N_63,In_253);
xor U201 (N_201,N_36,In_135);
nor U202 (N_202,In_191,In_265);
xor U203 (N_203,In_2,In_358);
nor U204 (N_204,N_23,N_68);
or U205 (N_205,N_30,In_125);
nor U206 (N_206,N_88,N_148);
and U207 (N_207,In_136,N_102);
nand U208 (N_208,N_66,In_67);
nand U209 (N_209,In_351,N_38);
nor U210 (N_210,In_418,N_51);
xnor U211 (N_211,In_172,N_84);
nor U212 (N_212,In_360,In_223);
or U213 (N_213,In_113,N_86);
nand U214 (N_214,N_107,In_44);
and U215 (N_215,In_370,N_90);
or U216 (N_216,In_66,In_495);
nor U217 (N_217,In_34,N_145);
or U218 (N_218,In_22,In_440);
xor U219 (N_219,In_252,N_52);
nor U220 (N_220,In_180,In_17);
nor U221 (N_221,In_255,In_423);
nor U222 (N_222,In_230,N_96);
nor U223 (N_223,N_123,In_359);
or U224 (N_224,In_145,N_134);
or U225 (N_225,N_217,N_176);
or U226 (N_226,N_19,In_369);
and U227 (N_227,N_116,In_178);
nand U228 (N_228,In_483,In_271);
and U229 (N_229,N_163,In_157);
or U230 (N_230,In_365,N_14);
or U231 (N_231,In_385,In_386);
or U232 (N_232,N_216,In_346);
or U233 (N_233,In_89,N_64);
xnor U234 (N_234,N_140,N_109);
nor U235 (N_235,In_339,In_406);
and U236 (N_236,N_146,In_484);
and U237 (N_237,N_208,In_304);
or U238 (N_238,N_77,N_93);
nor U239 (N_239,In_193,In_405);
nor U240 (N_240,In_70,N_141);
nand U241 (N_241,In_92,In_393);
or U242 (N_242,N_224,In_414);
and U243 (N_243,In_364,N_189);
nor U244 (N_244,N_58,In_347);
nor U245 (N_245,In_11,N_158);
or U246 (N_246,N_206,N_215);
nand U247 (N_247,N_33,In_35);
nor U248 (N_248,In_270,N_121);
or U249 (N_249,N_188,N_143);
or U250 (N_250,In_105,In_368);
nand U251 (N_251,In_475,N_157);
nor U252 (N_252,N_185,In_226);
and U253 (N_253,N_25,In_213);
nand U254 (N_254,In_444,In_171);
nand U255 (N_255,N_207,N_67);
and U256 (N_256,In_326,N_172);
nand U257 (N_257,N_194,In_488);
xor U258 (N_258,N_131,N_203);
or U259 (N_259,In_308,N_155);
nor U260 (N_260,In_139,N_39);
or U261 (N_261,N_13,In_98);
nand U262 (N_262,N_149,N_59);
or U263 (N_263,N_182,In_464);
and U264 (N_264,N_159,In_256);
xor U265 (N_265,N_132,In_401);
nor U266 (N_266,N_166,In_496);
or U267 (N_267,N_75,N_150);
and U268 (N_268,In_494,N_113);
nor U269 (N_269,N_184,In_285);
or U270 (N_270,In_195,N_101);
and U271 (N_271,N_222,In_104);
nand U272 (N_272,N_178,In_331);
or U273 (N_273,In_482,N_127);
nor U274 (N_274,N_95,N_156);
nand U275 (N_275,N_164,In_176);
and U276 (N_276,In_327,N_175);
nor U277 (N_277,In_118,In_122);
xnor U278 (N_278,N_169,N_69);
nand U279 (N_279,N_171,In_65);
nor U280 (N_280,N_192,In_15);
nand U281 (N_281,In_314,N_118);
and U282 (N_282,In_470,N_209);
or U283 (N_283,In_408,N_7);
nand U284 (N_284,N_204,N_125);
and U285 (N_285,N_223,N_186);
nor U286 (N_286,In_388,N_35);
nor U287 (N_287,N_151,In_119);
or U288 (N_288,N_167,N_133);
or U289 (N_289,N_218,N_136);
nor U290 (N_290,N_180,N_154);
or U291 (N_291,N_221,N_15);
and U292 (N_292,In_485,N_106);
nor U293 (N_293,In_318,In_426);
nor U294 (N_294,N_27,N_193);
and U295 (N_295,N_200,In_56);
or U296 (N_296,N_162,N_161);
nor U297 (N_297,In_443,In_383);
nor U298 (N_298,N_119,In_476);
nand U299 (N_299,In_362,N_6);
or U300 (N_300,N_233,N_268);
nor U301 (N_301,In_274,N_257);
nor U302 (N_302,N_235,N_201);
or U303 (N_303,N_10,N_263);
or U304 (N_304,N_237,In_349);
nor U305 (N_305,N_280,N_135);
or U306 (N_306,In_384,N_295);
xor U307 (N_307,In_91,N_274);
or U308 (N_308,N_168,N_275);
and U309 (N_309,In_190,In_305);
nand U310 (N_310,N_241,In_162);
and U311 (N_311,N_259,N_8);
and U312 (N_312,In_338,In_49);
nand U313 (N_313,In_292,N_214);
or U314 (N_314,In_487,N_244);
or U315 (N_315,N_247,N_297);
nand U316 (N_316,In_220,In_432);
xor U317 (N_317,N_254,N_115);
and U318 (N_318,In_284,N_71);
or U319 (N_319,In_478,N_279);
nor U320 (N_320,In_233,In_250);
and U321 (N_321,N_291,N_212);
and U322 (N_322,N_179,N_210);
nand U323 (N_323,N_177,N_174);
nand U324 (N_324,N_197,In_90);
xnor U325 (N_325,N_284,N_41);
and U326 (N_326,N_99,In_99);
and U327 (N_327,N_242,N_74);
nor U328 (N_328,N_205,In_24);
nor U329 (N_329,N_271,N_281);
nand U330 (N_330,N_190,N_225);
nand U331 (N_331,N_260,N_298);
nand U332 (N_332,N_264,N_296);
and U333 (N_333,In_454,N_20);
and U334 (N_334,In_325,In_174);
nor U335 (N_335,N_255,N_85);
or U336 (N_336,N_211,N_272);
nor U337 (N_337,In_288,In_55);
and U338 (N_338,N_165,N_292);
nand U339 (N_339,In_430,N_262);
or U340 (N_340,N_18,N_273);
or U341 (N_341,In_138,N_170);
xor U342 (N_342,In_154,N_103);
nand U343 (N_343,In_212,N_267);
nand U344 (N_344,In_6,N_258);
nor U345 (N_345,N_72,N_202);
and U346 (N_346,In_473,In_399);
nor U347 (N_347,In_391,N_61);
nand U348 (N_348,N_243,N_266);
and U349 (N_349,N_246,N_277);
nand U350 (N_350,N_94,In_187);
xor U351 (N_351,N_249,N_230);
nor U352 (N_352,N_276,In_382);
nand U353 (N_353,N_105,N_181);
nor U354 (N_354,N_245,N_110);
nand U355 (N_355,In_123,N_228);
nand U356 (N_356,N_238,N_229);
nand U357 (N_357,In_421,N_261);
and U358 (N_358,N_219,N_285);
or U359 (N_359,In_26,In_266);
nor U360 (N_360,N_152,N_282);
nand U361 (N_361,N_139,N_251);
nand U362 (N_362,In_77,In_170);
or U363 (N_363,In_336,N_252);
nand U364 (N_364,N_278,In_435);
or U365 (N_365,In_434,N_294);
nor U366 (N_366,N_234,N_270);
and U367 (N_367,N_226,N_78);
and U368 (N_368,N_213,N_195);
nor U369 (N_369,N_293,In_381);
nor U370 (N_370,N_80,N_265);
xor U371 (N_371,N_111,In_199);
nand U372 (N_372,N_287,In_455);
nand U373 (N_373,N_53,In_153);
or U374 (N_374,N_142,In_458);
and U375 (N_375,N_358,N_356);
xor U376 (N_376,N_334,N_26);
nand U377 (N_377,N_196,N_324);
xnor U378 (N_378,N_240,N_310);
or U379 (N_379,N_302,N_372);
and U380 (N_380,N_220,N_288);
and U381 (N_381,N_374,N_250);
and U382 (N_382,In_85,N_239);
and U383 (N_383,N_114,N_349);
nand U384 (N_384,N_333,N_81);
and U385 (N_385,N_339,N_327);
and U386 (N_386,N_368,N_191);
nand U387 (N_387,N_236,In_337);
nor U388 (N_388,In_471,N_325);
nand U389 (N_389,N_364,N_76);
and U390 (N_390,N_283,N_231);
nand U391 (N_391,N_343,N_361);
or U392 (N_392,N_269,N_304);
nand U393 (N_393,N_329,N_352);
or U394 (N_394,In_224,N_306);
nor U395 (N_395,N_335,N_346);
nand U396 (N_396,In_197,N_301);
and U397 (N_397,N_47,In_217);
xor U398 (N_398,N_316,N_332);
and U399 (N_399,N_313,N_227);
xor U400 (N_400,N_303,In_479);
nor U401 (N_401,N_299,N_183);
or U402 (N_402,N_365,In_177);
or U403 (N_403,N_286,N_232);
nor U404 (N_404,N_371,N_320);
nand U405 (N_405,N_347,N_338);
and U406 (N_406,N_363,N_342);
nor U407 (N_407,N_21,N_351);
nor U408 (N_408,N_305,N_198);
and U409 (N_409,N_323,N_354);
and U410 (N_410,N_348,N_307);
nand U411 (N_411,N_341,N_199);
nand U412 (N_412,In_324,N_367);
nand U413 (N_413,N_340,N_289);
and U414 (N_414,N_300,N_330);
or U415 (N_415,N_359,N_187);
xor U416 (N_416,N_248,N_253);
nand U417 (N_417,In_4,N_326);
and U418 (N_418,N_357,N_120);
or U419 (N_419,N_331,In_179);
or U420 (N_420,N_311,N_312);
and U421 (N_421,N_355,N_328);
xnor U422 (N_422,N_319,N_336);
nand U423 (N_423,N_337,N_317);
and U424 (N_424,N_362,In_239);
nor U425 (N_425,N_373,N_370);
or U426 (N_426,N_366,N_315);
xnor U427 (N_427,In_229,N_345);
and U428 (N_428,N_314,N_318);
nor U429 (N_429,N_308,N_369);
and U430 (N_430,N_344,N_160);
or U431 (N_431,N_353,N_322);
nand U432 (N_432,In_120,N_309);
nor U433 (N_433,N_290,N_321);
nor U434 (N_434,N_350,N_87);
or U435 (N_435,N_360,In_497);
or U436 (N_436,N_256,N_173);
nor U437 (N_437,N_153,N_191);
or U438 (N_438,N_354,N_199);
nand U439 (N_439,N_340,N_240);
nor U440 (N_440,N_370,N_310);
nand U441 (N_441,N_356,N_290);
nor U442 (N_442,N_250,In_177);
nand U443 (N_443,N_339,N_361);
and U444 (N_444,N_198,In_229);
or U445 (N_445,N_327,N_322);
or U446 (N_446,In_497,N_351);
or U447 (N_447,In_324,N_220);
and U448 (N_448,N_321,In_324);
and U449 (N_449,N_312,N_303);
or U450 (N_450,N_407,N_393);
xor U451 (N_451,N_421,N_402);
and U452 (N_452,N_403,N_446);
nor U453 (N_453,N_422,N_417);
and U454 (N_454,N_433,N_382);
nand U455 (N_455,N_391,N_389);
nand U456 (N_456,N_376,N_384);
nor U457 (N_457,N_434,N_396);
or U458 (N_458,N_442,N_423);
nand U459 (N_459,N_430,N_381);
xor U460 (N_460,N_420,N_408);
xor U461 (N_461,N_414,N_444);
nor U462 (N_462,N_385,N_448);
nor U463 (N_463,N_390,N_418);
or U464 (N_464,N_375,N_410);
and U465 (N_465,N_445,N_427);
and U466 (N_466,N_419,N_412);
nor U467 (N_467,N_438,N_425);
or U468 (N_468,N_441,N_401);
nand U469 (N_469,N_426,N_424);
nand U470 (N_470,N_394,N_437);
xnor U471 (N_471,N_447,N_428);
nand U472 (N_472,N_377,N_432);
nand U473 (N_473,N_380,N_397);
xnor U474 (N_474,N_406,N_411);
or U475 (N_475,N_409,N_443);
xor U476 (N_476,N_398,N_439);
nand U477 (N_477,N_379,N_388);
nand U478 (N_478,N_449,N_431);
or U479 (N_479,N_404,N_413);
and U480 (N_480,N_405,N_386);
or U481 (N_481,N_395,N_435);
nand U482 (N_482,N_378,N_399);
or U483 (N_483,N_392,N_440);
or U484 (N_484,N_387,N_415);
nor U485 (N_485,N_429,N_416);
and U486 (N_486,N_436,N_383);
nand U487 (N_487,N_400,N_424);
or U488 (N_488,N_440,N_428);
nand U489 (N_489,N_397,N_394);
nor U490 (N_490,N_386,N_389);
or U491 (N_491,N_378,N_442);
nand U492 (N_492,N_440,N_414);
or U493 (N_493,N_425,N_449);
nor U494 (N_494,N_384,N_447);
nand U495 (N_495,N_449,N_432);
nor U496 (N_496,N_377,N_395);
and U497 (N_497,N_393,N_428);
or U498 (N_498,N_444,N_418);
or U499 (N_499,N_449,N_444);
nor U500 (N_500,N_390,N_439);
and U501 (N_501,N_435,N_394);
and U502 (N_502,N_387,N_375);
nand U503 (N_503,N_413,N_436);
nand U504 (N_504,N_399,N_386);
or U505 (N_505,N_380,N_423);
xnor U506 (N_506,N_404,N_411);
and U507 (N_507,N_431,N_377);
nand U508 (N_508,N_424,N_441);
or U509 (N_509,N_444,N_427);
nand U510 (N_510,N_380,N_401);
and U511 (N_511,N_431,N_376);
nand U512 (N_512,N_425,N_390);
or U513 (N_513,N_404,N_408);
or U514 (N_514,N_438,N_429);
and U515 (N_515,N_419,N_388);
and U516 (N_516,N_386,N_387);
and U517 (N_517,N_378,N_382);
and U518 (N_518,N_391,N_381);
nor U519 (N_519,N_389,N_396);
nand U520 (N_520,N_386,N_402);
xor U521 (N_521,N_441,N_386);
or U522 (N_522,N_440,N_379);
nor U523 (N_523,N_410,N_396);
or U524 (N_524,N_412,N_414);
xnor U525 (N_525,N_480,N_472);
nand U526 (N_526,N_515,N_514);
and U527 (N_527,N_490,N_484);
nor U528 (N_528,N_499,N_462);
nand U529 (N_529,N_498,N_475);
and U530 (N_530,N_477,N_493);
nor U531 (N_531,N_459,N_521);
or U532 (N_532,N_512,N_479);
nor U533 (N_533,N_518,N_452);
nor U534 (N_534,N_473,N_471);
and U535 (N_535,N_482,N_467);
nand U536 (N_536,N_497,N_502);
xor U537 (N_537,N_491,N_513);
and U538 (N_538,N_517,N_465);
nand U539 (N_539,N_500,N_509);
nor U540 (N_540,N_451,N_496);
or U541 (N_541,N_481,N_501);
and U542 (N_542,N_495,N_463);
or U543 (N_543,N_474,N_511);
nor U544 (N_544,N_487,N_516);
nor U545 (N_545,N_464,N_469);
nor U546 (N_546,N_503,N_508);
and U547 (N_547,N_505,N_456);
nor U548 (N_548,N_519,N_476);
nand U549 (N_549,N_455,N_520);
and U550 (N_550,N_453,N_523);
nor U551 (N_551,N_457,N_461);
nor U552 (N_552,N_489,N_486);
nand U553 (N_553,N_524,N_483);
xnor U554 (N_554,N_470,N_466);
xor U555 (N_555,N_450,N_522);
and U556 (N_556,N_478,N_458);
nand U557 (N_557,N_506,N_460);
or U558 (N_558,N_468,N_488);
or U559 (N_559,N_504,N_510);
or U560 (N_560,N_494,N_492);
and U561 (N_561,N_454,N_485);
or U562 (N_562,N_507,N_463);
nand U563 (N_563,N_502,N_493);
nand U564 (N_564,N_487,N_503);
and U565 (N_565,N_520,N_451);
and U566 (N_566,N_522,N_490);
nor U567 (N_567,N_490,N_488);
xor U568 (N_568,N_487,N_519);
nand U569 (N_569,N_457,N_496);
or U570 (N_570,N_453,N_500);
nand U571 (N_571,N_524,N_486);
xor U572 (N_572,N_469,N_457);
nor U573 (N_573,N_452,N_498);
nor U574 (N_574,N_459,N_468);
xnor U575 (N_575,N_469,N_461);
nor U576 (N_576,N_487,N_511);
nor U577 (N_577,N_455,N_504);
xor U578 (N_578,N_462,N_498);
or U579 (N_579,N_454,N_507);
nor U580 (N_580,N_471,N_456);
nand U581 (N_581,N_464,N_521);
xor U582 (N_582,N_520,N_474);
and U583 (N_583,N_484,N_461);
nand U584 (N_584,N_478,N_480);
nand U585 (N_585,N_507,N_498);
nand U586 (N_586,N_485,N_460);
nand U587 (N_587,N_506,N_483);
or U588 (N_588,N_464,N_513);
or U589 (N_589,N_487,N_510);
and U590 (N_590,N_510,N_454);
and U591 (N_591,N_451,N_467);
nor U592 (N_592,N_518,N_489);
nor U593 (N_593,N_494,N_493);
nand U594 (N_594,N_521,N_497);
nor U595 (N_595,N_484,N_460);
nor U596 (N_596,N_517,N_481);
and U597 (N_597,N_453,N_481);
xnor U598 (N_598,N_472,N_496);
and U599 (N_599,N_519,N_455);
nor U600 (N_600,N_534,N_554);
or U601 (N_601,N_568,N_549);
or U602 (N_602,N_565,N_563);
or U603 (N_603,N_572,N_584);
xnor U604 (N_604,N_560,N_547);
nor U605 (N_605,N_594,N_528);
or U606 (N_606,N_585,N_544);
xnor U607 (N_607,N_527,N_589);
xnor U608 (N_608,N_580,N_575);
and U609 (N_609,N_579,N_593);
or U610 (N_610,N_536,N_599);
xor U611 (N_611,N_587,N_535);
nand U612 (N_612,N_533,N_541);
nand U613 (N_613,N_542,N_596);
or U614 (N_614,N_537,N_551);
or U615 (N_615,N_558,N_550);
or U616 (N_616,N_543,N_586);
and U617 (N_617,N_555,N_574);
nand U618 (N_618,N_530,N_578);
nor U619 (N_619,N_557,N_525);
and U620 (N_620,N_564,N_529);
and U621 (N_621,N_598,N_539);
and U622 (N_622,N_570,N_567);
xor U623 (N_623,N_591,N_569);
nand U624 (N_624,N_540,N_571);
nand U625 (N_625,N_546,N_588);
nor U626 (N_626,N_582,N_595);
and U627 (N_627,N_590,N_581);
nor U628 (N_628,N_526,N_545);
xnor U629 (N_629,N_573,N_532);
and U630 (N_630,N_559,N_562);
nor U631 (N_631,N_597,N_577);
xnor U632 (N_632,N_556,N_531);
nor U633 (N_633,N_548,N_553);
nor U634 (N_634,N_576,N_552);
nand U635 (N_635,N_566,N_592);
and U636 (N_636,N_583,N_561);
nor U637 (N_637,N_538,N_564);
nor U638 (N_638,N_555,N_593);
and U639 (N_639,N_576,N_526);
nor U640 (N_640,N_591,N_576);
nand U641 (N_641,N_589,N_554);
or U642 (N_642,N_543,N_549);
or U643 (N_643,N_555,N_537);
nand U644 (N_644,N_532,N_565);
nand U645 (N_645,N_538,N_525);
xor U646 (N_646,N_547,N_581);
nand U647 (N_647,N_556,N_588);
or U648 (N_648,N_548,N_535);
nand U649 (N_649,N_571,N_567);
nand U650 (N_650,N_549,N_596);
nand U651 (N_651,N_537,N_539);
or U652 (N_652,N_557,N_573);
nor U653 (N_653,N_546,N_592);
nand U654 (N_654,N_590,N_536);
xor U655 (N_655,N_584,N_598);
nor U656 (N_656,N_587,N_536);
xnor U657 (N_657,N_543,N_554);
xnor U658 (N_658,N_558,N_540);
nand U659 (N_659,N_586,N_588);
and U660 (N_660,N_561,N_575);
nand U661 (N_661,N_572,N_555);
nor U662 (N_662,N_587,N_569);
or U663 (N_663,N_541,N_599);
and U664 (N_664,N_539,N_592);
and U665 (N_665,N_570,N_550);
and U666 (N_666,N_554,N_576);
nand U667 (N_667,N_594,N_591);
nand U668 (N_668,N_570,N_528);
or U669 (N_669,N_551,N_546);
xor U670 (N_670,N_589,N_588);
nand U671 (N_671,N_593,N_526);
nand U672 (N_672,N_588,N_555);
nor U673 (N_673,N_534,N_545);
nor U674 (N_674,N_525,N_573);
or U675 (N_675,N_641,N_661);
nand U676 (N_676,N_637,N_640);
xor U677 (N_677,N_643,N_652);
nor U678 (N_678,N_621,N_602);
nor U679 (N_679,N_633,N_611);
or U680 (N_680,N_658,N_667);
nand U681 (N_681,N_620,N_651);
and U682 (N_682,N_638,N_673);
or U683 (N_683,N_659,N_657);
or U684 (N_684,N_625,N_606);
nand U685 (N_685,N_655,N_648);
or U686 (N_686,N_624,N_668);
nand U687 (N_687,N_627,N_618);
xor U688 (N_688,N_636,N_662);
or U689 (N_689,N_600,N_647);
or U690 (N_690,N_665,N_629);
nor U691 (N_691,N_674,N_639);
and U692 (N_692,N_615,N_650);
nand U693 (N_693,N_634,N_604);
nor U694 (N_694,N_644,N_619);
or U695 (N_695,N_663,N_646);
xor U696 (N_696,N_608,N_626);
nor U697 (N_697,N_664,N_669);
xnor U698 (N_698,N_666,N_610);
xnor U699 (N_699,N_613,N_614);
xor U700 (N_700,N_660,N_656);
xor U701 (N_701,N_603,N_623);
nor U702 (N_702,N_654,N_645);
xor U703 (N_703,N_649,N_628);
nor U704 (N_704,N_605,N_672);
nor U705 (N_705,N_617,N_635);
nand U706 (N_706,N_630,N_642);
nor U707 (N_707,N_601,N_612);
and U708 (N_708,N_622,N_670);
and U709 (N_709,N_653,N_609);
or U710 (N_710,N_607,N_671);
nor U711 (N_711,N_631,N_616);
nor U712 (N_712,N_632,N_622);
nor U713 (N_713,N_664,N_612);
nand U714 (N_714,N_635,N_674);
and U715 (N_715,N_628,N_601);
and U716 (N_716,N_619,N_669);
and U717 (N_717,N_603,N_673);
or U718 (N_718,N_644,N_635);
xnor U719 (N_719,N_617,N_652);
nand U720 (N_720,N_617,N_615);
nor U721 (N_721,N_649,N_608);
xnor U722 (N_722,N_639,N_625);
and U723 (N_723,N_613,N_642);
and U724 (N_724,N_625,N_635);
or U725 (N_725,N_672,N_614);
xnor U726 (N_726,N_616,N_647);
or U727 (N_727,N_642,N_601);
nand U728 (N_728,N_671,N_618);
and U729 (N_729,N_626,N_617);
xnor U730 (N_730,N_619,N_674);
or U731 (N_731,N_603,N_633);
nand U732 (N_732,N_658,N_635);
nor U733 (N_733,N_608,N_643);
and U734 (N_734,N_637,N_670);
nor U735 (N_735,N_648,N_651);
nand U736 (N_736,N_610,N_608);
and U737 (N_737,N_666,N_642);
nor U738 (N_738,N_659,N_603);
nor U739 (N_739,N_654,N_630);
nor U740 (N_740,N_618,N_641);
or U741 (N_741,N_664,N_649);
or U742 (N_742,N_648,N_641);
or U743 (N_743,N_659,N_653);
nor U744 (N_744,N_628,N_632);
or U745 (N_745,N_620,N_618);
nor U746 (N_746,N_603,N_661);
nand U747 (N_747,N_618,N_660);
or U748 (N_748,N_603,N_650);
nand U749 (N_749,N_658,N_632);
and U750 (N_750,N_700,N_680);
nor U751 (N_751,N_742,N_709);
or U752 (N_752,N_744,N_676);
xnor U753 (N_753,N_719,N_717);
xor U754 (N_754,N_683,N_696);
and U755 (N_755,N_732,N_746);
nor U756 (N_756,N_737,N_692);
nor U757 (N_757,N_728,N_722);
and U758 (N_758,N_749,N_684);
nand U759 (N_759,N_715,N_724);
or U760 (N_760,N_706,N_699);
nand U761 (N_761,N_714,N_747);
nor U762 (N_762,N_723,N_731);
nor U763 (N_763,N_698,N_687);
and U764 (N_764,N_741,N_738);
or U765 (N_765,N_739,N_718);
nor U766 (N_766,N_678,N_734);
nand U767 (N_767,N_691,N_694);
or U768 (N_768,N_711,N_729);
nor U769 (N_769,N_688,N_695);
or U770 (N_770,N_710,N_685);
nand U771 (N_771,N_701,N_682);
and U772 (N_772,N_708,N_735);
nand U773 (N_773,N_677,N_725);
nand U774 (N_774,N_727,N_740);
or U775 (N_775,N_736,N_726);
xor U776 (N_776,N_681,N_748);
nor U777 (N_777,N_743,N_689);
or U778 (N_778,N_730,N_675);
and U779 (N_779,N_703,N_704);
and U780 (N_780,N_712,N_720);
and U781 (N_781,N_686,N_733);
nor U782 (N_782,N_679,N_697);
or U783 (N_783,N_716,N_713);
xnor U784 (N_784,N_690,N_693);
and U785 (N_785,N_705,N_721);
or U786 (N_786,N_745,N_707);
nor U787 (N_787,N_702,N_745);
or U788 (N_788,N_718,N_712);
and U789 (N_789,N_686,N_701);
and U790 (N_790,N_680,N_736);
nand U791 (N_791,N_724,N_710);
nor U792 (N_792,N_726,N_732);
nand U793 (N_793,N_698,N_709);
nand U794 (N_794,N_716,N_690);
nor U795 (N_795,N_749,N_718);
xnor U796 (N_796,N_699,N_726);
nor U797 (N_797,N_679,N_726);
or U798 (N_798,N_698,N_737);
and U799 (N_799,N_731,N_716);
or U800 (N_800,N_700,N_677);
nor U801 (N_801,N_737,N_741);
nor U802 (N_802,N_701,N_734);
xor U803 (N_803,N_695,N_722);
nor U804 (N_804,N_715,N_728);
or U805 (N_805,N_709,N_728);
and U806 (N_806,N_732,N_744);
and U807 (N_807,N_709,N_688);
nand U808 (N_808,N_729,N_697);
or U809 (N_809,N_749,N_681);
nor U810 (N_810,N_716,N_681);
xnor U811 (N_811,N_702,N_710);
and U812 (N_812,N_687,N_728);
xor U813 (N_813,N_685,N_741);
nand U814 (N_814,N_745,N_714);
and U815 (N_815,N_691,N_714);
nor U816 (N_816,N_728,N_723);
xor U817 (N_817,N_736,N_679);
nand U818 (N_818,N_728,N_736);
or U819 (N_819,N_739,N_735);
nor U820 (N_820,N_714,N_730);
or U821 (N_821,N_699,N_698);
nand U822 (N_822,N_736,N_676);
xnor U823 (N_823,N_680,N_743);
and U824 (N_824,N_702,N_747);
or U825 (N_825,N_820,N_819);
or U826 (N_826,N_774,N_782);
nor U827 (N_827,N_802,N_810);
and U828 (N_828,N_800,N_784);
nor U829 (N_829,N_812,N_777);
nand U830 (N_830,N_788,N_765);
nor U831 (N_831,N_821,N_773);
xor U832 (N_832,N_796,N_778);
nand U833 (N_833,N_791,N_756);
and U834 (N_834,N_775,N_760);
nand U835 (N_835,N_792,N_768);
nand U836 (N_836,N_799,N_793);
and U837 (N_837,N_813,N_779);
nand U838 (N_838,N_798,N_789);
and U839 (N_839,N_761,N_815);
nor U840 (N_840,N_824,N_783);
nand U841 (N_841,N_759,N_794);
nand U842 (N_842,N_772,N_797);
nor U843 (N_843,N_807,N_767);
and U844 (N_844,N_771,N_806);
xor U845 (N_845,N_795,N_804);
or U846 (N_846,N_751,N_808);
nor U847 (N_847,N_818,N_776);
nor U848 (N_848,N_757,N_780);
nand U849 (N_849,N_803,N_823);
or U850 (N_850,N_801,N_814);
or U851 (N_851,N_805,N_769);
or U852 (N_852,N_822,N_781);
xor U853 (N_853,N_763,N_764);
nand U854 (N_854,N_785,N_811);
nand U855 (N_855,N_809,N_766);
and U856 (N_856,N_790,N_753);
or U857 (N_857,N_755,N_787);
nand U858 (N_858,N_754,N_758);
nand U859 (N_859,N_762,N_817);
and U860 (N_860,N_786,N_752);
nor U861 (N_861,N_770,N_816);
and U862 (N_862,N_750,N_798);
nand U863 (N_863,N_803,N_756);
nor U864 (N_864,N_824,N_796);
and U865 (N_865,N_754,N_796);
or U866 (N_866,N_777,N_774);
or U867 (N_867,N_812,N_820);
nand U868 (N_868,N_789,N_810);
and U869 (N_869,N_811,N_821);
nand U870 (N_870,N_799,N_822);
or U871 (N_871,N_787,N_754);
or U872 (N_872,N_765,N_777);
nor U873 (N_873,N_809,N_759);
or U874 (N_874,N_810,N_824);
xor U875 (N_875,N_805,N_793);
nand U876 (N_876,N_819,N_823);
nor U877 (N_877,N_806,N_773);
or U878 (N_878,N_813,N_757);
or U879 (N_879,N_750,N_764);
nor U880 (N_880,N_767,N_815);
or U881 (N_881,N_804,N_811);
or U882 (N_882,N_816,N_765);
nand U883 (N_883,N_814,N_784);
and U884 (N_884,N_773,N_812);
nand U885 (N_885,N_756,N_802);
and U886 (N_886,N_769,N_817);
nor U887 (N_887,N_816,N_811);
nor U888 (N_888,N_785,N_809);
nor U889 (N_889,N_762,N_798);
nor U890 (N_890,N_800,N_768);
nor U891 (N_891,N_752,N_764);
nand U892 (N_892,N_817,N_824);
or U893 (N_893,N_755,N_784);
or U894 (N_894,N_775,N_784);
or U895 (N_895,N_787,N_758);
nand U896 (N_896,N_752,N_765);
nor U897 (N_897,N_763,N_802);
and U898 (N_898,N_816,N_787);
or U899 (N_899,N_755,N_763);
nand U900 (N_900,N_874,N_834);
or U901 (N_901,N_835,N_887);
nand U902 (N_902,N_852,N_876);
nand U903 (N_903,N_895,N_869);
nand U904 (N_904,N_898,N_896);
and U905 (N_905,N_826,N_854);
nand U906 (N_906,N_846,N_866);
or U907 (N_907,N_883,N_880);
or U908 (N_908,N_829,N_899);
nor U909 (N_909,N_837,N_891);
nand U910 (N_910,N_838,N_879);
nand U911 (N_911,N_830,N_884);
or U912 (N_912,N_890,N_831);
and U913 (N_913,N_888,N_855);
and U914 (N_914,N_863,N_882);
or U915 (N_915,N_847,N_870);
or U916 (N_916,N_864,N_881);
and U917 (N_917,N_860,N_853);
nor U918 (N_918,N_839,N_825);
nand U919 (N_919,N_845,N_892);
nand U920 (N_920,N_844,N_842);
or U921 (N_921,N_872,N_877);
and U922 (N_922,N_867,N_865);
nor U923 (N_923,N_862,N_828);
xor U924 (N_924,N_836,N_861);
nand U925 (N_925,N_851,N_868);
nor U926 (N_926,N_849,N_841);
and U927 (N_927,N_833,N_885);
or U928 (N_928,N_878,N_875);
nand U929 (N_929,N_889,N_873);
nor U930 (N_930,N_886,N_897);
and U931 (N_931,N_832,N_843);
or U932 (N_932,N_858,N_827);
and U933 (N_933,N_840,N_859);
nor U934 (N_934,N_848,N_856);
nor U935 (N_935,N_894,N_871);
and U936 (N_936,N_857,N_850);
nand U937 (N_937,N_893,N_843);
or U938 (N_938,N_886,N_869);
or U939 (N_939,N_851,N_883);
and U940 (N_940,N_897,N_865);
nand U941 (N_941,N_839,N_857);
nor U942 (N_942,N_837,N_873);
nand U943 (N_943,N_861,N_859);
nor U944 (N_944,N_826,N_896);
or U945 (N_945,N_866,N_894);
nor U946 (N_946,N_834,N_848);
xor U947 (N_947,N_825,N_860);
and U948 (N_948,N_837,N_888);
or U949 (N_949,N_874,N_844);
xnor U950 (N_950,N_870,N_887);
nand U951 (N_951,N_826,N_843);
and U952 (N_952,N_836,N_825);
xnor U953 (N_953,N_899,N_890);
or U954 (N_954,N_871,N_895);
and U955 (N_955,N_874,N_848);
or U956 (N_956,N_827,N_834);
or U957 (N_957,N_882,N_853);
nand U958 (N_958,N_852,N_892);
and U959 (N_959,N_853,N_896);
and U960 (N_960,N_869,N_836);
nand U961 (N_961,N_881,N_885);
nor U962 (N_962,N_835,N_850);
or U963 (N_963,N_865,N_838);
and U964 (N_964,N_831,N_893);
nor U965 (N_965,N_874,N_898);
or U966 (N_966,N_867,N_886);
and U967 (N_967,N_885,N_870);
nand U968 (N_968,N_896,N_847);
or U969 (N_969,N_836,N_841);
nand U970 (N_970,N_846,N_849);
nand U971 (N_971,N_843,N_866);
or U972 (N_972,N_846,N_877);
or U973 (N_973,N_831,N_871);
and U974 (N_974,N_832,N_853);
nand U975 (N_975,N_919,N_953);
and U976 (N_976,N_965,N_974);
nor U977 (N_977,N_942,N_923);
nor U978 (N_978,N_971,N_944);
or U979 (N_979,N_949,N_914);
nor U980 (N_980,N_972,N_932);
nor U981 (N_981,N_909,N_920);
nor U982 (N_982,N_943,N_946);
nand U983 (N_983,N_903,N_931);
nand U984 (N_984,N_966,N_901);
or U985 (N_985,N_957,N_964);
nor U986 (N_986,N_959,N_963);
and U987 (N_987,N_910,N_973);
or U988 (N_988,N_938,N_945);
nand U989 (N_989,N_956,N_913);
and U990 (N_990,N_940,N_904);
nor U991 (N_991,N_900,N_926);
and U992 (N_992,N_939,N_907);
and U993 (N_993,N_924,N_934);
or U994 (N_994,N_935,N_960);
and U995 (N_995,N_951,N_918);
or U996 (N_996,N_958,N_941);
xor U997 (N_997,N_962,N_917);
or U998 (N_998,N_908,N_955);
or U999 (N_999,N_961,N_922);
and U1000 (N_1000,N_916,N_948);
nor U1001 (N_1001,N_911,N_928);
nand U1002 (N_1002,N_947,N_929);
or U1003 (N_1003,N_902,N_930);
or U1004 (N_1004,N_954,N_970);
or U1005 (N_1005,N_925,N_969);
xor U1006 (N_1006,N_906,N_967);
or U1007 (N_1007,N_927,N_936);
nand U1008 (N_1008,N_905,N_912);
nand U1009 (N_1009,N_921,N_952);
nand U1010 (N_1010,N_968,N_915);
or U1011 (N_1011,N_937,N_950);
nor U1012 (N_1012,N_933,N_904);
nor U1013 (N_1013,N_937,N_955);
or U1014 (N_1014,N_912,N_965);
or U1015 (N_1015,N_968,N_906);
or U1016 (N_1016,N_958,N_942);
and U1017 (N_1017,N_943,N_972);
xnor U1018 (N_1018,N_934,N_967);
or U1019 (N_1019,N_935,N_973);
nor U1020 (N_1020,N_972,N_957);
xnor U1021 (N_1021,N_959,N_902);
nor U1022 (N_1022,N_971,N_948);
nor U1023 (N_1023,N_919,N_918);
nor U1024 (N_1024,N_961,N_970);
nand U1025 (N_1025,N_952,N_938);
nor U1026 (N_1026,N_919,N_924);
or U1027 (N_1027,N_903,N_900);
and U1028 (N_1028,N_972,N_911);
xor U1029 (N_1029,N_911,N_938);
nand U1030 (N_1030,N_947,N_941);
or U1031 (N_1031,N_959,N_973);
nor U1032 (N_1032,N_922,N_932);
nor U1033 (N_1033,N_916,N_957);
xor U1034 (N_1034,N_952,N_948);
and U1035 (N_1035,N_920,N_923);
and U1036 (N_1036,N_967,N_951);
or U1037 (N_1037,N_928,N_967);
xnor U1038 (N_1038,N_902,N_925);
or U1039 (N_1039,N_934,N_942);
xnor U1040 (N_1040,N_946,N_904);
nor U1041 (N_1041,N_965,N_901);
nor U1042 (N_1042,N_972,N_903);
nand U1043 (N_1043,N_939,N_938);
and U1044 (N_1044,N_945,N_937);
nor U1045 (N_1045,N_910,N_918);
nand U1046 (N_1046,N_955,N_960);
and U1047 (N_1047,N_937,N_939);
nor U1048 (N_1048,N_933,N_972);
or U1049 (N_1049,N_933,N_950);
nor U1050 (N_1050,N_1033,N_1035);
or U1051 (N_1051,N_1040,N_1010);
nand U1052 (N_1052,N_979,N_1008);
nand U1053 (N_1053,N_1031,N_1018);
nand U1054 (N_1054,N_985,N_1039);
or U1055 (N_1055,N_999,N_1002);
nand U1056 (N_1056,N_1014,N_1025);
or U1057 (N_1057,N_1034,N_1003);
nand U1058 (N_1058,N_997,N_1045);
nor U1059 (N_1059,N_1021,N_1001);
and U1060 (N_1060,N_994,N_1043);
xor U1061 (N_1061,N_1048,N_1046);
or U1062 (N_1062,N_987,N_983);
and U1063 (N_1063,N_992,N_988);
nor U1064 (N_1064,N_1022,N_996);
nand U1065 (N_1065,N_1020,N_976);
nand U1066 (N_1066,N_1036,N_995);
xnor U1067 (N_1067,N_1012,N_1042);
nand U1068 (N_1068,N_1044,N_1024);
or U1069 (N_1069,N_1049,N_980);
nand U1070 (N_1070,N_1047,N_1017);
nand U1071 (N_1071,N_998,N_981);
nor U1072 (N_1072,N_977,N_1037);
nand U1073 (N_1073,N_1038,N_1030);
and U1074 (N_1074,N_1019,N_1005);
nand U1075 (N_1075,N_1011,N_1004);
xnor U1076 (N_1076,N_991,N_984);
nand U1077 (N_1077,N_989,N_1013);
nand U1078 (N_1078,N_982,N_1016);
or U1079 (N_1079,N_1028,N_986);
nor U1080 (N_1080,N_993,N_1029);
nand U1081 (N_1081,N_990,N_1007);
and U1082 (N_1082,N_1000,N_1041);
nor U1083 (N_1083,N_1023,N_978);
nor U1084 (N_1084,N_975,N_1026);
and U1085 (N_1085,N_1015,N_1032);
or U1086 (N_1086,N_1027,N_1006);
xor U1087 (N_1087,N_1009,N_1020);
and U1088 (N_1088,N_1004,N_981);
nor U1089 (N_1089,N_1003,N_1000);
or U1090 (N_1090,N_986,N_1034);
xnor U1091 (N_1091,N_985,N_999);
nor U1092 (N_1092,N_982,N_979);
nor U1093 (N_1093,N_1015,N_995);
nand U1094 (N_1094,N_1030,N_998);
or U1095 (N_1095,N_995,N_988);
xnor U1096 (N_1096,N_1018,N_1043);
or U1097 (N_1097,N_985,N_1004);
nor U1098 (N_1098,N_1021,N_1047);
and U1099 (N_1099,N_1049,N_977);
nand U1100 (N_1100,N_1039,N_994);
and U1101 (N_1101,N_1025,N_1042);
nor U1102 (N_1102,N_979,N_1011);
or U1103 (N_1103,N_1019,N_1041);
nand U1104 (N_1104,N_996,N_1000);
nand U1105 (N_1105,N_1028,N_983);
and U1106 (N_1106,N_1031,N_1048);
nor U1107 (N_1107,N_993,N_1025);
nand U1108 (N_1108,N_990,N_1021);
or U1109 (N_1109,N_997,N_979);
nand U1110 (N_1110,N_982,N_998);
and U1111 (N_1111,N_1039,N_979);
and U1112 (N_1112,N_1039,N_1030);
nor U1113 (N_1113,N_990,N_994);
and U1114 (N_1114,N_1010,N_980);
and U1115 (N_1115,N_1033,N_1006);
nand U1116 (N_1116,N_992,N_1046);
and U1117 (N_1117,N_1010,N_1026);
xor U1118 (N_1118,N_1016,N_981);
and U1119 (N_1119,N_1028,N_1027);
xnor U1120 (N_1120,N_994,N_980);
nand U1121 (N_1121,N_989,N_1028);
nand U1122 (N_1122,N_1033,N_1034);
nand U1123 (N_1123,N_1035,N_1030);
nand U1124 (N_1124,N_1011,N_984);
and U1125 (N_1125,N_1083,N_1124);
and U1126 (N_1126,N_1096,N_1122);
nor U1127 (N_1127,N_1088,N_1075);
and U1128 (N_1128,N_1095,N_1058);
or U1129 (N_1129,N_1100,N_1114);
nor U1130 (N_1130,N_1107,N_1067);
nand U1131 (N_1131,N_1089,N_1117);
or U1132 (N_1132,N_1066,N_1105);
and U1133 (N_1133,N_1052,N_1073);
and U1134 (N_1134,N_1104,N_1102);
or U1135 (N_1135,N_1090,N_1069);
nor U1136 (N_1136,N_1119,N_1099);
or U1137 (N_1137,N_1079,N_1068);
or U1138 (N_1138,N_1118,N_1123);
and U1139 (N_1139,N_1059,N_1086);
xor U1140 (N_1140,N_1094,N_1054);
nor U1141 (N_1141,N_1057,N_1093);
xor U1142 (N_1142,N_1098,N_1106);
nor U1143 (N_1143,N_1082,N_1078);
xor U1144 (N_1144,N_1056,N_1063);
nand U1145 (N_1145,N_1112,N_1081);
or U1146 (N_1146,N_1103,N_1108);
and U1147 (N_1147,N_1092,N_1055);
xnor U1148 (N_1148,N_1084,N_1072);
or U1149 (N_1149,N_1053,N_1065);
nor U1150 (N_1150,N_1087,N_1091);
nor U1151 (N_1151,N_1080,N_1074);
nor U1152 (N_1152,N_1116,N_1061);
or U1153 (N_1153,N_1121,N_1050);
and U1154 (N_1154,N_1051,N_1113);
and U1155 (N_1155,N_1070,N_1110);
and U1156 (N_1156,N_1077,N_1101);
nand U1157 (N_1157,N_1076,N_1115);
nor U1158 (N_1158,N_1062,N_1064);
and U1159 (N_1159,N_1060,N_1097);
or U1160 (N_1160,N_1085,N_1071);
or U1161 (N_1161,N_1111,N_1120);
xor U1162 (N_1162,N_1109,N_1107);
nor U1163 (N_1163,N_1062,N_1069);
nor U1164 (N_1164,N_1090,N_1105);
nand U1165 (N_1165,N_1071,N_1083);
and U1166 (N_1166,N_1080,N_1066);
and U1167 (N_1167,N_1079,N_1056);
nor U1168 (N_1168,N_1112,N_1098);
nor U1169 (N_1169,N_1096,N_1056);
nor U1170 (N_1170,N_1120,N_1112);
xnor U1171 (N_1171,N_1091,N_1118);
nand U1172 (N_1172,N_1053,N_1094);
or U1173 (N_1173,N_1050,N_1084);
nor U1174 (N_1174,N_1082,N_1052);
or U1175 (N_1175,N_1103,N_1079);
nor U1176 (N_1176,N_1053,N_1123);
or U1177 (N_1177,N_1093,N_1087);
and U1178 (N_1178,N_1088,N_1052);
nand U1179 (N_1179,N_1090,N_1100);
or U1180 (N_1180,N_1115,N_1123);
nand U1181 (N_1181,N_1103,N_1085);
nor U1182 (N_1182,N_1063,N_1095);
nand U1183 (N_1183,N_1116,N_1084);
xnor U1184 (N_1184,N_1099,N_1096);
and U1185 (N_1185,N_1097,N_1116);
and U1186 (N_1186,N_1119,N_1071);
nand U1187 (N_1187,N_1070,N_1067);
and U1188 (N_1188,N_1061,N_1068);
nor U1189 (N_1189,N_1085,N_1069);
or U1190 (N_1190,N_1108,N_1107);
xor U1191 (N_1191,N_1117,N_1083);
nand U1192 (N_1192,N_1106,N_1066);
and U1193 (N_1193,N_1054,N_1091);
nand U1194 (N_1194,N_1061,N_1102);
and U1195 (N_1195,N_1090,N_1061);
and U1196 (N_1196,N_1106,N_1112);
nand U1197 (N_1197,N_1055,N_1088);
nand U1198 (N_1198,N_1057,N_1110);
and U1199 (N_1199,N_1116,N_1086);
or U1200 (N_1200,N_1135,N_1153);
and U1201 (N_1201,N_1166,N_1129);
and U1202 (N_1202,N_1160,N_1150);
nand U1203 (N_1203,N_1183,N_1187);
xnor U1204 (N_1204,N_1145,N_1170);
nand U1205 (N_1205,N_1140,N_1161);
and U1206 (N_1206,N_1192,N_1142);
nand U1207 (N_1207,N_1156,N_1174);
or U1208 (N_1208,N_1185,N_1189);
and U1209 (N_1209,N_1163,N_1152);
or U1210 (N_1210,N_1193,N_1151);
or U1211 (N_1211,N_1154,N_1136);
or U1212 (N_1212,N_1191,N_1190);
or U1213 (N_1213,N_1172,N_1167);
or U1214 (N_1214,N_1141,N_1128);
or U1215 (N_1215,N_1175,N_1178);
or U1216 (N_1216,N_1147,N_1158);
nor U1217 (N_1217,N_1176,N_1188);
nor U1218 (N_1218,N_1162,N_1126);
and U1219 (N_1219,N_1139,N_1195);
xor U1220 (N_1220,N_1125,N_1157);
nor U1221 (N_1221,N_1127,N_1155);
and U1222 (N_1222,N_1194,N_1143);
nor U1223 (N_1223,N_1196,N_1134);
nor U1224 (N_1224,N_1197,N_1137);
xnor U1225 (N_1225,N_1130,N_1164);
or U1226 (N_1226,N_1177,N_1149);
xnor U1227 (N_1227,N_1186,N_1168);
or U1228 (N_1228,N_1169,N_1179);
and U1229 (N_1229,N_1138,N_1198);
or U1230 (N_1230,N_1165,N_1199);
and U1231 (N_1231,N_1133,N_1184);
or U1232 (N_1232,N_1181,N_1148);
nor U1233 (N_1233,N_1182,N_1180);
nor U1234 (N_1234,N_1132,N_1173);
nand U1235 (N_1235,N_1159,N_1144);
nand U1236 (N_1236,N_1171,N_1131);
nor U1237 (N_1237,N_1146,N_1194);
xnor U1238 (N_1238,N_1177,N_1129);
and U1239 (N_1239,N_1173,N_1163);
nand U1240 (N_1240,N_1138,N_1141);
or U1241 (N_1241,N_1128,N_1195);
or U1242 (N_1242,N_1195,N_1150);
nand U1243 (N_1243,N_1136,N_1184);
and U1244 (N_1244,N_1148,N_1136);
and U1245 (N_1245,N_1143,N_1135);
and U1246 (N_1246,N_1141,N_1142);
nor U1247 (N_1247,N_1157,N_1138);
and U1248 (N_1248,N_1143,N_1171);
and U1249 (N_1249,N_1128,N_1135);
or U1250 (N_1250,N_1160,N_1126);
and U1251 (N_1251,N_1163,N_1136);
and U1252 (N_1252,N_1139,N_1129);
nand U1253 (N_1253,N_1160,N_1147);
or U1254 (N_1254,N_1195,N_1161);
xnor U1255 (N_1255,N_1125,N_1178);
and U1256 (N_1256,N_1174,N_1197);
and U1257 (N_1257,N_1158,N_1148);
or U1258 (N_1258,N_1186,N_1187);
and U1259 (N_1259,N_1165,N_1171);
xor U1260 (N_1260,N_1155,N_1181);
nand U1261 (N_1261,N_1194,N_1195);
xor U1262 (N_1262,N_1145,N_1199);
nand U1263 (N_1263,N_1191,N_1176);
or U1264 (N_1264,N_1160,N_1144);
xor U1265 (N_1265,N_1193,N_1129);
nand U1266 (N_1266,N_1178,N_1153);
nand U1267 (N_1267,N_1143,N_1129);
or U1268 (N_1268,N_1190,N_1198);
or U1269 (N_1269,N_1130,N_1158);
xor U1270 (N_1270,N_1138,N_1176);
and U1271 (N_1271,N_1166,N_1195);
or U1272 (N_1272,N_1143,N_1142);
xnor U1273 (N_1273,N_1171,N_1156);
or U1274 (N_1274,N_1186,N_1151);
and U1275 (N_1275,N_1207,N_1233);
nor U1276 (N_1276,N_1228,N_1263);
xor U1277 (N_1277,N_1223,N_1244);
nor U1278 (N_1278,N_1246,N_1220);
or U1279 (N_1279,N_1250,N_1236);
or U1280 (N_1280,N_1201,N_1259);
or U1281 (N_1281,N_1221,N_1219);
xor U1282 (N_1282,N_1272,N_1249);
or U1283 (N_1283,N_1203,N_1206);
nor U1284 (N_1284,N_1208,N_1231);
and U1285 (N_1285,N_1204,N_1270);
and U1286 (N_1286,N_1258,N_1260);
nor U1287 (N_1287,N_1253,N_1248);
or U1288 (N_1288,N_1224,N_1229);
nor U1289 (N_1289,N_1209,N_1247);
and U1290 (N_1290,N_1211,N_1266);
xor U1291 (N_1291,N_1235,N_1227);
nor U1292 (N_1292,N_1226,N_1218);
nand U1293 (N_1293,N_1257,N_1267);
or U1294 (N_1294,N_1269,N_1252);
and U1295 (N_1295,N_1212,N_1241);
or U1296 (N_1296,N_1232,N_1243);
or U1297 (N_1297,N_1245,N_1202);
nand U1298 (N_1298,N_1238,N_1254);
nor U1299 (N_1299,N_1251,N_1214);
or U1300 (N_1300,N_1200,N_1234);
nand U1301 (N_1301,N_1256,N_1255);
and U1302 (N_1302,N_1261,N_1274);
and U1303 (N_1303,N_1237,N_1271);
nand U1304 (N_1304,N_1217,N_1273);
nor U1305 (N_1305,N_1210,N_1264);
nor U1306 (N_1306,N_1240,N_1215);
or U1307 (N_1307,N_1222,N_1230);
or U1308 (N_1308,N_1268,N_1213);
xnor U1309 (N_1309,N_1225,N_1262);
or U1310 (N_1310,N_1242,N_1239);
or U1311 (N_1311,N_1216,N_1265);
nand U1312 (N_1312,N_1205,N_1211);
nand U1313 (N_1313,N_1231,N_1229);
nor U1314 (N_1314,N_1243,N_1238);
xnor U1315 (N_1315,N_1245,N_1214);
and U1316 (N_1316,N_1269,N_1259);
or U1317 (N_1317,N_1227,N_1204);
nor U1318 (N_1318,N_1205,N_1200);
nor U1319 (N_1319,N_1274,N_1221);
nor U1320 (N_1320,N_1234,N_1247);
nand U1321 (N_1321,N_1207,N_1223);
nor U1322 (N_1322,N_1215,N_1202);
and U1323 (N_1323,N_1254,N_1252);
nand U1324 (N_1324,N_1233,N_1223);
nand U1325 (N_1325,N_1213,N_1220);
and U1326 (N_1326,N_1236,N_1251);
xor U1327 (N_1327,N_1210,N_1247);
nor U1328 (N_1328,N_1212,N_1219);
and U1329 (N_1329,N_1202,N_1248);
nor U1330 (N_1330,N_1255,N_1239);
and U1331 (N_1331,N_1259,N_1236);
and U1332 (N_1332,N_1249,N_1215);
and U1333 (N_1333,N_1225,N_1272);
or U1334 (N_1334,N_1267,N_1233);
and U1335 (N_1335,N_1263,N_1229);
nand U1336 (N_1336,N_1245,N_1268);
or U1337 (N_1337,N_1237,N_1243);
and U1338 (N_1338,N_1251,N_1221);
or U1339 (N_1339,N_1246,N_1206);
nor U1340 (N_1340,N_1244,N_1222);
and U1341 (N_1341,N_1223,N_1200);
nand U1342 (N_1342,N_1231,N_1244);
nor U1343 (N_1343,N_1237,N_1252);
nand U1344 (N_1344,N_1242,N_1200);
or U1345 (N_1345,N_1230,N_1251);
xor U1346 (N_1346,N_1266,N_1208);
nor U1347 (N_1347,N_1208,N_1200);
or U1348 (N_1348,N_1227,N_1224);
and U1349 (N_1349,N_1214,N_1234);
or U1350 (N_1350,N_1338,N_1275);
nand U1351 (N_1351,N_1316,N_1319);
nand U1352 (N_1352,N_1333,N_1304);
nor U1353 (N_1353,N_1280,N_1299);
nand U1354 (N_1354,N_1308,N_1335);
and U1355 (N_1355,N_1285,N_1324);
and U1356 (N_1356,N_1348,N_1289);
xnor U1357 (N_1357,N_1347,N_1276);
nor U1358 (N_1358,N_1314,N_1321);
xnor U1359 (N_1359,N_1296,N_1309);
or U1360 (N_1360,N_1290,N_1291);
and U1361 (N_1361,N_1323,N_1294);
or U1362 (N_1362,N_1320,N_1302);
or U1363 (N_1363,N_1337,N_1334);
or U1364 (N_1364,N_1342,N_1293);
and U1365 (N_1365,N_1318,N_1330);
and U1366 (N_1366,N_1349,N_1288);
xnor U1367 (N_1367,N_1339,N_1282);
or U1368 (N_1368,N_1328,N_1277);
nor U1369 (N_1369,N_1327,N_1305);
nor U1370 (N_1370,N_1341,N_1315);
xnor U1371 (N_1371,N_1332,N_1346);
nor U1372 (N_1372,N_1307,N_1298);
nor U1373 (N_1373,N_1278,N_1343);
and U1374 (N_1374,N_1281,N_1340);
nand U1375 (N_1375,N_1303,N_1331);
nand U1376 (N_1376,N_1317,N_1279);
nor U1377 (N_1377,N_1325,N_1322);
nand U1378 (N_1378,N_1311,N_1286);
nor U1379 (N_1379,N_1329,N_1295);
and U1380 (N_1380,N_1312,N_1344);
and U1381 (N_1381,N_1292,N_1306);
xnor U1382 (N_1382,N_1310,N_1297);
or U1383 (N_1383,N_1287,N_1300);
and U1384 (N_1384,N_1345,N_1313);
and U1385 (N_1385,N_1326,N_1283);
nand U1386 (N_1386,N_1284,N_1336);
xnor U1387 (N_1387,N_1301,N_1284);
nor U1388 (N_1388,N_1347,N_1315);
nor U1389 (N_1389,N_1338,N_1310);
and U1390 (N_1390,N_1337,N_1308);
or U1391 (N_1391,N_1344,N_1299);
or U1392 (N_1392,N_1289,N_1323);
and U1393 (N_1393,N_1349,N_1335);
nor U1394 (N_1394,N_1336,N_1334);
nand U1395 (N_1395,N_1282,N_1330);
nand U1396 (N_1396,N_1332,N_1314);
nor U1397 (N_1397,N_1319,N_1312);
nand U1398 (N_1398,N_1340,N_1345);
or U1399 (N_1399,N_1292,N_1287);
xnor U1400 (N_1400,N_1304,N_1283);
xnor U1401 (N_1401,N_1283,N_1307);
or U1402 (N_1402,N_1281,N_1314);
nand U1403 (N_1403,N_1283,N_1329);
nand U1404 (N_1404,N_1306,N_1325);
nand U1405 (N_1405,N_1313,N_1309);
and U1406 (N_1406,N_1343,N_1314);
nand U1407 (N_1407,N_1308,N_1288);
nand U1408 (N_1408,N_1289,N_1282);
nor U1409 (N_1409,N_1316,N_1322);
nand U1410 (N_1410,N_1339,N_1327);
nor U1411 (N_1411,N_1280,N_1276);
xnor U1412 (N_1412,N_1297,N_1335);
or U1413 (N_1413,N_1327,N_1349);
and U1414 (N_1414,N_1347,N_1321);
and U1415 (N_1415,N_1292,N_1290);
nor U1416 (N_1416,N_1326,N_1323);
and U1417 (N_1417,N_1333,N_1284);
and U1418 (N_1418,N_1326,N_1291);
and U1419 (N_1419,N_1276,N_1284);
xnor U1420 (N_1420,N_1277,N_1299);
and U1421 (N_1421,N_1301,N_1327);
or U1422 (N_1422,N_1337,N_1300);
nand U1423 (N_1423,N_1347,N_1340);
nand U1424 (N_1424,N_1290,N_1330);
and U1425 (N_1425,N_1360,N_1354);
nor U1426 (N_1426,N_1420,N_1375);
or U1427 (N_1427,N_1410,N_1388);
and U1428 (N_1428,N_1412,N_1407);
or U1429 (N_1429,N_1364,N_1422);
nor U1430 (N_1430,N_1421,N_1395);
nor U1431 (N_1431,N_1369,N_1386);
or U1432 (N_1432,N_1351,N_1361);
nand U1433 (N_1433,N_1376,N_1384);
xnor U1434 (N_1434,N_1385,N_1409);
nand U1435 (N_1435,N_1366,N_1380);
nand U1436 (N_1436,N_1411,N_1401);
and U1437 (N_1437,N_1374,N_1416);
nand U1438 (N_1438,N_1350,N_1377);
nand U1439 (N_1439,N_1415,N_1413);
and U1440 (N_1440,N_1391,N_1408);
xor U1441 (N_1441,N_1363,N_1397);
or U1442 (N_1442,N_1399,N_1414);
or U1443 (N_1443,N_1359,N_1362);
nor U1444 (N_1444,N_1358,N_1368);
and U1445 (N_1445,N_1370,N_1423);
nand U1446 (N_1446,N_1352,N_1405);
or U1447 (N_1447,N_1383,N_1382);
xor U1448 (N_1448,N_1404,N_1365);
or U1449 (N_1449,N_1417,N_1356);
nand U1450 (N_1450,N_1378,N_1419);
and U1451 (N_1451,N_1357,N_1424);
nor U1452 (N_1452,N_1371,N_1394);
nor U1453 (N_1453,N_1355,N_1389);
nor U1454 (N_1454,N_1381,N_1373);
or U1455 (N_1455,N_1403,N_1396);
nor U1456 (N_1456,N_1418,N_1400);
nor U1457 (N_1457,N_1402,N_1367);
nor U1458 (N_1458,N_1372,N_1393);
or U1459 (N_1459,N_1390,N_1398);
and U1460 (N_1460,N_1379,N_1387);
nand U1461 (N_1461,N_1392,N_1353);
nor U1462 (N_1462,N_1406,N_1398);
or U1463 (N_1463,N_1383,N_1365);
or U1464 (N_1464,N_1398,N_1412);
nand U1465 (N_1465,N_1382,N_1360);
nand U1466 (N_1466,N_1398,N_1407);
or U1467 (N_1467,N_1378,N_1410);
nor U1468 (N_1468,N_1382,N_1397);
xnor U1469 (N_1469,N_1388,N_1363);
nor U1470 (N_1470,N_1380,N_1417);
nor U1471 (N_1471,N_1410,N_1372);
and U1472 (N_1472,N_1357,N_1386);
xnor U1473 (N_1473,N_1358,N_1381);
and U1474 (N_1474,N_1370,N_1358);
or U1475 (N_1475,N_1385,N_1414);
nand U1476 (N_1476,N_1394,N_1352);
and U1477 (N_1477,N_1368,N_1398);
or U1478 (N_1478,N_1415,N_1395);
and U1479 (N_1479,N_1350,N_1352);
or U1480 (N_1480,N_1408,N_1418);
nand U1481 (N_1481,N_1363,N_1376);
and U1482 (N_1482,N_1375,N_1360);
nand U1483 (N_1483,N_1389,N_1403);
nand U1484 (N_1484,N_1358,N_1396);
and U1485 (N_1485,N_1381,N_1407);
or U1486 (N_1486,N_1411,N_1375);
or U1487 (N_1487,N_1376,N_1371);
nand U1488 (N_1488,N_1382,N_1384);
nor U1489 (N_1489,N_1421,N_1371);
xnor U1490 (N_1490,N_1371,N_1419);
or U1491 (N_1491,N_1402,N_1356);
and U1492 (N_1492,N_1391,N_1405);
xor U1493 (N_1493,N_1411,N_1396);
or U1494 (N_1494,N_1381,N_1410);
nor U1495 (N_1495,N_1357,N_1368);
and U1496 (N_1496,N_1369,N_1368);
nor U1497 (N_1497,N_1416,N_1393);
nor U1498 (N_1498,N_1350,N_1404);
or U1499 (N_1499,N_1366,N_1370);
xnor U1500 (N_1500,N_1434,N_1491);
and U1501 (N_1501,N_1452,N_1489);
or U1502 (N_1502,N_1455,N_1479);
nand U1503 (N_1503,N_1444,N_1493);
nand U1504 (N_1504,N_1430,N_1461);
nor U1505 (N_1505,N_1473,N_1447);
and U1506 (N_1506,N_1459,N_1441);
or U1507 (N_1507,N_1435,N_1480);
or U1508 (N_1508,N_1437,N_1443);
or U1509 (N_1509,N_1467,N_1497);
nor U1510 (N_1510,N_1427,N_1490);
nand U1511 (N_1511,N_1478,N_1431);
or U1512 (N_1512,N_1474,N_1492);
or U1513 (N_1513,N_1429,N_1440);
and U1514 (N_1514,N_1458,N_1494);
nand U1515 (N_1515,N_1469,N_1476);
or U1516 (N_1516,N_1445,N_1472);
or U1517 (N_1517,N_1471,N_1454);
nand U1518 (N_1518,N_1498,N_1442);
xnor U1519 (N_1519,N_1448,N_1464);
or U1520 (N_1520,N_1470,N_1425);
and U1521 (N_1521,N_1486,N_1468);
and U1522 (N_1522,N_1446,N_1488);
and U1523 (N_1523,N_1456,N_1438);
or U1524 (N_1524,N_1433,N_1457);
or U1525 (N_1525,N_1481,N_1439);
and U1526 (N_1526,N_1484,N_1449);
or U1527 (N_1527,N_1436,N_1465);
nor U1528 (N_1528,N_1483,N_1487);
nor U1529 (N_1529,N_1451,N_1495);
or U1530 (N_1530,N_1499,N_1450);
nor U1531 (N_1531,N_1426,N_1462);
nor U1532 (N_1532,N_1485,N_1477);
nor U1533 (N_1533,N_1460,N_1463);
and U1534 (N_1534,N_1453,N_1466);
nand U1535 (N_1535,N_1428,N_1432);
nand U1536 (N_1536,N_1496,N_1475);
nor U1537 (N_1537,N_1482,N_1467);
and U1538 (N_1538,N_1457,N_1497);
and U1539 (N_1539,N_1490,N_1428);
xnor U1540 (N_1540,N_1479,N_1429);
nand U1541 (N_1541,N_1477,N_1431);
or U1542 (N_1542,N_1454,N_1433);
and U1543 (N_1543,N_1459,N_1466);
nor U1544 (N_1544,N_1475,N_1476);
and U1545 (N_1545,N_1474,N_1428);
and U1546 (N_1546,N_1472,N_1487);
nand U1547 (N_1547,N_1466,N_1492);
or U1548 (N_1548,N_1477,N_1448);
nor U1549 (N_1549,N_1466,N_1474);
or U1550 (N_1550,N_1490,N_1480);
and U1551 (N_1551,N_1433,N_1443);
and U1552 (N_1552,N_1439,N_1468);
and U1553 (N_1553,N_1482,N_1442);
nor U1554 (N_1554,N_1483,N_1446);
xnor U1555 (N_1555,N_1488,N_1486);
nand U1556 (N_1556,N_1483,N_1498);
and U1557 (N_1557,N_1451,N_1498);
nor U1558 (N_1558,N_1474,N_1435);
or U1559 (N_1559,N_1468,N_1436);
and U1560 (N_1560,N_1476,N_1457);
nand U1561 (N_1561,N_1446,N_1436);
or U1562 (N_1562,N_1427,N_1493);
nor U1563 (N_1563,N_1433,N_1479);
nand U1564 (N_1564,N_1454,N_1448);
or U1565 (N_1565,N_1426,N_1441);
nor U1566 (N_1566,N_1480,N_1453);
nand U1567 (N_1567,N_1496,N_1491);
nor U1568 (N_1568,N_1484,N_1438);
nor U1569 (N_1569,N_1497,N_1441);
and U1570 (N_1570,N_1456,N_1485);
xor U1571 (N_1571,N_1482,N_1479);
and U1572 (N_1572,N_1463,N_1461);
or U1573 (N_1573,N_1480,N_1463);
nor U1574 (N_1574,N_1466,N_1467);
nor U1575 (N_1575,N_1527,N_1535);
and U1576 (N_1576,N_1538,N_1506);
nor U1577 (N_1577,N_1522,N_1518);
or U1578 (N_1578,N_1551,N_1547);
nor U1579 (N_1579,N_1563,N_1560);
or U1580 (N_1580,N_1520,N_1531);
and U1581 (N_1581,N_1523,N_1532);
and U1582 (N_1582,N_1524,N_1504);
and U1583 (N_1583,N_1572,N_1521);
or U1584 (N_1584,N_1546,N_1541);
nor U1585 (N_1585,N_1509,N_1544);
or U1586 (N_1586,N_1505,N_1569);
nand U1587 (N_1587,N_1530,N_1565);
nand U1588 (N_1588,N_1537,N_1558);
nor U1589 (N_1589,N_1528,N_1556);
and U1590 (N_1590,N_1514,N_1512);
nand U1591 (N_1591,N_1543,N_1502);
and U1592 (N_1592,N_1510,N_1542);
nor U1593 (N_1593,N_1540,N_1574);
and U1594 (N_1594,N_1508,N_1525);
nor U1595 (N_1595,N_1503,N_1526);
or U1596 (N_1596,N_1549,N_1536);
nand U1597 (N_1597,N_1570,N_1500);
xnor U1598 (N_1598,N_1513,N_1511);
nand U1599 (N_1599,N_1545,N_1559);
or U1600 (N_1600,N_1573,N_1539);
nor U1601 (N_1601,N_1567,N_1552);
and U1602 (N_1602,N_1534,N_1571);
nor U1603 (N_1603,N_1529,N_1561);
nor U1604 (N_1604,N_1507,N_1548);
nor U1605 (N_1605,N_1566,N_1533);
nor U1606 (N_1606,N_1501,N_1555);
xor U1607 (N_1607,N_1519,N_1564);
and U1608 (N_1608,N_1550,N_1516);
nor U1609 (N_1609,N_1515,N_1557);
or U1610 (N_1610,N_1568,N_1562);
nor U1611 (N_1611,N_1517,N_1554);
and U1612 (N_1612,N_1553,N_1523);
nor U1613 (N_1613,N_1512,N_1553);
nand U1614 (N_1614,N_1567,N_1554);
and U1615 (N_1615,N_1569,N_1563);
nor U1616 (N_1616,N_1536,N_1537);
nor U1617 (N_1617,N_1548,N_1557);
nor U1618 (N_1618,N_1518,N_1531);
or U1619 (N_1619,N_1528,N_1516);
and U1620 (N_1620,N_1544,N_1569);
nor U1621 (N_1621,N_1557,N_1518);
and U1622 (N_1622,N_1536,N_1503);
nand U1623 (N_1623,N_1542,N_1503);
nand U1624 (N_1624,N_1513,N_1538);
nor U1625 (N_1625,N_1526,N_1525);
or U1626 (N_1626,N_1540,N_1553);
nor U1627 (N_1627,N_1518,N_1565);
nand U1628 (N_1628,N_1545,N_1521);
and U1629 (N_1629,N_1555,N_1524);
and U1630 (N_1630,N_1529,N_1508);
or U1631 (N_1631,N_1564,N_1500);
or U1632 (N_1632,N_1542,N_1507);
or U1633 (N_1633,N_1558,N_1571);
or U1634 (N_1634,N_1550,N_1527);
and U1635 (N_1635,N_1523,N_1506);
nor U1636 (N_1636,N_1555,N_1546);
xor U1637 (N_1637,N_1516,N_1562);
nor U1638 (N_1638,N_1513,N_1544);
or U1639 (N_1639,N_1568,N_1564);
nand U1640 (N_1640,N_1504,N_1569);
nand U1641 (N_1641,N_1549,N_1514);
and U1642 (N_1642,N_1510,N_1537);
and U1643 (N_1643,N_1504,N_1511);
and U1644 (N_1644,N_1541,N_1522);
xor U1645 (N_1645,N_1501,N_1517);
and U1646 (N_1646,N_1531,N_1516);
nor U1647 (N_1647,N_1538,N_1525);
and U1648 (N_1648,N_1524,N_1515);
nand U1649 (N_1649,N_1538,N_1543);
nand U1650 (N_1650,N_1623,N_1621);
nor U1651 (N_1651,N_1639,N_1588);
or U1652 (N_1652,N_1611,N_1577);
or U1653 (N_1653,N_1595,N_1584);
or U1654 (N_1654,N_1583,N_1609);
or U1655 (N_1655,N_1632,N_1590);
nand U1656 (N_1656,N_1585,N_1643);
nor U1657 (N_1657,N_1635,N_1630);
nand U1658 (N_1658,N_1637,N_1616);
xor U1659 (N_1659,N_1606,N_1582);
nand U1660 (N_1660,N_1642,N_1624);
and U1661 (N_1661,N_1605,N_1598);
and U1662 (N_1662,N_1645,N_1586);
nor U1663 (N_1663,N_1618,N_1581);
nor U1664 (N_1664,N_1612,N_1633);
nand U1665 (N_1665,N_1640,N_1603);
nand U1666 (N_1666,N_1626,N_1625);
nand U1667 (N_1667,N_1649,N_1576);
nor U1668 (N_1668,N_1620,N_1575);
nor U1669 (N_1669,N_1641,N_1614);
and U1670 (N_1670,N_1644,N_1619);
xnor U1671 (N_1671,N_1648,N_1601);
nand U1672 (N_1672,N_1600,N_1593);
nand U1673 (N_1673,N_1579,N_1628);
or U1674 (N_1674,N_1580,N_1629);
nor U1675 (N_1675,N_1610,N_1631);
xnor U1676 (N_1676,N_1599,N_1592);
nor U1677 (N_1677,N_1647,N_1638);
or U1678 (N_1678,N_1591,N_1622);
and U1679 (N_1679,N_1578,N_1597);
nor U1680 (N_1680,N_1607,N_1596);
and U1681 (N_1681,N_1615,N_1608);
and U1682 (N_1682,N_1594,N_1627);
nor U1683 (N_1683,N_1604,N_1589);
or U1684 (N_1684,N_1613,N_1602);
nor U1685 (N_1685,N_1636,N_1646);
or U1686 (N_1686,N_1634,N_1617);
and U1687 (N_1687,N_1587,N_1612);
or U1688 (N_1688,N_1616,N_1590);
and U1689 (N_1689,N_1577,N_1627);
and U1690 (N_1690,N_1609,N_1603);
nor U1691 (N_1691,N_1649,N_1601);
nand U1692 (N_1692,N_1611,N_1647);
nand U1693 (N_1693,N_1606,N_1610);
nand U1694 (N_1694,N_1647,N_1624);
or U1695 (N_1695,N_1642,N_1599);
or U1696 (N_1696,N_1646,N_1596);
nand U1697 (N_1697,N_1605,N_1602);
or U1698 (N_1698,N_1579,N_1577);
nand U1699 (N_1699,N_1615,N_1580);
and U1700 (N_1700,N_1621,N_1647);
or U1701 (N_1701,N_1642,N_1634);
and U1702 (N_1702,N_1589,N_1586);
and U1703 (N_1703,N_1612,N_1589);
nor U1704 (N_1704,N_1603,N_1638);
and U1705 (N_1705,N_1611,N_1621);
xor U1706 (N_1706,N_1645,N_1591);
xnor U1707 (N_1707,N_1629,N_1649);
nor U1708 (N_1708,N_1583,N_1648);
and U1709 (N_1709,N_1640,N_1634);
xor U1710 (N_1710,N_1605,N_1619);
nand U1711 (N_1711,N_1582,N_1577);
nand U1712 (N_1712,N_1577,N_1581);
nand U1713 (N_1713,N_1593,N_1589);
nand U1714 (N_1714,N_1643,N_1618);
or U1715 (N_1715,N_1603,N_1587);
nor U1716 (N_1716,N_1584,N_1593);
or U1717 (N_1717,N_1646,N_1648);
nand U1718 (N_1718,N_1648,N_1616);
nor U1719 (N_1719,N_1622,N_1606);
nor U1720 (N_1720,N_1593,N_1578);
and U1721 (N_1721,N_1583,N_1596);
and U1722 (N_1722,N_1616,N_1595);
nor U1723 (N_1723,N_1630,N_1641);
or U1724 (N_1724,N_1636,N_1575);
or U1725 (N_1725,N_1697,N_1716);
nand U1726 (N_1726,N_1684,N_1664);
and U1727 (N_1727,N_1724,N_1701);
nor U1728 (N_1728,N_1654,N_1653);
nand U1729 (N_1729,N_1702,N_1671);
and U1730 (N_1730,N_1667,N_1696);
nand U1731 (N_1731,N_1699,N_1718);
nand U1732 (N_1732,N_1666,N_1717);
and U1733 (N_1733,N_1707,N_1659);
nand U1734 (N_1734,N_1721,N_1657);
nor U1735 (N_1735,N_1651,N_1709);
or U1736 (N_1736,N_1705,N_1656);
and U1737 (N_1737,N_1675,N_1713);
nand U1738 (N_1738,N_1680,N_1686);
nand U1739 (N_1739,N_1690,N_1681);
xor U1740 (N_1740,N_1694,N_1685);
nor U1741 (N_1741,N_1688,N_1692);
and U1742 (N_1742,N_1691,N_1710);
nand U1743 (N_1743,N_1708,N_1695);
and U1744 (N_1744,N_1720,N_1712);
nand U1745 (N_1745,N_1698,N_1703);
xor U1746 (N_1746,N_1668,N_1660);
nand U1747 (N_1747,N_1683,N_1669);
and U1748 (N_1748,N_1662,N_1719);
or U1749 (N_1749,N_1650,N_1723);
or U1750 (N_1750,N_1706,N_1652);
xor U1751 (N_1751,N_1672,N_1700);
or U1752 (N_1752,N_1655,N_1678);
or U1753 (N_1753,N_1687,N_1674);
nor U1754 (N_1754,N_1714,N_1682);
and U1755 (N_1755,N_1663,N_1665);
or U1756 (N_1756,N_1679,N_1676);
nand U1757 (N_1757,N_1711,N_1677);
xor U1758 (N_1758,N_1661,N_1658);
xnor U1759 (N_1759,N_1693,N_1704);
nor U1760 (N_1760,N_1715,N_1673);
or U1761 (N_1761,N_1722,N_1689);
nand U1762 (N_1762,N_1670,N_1703);
nor U1763 (N_1763,N_1719,N_1653);
or U1764 (N_1764,N_1720,N_1724);
or U1765 (N_1765,N_1663,N_1672);
xnor U1766 (N_1766,N_1707,N_1721);
nor U1767 (N_1767,N_1683,N_1675);
nand U1768 (N_1768,N_1721,N_1651);
or U1769 (N_1769,N_1657,N_1653);
or U1770 (N_1770,N_1655,N_1665);
or U1771 (N_1771,N_1716,N_1685);
xnor U1772 (N_1772,N_1679,N_1720);
and U1773 (N_1773,N_1679,N_1668);
nand U1774 (N_1774,N_1706,N_1711);
nand U1775 (N_1775,N_1713,N_1664);
nand U1776 (N_1776,N_1683,N_1658);
or U1777 (N_1777,N_1656,N_1659);
xnor U1778 (N_1778,N_1719,N_1687);
nor U1779 (N_1779,N_1658,N_1654);
nor U1780 (N_1780,N_1723,N_1660);
nor U1781 (N_1781,N_1657,N_1650);
nand U1782 (N_1782,N_1672,N_1710);
nor U1783 (N_1783,N_1685,N_1702);
nand U1784 (N_1784,N_1657,N_1707);
nor U1785 (N_1785,N_1682,N_1661);
or U1786 (N_1786,N_1717,N_1685);
nand U1787 (N_1787,N_1685,N_1661);
xnor U1788 (N_1788,N_1708,N_1653);
or U1789 (N_1789,N_1694,N_1712);
nor U1790 (N_1790,N_1683,N_1696);
xnor U1791 (N_1791,N_1650,N_1677);
and U1792 (N_1792,N_1697,N_1724);
or U1793 (N_1793,N_1662,N_1720);
or U1794 (N_1794,N_1655,N_1671);
or U1795 (N_1795,N_1661,N_1705);
xnor U1796 (N_1796,N_1694,N_1688);
or U1797 (N_1797,N_1705,N_1691);
xor U1798 (N_1798,N_1681,N_1722);
or U1799 (N_1799,N_1651,N_1670);
or U1800 (N_1800,N_1728,N_1778);
or U1801 (N_1801,N_1726,N_1797);
nand U1802 (N_1802,N_1751,N_1744);
nand U1803 (N_1803,N_1784,N_1736);
nor U1804 (N_1804,N_1787,N_1789);
and U1805 (N_1805,N_1753,N_1746);
and U1806 (N_1806,N_1796,N_1766);
nand U1807 (N_1807,N_1742,N_1750);
or U1808 (N_1808,N_1779,N_1741);
and U1809 (N_1809,N_1792,N_1757);
nor U1810 (N_1810,N_1756,N_1799);
xnor U1811 (N_1811,N_1782,N_1762);
and U1812 (N_1812,N_1775,N_1737);
and U1813 (N_1813,N_1745,N_1776);
nand U1814 (N_1814,N_1738,N_1783);
nand U1815 (N_1815,N_1786,N_1785);
or U1816 (N_1816,N_1767,N_1732);
nor U1817 (N_1817,N_1759,N_1740);
nor U1818 (N_1818,N_1770,N_1725);
nand U1819 (N_1819,N_1795,N_1733);
and U1820 (N_1820,N_1790,N_1772);
nor U1821 (N_1821,N_1771,N_1747);
nand U1822 (N_1822,N_1774,N_1769);
nand U1823 (N_1823,N_1761,N_1739);
xnor U1824 (N_1824,N_1729,N_1793);
nand U1825 (N_1825,N_1760,N_1749);
or U1826 (N_1826,N_1768,N_1781);
xor U1827 (N_1827,N_1763,N_1773);
nand U1828 (N_1828,N_1794,N_1727);
nand U1829 (N_1829,N_1791,N_1752);
or U1830 (N_1830,N_1748,N_1734);
nor U1831 (N_1831,N_1754,N_1758);
and U1832 (N_1832,N_1780,N_1730);
or U1833 (N_1833,N_1743,N_1777);
or U1834 (N_1834,N_1755,N_1788);
nand U1835 (N_1835,N_1735,N_1765);
nand U1836 (N_1836,N_1764,N_1731);
nor U1837 (N_1837,N_1798,N_1775);
or U1838 (N_1838,N_1732,N_1735);
nor U1839 (N_1839,N_1742,N_1791);
or U1840 (N_1840,N_1741,N_1735);
xor U1841 (N_1841,N_1762,N_1789);
or U1842 (N_1842,N_1752,N_1731);
nand U1843 (N_1843,N_1767,N_1788);
nand U1844 (N_1844,N_1780,N_1751);
nor U1845 (N_1845,N_1738,N_1763);
nand U1846 (N_1846,N_1759,N_1796);
and U1847 (N_1847,N_1742,N_1726);
nor U1848 (N_1848,N_1749,N_1752);
nor U1849 (N_1849,N_1726,N_1772);
nand U1850 (N_1850,N_1777,N_1765);
or U1851 (N_1851,N_1729,N_1754);
nand U1852 (N_1852,N_1761,N_1742);
or U1853 (N_1853,N_1797,N_1742);
nand U1854 (N_1854,N_1786,N_1790);
nor U1855 (N_1855,N_1750,N_1792);
nand U1856 (N_1856,N_1783,N_1782);
nand U1857 (N_1857,N_1741,N_1762);
xor U1858 (N_1858,N_1796,N_1736);
nand U1859 (N_1859,N_1743,N_1754);
or U1860 (N_1860,N_1789,N_1794);
and U1861 (N_1861,N_1748,N_1751);
and U1862 (N_1862,N_1735,N_1767);
nand U1863 (N_1863,N_1747,N_1754);
or U1864 (N_1864,N_1794,N_1772);
nor U1865 (N_1865,N_1747,N_1791);
and U1866 (N_1866,N_1733,N_1725);
and U1867 (N_1867,N_1742,N_1776);
nand U1868 (N_1868,N_1762,N_1745);
nand U1869 (N_1869,N_1745,N_1784);
nand U1870 (N_1870,N_1734,N_1733);
nor U1871 (N_1871,N_1737,N_1749);
or U1872 (N_1872,N_1784,N_1737);
xor U1873 (N_1873,N_1779,N_1790);
nor U1874 (N_1874,N_1746,N_1793);
xnor U1875 (N_1875,N_1806,N_1844);
and U1876 (N_1876,N_1817,N_1831);
nand U1877 (N_1877,N_1873,N_1849);
nor U1878 (N_1878,N_1864,N_1848);
or U1879 (N_1879,N_1816,N_1824);
and U1880 (N_1880,N_1805,N_1859);
or U1881 (N_1881,N_1820,N_1851);
nor U1882 (N_1882,N_1815,N_1862);
or U1883 (N_1883,N_1872,N_1860);
and U1884 (N_1884,N_1865,N_1821);
xnor U1885 (N_1885,N_1874,N_1841);
or U1886 (N_1886,N_1866,N_1842);
nor U1887 (N_1887,N_1858,N_1861);
nand U1888 (N_1888,N_1830,N_1818);
nor U1889 (N_1889,N_1856,N_1809);
nand U1890 (N_1890,N_1843,N_1863);
nand U1891 (N_1891,N_1854,N_1835);
nor U1892 (N_1892,N_1828,N_1803);
or U1893 (N_1893,N_1804,N_1833);
or U1894 (N_1894,N_1847,N_1870);
or U1895 (N_1895,N_1868,N_1838);
or U1896 (N_1896,N_1813,N_1802);
and U1897 (N_1897,N_1822,N_1808);
xor U1898 (N_1898,N_1840,N_1845);
and U1899 (N_1899,N_1846,N_1807);
or U1900 (N_1900,N_1837,N_1850);
or U1901 (N_1901,N_1825,N_1811);
nand U1902 (N_1902,N_1867,N_1801);
nand U1903 (N_1903,N_1826,N_1829);
or U1904 (N_1904,N_1834,N_1839);
or U1905 (N_1905,N_1855,N_1827);
nand U1906 (N_1906,N_1810,N_1852);
and U1907 (N_1907,N_1819,N_1800);
nand U1908 (N_1908,N_1823,N_1814);
xnor U1909 (N_1909,N_1832,N_1812);
xor U1910 (N_1910,N_1857,N_1836);
or U1911 (N_1911,N_1869,N_1853);
nand U1912 (N_1912,N_1871,N_1821);
or U1913 (N_1913,N_1825,N_1846);
nand U1914 (N_1914,N_1803,N_1852);
nand U1915 (N_1915,N_1853,N_1840);
nand U1916 (N_1916,N_1816,N_1858);
nor U1917 (N_1917,N_1833,N_1827);
nor U1918 (N_1918,N_1824,N_1814);
nor U1919 (N_1919,N_1818,N_1807);
and U1920 (N_1920,N_1834,N_1805);
or U1921 (N_1921,N_1861,N_1811);
xnor U1922 (N_1922,N_1872,N_1841);
and U1923 (N_1923,N_1815,N_1864);
xor U1924 (N_1924,N_1819,N_1822);
nor U1925 (N_1925,N_1850,N_1867);
nor U1926 (N_1926,N_1862,N_1842);
nor U1927 (N_1927,N_1813,N_1871);
and U1928 (N_1928,N_1853,N_1859);
nor U1929 (N_1929,N_1804,N_1816);
or U1930 (N_1930,N_1823,N_1805);
xnor U1931 (N_1931,N_1826,N_1870);
or U1932 (N_1932,N_1821,N_1869);
xnor U1933 (N_1933,N_1853,N_1862);
xnor U1934 (N_1934,N_1821,N_1852);
nor U1935 (N_1935,N_1854,N_1847);
xnor U1936 (N_1936,N_1854,N_1867);
nor U1937 (N_1937,N_1816,N_1815);
nor U1938 (N_1938,N_1807,N_1839);
nand U1939 (N_1939,N_1858,N_1871);
nand U1940 (N_1940,N_1803,N_1804);
xnor U1941 (N_1941,N_1824,N_1858);
nor U1942 (N_1942,N_1846,N_1827);
or U1943 (N_1943,N_1852,N_1854);
or U1944 (N_1944,N_1871,N_1855);
nand U1945 (N_1945,N_1847,N_1856);
and U1946 (N_1946,N_1856,N_1874);
nor U1947 (N_1947,N_1840,N_1838);
and U1948 (N_1948,N_1869,N_1842);
nand U1949 (N_1949,N_1818,N_1810);
nand U1950 (N_1950,N_1910,N_1918);
xnor U1951 (N_1951,N_1905,N_1908);
or U1952 (N_1952,N_1878,N_1925);
and U1953 (N_1953,N_1916,N_1897);
and U1954 (N_1954,N_1913,N_1893);
nor U1955 (N_1955,N_1880,N_1892);
nand U1956 (N_1956,N_1909,N_1887);
or U1957 (N_1957,N_1920,N_1900);
and U1958 (N_1958,N_1876,N_1895);
or U1959 (N_1959,N_1902,N_1935);
and U1960 (N_1960,N_1923,N_1932);
xor U1961 (N_1961,N_1930,N_1942);
nor U1962 (N_1962,N_1883,N_1943);
nand U1963 (N_1963,N_1924,N_1927);
xor U1964 (N_1964,N_1945,N_1933);
and U1965 (N_1965,N_1946,N_1901);
nand U1966 (N_1966,N_1904,N_1934);
nor U1967 (N_1967,N_1907,N_1899);
xnor U1968 (N_1968,N_1915,N_1884);
nand U1969 (N_1969,N_1898,N_1877);
and U1970 (N_1970,N_1882,N_1888);
and U1971 (N_1971,N_1890,N_1903);
or U1972 (N_1972,N_1937,N_1875);
nor U1973 (N_1973,N_1947,N_1948);
nor U1974 (N_1974,N_1938,N_1896);
and U1975 (N_1975,N_1940,N_1889);
or U1976 (N_1976,N_1906,N_1891);
and U1977 (N_1977,N_1881,N_1921);
nand U1978 (N_1978,N_1879,N_1914);
nor U1979 (N_1979,N_1885,N_1922);
xor U1980 (N_1980,N_1936,N_1949);
or U1981 (N_1981,N_1911,N_1928);
nor U1982 (N_1982,N_1894,N_1912);
or U1983 (N_1983,N_1939,N_1926);
or U1984 (N_1984,N_1917,N_1944);
nor U1985 (N_1985,N_1941,N_1919);
xnor U1986 (N_1986,N_1929,N_1931);
nand U1987 (N_1987,N_1886,N_1904);
and U1988 (N_1988,N_1933,N_1947);
or U1989 (N_1989,N_1883,N_1905);
nor U1990 (N_1990,N_1945,N_1901);
and U1991 (N_1991,N_1929,N_1899);
nand U1992 (N_1992,N_1936,N_1902);
and U1993 (N_1993,N_1944,N_1927);
and U1994 (N_1994,N_1906,N_1918);
or U1995 (N_1995,N_1934,N_1876);
or U1996 (N_1996,N_1896,N_1884);
nor U1997 (N_1997,N_1912,N_1942);
xor U1998 (N_1998,N_1921,N_1945);
or U1999 (N_1999,N_1932,N_1944);
or U2000 (N_2000,N_1887,N_1937);
nand U2001 (N_2001,N_1877,N_1928);
or U2002 (N_2002,N_1939,N_1902);
and U2003 (N_2003,N_1916,N_1924);
nor U2004 (N_2004,N_1933,N_1920);
nor U2005 (N_2005,N_1907,N_1919);
or U2006 (N_2006,N_1896,N_1892);
nand U2007 (N_2007,N_1937,N_1905);
nand U2008 (N_2008,N_1921,N_1888);
and U2009 (N_2009,N_1877,N_1885);
nand U2010 (N_2010,N_1887,N_1915);
nand U2011 (N_2011,N_1914,N_1892);
and U2012 (N_2012,N_1931,N_1910);
or U2013 (N_2013,N_1901,N_1893);
and U2014 (N_2014,N_1911,N_1922);
and U2015 (N_2015,N_1895,N_1878);
and U2016 (N_2016,N_1877,N_1881);
and U2017 (N_2017,N_1929,N_1939);
and U2018 (N_2018,N_1911,N_1926);
or U2019 (N_2019,N_1909,N_1903);
nand U2020 (N_2020,N_1936,N_1891);
nor U2021 (N_2021,N_1879,N_1935);
nor U2022 (N_2022,N_1915,N_1892);
or U2023 (N_2023,N_1923,N_1893);
and U2024 (N_2024,N_1934,N_1882);
and U2025 (N_2025,N_1953,N_2019);
nand U2026 (N_2026,N_1970,N_2023);
nor U2027 (N_2027,N_1967,N_1977);
nor U2028 (N_2028,N_1957,N_1988);
xnor U2029 (N_2029,N_1976,N_1954);
or U2030 (N_2030,N_2005,N_2018);
nor U2031 (N_2031,N_2004,N_1955);
nor U2032 (N_2032,N_1983,N_2001);
nor U2033 (N_2033,N_1972,N_1965);
xor U2034 (N_2034,N_1962,N_1996);
and U2035 (N_2035,N_1979,N_2021);
or U2036 (N_2036,N_2013,N_1987);
xor U2037 (N_2037,N_1956,N_1999);
nand U2038 (N_2038,N_2017,N_1978);
nor U2039 (N_2039,N_1994,N_2015);
and U2040 (N_2040,N_2011,N_1980);
or U2041 (N_2041,N_1992,N_1986);
or U2042 (N_2042,N_1991,N_2006);
nor U2043 (N_2043,N_1958,N_1974);
nand U2044 (N_2044,N_1989,N_1961);
or U2045 (N_2045,N_1968,N_2014);
nand U2046 (N_2046,N_1997,N_1951);
or U2047 (N_2047,N_2010,N_1950);
and U2048 (N_2048,N_1971,N_2008);
nor U2049 (N_2049,N_1960,N_2000);
or U2050 (N_2050,N_2009,N_1964);
nor U2051 (N_2051,N_1993,N_2016);
and U2052 (N_2052,N_1995,N_1973);
or U2053 (N_2053,N_2007,N_2020);
nand U2054 (N_2054,N_1984,N_1952);
or U2055 (N_2055,N_1998,N_1966);
and U2056 (N_2056,N_1982,N_1981);
nand U2057 (N_2057,N_1990,N_2022);
or U2058 (N_2058,N_2012,N_2003);
or U2059 (N_2059,N_2002,N_1959);
and U2060 (N_2060,N_1969,N_2024);
or U2061 (N_2061,N_1985,N_1975);
and U2062 (N_2062,N_1963,N_1953);
and U2063 (N_2063,N_2002,N_2021);
or U2064 (N_2064,N_1955,N_2013);
or U2065 (N_2065,N_1969,N_2004);
or U2066 (N_2066,N_1953,N_1974);
nor U2067 (N_2067,N_2021,N_1985);
nor U2068 (N_2068,N_1966,N_1986);
nor U2069 (N_2069,N_1978,N_1979);
nand U2070 (N_2070,N_1974,N_1989);
or U2071 (N_2071,N_1961,N_2000);
or U2072 (N_2072,N_2001,N_1995);
nand U2073 (N_2073,N_1958,N_2001);
nor U2074 (N_2074,N_1966,N_2016);
and U2075 (N_2075,N_2005,N_1961);
or U2076 (N_2076,N_1956,N_1955);
nand U2077 (N_2077,N_1977,N_1968);
nor U2078 (N_2078,N_1962,N_1954);
nand U2079 (N_2079,N_1966,N_1989);
nand U2080 (N_2080,N_1997,N_2000);
nand U2081 (N_2081,N_1994,N_2008);
xnor U2082 (N_2082,N_2014,N_2006);
nand U2083 (N_2083,N_2020,N_2018);
and U2084 (N_2084,N_2014,N_1969);
nand U2085 (N_2085,N_1995,N_1989);
or U2086 (N_2086,N_1965,N_1953);
or U2087 (N_2087,N_1995,N_2018);
nand U2088 (N_2088,N_2006,N_1982);
nor U2089 (N_2089,N_1973,N_1988);
or U2090 (N_2090,N_1950,N_1967);
or U2091 (N_2091,N_2016,N_1955);
nand U2092 (N_2092,N_2011,N_1991);
nor U2093 (N_2093,N_1974,N_1985);
nand U2094 (N_2094,N_1991,N_1962);
nand U2095 (N_2095,N_1993,N_2015);
nand U2096 (N_2096,N_2005,N_1957);
or U2097 (N_2097,N_2008,N_2021);
and U2098 (N_2098,N_1985,N_1966);
or U2099 (N_2099,N_2004,N_1979);
nand U2100 (N_2100,N_2098,N_2049);
and U2101 (N_2101,N_2054,N_2025);
and U2102 (N_2102,N_2080,N_2090);
and U2103 (N_2103,N_2036,N_2057);
nand U2104 (N_2104,N_2067,N_2047);
or U2105 (N_2105,N_2081,N_2092);
and U2106 (N_2106,N_2071,N_2091);
and U2107 (N_2107,N_2060,N_2074);
xnor U2108 (N_2108,N_2097,N_2072);
xnor U2109 (N_2109,N_2038,N_2093);
and U2110 (N_2110,N_2084,N_2037);
nand U2111 (N_2111,N_2095,N_2064);
or U2112 (N_2112,N_2035,N_2089);
nand U2113 (N_2113,N_2086,N_2056);
nand U2114 (N_2114,N_2042,N_2033);
and U2115 (N_2115,N_2055,N_2050);
xor U2116 (N_2116,N_2045,N_2039);
xnor U2117 (N_2117,N_2066,N_2068);
or U2118 (N_2118,N_2051,N_2079);
or U2119 (N_2119,N_2034,N_2048);
nor U2120 (N_2120,N_2063,N_2077);
nor U2121 (N_2121,N_2026,N_2076);
and U2122 (N_2122,N_2099,N_2032);
and U2123 (N_2123,N_2043,N_2052);
or U2124 (N_2124,N_2053,N_2094);
nand U2125 (N_2125,N_2069,N_2082);
nor U2126 (N_2126,N_2096,N_2046);
and U2127 (N_2127,N_2040,N_2078);
nor U2128 (N_2128,N_2065,N_2087);
or U2129 (N_2129,N_2059,N_2031);
xnor U2130 (N_2130,N_2070,N_2041);
xnor U2131 (N_2131,N_2061,N_2083);
nand U2132 (N_2132,N_2058,N_2029);
nor U2133 (N_2133,N_2073,N_2027);
and U2134 (N_2134,N_2062,N_2030);
or U2135 (N_2135,N_2044,N_2028);
or U2136 (N_2136,N_2085,N_2075);
or U2137 (N_2137,N_2088,N_2035);
nor U2138 (N_2138,N_2025,N_2092);
xor U2139 (N_2139,N_2052,N_2078);
or U2140 (N_2140,N_2044,N_2050);
nor U2141 (N_2141,N_2066,N_2071);
nand U2142 (N_2142,N_2078,N_2087);
xnor U2143 (N_2143,N_2096,N_2084);
nor U2144 (N_2144,N_2087,N_2070);
nor U2145 (N_2145,N_2090,N_2082);
xor U2146 (N_2146,N_2078,N_2051);
nand U2147 (N_2147,N_2062,N_2074);
and U2148 (N_2148,N_2093,N_2042);
nand U2149 (N_2149,N_2046,N_2075);
or U2150 (N_2150,N_2072,N_2092);
nand U2151 (N_2151,N_2069,N_2081);
or U2152 (N_2152,N_2064,N_2074);
or U2153 (N_2153,N_2028,N_2050);
xor U2154 (N_2154,N_2045,N_2082);
or U2155 (N_2155,N_2031,N_2041);
xnor U2156 (N_2156,N_2028,N_2036);
nor U2157 (N_2157,N_2091,N_2083);
or U2158 (N_2158,N_2096,N_2038);
xnor U2159 (N_2159,N_2099,N_2097);
nand U2160 (N_2160,N_2051,N_2093);
nand U2161 (N_2161,N_2051,N_2085);
or U2162 (N_2162,N_2068,N_2072);
nand U2163 (N_2163,N_2060,N_2030);
nor U2164 (N_2164,N_2060,N_2077);
or U2165 (N_2165,N_2063,N_2081);
nor U2166 (N_2166,N_2036,N_2082);
xor U2167 (N_2167,N_2062,N_2027);
nor U2168 (N_2168,N_2077,N_2038);
nand U2169 (N_2169,N_2061,N_2088);
and U2170 (N_2170,N_2071,N_2085);
xnor U2171 (N_2171,N_2078,N_2045);
or U2172 (N_2172,N_2056,N_2045);
nor U2173 (N_2173,N_2027,N_2042);
or U2174 (N_2174,N_2027,N_2057);
or U2175 (N_2175,N_2122,N_2123);
and U2176 (N_2176,N_2127,N_2124);
nand U2177 (N_2177,N_2152,N_2161);
xor U2178 (N_2178,N_2113,N_2119);
nor U2179 (N_2179,N_2157,N_2126);
nor U2180 (N_2180,N_2112,N_2118);
nand U2181 (N_2181,N_2141,N_2132);
nand U2182 (N_2182,N_2131,N_2163);
nor U2183 (N_2183,N_2162,N_2135);
nor U2184 (N_2184,N_2108,N_2101);
nand U2185 (N_2185,N_2153,N_2109);
or U2186 (N_2186,N_2154,N_2147);
or U2187 (N_2187,N_2144,N_2130);
and U2188 (N_2188,N_2160,N_2146);
or U2189 (N_2189,N_2138,N_2174);
xor U2190 (N_2190,N_2120,N_2167);
or U2191 (N_2191,N_2100,N_2142);
and U2192 (N_2192,N_2103,N_2164);
nand U2193 (N_2193,N_2125,N_2102);
nor U2194 (N_2194,N_2143,N_2114);
nand U2195 (N_2195,N_2121,N_2106);
xor U2196 (N_2196,N_2145,N_2137);
nand U2197 (N_2197,N_2173,N_2140);
nand U2198 (N_2198,N_2117,N_2165);
xnor U2199 (N_2199,N_2139,N_2110);
nand U2200 (N_2200,N_2148,N_2169);
and U2201 (N_2201,N_2159,N_2171);
xnor U2202 (N_2202,N_2128,N_2133);
or U2203 (N_2203,N_2170,N_2166);
nand U2204 (N_2204,N_2136,N_2156);
xnor U2205 (N_2205,N_2172,N_2155);
nor U2206 (N_2206,N_2105,N_2129);
nor U2207 (N_2207,N_2149,N_2111);
or U2208 (N_2208,N_2168,N_2150);
nor U2209 (N_2209,N_2115,N_2116);
and U2210 (N_2210,N_2104,N_2107);
nand U2211 (N_2211,N_2151,N_2134);
nor U2212 (N_2212,N_2158,N_2144);
and U2213 (N_2213,N_2115,N_2156);
or U2214 (N_2214,N_2111,N_2114);
nor U2215 (N_2215,N_2127,N_2133);
nand U2216 (N_2216,N_2147,N_2153);
nand U2217 (N_2217,N_2144,N_2173);
nor U2218 (N_2218,N_2141,N_2161);
and U2219 (N_2219,N_2173,N_2129);
or U2220 (N_2220,N_2145,N_2109);
or U2221 (N_2221,N_2112,N_2119);
nor U2222 (N_2222,N_2108,N_2146);
and U2223 (N_2223,N_2171,N_2167);
nand U2224 (N_2224,N_2135,N_2141);
nand U2225 (N_2225,N_2151,N_2111);
and U2226 (N_2226,N_2109,N_2139);
and U2227 (N_2227,N_2165,N_2141);
nor U2228 (N_2228,N_2101,N_2110);
nor U2229 (N_2229,N_2145,N_2104);
nand U2230 (N_2230,N_2106,N_2169);
nor U2231 (N_2231,N_2172,N_2163);
or U2232 (N_2232,N_2173,N_2109);
or U2233 (N_2233,N_2124,N_2145);
and U2234 (N_2234,N_2109,N_2168);
and U2235 (N_2235,N_2151,N_2118);
or U2236 (N_2236,N_2129,N_2107);
nand U2237 (N_2237,N_2169,N_2162);
or U2238 (N_2238,N_2127,N_2137);
and U2239 (N_2239,N_2162,N_2123);
nand U2240 (N_2240,N_2105,N_2120);
or U2241 (N_2241,N_2146,N_2140);
or U2242 (N_2242,N_2110,N_2137);
or U2243 (N_2243,N_2108,N_2141);
nor U2244 (N_2244,N_2143,N_2125);
nor U2245 (N_2245,N_2143,N_2173);
and U2246 (N_2246,N_2166,N_2143);
nor U2247 (N_2247,N_2122,N_2142);
nor U2248 (N_2248,N_2107,N_2159);
nand U2249 (N_2249,N_2118,N_2115);
xor U2250 (N_2250,N_2187,N_2209);
and U2251 (N_2251,N_2228,N_2198);
and U2252 (N_2252,N_2248,N_2207);
and U2253 (N_2253,N_2223,N_2201);
xor U2254 (N_2254,N_2175,N_2217);
xnor U2255 (N_2255,N_2224,N_2238);
nand U2256 (N_2256,N_2216,N_2243);
nand U2257 (N_2257,N_2194,N_2179);
and U2258 (N_2258,N_2239,N_2210);
nor U2259 (N_2259,N_2176,N_2190);
nor U2260 (N_2260,N_2191,N_2204);
nand U2261 (N_2261,N_2213,N_2202);
xnor U2262 (N_2262,N_2180,N_2195);
nand U2263 (N_2263,N_2181,N_2214);
and U2264 (N_2264,N_2203,N_2222);
and U2265 (N_2265,N_2232,N_2233);
or U2266 (N_2266,N_2184,N_2226);
and U2267 (N_2267,N_2246,N_2177);
xor U2268 (N_2268,N_2197,N_2247);
nand U2269 (N_2269,N_2241,N_2189);
and U2270 (N_2270,N_2242,N_2249);
xnor U2271 (N_2271,N_2188,N_2225);
nor U2272 (N_2272,N_2211,N_2205);
or U2273 (N_2273,N_2245,N_2185);
or U2274 (N_2274,N_2178,N_2219);
and U2275 (N_2275,N_2182,N_2221);
xor U2276 (N_2276,N_2230,N_2240);
or U2277 (N_2277,N_2186,N_2196);
nor U2278 (N_2278,N_2218,N_2183);
nand U2279 (N_2279,N_2237,N_2220);
nand U2280 (N_2280,N_2192,N_2227);
nor U2281 (N_2281,N_2200,N_2215);
xnor U2282 (N_2282,N_2231,N_2199);
nor U2283 (N_2283,N_2193,N_2236);
or U2284 (N_2284,N_2212,N_2208);
xor U2285 (N_2285,N_2229,N_2234);
or U2286 (N_2286,N_2206,N_2244);
and U2287 (N_2287,N_2235,N_2248);
nor U2288 (N_2288,N_2245,N_2247);
xnor U2289 (N_2289,N_2209,N_2208);
nor U2290 (N_2290,N_2246,N_2179);
nor U2291 (N_2291,N_2200,N_2232);
nand U2292 (N_2292,N_2181,N_2236);
and U2293 (N_2293,N_2226,N_2210);
and U2294 (N_2294,N_2196,N_2235);
and U2295 (N_2295,N_2196,N_2190);
nand U2296 (N_2296,N_2205,N_2226);
nand U2297 (N_2297,N_2181,N_2188);
and U2298 (N_2298,N_2249,N_2191);
or U2299 (N_2299,N_2183,N_2217);
xnor U2300 (N_2300,N_2235,N_2240);
and U2301 (N_2301,N_2227,N_2183);
nand U2302 (N_2302,N_2183,N_2235);
or U2303 (N_2303,N_2199,N_2228);
or U2304 (N_2304,N_2233,N_2192);
nand U2305 (N_2305,N_2199,N_2216);
or U2306 (N_2306,N_2233,N_2211);
and U2307 (N_2307,N_2185,N_2240);
or U2308 (N_2308,N_2192,N_2207);
or U2309 (N_2309,N_2242,N_2212);
and U2310 (N_2310,N_2218,N_2178);
and U2311 (N_2311,N_2201,N_2202);
nor U2312 (N_2312,N_2198,N_2210);
nor U2313 (N_2313,N_2247,N_2240);
or U2314 (N_2314,N_2214,N_2249);
and U2315 (N_2315,N_2216,N_2234);
nor U2316 (N_2316,N_2213,N_2187);
and U2317 (N_2317,N_2184,N_2215);
nor U2318 (N_2318,N_2235,N_2229);
nand U2319 (N_2319,N_2179,N_2176);
or U2320 (N_2320,N_2242,N_2178);
nor U2321 (N_2321,N_2181,N_2231);
and U2322 (N_2322,N_2241,N_2235);
nor U2323 (N_2323,N_2207,N_2191);
xor U2324 (N_2324,N_2221,N_2247);
nor U2325 (N_2325,N_2299,N_2281);
nor U2326 (N_2326,N_2262,N_2291);
nand U2327 (N_2327,N_2276,N_2277);
nor U2328 (N_2328,N_2319,N_2305);
and U2329 (N_2329,N_2298,N_2293);
and U2330 (N_2330,N_2313,N_2316);
and U2331 (N_2331,N_2275,N_2321);
nand U2332 (N_2332,N_2278,N_2280);
nor U2333 (N_2333,N_2263,N_2315);
nor U2334 (N_2334,N_2297,N_2270);
nand U2335 (N_2335,N_2282,N_2308);
nor U2336 (N_2336,N_2260,N_2311);
nor U2337 (N_2337,N_2286,N_2296);
or U2338 (N_2338,N_2252,N_2307);
and U2339 (N_2339,N_2258,N_2273);
and U2340 (N_2340,N_2324,N_2292);
nand U2341 (N_2341,N_2322,N_2283);
and U2342 (N_2342,N_2250,N_2279);
nor U2343 (N_2343,N_2253,N_2269);
or U2344 (N_2344,N_2302,N_2295);
and U2345 (N_2345,N_2267,N_2301);
nor U2346 (N_2346,N_2310,N_2287);
and U2347 (N_2347,N_2266,N_2264);
and U2348 (N_2348,N_2290,N_2318);
nor U2349 (N_2349,N_2256,N_2323);
or U2350 (N_2350,N_2303,N_2317);
nand U2351 (N_2351,N_2309,N_2314);
xnor U2352 (N_2352,N_2288,N_2274);
nand U2353 (N_2353,N_2272,N_2320);
nand U2354 (N_2354,N_2251,N_2294);
or U2355 (N_2355,N_2257,N_2306);
and U2356 (N_2356,N_2271,N_2285);
nand U2357 (N_2357,N_2255,N_2284);
and U2358 (N_2358,N_2300,N_2289);
and U2359 (N_2359,N_2265,N_2261);
or U2360 (N_2360,N_2304,N_2312);
and U2361 (N_2361,N_2259,N_2254);
and U2362 (N_2362,N_2268,N_2271);
and U2363 (N_2363,N_2300,N_2294);
or U2364 (N_2364,N_2255,N_2278);
or U2365 (N_2365,N_2307,N_2259);
or U2366 (N_2366,N_2260,N_2276);
and U2367 (N_2367,N_2253,N_2264);
and U2368 (N_2368,N_2259,N_2293);
nor U2369 (N_2369,N_2301,N_2269);
nand U2370 (N_2370,N_2250,N_2308);
xor U2371 (N_2371,N_2313,N_2261);
and U2372 (N_2372,N_2321,N_2310);
or U2373 (N_2373,N_2255,N_2252);
nor U2374 (N_2374,N_2303,N_2286);
or U2375 (N_2375,N_2317,N_2311);
nor U2376 (N_2376,N_2316,N_2291);
nand U2377 (N_2377,N_2267,N_2299);
and U2378 (N_2378,N_2323,N_2262);
nand U2379 (N_2379,N_2309,N_2271);
nand U2380 (N_2380,N_2324,N_2322);
and U2381 (N_2381,N_2261,N_2255);
and U2382 (N_2382,N_2280,N_2272);
and U2383 (N_2383,N_2298,N_2268);
and U2384 (N_2384,N_2313,N_2257);
nor U2385 (N_2385,N_2309,N_2307);
or U2386 (N_2386,N_2314,N_2300);
and U2387 (N_2387,N_2284,N_2253);
nor U2388 (N_2388,N_2307,N_2267);
and U2389 (N_2389,N_2286,N_2324);
and U2390 (N_2390,N_2324,N_2284);
and U2391 (N_2391,N_2307,N_2293);
and U2392 (N_2392,N_2267,N_2273);
and U2393 (N_2393,N_2265,N_2275);
or U2394 (N_2394,N_2268,N_2302);
nor U2395 (N_2395,N_2253,N_2321);
and U2396 (N_2396,N_2250,N_2301);
nand U2397 (N_2397,N_2311,N_2323);
and U2398 (N_2398,N_2275,N_2303);
xor U2399 (N_2399,N_2308,N_2260);
or U2400 (N_2400,N_2389,N_2339);
and U2401 (N_2401,N_2377,N_2364);
and U2402 (N_2402,N_2327,N_2382);
or U2403 (N_2403,N_2385,N_2340);
and U2404 (N_2404,N_2390,N_2370);
or U2405 (N_2405,N_2345,N_2365);
nor U2406 (N_2406,N_2380,N_2337);
nor U2407 (N_2407,N_2394,N_2343);
or U2408 (N_2408,N_2393,N_2352);
or U2409 (N_2409,N_2354,N_2346);
nor U2410 (N_2410,N_2330,N_2384);
and U2411 (N_2411,N_2342,N_2399);
nor U2412 (N_2412,N_2332,N_2387);
or U2413 (N_2413,N_2328,N_2341);
or U2414 (N_2414,N_2361,N_2347);
nand U2415 (N_2415,N_2386,N_2325);
nand U2416 (N_2416,N_2391,N_2392);
nand U2417 (N_2417,N_2355,N_2326);
and U2418 (N_2418,N_2388,N_2398);
nand U2419 (N_2419,N_2378,N_2333);
nand U2420 (N_2420,N_2397,N_2338);
nand U2421 (N_2421,N_2369,N_2350);
nor U2422 (N_2422,N_2334,N_2396);
nand U2423 (N_2423,N_2395,N_2372);
or U2424 (N_2424,N_2381,N_2331);
nor U2425 (N_2425,N_2351,N_2360);
or U2426 (N_2426,N_2358,N_2367);
or U2427 (N_2427,N_2348,N_2375);
or U2428 (N_2428,N_2359,N_2383);
or U2429 (N_2429,N_2373,N_2368);
xor U2430 (N_2430,N_2336,N_2379);
or U2431 (N_2431,N_2349,N_2362);
xor U2432 (N_2432,N_2371,N_2363);
or U2433 (N_2433,N_2329,N_2357);
xnor U2434 (N_2434,N_2344,N_2335);
and U2435 (N_2435,N_2374,N_2353);
and U2436 (N_2436,N_2366,N_2356);
or U2437 (N_2437,N_2376,N_2331);
or U2438 (N_2438,N_2344,N_2327);
and U2439 (N_2439,N_2377,N_2358);
nand U2440 (N_2440,N_2371,N_2358);
or U2441 (N_2441,N_2353,N_2351);
nand U2442 (N_2442,N_2369,N_2372);
nor U2443 (N_2443,N_2333,N_2393);
or U2444 (N_2444,N_2347,N_2337);
xor U2445 (N_2445,N_2372,N_2381);
nand U2446 (N_2446,N_2379,N_2359);
nor U2447 (N_2447,N_2334,N_2343);
nor U2448 (N_2448,N_2350,N_2393);
or U2449 (N_2449,N_2361,N_2350);
and U2450 (N_2450,N_2326,N_2344);
or U2451 (N_2451,N_2384,N_2390);
and U2452 (N_2452,N_2399,N_2398);
or U2453 (N_2453,N_2378,N_2385);
nand U2454 (N_2454,N_2340,N_2363);
xnor U2455 (N_2455,N_2371,N_2356);
nand U2456 (N_2456,N_2394,N_2326);
nand U2457 (N_2457,N_2372,N_2385);
or U2458 (N_2458,N_2346,N_2366);
nor U2459 (N_2459,N_2333,N_2372);
nand U2460 (N_2460,N_2366,N_2344);
nor U2461 (N_2461,N_2355,N_2348);
nor U2462 (N_2462,N_2393,N_2381);
xor U2463 (N_2463,N_2386,N_2377);
nand U2464 (N_2464,N_2370,N_2389);
nand U2465 (N_2465,N_2390,N_2392);
or U2466 (N_2466,N_2391,N_2396);
and U2467 (N_2467,N_2383,N_2335);
nor U2468 (N_2468,N_2380,N_2395);
nand U2469 (N_2469,N_2381,N_2339);
and U2470 (N_2470,N_2342,N_2388);
nor U2471 (N_2471,N_2393,N_2347);
nor U2472 (N_2472,N_2327,N_2389);
nand U2473 (N_2473,N_2355,N_2360);
and U2474 (N_2474,N_2388,N_2365);
xor U2475 (N_2475,N_2474,N_2444);
nor U2476 (N_2476,N_2407,N_2471);
or U2477 (N_2477,N_2456,N_2459);
and U2478 (N_2478,N_2417,N_2401);
nand U2479 (N_2479,N_2426,N_2422);
nor U2480 (N_2480,N_2441,N_2410);
nor U2481 (N_2481,N_2433,N_2458);
nand U2482 (N_2482,N_2466,N_2447);
nor U2483 (N_2483,N_2429,N_2430);
and U2484 (N_2484,N_2468,N_2420);
nor U2485 (N_2485,N_2415,N_2469);
nor U2486 (N_2486,N_2473,N_2409);
nand U2487 (N_2487,N_2438,N_2428);
or U2488 (N_2488,N_2434,N_2465);
xor U2489 (N_2489,N_2463,N_2431);
nand U2490 (N_2490,N_2436,N_2424);
nor U2491 (N_2491,N_2450,N_2413);
or U2492 (N_2492,N_2451,N_2427);
nand U2493 (N_2493,N_2455,N_2400);
and U2494 (N_2494,N_2404,N_2439);
or U2495 (N_2495,N_2425,N_2443);
nand U2496 (N_2496,N_2402,N_2449);
nand U2497 (N_2497,N_2472,N_2421);
xor U2498 (N_2498,N_2414,N_2446);
or U2499 (N_2499,N_2453,N_2452);
or U2500 (N_2500,N_2435,N_2462);
nor U2501 (N_2501,N_2423,N_2437);
nor U2502 (N_2502,N_2416,N_2467);
or U2503 (N_2503,N_2406,N_2403);
xor U2504 (N_2504,N_2448,N_2411);
nand U2505 (N_2505,N_2461,N_2460);
nand U2506 (N_2506,N_2457,N_2432);
or U2507 (N_2507,N_2442,N_2405);
or U2508 (N_2508,N_2408,N_2412);
or U2509 (N_2509,N_2418,N_2440);
nor U2510 (N_2510,N_2419,N_2445);
or U2511 (N_2511,N_2470,N_2464);
nor U2512 (N_2512,N_2454,N_2447);
and U2513 (N_2513,N_2460,N_2455);
nand U2514 (N_2514,N_2467,N_2460);
nand U2515 (N_2515,N_2411,N_2473);
and U2516 (N_2516,N_2404,N_2460);
or U2517 (N_2517,N_2420,N_2418);
nand U2518 (N_2518,N_2435,N_2429);
or U2519 (N_2519,N_2414,N_2402);
or U2520 (N_2520,N_2405,N_2454);
and U2521 (N_2521,N_2403,N_2471);
and U2522 (N_2522,N_2454,N_2421);
or U2523 (N_2523,N_2473,N_2459);
nand U2524 (N_2524,N_2468,N_2432);
nand U2525 (N_2525,N_2409,N_2449);
and U2526 (N_2526,N_2405,N_2425);
nand U2527 (N_2527,N_2419,N_2420);
xor U2528 (N_2528,N_2456,N_2442);
or U2529 (N_2529,N_2410,N_2412);
nand U2530 (N_2530,N_2427,N_2430);
or U2531 (N_2531,N_2446,N_2440);
nand U2532 (N_2532,N_2463,N_2411);
xor U2533 (N_2533,N_2433,N_2421);
or U2534 (N_2534,N_2471,N_2433);
nand U2535 (N_2535,N_2450,N_2462);
or U2536 (N_2536,N_2466,N_2471);
nand U2537 (N_2537,N_2429,N_2436);
or U2538 (N_2538,N_2432,N_2404);
and U2539 (N_2539,N_2457,N_2442);
xor U2540 (N_2540,N_2467,N_2472);
and U2541 (N_2541,N_2404,N_2437);
nand U2542 (N_2542,N_2471,N_2467);
nor U2543 (N_2543,N_2415,N_2444);
nor U2544 (N_2544,N_2428,N_2465);
and U2545 (N_2545,N_2438,N_2459);
and U2546 (N_2546,N_2407,N_2453);
nand U2547 (N_2547,N_2428,N_2441);
and U2548 (N_2548,N_2435,N_2421);
nor U2549 (N_2549,N_2427,N_2406);
nand U2550 (N_2550,N_2542,N_2526);
and U2551 (N_2551,N_2499,N_2528);
or U2552 (N_2552,N_2508,N_2490);
or U2553 (N_2553,N_2529,N_2519);
and U2554 (N_2554,N_2532,N_2516);
and U2555 (N_2555,N_2505,N_2481);
and U2556 (N_2556,N_2483,N_2494);
nor U2557 (N_2557,N_2515,N_2502);
or U2558 (N_2558,N_2524,N_2537);
nor U2559 (N_2559,N_2535,N_2534);
nor U2560 (N_2560,N_2531,N_2491);
nand U2561 (N_2561,N_2530,N_2545);
or U2562 (N_2562,N_2547,N_2496);
nand U2563 (N_2563,N_2500,N_2512);
or U2564 (N_2564,N_2541,N_2488);
and U2565 (N_2565,N_2540,N_2489);
nor U2566 (N_2566,N_2475,N_2478);
or U2567 (N_2567,N_2523,N_2476);
xnor U2568 (N_2568,N_2484,N_2503);
nor U2569 (N_2569,N_2521,N_2527);
or U2570 (N_2570,N_2486,N_2477);
nor U2571 (N_2571,N_2513,N_2504);
nor U2572 (N_2572,N_2522,N_2479);
nor U2573 (N_2573,N_2517,N_2510);
or U2574 (N_2574,N_2487,N_2501);
xor U2575 (N_2575,N_2482,N_2525);
nor U2576 (N_2576,N_2533,N_2546);
nor U2577 (N_2577,N_2520,N_2493);
nand U2578 (N_2578,N_2536,N_2544);
nand U2579 (N_2579,N_2495,N_2543);
nand U2580 (N_2580,N_2485,N_2514);
nand U2581 (N_2581,N_2548,N_2511);
nand U2582 (N_2582,N_2506,N_2538);
xnor U2583 (N_2583,N_2480,N_2509);
and U2584 (N_2584,N_2497,N_2549);
nor U2585 (N_2585,N_2539,N_2518);
nand U2586 (N_2586,N_2492,N_2498);
and U2587 (N_2587,N_2507,N_2496);
or U2588 (N_2588,N_2480,N_2483);
and U2589 (N_2589,N_2493,N_2534);
nand U2590 (N_2590,N_2487,N_2519);
and U2591 (N_2591,N_2535,N_2514);
and U2592 (N_2592,N_2514,N_2500);
nand U2593 (N_2593,N_2520,N_2524);
nand U2594 (N_2594,N_2513,N_2520);
nor U2595 (N_2595,N_2506,N_2508);
or U2596 (N_2596,N_2498,N_2507);
or U2597 (N_2597,N_2521,N_2485);
or U2598 (N_2598,N_2490,N_2517);
nor U2599 (N_2599,N_2482,N_2541);
and U2600 (N_2600,N_2499,N_2530);
nand U2601 (N_2601,N_2482,N_2537);
and U2602 (N_2602,N_2491,N_2546);
or U2603 (N_2603,N_2513,N_2485);
and U2604 (N_2604,N_2510,N_2505);
nand U2605 (N_2605,N_2523,N_2487);
xnor U2606 (N_2606,N_2535,N_2523);
nand U2607 (N_2607,N_2508,N_2477);
nor U2608 (N_2608,N_2484,N_2521);
xor U2609 (N_2609,N_2493,N_2523);
xnor U2610 (N_2610,N_2492,N_2507);
or U2611 (N_2611,N_2538,N_2541);
nand U2612 (N_2612,N_2513,N_2549);
nor U2613 (N_2613,N_2483,N_2501);
or U2614 (N_2614,N_2499,N_2548);
or U2615 (N_2615,N_2501,N_2549);
nor U2616 (N_2616,N_2543,N_2483);
nand U2617 (N_2617,N_2546,N_2534);
nor U2618 (N_2618,N_2531,N_2523);
nand U2619 (N_2619,N_2499,N_2531);
nand U2620 (N_2620,N_2504,N_2522);
xnor U2621 (N_2621,N_2501,N_2507);
and U2622 (N_2622,N_2478,N_2515);
nor U2623 (N_2623,N_2518,N_2478);
or U2624 (N_2624,N_2476,N_2528);
or U2625 (N_2625,N_2616,N_2622);
or U2626 (N_2626,N_2569,N_2623);
nand U2627 (N_2627,N_2559,N_2568);
nand U2628 (N_2628,N_2605,N_2586);
and U2629 (N_2629,N_2593,N_2567);
or U2630 (N_2630,N_2587,N_2610);
and U2631 (N_2631,N_2582,N_2584);
and U2632 (N_2632,N_2561,N_2600);
nor U2633 (N_2633,N_2556,N_2573);
and U2634 (N_2634,N_2574,N_2617);
or U2635 (N_2635,N_2591,N_2604);
nand U2636 (N_2636,N_2560,N_2585);
nor U2637 (N_2637,N_2598,N_2583);
nor U2638 (N_2638,N_2589,N_2555);
xor U2639 (N_2639,N_2612,N_2603);
nor U2640 (N_2640,N_2613,N_2594);
xnor U2641 (N_2641,N_2565,N_2608);
and U2642 (N_2642,N_2624,N_2551);
nor U2643 (N_2643,N_2621,N_2619);
and U2644 (N_2644,N_2578,N_2557);
nand U2645 (N_2645,N_2597,N_2579);
nor U2646 (N_2646,N_2558,N_2577);
nor U2647 (N_2647,N_2602,N_2570);
xnor U2648 (N_2648,N_2580,N_2611);
and U2649 (N_2649,N_2562,N_2607);
nor U2650 (N_2650,N_2601,N_2592);
nor U2651 (N_2651,N_2571,N_2618);
or U2652 (N_2652,N_2596,N_2614);
xnor U2653 (N_2653,N_2554,N_2599);
or U2654 (N_2654,N_2595,N_2588);
nand U2655 (N_2655,N_2553,N_2615);
nor U2656 (N_2656,N_2572,N_2566);
nor U2657 (N_2657,N_2563,N_2564);
and U2658 (N_2658,N_2581,N_2609);
nand U2659 (N_2659,N_2590,N_2552);
nand U2660 (N_2660,N_2575,N_2550);
and U2661 (N_2661,N_2576,N_2620);
nor U2662 (N_2662,N_2606,N_2610);
or U2663 (N_2663,N_2565,N_2580);
and U2664 (N_2664,N_2557,N_2623);
nor U2665 (N_2665,N_2594,N_2611);
nor U2666 (N_2666,N_2615,N_2621);
nand U2667 (N_2667,N_2605,N_2614);
and U2668 (N_2668,N_2603,N_2597);
and U2669 (N_2669,N_2590,N_2562);
nor U2670 (N_2670,N_2597,N_2604);
nor U2671 (N_2671,N_2604,N_2568);
nand U2672 (N_2672,N_2608,N_2613);
or U2673 (N_2673,N_2609,N_2616);
nand U2674 (N_2674,N_2613,N_2582);
nor U2675 (N_2675,N_2576,N_2581);
or U2676 (N_2676,N_2595,N_2585);
and U2677 (N_2677,N_2580,N_2560);
nor U2678 (N_2678,N_2624,N_2596);
xnor U2679 (N_2679,N_2552,N_2563);
nor U2680 (N_2680,N_2578,N_2617);
nor U2681 (N_2681,N_2597,N_2573);
xor U2682 (N_2682,N_2601,N_2562);
nor U2683 (N_2683,N_2606,N_2583);
nand U2684 (N_2684,N_2580,N_2595);
and U2685 (N_2685,N_2623,N_2572);
and U2686 (N_2686,N_2565,N_2561);
or U2687 (N_2687,N_2552,N_2569);
xnor U2688 (N_2688,N_2563,N_2557);
nor U2689 (N_2689,N_2580,N_2608);
or U2690 (N_2690,N_2562,N_2589);
nor U2691 (N_2691,N_2570,N_2613);
xor U2692 (N_2692,N_2551,N_2594);
nand U2693 (N_2693,N_2559,N_2585);
or U2694 (N_2694,N_2598,N_2593);
or U2695 (N_2695,N_2591,N_2603);
and U2696 (N_2696,N_2602,N_2559);
nor U2697 (N_2697,N_2587,N_2588);
and U2698 (N_2698,N_2615,N_2572);
nand U2699 (N_2699,N_2579,N_2601);
or U2700 (N_2700,N_2641,N_2685);
and U2701 (N_2701,N_2686,N_2664);
nand U2702 (N_2702,N_2662,N_2693);
nand U2703 (N_2703,N_2654,N_2667);
nor U2704 (N_2704,N_2680,N_2630);
and U2705 (N_2705,N_2679,N_2647);
nand U2706 (N_2706,N_2663,N_2639);
nor U2707 (N_2707,N_2690,N_2656);
nor U2708 (N_2708,N_2666,N_2650);
or U2709 (N_2709,N_2653,N_2668);
and U2710 (N_2710,N_2687,N_2655);
nor U2711 (N_2711,N_2683,N_2644);
and U2712 (N_2712,N_2696,N_2681);
or U2713 (N_2713,N_2633,N_2670);
nand U2714 (N_2714,N_2637,N_2682);
and U2715 (N_2715,N_2645,N_2657);
or U2716 (N_2716,N_2634,N_2632);
or U2717 (N_2717,N_2676,N_2661);
or U2718 (N_2718,N_2660,N_2675);
and U2719 (N_2719,N_2671,N_2699);
and U2720 (N_2720,N_2658,N_2646);
or U2721 (N_2721,N_2649,N_2692);
and U2722 (N_2722,N_2665,N_2694);
or U2723 (N_2723,N_2628,N_2673);
xnor U2724 (N_2724,N_2652,N_2678);
and U2725 (N_2725,N_2688,N_2629);
nor U2726 (N_2726,N_2684,N_2631);
nand U2727 (N_2727,N_2627,N_2695);
nor U2728 (N_2728,N_2638,N_2651);
nor U2729 (N_2729,N_2642,N_2689);
and U2730 (N_2730,N_2669,N_2625);
nor U2731 (N_2731,N_2643,N_2698);
nand U2732 (N_2732,N_2648,N_2674);
or U2733 (N_2733,N_2635,N_2691);
or U2734 (N_2734,N_2672,N_2640);
nor U2735 (N_2735,N_2677,N_2636);
nand U2736 (N_2736,N_2659,N_2626);
or U2737 (N_2737,N_2697,N_2645);
nor U2738 (N_2738,N_2656,N_2629);
nor U2739 (N_2739,N_2687,N_2662);
nor U2740 (N_2740,N_2691,N_2656);
nor U2741 (N_2741,N_2640,N_2678);
or U2742 (N_2742,N_2630,N_2675);
nand U2743 (N_2743,N_2645,N_2681);
or U2744 (N_2744,N_2696,N_2679);
nor U2745 (N_2745,N_2658,N_2627);
or U2746 (N_2746,N_2699,N_2640);
and U2747 (N_2747,N_2689,N_2648);
or U2748 (N_2748,N_2631,N_2654);
nor U2749 (N_2749,N_2648,N_2694);
or U2750 (N_2750,N_2693,N_2687);
and U2751 (N_2751,N_2641,N_2661);
nor U2752 (N_2752,N_2668,N_2666);
nor U2753 (N_2753,N_2647,N_2689);
or U2754 (N_2754,N_2652,N_2653);
nand U2755 (N_2755,N_2657,N_2640);
nor U2756 (N_2756,N_2678,N_2644);
or U2757 (N_2757,N_2633,N_2674);
nand U2758 (N_2758,N_2657,N_2698);
and U2759 (N_2759,N_2657,N_2667);
and U2760 (N_2760,N_2680,N_2679);
or U2761 (N_2761,N_2636,N_2652);
or U2762 (N_2762,N_2632,N_2675);
and U2763 (N_2763,N_2631,N_2650);
nor U2764 (N_2764,N_2676,N_2666);
nor U2765 (N_2765,N_2675,N_2646);
and U2766 (N_2766,N_2648,N_2625);
and U2767 (N_2767,N_2665,N_2629);
nor U2768 (N_2768,N_2646,N_2689);
and U2769 (N_2769,N_2637,N_2695);
and U2770 (N_2770,N_2639,N_2678);
and U2771 (N_2771,N_2656,N_2670);
nor U2772 (N_2772,N_2641,N_2683);
or U2773 (N_2773,N_2679,N_2644);
xnor U2774 (N_2774,N_2657,N_2632);
and U2775 (N_2775,N_2716,N_2703);
and U2776 (N_2776,N_2771,N_2700);
xnor U2777 (N_2777,N_2718,N_2752);
xor U2778 (N_2778,N_2763,N_2770);
nor U2779 (N_2779,N_2740,N_2746);
xor U2780 (N_2780,N_2760,N_2721);
nor U2781 (N_2781,N_2745,N_2757);
and U2782 (N_2782,N_2733,N_2710);
nand U2783 (N_2783,N_2758,N_2762);
or U2784 (N_2784,N_2769,N_2720);
or U2785 (N_2785,N_2773,N_2730);
xor U2786 (N_2786,N_2724,N_2722);
nand U2787 (N_2787,N_2728,N_2756);
nor U2788 (N_2788,N_2737,N_2748);
nand U2789 (N_2789,N_2725,N_2706);
and U2790 (N_2790,N_2704,N_2747);
nand U2791 (N_2791,N_2755,N_2749);
nand U2792 (N_2792,N_2712,N_2738);
nand U2793 (N_2793,N_2734,N_2729);
nand U2794 (N_2794,N_2736,N_2727);
and U2795 (N_2795,N_2709,N_2715);
nand U2796 (N_2796,N_2735,N_2711);
nor U2797 (N_2797,N_2759,N_2707);
nand U2798 (N_2798,N_2753,N_2742);
nor U2799 (N_2799,N_2726,N_2732);
and U2800 (N_2800,N_2766,N_2719);
or U2801 (N_2801,N_2705,N_2713);
nand U2802 (N_2802,N_2765,N_2743);
and U2803 (N_2803,N_2741,N_2717);
and U2804 (N_2804,N_2739,N_2772);
or U2805 (N_2805,N_2714,N_2767);
nand U2806 (N_2806,N_2701,N_2764);
or U2807 (N_2807,N_2754,N_2723);
nor U2808 (N_2808,N_2731,N_2750);
or U2809 (N_2809,N_2774,N_2744);
xnor U2810 (N_2810,N_2761,N_2708);
nand U2811 (N_2811,N_2768,N_2751);
or U2812 (N_2812,N_2702,N_2748);
nor U2813 (N_2813,N_2772,N_2759);
nand U2814 (N_2814,N_2754,N_2756);
nor U2815 (N_2815,N_2716,N_2729);
and U2816 (N_2816,N_2701,N_2708);
nor U2817 (N_2817,N_2712,N_2734);
and U2818 (N_2818,N_2706,N_2772);
nor U2819 (N_2819,N_2767,N_2720);
and U2820 (N_2820,N_2720,N_2748);
and U2821 (N_2821,N_2719,N_2724);
nand U2822 (N_2822,N_2736,N_2706);
and U2823 (N_2823,N_2764,N_2763);
nand U2824 (N_2824,N_2701,N_2745);
and U2825 (N_2825,N_2745,N_2719);
nand U2826 (N_2826,N_2700,N_2742);
or U2827 (N_2827,N_2770,N_2764);
and U2828 (N_2828,N_2740,N_2763);
or U2829 (N_2829,N_2711,N_2768);
or U2830 (N_2830,N_2749,N_2724);
xnor U2831 (N_2831,N_2750,N_2756);
or U2832 (N_2832,N_2745,N_2711);
nand U2833 (N_2833,N_2709,N_2704);
nand U2834 (N_2834,N_2753,N_2723);
nand U2835 (N_2835,N_2762,N_2705);
nand U2836 (N_2836,N_2700,N_2762);
nand U2837 (N_2837,N_2709,N_2748);
nor U2838 (N_2838,N_2709,N_2753);
or U2839 (N_2839,N_2768,N_2762);
or U2840 (N_2840,N_2771,N_2741);
nand U2841 (N_2841,N_2734,N_2767);
and U2842 (N_2842,N_2730,N_2740);
nor U2843 (N_2843,N_2768,N_2747);
xor U2844 (N_2844,N_2721,N_2715);
and U2845 (N_2845,N_2702,N_2731);
xor U2846 (N_2846,N_2772,N_2716);
nor U2847 (N_2847,N_2770,N_2769);
nor U2848 (N_2848,N_2727,N_2759);
or U2849 (N_2849,N_2715,N_2767);
or U2850 (N_2850,N_2822,N_2778);
nand U2851 (N_2851,N_2834,N_2805);
or U2852 (N_2852,N_2843,N_2821);
and U2853 (N_2853,N_2798,N_2813);
or U2854 (N_2854,N_2832,N_2787);
or U2855 (N_2855,N_2783,N_2841);
nand U2856 (N_2856,N_2808,N_2817);
nand U2857 (N_2857,N_2831,N_2780);
and U2858 (N_2858,N_2802,N_2838);
nand U2859 (N_2859,N_2803,N_2825);
nor U2860 (N_2860,N_2835,N_2800);
or U2861 (N_2861,N_2788,N_2791);
nor U2862 (N_2862,N_2816,N_2796);
and U2863 (N_2863,N_2836,N_2775);
nand U2864 (N_2864,N_2777,N_2806);
nand U2865 (N_2865,N_2837,N_2776);
nand U2866 (N_2866,N_2840,N_2818);
nor U2867 (N_2867,N_2809,N_2785);
or U2868 (N_2868,N_2779,N_2799);
nand U2869 (N_2869,N_2795,N_2839);
xor U2870 (N_2870,N_2804,N_2849);
nand U2871 (N_2871,N_2827,N_2797);
xor U2872 (N_2872,N_2786,N_2793);
and U2873 (N_2873,N_2842,N_2807);
nand U2874 (N_2874,N_2790,N_2782);
and U2875 (N_2875,N_2830,N_2784);
nor U2876 (N_2876,N_2828,N_2844);
and U2877 (N_2877,N_2814,N_2819);
or U2878 (N_2878,N_2801,N_2829);
nand U2879 (N_2879,N_2789,N_2781);
and U2880 (N_2880,N_2833,N_2794);
or U2881 (N_2881,N_2847,N_2815);
or U2882 (N_2882,N_2823,N_2820);
and U2883 (N_2883,N_2845,N_2826);
xnor U2884 (N_2884,N_2824,N_2810);
nand U2885 (N_2885,N_2792,N_2812);
or U2886 (N_2886,N_2848,N_2811);
or U2887 (N_2887,N_2846,N_2779);
nand U2888 (N_2888,N_2806,N_2790);
xor U2889 (N_2889,N_2816,N_2809);
xor U2890 (N_2890,N_2813,N_2815);
and U2891 (N_2891,N_2808,N_2799);
nand U2892 (N_2892,N_2799,N_2849);
nand U2893 (N_2893,N_2823,N_2803);
or U2894 (N_2894,N_2793,N_2811);
xor U2895 (N_2895,N_2832,N_2807);
xnor U2896 (N_2896,N_2832,N_2829);
nor U2897 (N_2897,N_2816,N_2831);
xnor U2898 (N_2898,N_2831,N_2821);
and U2899 (N_2899,N_2786,N_2828);
nand U2900 (N_2900,N_2838,N_2834);
nand U2901 (N_2901,N_2845,N_2806);
or U2902 (N_2902,N_2820,N_2836);
and U2903 (N_2903,N_2799,N_2821);
nand U2904 (N_2904,N_2833,N_2822);
nand U2905 (N_2905,N_2845,N_2777);
or U2906 (N_2906,N_2795,N_2834);
nor U2907 (N_2907,N_2829,N_2778);
nor U2908 (N_2908,N_2777,N_2815);
and U2909 (N_2909,N_2832,N_2783);
nand U2910 (N_2910,N_2776,N_2819);
nand U2911 (N_2911,N_2847,N_2819);
and U2912 (N_2912,N_2788,N_2831);
nor U2913 (N_2913,N_2783,N_2844);
and U2914 (N_2914,N_2786,N_2803);
or U2915 (N_2915,N_2845,N_2808);
or U2916 (N_2916,N_2800,N_2814);
or U2917 (N_2917,N_2811,N_2802);
or U2918 (N_2918,N_2780,N_2787);
or U2919 (N_2919,N_2816,N_2810);
nand U2920 (N_2920,N_2808,N_2802);
xor U2921 (N_2921,N_2825,N_2838);
or U2922 (N_2922,N_2816,N_2782);
and U2923 (N_2923,N_2829,N_2775);
nand U2924 (N_2924,N_2787,N_2792);
or U2925 (N_2925,N_2918,N_2850);
and U2926 (N_2926,N_2862,N_2920);
nor U2927 (N_2927,N_2868,N_2855);
xor U2928 (N_2928,N_2897,N_2891);
nor U2929 (N_2929,N_2851,N_2856);
nor U2930 (N_2930,N_2860,N_2922);
and U2931 (N_2931,N_2854,N_2892);
and U2932 (N_2932,N_2905,N_2903);
nor U2933 (N_2933,N_2878,N_2881);
and U2934 (N_2934,N_2912,N_2916);
and U2935 (N_2935,N_2871,N_2877);
and U2936 (N_2936,N_2910,N_2884);
or U2937 (N_2937,N_2859,N_2882);
and U2938 (N_2938,N_2923,N_2909);
nand U2939 (N_2939,N_2901,N_2902);
xnor U2940 (N_2940,N_2924,N_2879);
and U2941 (N_2941,N_2870,N_2906);
nand U2942 (N_2942,N_2898,N_2886);
nor U2943 (N_2943,N_2904,N_2887);
nand U2944 (N_2944,N_2883,N_2895);
and U2945 (N_2945,N_2872,N_2894);
nand U2946 (N_2946,N_2911,N_2858);
xor U2947 (N_2947,N_2861,N_2893);
and U2948 (N_2948,N_2913,N_2885);
and U2949 (N_2949,N_2869,N_2899);
or U2950 (N_2950,N_2863,N_2890);
nand U2951 (N_2951,N_2874,N_2888);
and U2952 (N_2952,N_2857,N_2900);
nor U2953 (N_2953,N_2880,N_2865);
or U2954 (N_2954,N_2907,N_2875);
nor U2955 (N_2955,N_2864,N_2917);
nor U2956 (N_2956,N_2852,N_2889);
or U2957 (N_2957,N_2908,N_2914);
or U2958 (N_2958,N_2919,N_2867);
nand U2959 (N_2959,N_2853,N_2915);
nand U2960 (N_2960,N_2866,N_2873);
xnor U2961 (N_2961,N_2896,N_2921);
and U2962 (N_2962,N_2876,N_2852);
nand U2963 (N_2963,N_2919,N_2880);
and U2964 (N_2964,N_2892,N_2873);
nor U2965 (N_2965,N_2865,N_2860);
nand U2966 (N_2966,N_2888,N_2903);
nand U2967 (N_2967,N_2880,N_2924);
or U2968 (N_2968,N_2864,N_2889);
and U2969 (N_2969,N_2899,N_2856);
and U2970 (N_2970,N_2909,N_2884);
and U2971 (N_2971,N_2913,N_2908);
xor U2972 (N_2972,N_2904,N_2862);
nor U2973 (N_2973,N_2877,N_2865);
or U2974 (N_2974,N_2892,N_2922);
and U2975 (N_2975,N_2872,N_2870);
nor U2976 (N_2976,N_2866,N_2861);
nor U2977 (N_2977,N_2916,N_2876);
nand U2978 (N_2978,N_2868,N_2908);
and U2979 (N_2979,N_2908,N_2901);
or U2980 (N_2980,N_2888,N_2873);
nor U2981 (N_2981,N_2883,N_2864);
and U2982 (N_2982,N_2870,N_2873);
or U2983 (N_2983,N_2852,N_2875);
nand U2984 (N_2984,N_2880,N_2915);
or U2985 (N_2985,N_2920,N_2922);
nand U2986 (N_2986,N_2853,N_2867);
nand U2987 (N_2987,N_2866,N_2885);
nor U2988 (N_2988,N_2874,N_2865);
or U2989 (N_2989,N_2881,N_2863);
or U2990 (N_2990,N_2868,N_2876);
nand U2991 (N_2991,N_2859,N_2916);
nor U2992 (N_2992,N_2914,N_2891);
nor U2993 (N_2993,N_2854,N_2899);
nand U2994 (N_2994,N_2852,N_2891);
nor U2995 (N_2995,N_2865,N_2908);
and U2996 (N_2996,N_2909,N_2910);
nor U2997 (N_2997,N_2902,N_2862);
or U2998 (N_2998,N_2868,N_2872);
and U2999 (N_2999,N_2867,N_2875);
nor UO_0 (O_0,N_2976,N_2934);
nand UO_1 (O_1,N_2968,N_2967);
or UO_2 (O_2,N_2956,N_2944);
nor UO_3 (O_3,N_2999,N_2927);
nand UO_4 (O_4,N_2992,N_2978);
or UO_5 (O_5,N_2989,N_2955);
xnor UO_6 (O_6,N_2943,N_2986);
nor UO_7 (O_7,N_2925,N_2926);
nand UO_8 (O_8,N_2946,N_2939);
nor UO_9 (O_9,N_2952,N_2979);
nor UO_10 (O_10,N_2932,N_2940);
and UO_11 (O_11,N_2997,N_2998);
xor UO_12 (O_12,N_2958,N_2987);
nor UO_13 (O_13,N_2938,N_2991);
nand UO_14 (O_14,N_2959,N_2961);
xor UO_15 (O_15,N_2974,N_2970);
and UO_16 (O_16,N_2941,N_2953);
nand UO_17 (O_17,N_2936,N_2996);
nand UO_18 (O_18,N_2984,N_2957);
xor UO_19 (O_19,N_2972,N_2930);
or UO_20 (O_20,N_2950,N_2928);
and UO_21 (O_21,N_2990,N_2973);
or UO_22 (O_22,N_2937,N_2983);
and UO_23 (O_23,N_2980,N_2994);
or UO_24 (O_24,N_2949,N_2963);
nor UO_25 (O_25,N_2971,N_2951);
nand UO_26 (O_26,N_2962,N_2929);
or UO_27 (O_27,N_2945,N_2988);
nand UO_28 (O_28,N_2995,N_2933);
nand UO_29 (O_29,N_2982,N_2966);
xor UO_30 (O_30,N_2993,N_2969);
nor UO_31 (O_31,N_2948,N_2954);
or UO_32 (O_32,N_2947,N_2965);
nor UO_33 (O_33,N_2942,N_2960);
or UO_34 (O_34,N_2985,N_2935);
or UO_35 (O_35,N_2931,N_2977);
and UO_36 (O_36,N_2964,N_2981);
nor UO_37 (O_37,N_2975,N_2992);
or UO_38 (O_38,N_2933,N_2939);
or UO_39 (O_39,N_2942,N_2959);
and UO_40 (O_40,N_2965,N_2987);
nand UO_41 (O_41,N_2963,N_2959);
nor UO_42 (O_42,N_2996,N_2934);
and UO_43 (O_43,N_2927,N_2935);
or UO_44 (O_44,N_2973,N_2964);
and UO_45 (O_45,N_2957,N_2985);
nor UO_46 (O_46,N_2963,N_2929);
xnor UO_47 (O_47,N_2941,N_2929);
or UO_48 (O_48,N_2968,N_2944);
and UO_49 (O_49,N_2966,N_2999);
and UO_50 (O_50,N_2970,N_2933);
or UO_51 (O_51,N_2976,N_2983);
and UO_52 (O_52,N_2978,N_2926);
and UO_53 (O_53,N_2978,N_2971);
and UO_54 (O_54,N_2946,N_2947);
and UO_55 (O_55,N_2988,N_2961);
or UO_56 (O_56,N_2969,N_2965);
and UO_57 (O_57,N_2932,N_2947);
nand UO_58 (O_58,N_2948,N_2991);
nor UO_59 (O_59,N_2934,N_2978);
or UO_60 (O_60,N_2951,N_2952);
nand UO_61 (O_61,N_2986,N_2999);
nor UO_62 (O_62,N_2977,N_2972);
nor UO_63 (O_63,N_2983,N_2941);
nor UO_64 (O_64,N_2973,N_2984);
and UO_65 (O_65,N_2965,N_2943);
or UO_66 (O_66,N_2967,N_2940);
or UO_67 (O_67,N_2940,N_2925);
and UO_68 (O_68,N_2941,N_2996);
or UO_69 (O_69,N_2974,N_2943);
and UO_70 (O_70,N_2930,N_2971);
or UO_71 (O_71,N_2939,N_2930);
nand UO_72 (O_72,N_2942,N_2966);
xor UO_73 (O_73,N_2979,N_2949);
or UO_74 (O_74,N_2950,N_2968);
xor UO_75 (O_75,N_2961,N_2932);
xor UO_76 (O_76,N_2949,N_2948);
nor UO_77 (O_77,N_2957,N_2959);
or UO_78 (O_78,N_2957,N_2955);
nor UO_79 (O_79,N_2965,N_2975);
or UO_80 (O_80,N_2957,N_2999);
nand UO_81 (O_81,N_2969,N_2927);
or UO_82 (O_82,N_2939,N_2937);
and UO_83 (O_83,N_2970,N_2932);
and UO_84 (O_84,N_2957,N_2963);
nand UO_85 (O_85,N_2936,N_2979);
and UO_86 (O_86,N_2999,N_2935);
nor UO_87 (O_87,N_2939,N_2952);
or UO_88 (O_88,N_2987,N_2989);
xnor UO_89 (O_89,N_2938,N_2927);
nor UO_90 (O_90,N_2990,N_2996);
nand UO_91 (O_91,N_2994,N_2962);
nor UO_92 (O_92,N_2985,N_2955);
xor UO_93 (O_93,N_2937,N_2975);
nand UO_94 (O_94,N_2926,N_2977);
nor UO_95 (O_95,N_2976,N_2938);
nand UO_96 (O_96,N_2982,N_2976);
or UO_97 (O_97,N_2947,N_2978);
nand UO_98 (O_98,N_2960,N_2948);
and UO_99 (O_99,N_2995,N_2959);
or UO_100 (O_100,N_2925,N_2994);
and UO_101 (O_101,N_2980,N_2946);
nand UO_102 (O_102,N_2932,N_2942);
and UO_103 (O_103,N_2946,N_2953);
and UO_104 (O_104,N_2953,N_2926);
or UO_105 (O_105,N_2977,N_2970);
nand UO_106 (O_106,N_2990,N_2999);
and UO_107 (O_107,N_2955,N_2993);
or UO_108 (O_108,N_2940,N_2995);
or UO_109 (O_109,N_2993,N_2943);
nor UO_110 (O_110,N_2930,N_2986);
nor UO_111 (O_111,N_2976,N_2970);
or UO_112 (O_112,N_2937,N_2979);
nor UO_113 (O_113,N_2927,N_2954);
nand UO_114 (O_114,N_2985,N_2939);
nand UO_115 (O_115,N_2960,N_2980);
nand UO_116 (O_116,N_2986,N_2965);
and UO_117 (O_117,N_2959,N_2996);
or UO_118 (O_118,N_2928,N_2981);
and UO_119 (O_119,N_2989,N_2973);
and UO_120 (O_120,N_2978,N_2997);
or UO_121 (O_121,N_2957,N_2938);
nor UO_122 (O_122,N_2941,N_2963);
xnor UO_123 (O_123,N_2982,N_2932);
or UO_124 (O_124,N_2998,N_2965);
and UO_125 (O_125,N_2964,N_2982);
or UO_126 (O_126,N_2939,N_2948);
or UO_127 (O_127,N_2938,N_2928);
nor UO_128 (O_128,N_2953,N_2982);
or UO_129 (O_129,N_2960,N_2966);
nor UO_130 (O_130,N_2952,N_2962);
or UO_131 (O_131,N_2939,N_2961);
or UO_132 (O_132,N_2992,N_2971);
and UO_133 (O_133,N_2974,N_2993);
and UO_134 (O_134,N_2967,N_2944);
nor UO_135 (O_135,N_2956,N_2952);
and UO_136 (O_136,N_2949,N_2951);
and UO_137 (O_137,N_2930,N_2926);
xnor UO_138 (O_138,N_2973,N_2983);
and UO_139 (O_139,N_2999,N_2964);
nand UO_140 (O_140,N_2965,N_2971);
or UO_141 (O_141,N_2997,N_2968);
xnor UO_142 (O_142,N_2930,N_2993);
and UO_143 (O_143,N_2965,N_2981);
and UO_144 (O_144,N_2998,N_2979);
and UO_145 (O_145,N_2996,N_2943);
or UO_146 (O_146,N_2945,N_2974);
and UO_147 (O_147,N_2970,N_2978);
and UO_148 (O_148,N_2950,N_2957);
nand UO_149 (O_149,N_2934,N_2995);
or UO_150 (O_150,N_2984,N_2988);
or UO_151 (O_151,N_2986,N_2975);
nand UO_152 (O_152,N_2953,N_2961);
xnor UO_153 (O_153,N_2962,N_2983);
xor UO_154 (O_154,N_2944,N_2950);
nor UO_155 (O_155,N_2960,N_2964);
and UO_156 (O_156,N_2958,N_2951);
and UO_157 (O_157,N_2981,N_2946);
and UO_158 (O_158,N_2977,N_2966);
or UO_159 (O_159,N_2994,N_2996);
and UO_160 (O_160,N_2962,N_2927);
and UO_161 (O_161,N_2968,N_2977);
or UO_162 (O_162,N_2945,N_2951);
nor UO_163 (O_163,N_2955,N_2966);
xnor UO_164 (O_164,N_2941,N_2995);
nor UO_165 (O_165,N_2941,N_2977);
or UO_166 (O_166,N_2926,N_2928);
or UO_167 (O_167,N_2933,N_2993);
or UO_168 (O_168,N_2982,N_2972);
xor UO_169 (O_169,N_2928,N_2996);
xnor UO_170 (O_170,N_2968,N_2960);
xnor UO_171 (O_171,N_2927,N_2930);
nand UO_172 (O_172,N_2990,N_2991);
xor UO_173 (O_173,N_2970,N_2975);
and UO_174 (O_174,N_2942,N_2969);
nand UO_175 (O_175,N_2939,N_2984);
or UO_176 (O_176,N_2970,N_2991);
nand UO_177 (O_177,N_2961,N_2957);
nor UO_178 (O_178,N_2975,N_2978);
and UO_179 (O_179,N_2937,N_2950);
or UO_180 (O_180,N_2946,N_2937);
and UO_181 (O_181,N_2929,N_2937);
nor UO_182 (O_182,N_2952,N_2989);
or UO_183 (O_183,N_2979,N_2972);
and UO_184 (O_184,N_2978,N_2980);
or UO_185 (O_185,N_2988,N_2927);
and UO_186 (O_186,N_2936,N_2971);
xnor UO_187 (O_187,N_2976,N_2946);
or UO_188 (O_188,N_2998,N_2988);
and UO_189 (O_189,N_2984,N_2981);
or UO_190 (O_190,N_2968,N_2975);
or UO_191 (O_191,N_2962,N_2970);
nor UO_192 (O_192,N_2941,N_2933);
or UO_193 (O_193,N_2932,N_2941);
nor UO_194 (O_194,N_2999,N_2960);
nor UO_195 (O_195,N_2959,N_2977);
nand UO_196 (O_196,N_2962,N_2974);
and UO_197 (O_197,N_2990,N_2931);
or UO_198 (O_198,N_2988,N_2959);
or UO_199 (O_199,N_2962,N_2938);
nand UO_200 (O_200,N_2936,N_2937);
nand UO_201 (O_201,N_2928,N_2991);
and UO_202 (O_202,N_2969,N_2935);
xnor UO_203 (O_203,N_2950,N_2979);
nand UO_204 (O_204,N_2963,N_2960);
and UO_205 (O_205,N_2938,N_2947);
nor UO_206 (O_206,N_2983,N_2959);
nand UO_207 (O_207,N_2977,N_2971);
nor UO_208 (O_208,N_2943,N_2968);
or UO_209 (O_209,N_2967,N_2980);
and UO_210 (O_210,N_2966,N_2954);
nor UO_211 (O_211,N_2959,N_2937);
or UO_212 (O_212,N_2949,N_2968);
and UO_213 (O_213,N_2970,N_2935);
nand UO_214 (O_214,N_2981,N_2954);
and UO_215 (O_215,N_2989,N_2956);
or UO_216 (O_216,N_2977,N_2942);
nand UO_217 (O_217,N_2979,N_2953);
nor UO_218 (O_218,N_2968,N_2964);
nor UO_219 (O_219,N_2981,N_2927);
or UO_220 (O_220,N_2953,N_2956);
nor UO_221 (O_221,N_2954,N_2965);
xor UO_222 (O_222,N_2976,N_2985);
and UO_223 (O_223,N_2969,N_2939);
nor UO_224 (O_224,N_2953,N_2958);
nand UO_225 (O_225,N_2998,N_2983);
and UO_226 (O_226,N_2999,N_2985);
and UO_227 (O_227,N_2979,N_2974);
xor UO_228 (O_228,N_2975,N_2973);
nand UO_229 (O_229,N_2989,N_2977);
nand UO_230 (O_230,N_2953,N_2968);
nand UO_231 (O_231,N_2945,N_2936);
or UO_232 (O_232,N_2966,N_2958);
and UO_233 (O_233,N_2958,N_2988);
nand UO_234 (O_234,N_2975,N_2929);
xnor UO_235 (O_235,N_2985,N_2972);
and UO_236 (O_236,N_2992,N_2970);
nor UO_237 (O_237,N_2946,N_2988);
nand UO_238 (O_238,N_2928,N_2946);
nor UO_239 (O_239,N_2982,N_2960);
and UO_240 (O_240,N_2940,N_2961);
and UO_241 (O_241,N_2963,N_2978);
or UO_242 (O_242,N_2989,N_2995);
and UO_243 (O_243,N_2936,N_2932);
and UO_244 (O_244,N_2997,N_2984);
nor UO_245 (O_245,N_2984,N_2949);
xnor UO_246 (O_246,N_2966,N_2934);
nand UO_247 (O_247,N_2939,N_2940);
nor UO_248 (O_248,N_2954,N_2999);
nand UO_249 (O_249,N_2935,N_2953);
and UO_250 (O_250,N_2976,N_2979);
xor UO_251 (O_251,N_2932,N_2925);
and UO_252 (O_252,N_2984,N_2977);
or UO_253 (O_253,N_2990,N_2997);
or UO_254 (O_254,N_2925,N_2939);
and UO_255 (O_255,N_2929,N_2969);
or UO_256 (O_256,N_2932,N_2976);
and UO_257 (O_257,N_2992,N_2969);
nor UO_258 (O_258,N_2951,N_2996);
nor UO_259 (O_259,N_2967,N_2986);
or UO_260 (O_260,N_2941,N_2930);
or UO_261 (O_261,N_2956,N_2942);
and UO_262 (O_262,N_2964,N_2934);
or UO_263 (O_263,N_2937,N_2974);
nand UO_264 (O_264,N_2945,N_2930);
and UO_265 (O_265,N_2958,N_2990);
nand UO_266 (O_266,N_2956,N_2931);
and UO_267 (O_267,N_2935,N_2987);
and UO_268 (O_268,N_2930,N_2934);
nor UO_269 (O_269,N_2965,N_2976);
or UO_270 (O_270,N_2978,N_2930);
nor UO_271 (O_271,N_2925,N_2965);
nor UO_272 (O_272,N_2972,N_2980);
and UO_273 (O_273,N_2959,N_2984);
nand UO_274 (O_274,N_2953,N_2972);
nor UO_275 (O_275,N_2945,N_2969);
and UO_276 (O_276,N_2994,N_2971);
nand UO_277 (O_277,N_2933,N_2936);
nor UO_278 (O_278,N_2971,N_2991);
nor UO_279 (O_279,N_2963,N_2950);
or UO_280 (O_280,N_2990,N_2967);
and UO_281 (O_281,N_2928,N_2976);
nand UO_282 (O_282,N_2985,N_2981);
nor UO_283 (O_283,N_2935,N_2929);
and UO_284 (O_284,N_2929,N_2998);
or UO_285 (O_285,N_2938,N_2956);
and UO_286 (O_286,N_2965,N_2992);
or UO_287 (O_287,N_2974,N_2954);
and UO_288 (O_288,N_2964,N_2944);
or UO_289 (O_289,N_2935,N_2966);
nand UO_290 (O_290,N_2990,N_2947);
and UO_291 (O_291,N_2982,N_2947);
and UO_292 (O_292,N_2940,N_2992);
nand UO_293 (O_293,N_2961,N_2990);
or UO_294 (O_294,N_2999,N_2943);
nor UO_295 (O_295,N_2964,N_2984);
nand UO_296 (O_296,N_2998,N_2973);
or UO_297 (O_297,N_2971,N_2943);
nand UO_298 (O_298,N_2941,N_2957);
xnor UO_299 (O_299,N_2982,N_2989);
and UO_300 (O_300,N_2965,N_2973);
nor UO_301 (O_301,N_2976,N_2957);
and UO_302 (O_302,N_2931,N_2993);
nand UO_303 (O_303,N_2954,N_2953);
and UO_304 (O_304,N_2958,N_2984);
nand UO_305 (O_305,N_2981,N_2953);
xor UO_306 (O_306,N_2968,N_2999);
nand UO_307 (O_307,N_2984,N_2935);
xor UO_308 (O_308,N_2966,N_2980);
and UO_309 (O_309,N_2956,N_2948);
nand UO_310 (O_310,N_2966,N_2988);
nor UO_311 (O_311,N_2947,N_2949);
nand UO_312 (O_312,N_2937,N_2952);
or UO_313 (O_313,N_2936,N_2927);
or UO_314 (O_314,N_2981,N_2951);
nor UO_315 (O_315,N_2960,N_2938);
or UO_316 (O_316,N_2970,N_2988);
nor UO_317 (O_317,N_2950,N_2961);
xor UO_318 (O_318,N_2927,N_2965);
or UO_319 (O_319,N_2976,N_2969);
and UO_320 (O_320,N_2931,N_2953);
and UO_321 (O_321,N_2955,N_2945);
nand UO_322 (O_322,N_2934,N_2940);
and UO_323 (O_323,N_2972,N_2929);
nor UO_324 (O_324,N_2959,N_2947);
nand UO_325 (O_325,N_2995,N_2974);
and UO_326 (O_326,N_2991,N_2936);
nor UO_327 (O_327,N_2995,N_2954);
and UO_328 (O_328,N_2964,N_2936);
nand UO_329 (O_329,N_2966,N_2929);
nand UO_330 (O_330,N_2932,N_2984);
or UO_331 (O_331,N_2988,N_2938);
and UO_332 (O_332,N_2967,N_2930);
and UO_333 (O_333,N_2993,N_2983);
and UO_334 (O_334,N_2988,N_2963);
or UO_335 (O_335,N_2942,N_2948);
nand UO_336 (O_336,N_2949,N_2936);
or UO_337 (O_337,N_2944,N_2943);
or UO_338 (O_338,N_2960,N_2931);
or UO_339 (O_339,N_2974,N_2971);
nand UO_340 (O_340,N_2993,N_2973);
nand UO_341 (O_341,N_2941,N_2951);
nor UO_342 (O_342,N_2968,N_2962);
or UO_343 (O_343,N_2984,N_2931);
xnor UO_344 (O_344,N_2948,N_2978);
nor UO_345 (O_345,N_2932,N_2977);
or UO_346 (O_346,N_2991,N_2956);
and UO_347 (O_347,N_2929,N_2973);
nand UO_348 (O_348,N_2970,N_2969);
nand UO_349 (O_349,N_2962,N_2926);
nor UO_350 (O_350,N_2926,N_2936);
or UO_351 (O_351,N_2975,N_2999);
nand UO_352 (O_352,N_2985,N_2930);
nand UO_353 (O_353,N_2977,N_2945);
nor UO_354 (O_354,N_2976,N_2944);
and UO_355 (O_355,N_2981,N_2988);
or UO_356 (O_356,N_2945,N_2989);
nor UO_357 (O_357,N_2938,N_2974);
and UO_358 (O_358,N_2969,N_2973);
nand UO_359 (O_359,N_2934,N_2983);
and UO_360 (O_360,N_2954,N_2941);
nor UO_361 (O_361,N_2992,N_2933);
nand UO_362 (O_362,N_2929,N_2971);
or UO_363 (O_363,N_2955,N_2979);
and UO_364 (O_364,N_2933,N_2935);
nand UO_365 (O_365,N_2928,N_2977);
and UO_366 (O_366,N_2961,N_2985);
or UO_367 (O_367,N_2990,N_2984);
and UO_368 (O_368,N_2983,N_2936);
or UO_369 (O_369,N_2983,N_2988);
nand UO_370 (O_370,N_2925,N_2997);
nand UO_371 (O_371,N_2992,N_2973);
and UO_372 (O_372,N_2932,N_2987);
nand UO_373 (O_373,N_2949,N_2953);
and UO_374 (O_374,N_2976,N_2974);
and UO_375 (O_375,N_2969,N_2982);
and UO_376 (O_376,N_2993,N_2926);
xor UO_377 (O_377,N_2950,N_2969);
and UO_378 (O_378,N_2989,N_2964);
or UO_379 (O_379,N_2975,N_2925);
nand UO_380 (O_380,N_2988,N_2997);
nor UO_381 (O_381,N_2943,N_2941);
or UO_382 (O_382,N_2928,N_2984);
or UO_383 (O_383,N_2989,N_2998);
xnor UO_384 (O_384,N_2951,N_2959);
xor UO_385 (O_385,N_2966,N_2986);
xor UO_386 (O_386,N_2938,N_2961);
or UO_387 (O_387,N_2941,N_2952);
nor UO_388 (O_388,N_2989,N_2930);
nand UO_389 (O_389,N_2926,N_2967);
and UO_390 (O_390,N_2942,N_2953);
or UO_391 (O_391,N_2974,N_2981);
nor UO_392 (O_392,N_2984,N_2983);
and UO_393 (O_393,N_2958,N_2972);
nor UO_394 (O_394,N_2994,N_2981);
or UO_395 (O_395,N_2952,N_2959);
nor UO_396 (O_396,N_2964,N_2990);
nor UO_397 (O_397,N_2937,N_2942);
xnor UO_398 (O_398,N_2948,N_2979);
and UO_399 (O_399,N_2977,N_2960);
xor UO_400 (O_400,N_2938,N_2959);
nor UO_401 (O_401,N_2970,N_2938);
and UO_402 (O_402,N_2940,N_2976);
or UO_403 (O_403,N_2957,N_2971);
nor UO_404 (O_404,N_2931,N_2965);
nor UO_405 (O_405,N_2959,N_2927);
nor UO_406 (O_406,N_2952,N_2970);
or UO_407 (O_407,N_2956,N_2965);
and UO_408 (O_408,N_2970,N_2966);
or UO_409 (O_409,N_2949,N_2989);
nand UO_410 (O_410,N_2980,N_2979);
and UO_411 (O_411,N_2987,N_2994);
xor UO_412 (O_412,N_2978,N_2929);
nand UO_413 (O_413,N_2976,N_2947);
or UO_414 (O_414,N_2933,N_2975);
nand UO_415 (O_415,N_2946,N_2966);
nor UO_416 (O_416,N_2962,N_2966);
nor UO_417 (O_417,N_2971,N_2993);
nand UO_418 (O_418,N_2973,N_2966);
or UO_419 (O_419,N_2973,N_2950);
nor UO_420 (O_420,N_2957,N_2936);
nand UO_421 (O_421,N_2952,N_2931);
nor UO_422 (O_422,N_2984,N_2930);
or UO_423 (O_423,N_2954,N_2987);
xnor UO_424 (O_424,N_2955,N_2967);
nor UO_425 (O_425,N_2987,N_2982);
nor UO_426 (O_426,N_2988,N_2928);
nor UO_427 (O_427,N_2954,N_2964);
or UO_428 (O_428,N_2930,N_2931);
nor UO_429 (O_429,N_2952,N_2994);
nand UO_430 (O_430,N_2934,N_2943);
or UO_431 (O_431,N_2951,N_2975);
nand UO_432 (O_432,N_2972,N_2969);
nor UO_433 (O_433,N_2991,N_2988);
nor UO_434 (O_434,N_2937,N_2978);
nand UO_435 (O_435,N_2950,N_2985);
and UO_436 (O_436,N_2971,N_2963);
nor UO_437 (O_437,N_2957,N_2926);
nor UO_438 (O_438,N_2927,N_2977);
xnor UO_439 (O_439,N_2959,N_2935);
xnor UO_440 (O_440,N_2969,N_2926);
nor UO_441 (O_441,N_2940,N_2972);
nand UO_442 (O_442,N_2935,N_2963);
xnor UO_443 (O_443,N_2926,N_2946);
xor UO_444 (O_444,N_2981,N_2968);
or UO_445 (O_445,N_2935,N_2937);
nor UO_446 (O_446,N_2977,N_2985);
nor UO_447 (O_447,N_2947,N_2931);
or UO_448 (O_448,N_2979,N_2981);
nor UO_449 (O_449,N_2964,N_2951);
nand UO_450 (O_450,N_2957,N_2948);
or UO_451 (O_451,N_2989,N_2974);
or UO_452 (O_452,N_2994,N_2926);
nor UO_453 (O_453,N_2981,N_2996);
or UO_454 (O_454,N_2930,N_2979);
or UO_455 (O_455,N_2981,N_2947);
or UO_456 (O_456,N_2977,N_2969);
nor UO_457 (O_457,N_2971,N_2983);
nand UO_458 (O_458,N_2941,N_2988);
nand UO_459 (O_459,N_2942,N_2964);
nor UO_460 (O_460,N_2949,N_2995);
nand UO_461 (O_461,N_2975,N_2931);
or UO_462 (O_462,N_2986,N_2959);
and UO_463 (O_463,N_2938,N_2950);
nand UO_464 (O_464,N_2937,N_2934);
and UO_465 (O_465,N_2926,N_2938);
and UO_466 (O_466,N_2925,N_2963);
or UO_467 (O_467,N_2975,N_2981);
nor UO_468 (O_468,N_2966,N_2969);
or UO_469 (O_469,N_2952,N_2987);
nand UO_470 (O_470,N_2963,N_2954);
nand UO_471 (O_471,N_2976,N_2950);
xor UO_472 (O_472,N_2942,N_2984);
xor UO_473 (O_473,N_2984,N_2991);
nor UO_474 (O_474,N_2981,N_2933);
nor UO_475 (O_475,N_2994,N_2989);
nand UO_476 (O_476,N_2955,N_2943);
or UO_477 (O_477,N_2997,N_2940);
nand UO_478 (O_478,N_2993,N_2992);
nor UO_479 (O_479,N_2989,N_2970);
or UO_480 (O_480,N_2993,N_2988);
nand UO_481 (O_481,N_2989,N_2953);
xor UO_482 (O_482,N_2926,N_2960);
or UO_483 (O_483,N_2980,N_2937);
xnor UO_484 (O_484,N_2992,N_2942);
nand UO_485 (O_485,N_2925,N_2971);
and UO_486 (O_486,N_2941,N_2974);
nor UO_487 (O_487,N_2955,N_2925);
xor UO_488 (O_488,N_2947,N_2979);
nand UO_489 (O_489,N_2954,N_2983);
and UO_490 (O_490,N_2974,N_2975);
nand UO_491 (O_491,N_2979,N_2957);
and UO_492 (O_492,N_2930,N_2981);
and UO_493 (O_493,N_2962,N_2949);
nor UO_494 (O_494,N_2954,N_2957);
or UO_495 (O_495,N_2935,N_2992);
and UO_496 (O_496,N_2996,N_2958);
nand UO_497 (O_497,N_2977,N_2992);
nand UO_498 (O_498,N_2960,N_2987);
nand UO_499 (O_499,N_2938,N_2982);
endmodule