module basic_2000_20000_2500_125_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_982,In_1606);
and U1 (N_1,In_1716,In_1832);
nand U2 (N_2,In_772,In_1996);
nand U3 (N_3,In_1933,In_420);
or U4 (N_4,In_911,In_1852);
nand U5 (N_5,In_493,In_1183);
xor U6 (N_6,In_517,In_133);
or U7 (N_7,In_1835,In_1316);
nor U8 (N_8,In_264,In_1690);
nand U9 (N_9,In_1007,In_435);
nand U10 (N_10,In_963,In_959);
nand U11 (N_11,In_1838,In_243);
and U12 (N_12,In_1611,In_1805);
nor U13 (N_13,In_85,In_977);
nor U14 (N_14,In_1775,In_478);
nor U15 (N_15,In_1024,In_1772);
and U16 (N_16,In_1502,In_1720);
xnor U17 (N_17,In_1175,In_438);
nor U18 (N_18,In_162,In_849);
nand U19 (N_19,In_1081,In_715);
and U20 (N_20,In_537,In_328);
nand U21 (N_21,In_1371,In_767);
or U22 (N_22,In_1721,In_1140);
and U23 (N_23,In_411,In_121);
or U24 (N_24,In_804,In_931);
and U25 (N_25,In_1416,In_1536);
and U26 (N_26,In_757,In_1356);
or U27 (N_27,In_1119,In_1985);
and U28 (N_28,In_437,In_1913);
and U29 (N_29,In_704,In_453);
nand U30 (N_30,In_111,In_1111);
or U31 (N_31,In_1281,In_1511);
nand U32 (N_32,In_1964,In_1914);
and U33 (N_33,In_131,In_204);
nor U34 (N_34,In_236,In_32);
nand U35 (N_35,In_1857,In_1643);
or U36 (N_36,In_895,In_1849);
nand U37 (N_37,In_1987,In_1702);
nor U38 (N_38,In_166,In_433);
and U39 (N_39,In_1032,In_344);
nand U40 (N_40,In_457,In_315);
and U41 (N_41,In_1198,In_1095);
nand U42 (N_42,In_614,In_1072);
nand U43 (N_43,In_153,In_1609);
or U44 (N_44,In_762,In_638);
nand U45 (N_45,In_365,In_1724);
nand U46 (N_46,In_1163,In_285);
nand U47 (N_47,In_717,In_316);
xnor U48 (N_48,In_975,In_317);
and U49 (N_49,In_774,In_802);
or U50 (N_50,In_1623,In_1937);
and U51 (N_51,In_1197,In_515);
or U52 (N_52,In_413,In_75);
or U53 (N_53,In_36,In_1470);
and U54 (N_54,In_401,In_539);
nand U55 (N_55,In_1120,In_334);
and U56 (N_56,In_469,In_944);
xor U57 (N_57,In_1559,In_1718);
nand U58 (N_58,In_1530,In_1206);
or U59 (N_59,In_1287,In_590);
and U60 (N_60,In_641,In_1742);
or U61 (N_61,In_1886,In_1621);
and U62 (N_62,In_42,In_817);
xnor U63 (N_63,In_1615,In_1193);
nand U64 (N_64,In_314,In_323);
and U65 (N_65,In_1863,In_1649);
nor U66 (N_66,In_630,In_547);
and U67 (N_67,In_1986,In_1541);
nand U68 (N_68,In_207,In_626);
and U69 (N_69,In_218,In_228);
nand U70 (N_70,In_11,In_492);
or U71 (N_71,In_138,In_68);
nor U72 (N_72,In_1504,In_1456);
or U73 (N_73,In_978,In_1491);
and U74 (N_74,In_289,In_499);
and U75 (N_75,In_1034,In_576);
nand U76 (N_76,In_1090,In_522);
nor U77 (N_77,In_789,In_1876);
xnor U78 (N_78,In_693,In_1570);
nor U79 (N_79,In_884,In_966);
nand U80 (N_80,In_1158,In_873);
and U81 (N_81,In_368,In_920);
nor U82 (N_82,In_1188,In_1247);
nand U83 (N_83,In_1887,In_1947);
nand U84 (N_84,In_70,In_1600);
and U85 (N_85,In_617,In_991);
nand U86 (N_86,In_439,In_1226);
or U87 (N_87,In_878,In_1178);
or U88 (N_88,In_1903,In_1804);
nand U89 (N_89,In_1415,In_1629);
nor U90 (N_90,In_970,In_1267);
nand U91 (N_91,In_839,In_1757);
or U92 (N_92,In_1413,In_1001);
nor U93 (N_93,In_1513,In_600);
and U94 (N_94,In_1301,In_19);
xnor U95 (N_95,In_612,In_950);
xnor U96 (N_96,In_562,In_1483);
and U97 (N_97,In_1362,In_685);
nand U98 (N_98,In_1668,In_737);
nand U99 (N_99,In_434,In_471);
and U100 (N_100,In_18,In_1822);
and U101 (N_101,In_376,In_1783);
nor U102 (N_102,In_1377,In_245);
and U103 (N_103,In_1018,In_1970);
nand U104 (N_104,In_548,In_1101);
nand U105 (N_105,In_649,In_89);
xnor U106 (N_106,In_0,In_1142);
and U107 (N_107,In_589,In_157);
nor U108 (N_108,In_136,In_1255);
or U109 (N_109,In_1225,In_1517);
xor U110 (N_110,In_1641,In_1029);
nand U111 (N_111,In_301,In_1363);
nor U112 (N_112,In_1153,In_1758);
and U113 (N_113,In_209,In_1931);
nor U114 (N_114,In_779,In_1813);
nor U115 (N_115,In_308,In_520);
nand U116 (N_116,In_1222,In_1786);
nor U117 (N_117,In_1418,In_467);
and U118 (N_118,In_350,In_838);
nand U119 (N_119,In_1350,In_303);
and U120 (N_120,In_417,In_431);
nand U121 (N_121,In_1793,In_1239);
and U122 (N_122,In_187,In_398);
and U123 (N_123,In_21,In_197);
nor U124 (N_124,In_1484,In_874);
and U125 (N_125,In_1573,In_1434);
nor U126 (N_126,In_4,In_1242);
nor U127 (N_127,In_940,In_102);
nand U128 (N_128,In_1639,In_1501);
or U129 (N_129,In_1698,In_900);
nor U130 (N_130,In_1278,In_465);
nand U131 (N_131,In_1166,In_930);
nor U132 (N_132,In_1447,In_700);
nand U133 (N_133,In_1408,In_1023);
nor U134 (N_134,In_9,In_1700);
xnor U135 (N_135,In_1842,In_828);
nor U136 (N_136,In_1531,In_917);
and U137 (N_137,In_72,In_1323);
nand U138 (N_138,In_577,In_1869);
nor U139 (N_139,In_1781,In_1788);
nor U140 (N_140,In_430,In_844);
nor U141 (N_141,In_559,In_958);
or U142 (N_142,In_1093,In_1157);
nor U143 (N_143,In_812,In_1848);
nor U144 (N_144,In_108,In_258);
and U145 (N_145,In_645,In_634);
nor U146 (N_146,In_999,In_485);
nor U147 (N_147,In_1170,In_646);
or U148 (N_148,In_856,In_1821);
nand U149 (N_149,In_1179,In_1542);
or U150 (N_150,In_824,In_945);
nand U151 (N_151,In_1610,In_27);
or U152 (N_152,In_295,In_1921);
xnor U153 (N_153,In_882,In_833);
and U154 (N_154,In_139,In_450);
or U155 (N_155,In_1823,In_1839);
xor U156 (N_156,In_126,In_1650);
or U157 (N_157,In_575,In_905);
xor U158 (N_158,In_1192,In_1122);
and U159 (N_159,In_897,In_568);
nor U160 (N_160,In_837,In_1398);
nor U161 (N_161,In_1113,N_155);
or U162 (N_162,In_470,In_148);
xor U163 (N_163,In_1597,In_355);
xnor U164 (N_164,In_146,In_1710);
and U165 (N_165,In_1490,In_821);
nor U166 (N_166,In_1164,In_830);
nand U167 (N_167,In_428,In_1548);
nor U168 (N_168,In_1176,In_132);
xnor U169 (N_169,In_644,In_775);
or U170 (N_170,In_163,In_1711);
or U171 (N_171,In_22,In_1952);
nand U172 (N_172,In_1445,In_1291);
or U173 (N_173,In_747,In_1558);
and U174 (N_174,In_707,In_1306);
or U175 (N_175,In_1011,In_114);
or U176 (N_176,N_61,In_642);
nand U177 (N_177,In_888,N_69);
xnor U178 (N_178,In_1732,In_956);
and U179 (N_179,In_1500,In_252);
xor U180 (N_180,In_1397,In_1833);
nor U181 (N_181,N_98,In_1201);
nor U182 (N_182,In_1046,In_1677);
nand U183 (N_183,In_1207,In_848);
and U184 (N_184,In_1393,In_402);
or U185 (N_185,In_486,In_765);
nand U186 (N_186,In_1475,In_1203);
xor U187 (N_187,In_134,In_455);
nor U188 (N_188,In_117,In_683);
or U189 (N_189,In_1594,N_149);
nor U190 (N_190,In_1519,In_1954);
and U191 (N_191,N_84,In_1796);
nor U192 (N_192,In_1695,In_1489);
nor U193 (N_193,In_1187,In_1130);
and U194 (N_194,In_1395,In_1552);
or U195 (N_195,In_1686,In_1068);
nor U196 (N_196,In_968,In_521);
nor U197 (N_197,In_1866,In_342);
nor U198 (N_198,In_1993,N_36);
and U199 (N_199,In_1902,N_146);
and U200 (N_200,In_198,N_153);
nand U201 (N_201,N_156,In_863);
nor U202 (N_202,In_362,In_508);
or U203 (N_203,In_395,In_302);
xnor U204 (N_204,N_118,In_1108);
nor U205 (N_205,In_1331,N_55);
nor U206 (N_206,In_1917,In_1488);
nand U207 (N_207,N_22,In_1992);
nand U208 (N_208,In_1053,In_660);
nor U209 (N_209,In_193,In_1737);
nor U210 (N_210,In_926,In_1874);
nand U211 (N_211,In_1890,N_103);
xnor U212 (N_212,In_173,In_1208);
nand U213 (N_213,In_384,In_290);
nand U214 (N_214,In_40,N_151);
or U215 (N_215,In_1043,In_281);
or U216 (N_216,In_1134,In_1476);
nand U217 (N_217,In_1858,In_908);
and U218 (N_218,In_175,N_76);
or U219 (N_219,In_1879,In_1384);
nand U220 (N_220,In_1738,In_1925);
or U221 (N_221,In_1274,In_1870);
and U222 (N_222,In_500,N_43);
nor U223 (N_223,In_1982,In_1588);
nand U224 (N_224,In_674,In_358);
and U225 (N_225,In_17,In_976);
nor U226 (N_226,In_1437,In_1676);
or U227 (N_227,In_116,In_377);
nor U228 (N_228,In_1620,N_62);
nor U229 (N_229,In_1486,In_1082);
and U230 (N_230,In_1927,In_661);
nand U231 (N_231,In_534,N_79);
or U232 (N_232,In_957,In_813);
nor U233 (N_233,In_1628,In_1094);
nand U234 (N_234,In_1314,In_1406);
nand U235 (N_235,In_92,In_1002);
nor U236 (N_236,In_454,In_1778);
xnor U237 (N_237,In_189,In_766);
nor U238 (N_238,In_185,In_123);
or U239 (N_239,In_1799,In_1181);
and U240 (N_240,In_1139,In_1260);
xor U241 (N_241,In_29,N_135);
nand U242 (N_242,In_423,N_0);
nor U243 (N_243,In_210,In_1782);
xnor U244 (N_244,In_1774,In_1599);
or U245 (N_245,In_1078,In_1521);
nand U246 (N_246,In_654,In_1978);
or U247 (N_247,In_896,In_341);
or U248 (N_248,In_300,In_800);
and U249 (N_249,In_1613,In_591);
nor U250 (N_250,In_129,In_1825);
xnor U251 (N_251,N_68,In_601);
and U252 (N_252,In_369,In_1304);
nand U253 (N_253,In_867,In_569);
or U254 (N_254,In_753,In_987);
nand U255 (N_255,In_578,In_152);
nor U256 (N_256,In_385,In_66);
or U257 (N_257,In_1177,In_1587);
or U258 (N_258,In_296,In_1348);
nand U259 (N_259,N_38,In_8);
nand U260 (N_260,In_983,In_1310);
nor U261 (N_261,In_980,In_53);
and U262 (N_262,In_406,In_158);
and U263 (N_263,In_1693,In_1336);
or U264 (N_264,In_781,N_40);
or U265 (N_265,In_597,In_1915);
and U266 (N_266,In_793,In_327);
or U267 (N_267,In_764,In_1000);
and U268 (N_268,N_37,In_827);
and U269 (N_269,In_1659,In_1216);
nor U270 (N_270,In_893,In_690);
nor U271 (N_271,In_866,In_1726);
and U272 (N_272,In_1419,In_546);
nand U273 (N_273,N_113,In_745);
or U274 (N_274,In_1012,In_1049);
nor U275 (N_275,In_1357,In_1539);
and U276 (N_276,In_1655,N_115);
or U277 (N_277,In_217,In_443);
nand U278 (N_278,In_914,In_835);
and U279 (N_279,In_30,In_906);
nor U280 (N_280,N_58,In_1067);
nand U281 (N_281,N_64,In_480);
or U282 (N_282,In_1494,In_555);
xnor U283 (N_283,In_865,In_106);
or U284 (N_284,In_1859,In_1753);
nor U285 (N_285,In_370,In_864);
or U286 (N_286,In_1872,In_63);
and U287 (N_287,In_1037,In_1471);
and U288 (N_288,In_935,In_843);
nor U289 (N_289,In_1967,In_1878);
or U290 (N_290,In_1524,In_1147);
and U291 (N_291,In_1069,In_609);
and U292 (N_292,In_672,In_585);
nor U293 (N_293,In_1123,In_840);
or U294 (N_294,In_1185,In_259);
and U295 (N_295,N_157,In_662);
and U296 (N_296,In_99,In_697);
xor U297 (N_297,In_1202,In_1723);
or U298 (N_298,In_1219,In_1920);
xnor U299 (N_299,In_86,In_1983);
or U300 (N_300,In_1048,In_599);
xor U301 (N_301,In_422,In_1057);
nor U302 (N_302,In_1309,In_1706);
nand U303 (N_303,In_795,In_1340);
and U304 (N_304,In_319,In_1972);
or U305 (N_305,In_588,In_616);
nor U306 (N_306,In_1891,In_1318);
or U307 (N_307,In_862,In_1560);
nand U308 (N_308,In_97,In_1420);
xor U309 (N_309,In_118,In_1104);
and U310 (N_310,N_45,In_1603);
or U311 (N_311,N_112,In_13);
and U312 (N_312,In_1767,In_1237);
or U313 (N_313,In_381,In_1929);
or U314 (N_314,In_229,In_785);
or U315 (N_315,In_321,In_1771);
nand U316 (N_316,In_593,In_141);
nor U317 (N_317,In_7,In_159);
or U318 (N_318,In_1214,In_771);
nand U319 (N_319,In_540,In_1060);
nand U320 (N_320,N_41,N_292);
or U321 (N_321,In_1780,In_1598);
and U322 (N_322,In_1211,In_1151);
and U323 (N_323,In_410,In_266);
and U324 (N_324,In_1819,In_203);
nand U325 (N_325,In_1422,In_240);
and U326 (N_326,In_657,N_178);
and U327 (N_327,In_233,In_792);
nor U328 (N_328,In_379,In_104);
nor U329 (N_329,In_244,N_199);
or U330 (N_330,In_1999,N_67);
nor U331 (N_331,In_985,In_992);
or U332 (N_332,In_1212,In_1453);
and U333 (N_333,In_819,In_798);
or U334 (N_334,N_121,N_229);
nand U335 (N_335,In_1820,In_489);
and U336 (N_336,In_1436,N_106);
or U337 (N_337,In_282,In_1035);
nor U338 (N_338,In_1343,In_586);
and U339 (N_339,In_552,In_543);
nor U340 (N_340,In_1468,In_1283);
nand U341 (N_341,In_1244,In_1697);
xor U342 (N_342,In_1339,In_199);
nor U343 (N_343,In_832,N_124);
nor U344 (N_344,N_265,In_1856);
nand U345 (N_345,In_359,In_1372);
or U346 (N_346,In_1342,In_1039);
or U347 (N_347,In_34,In_1110);
or U348 (N_348,In_214,In_1617);
nor U349 (N_349,In_698,N_92);
nand U350 (N_350,In_553,In_1425);
nor U351 (N_351,In_275,In_1694);
nand U352 (N_352,N_221,N_192);
and U353 (N_353,In_998,In_1990);
nor U354 (N_354,In_1064,In_556);
nor U355 (N_355,In_405,In_1292);
nand U356 (N_356,In_1546,In_1748);
nor U357 (N_357,In_1266,In_633);
and U358 (N_358,In_399,In_326);
and U359 (N_359,In_875,In_1322);
nor U360 (N_360,In_1658,N_96);
or U361 (N_361,In_857,In_720);
and U362 (N_362,In_1829,In_424);
and U363 (N_363,In_24,In_1457);
or U364 (N_364,In_1712,In_1544);
xor U365 (N_365,N_297,N_10);
and U366 (N_366,N_308,In_834);
nand U367 (N_367,In_1146,In_1405);
nor U368 (N_368,In_1683,N_268);
nor U369 (N_369,N_80,In_1124);
nor U370 (N_370,In_909,In_1351);
nor U371 (N_371,In_98,N_189);
nor U372 (N_372,N_148,N_218);
nor U373 (N_373,In_312,In_1750);
nand U374 (N_374,In_1785,In_1708);
nand U375 (N_375,In_1557,In_1382);
xor U376 (N_376,In_1112,In_338);
xnor U377 (N_377,In_995,In_572);
and U378 (N_378,In_1515,In_1107);
or U379 (N_379,In_1847,In_474);
or U380 (N_380,In_928,In_1640);
nand U381 (N_381,In_1387,In_31);
nor U382 (N_382,N_3,N_303);
nor U383 (N_383,In_1853,In_331);
nor U384 (N_384,In_1851,In_979);
and U385 (N_385,In_790,N_227);
or U386 (N_386,In_1366,N_168);
xor U387 (N_387,In_847,In_1654);
nand U388 (N_388,In_330,In_1298);
nor U389 (N_389,In_871,In_291);
and U390 (N_390,In_692,In_807);
or U391 (N_391,N_119,In_953);
nor U392 (N_392,In_1355,In_505);
and U393 (N_393,In_347,In_581);
and U394 (N_394,In_249,In_299);
and U395 (N_395,In_1026,In_1592);
nand U396 (N_396,In_712,In_531);
or U397 (N_397,In_570,In_1186);
or U398 (N_398,In_109,In_566);
nand U399 (N_399,N_109,N_26);
nand U400 (N_400,In_115,N_269);
and U401 (N_401,In_178,In_1830);
or U402 (N_402,In_339,In_1745);
and U403 (N_403,In_447,In_1579);
nand U404 (N_404,In_990,In_1624);
nand U405 (N_405,N_32,In_740);
nor U406 (N_406,N_78,In_1252);
and U407 (N_407,In_1066,In_969);
nor U408 (N_408,In_169,In_1794);
and U409 (N_409,In_748,In_797);
nand U410 (N_410,In_1747,In_1321);
or U411 (N_411,In_1052,In_1006);
nand U412 (N_412,In_845,In_1800);
nor U413 (N_413,In_216,In_254);
or U414 (N_414,In_1901,In_655);
and U415 (N_415,In_1379,In_1651);
and U416 (N_416,In_1271,In_542);
nand U417 (N_417,In_345,In_414);
and U418 (N_418,In_733,In_1296);
or U419 (N_419,In_76,In_293);
nand U420 (N_420,In_1086,N_313);
and U421 (N_421,In_647,In_1087);
and U422 (N_422,In_1446,In_1875);
or U423 (N_423,N_202,In_726);
nor U424 (N_424,N_83,In_1604);
or U425 (N_425,In_507,In_55);
and U426 (N_426,In_67,In_1596);
or U427 (N_427,N_250,In_127);
nand U428 (N_428,N_216,In_1098);
nor U429 (N_429,In_731,In_1062);
and U430 (N_430,In_1150,In_287);
or U431 (N_431,N_31,In_1294);
or U432 (N_432,In_898,In_1670);
xor U433 (N_433,In_62,In_391);
or U434 (N_434,In_113,In_90);
xnor U435 (N_435,In_786,In_686);
and U436 (N_436,In_260,In_1257);
and U437 (N_437,N_284,In_1602);
and U438 (N_438,In_309,In_1518);
nor U439 (N_439,N_140,In_622);
or U440 (N_440,In_1254,In_238);
or U441 (N_441,In_759,In_442);
xor U442 (N_442,In_1752,In_1189);
or U443 (N_443,In_596,In_333);
nand U444 (N_444,In_892,In_140);
or U445 (N_445,N_87,In_1565);
and U446 (N_446,In_1516,In_1563);
or U447 (N_447,In_755,In_663);
nor U448 (N_448,N_27,In_1288);
xor U449 (N_449,N_104,In_1662);
nor U450 (N_450,N_196,In_1469);
nand U451 (N_451,N_253,In_964);
or U452 (N_452,In_1477,N_95);
and U453 (N_453,In_1664,In_924);
or U454 (N_454,N_274,In_1191);
xnor U455 (N_455,In_1918,In_1884);
and U456 (N_456,In_533,N_160);
and U457 (N_457,In_853,In_814);
nor U458 (N_458,In_1691,N_137);
nor U459 (N_459,In_1367,In_46);
and U460 (N_460,In_611,In_1441);
nand U461 (N_461,In_605,N_169);
or U462 (N_462,In_294,N_131);
nand U463 (N_463,In_1582,In_1289);
nor U464 (N_464,In_1850,In_1860);
or U465 (N_465,N_288,In_1689);
or U466 (N_466,In_984,In_512);
and U467 (N_467,In_364,In_497);
or U468 (N_468,N_215,In_170);
nand U469 (N_469,In_224,In_318);
and U470 (N_470,In_514,In_241);
and U471 (N_471,N_277,In_1159);
nand U472 (N_472,In_903,In_818);
and U473 (N_473,N_319,In_1899);
nand U474 (N_474,In_110,N_54);
xnor U475 (N_475,In_380,In_322);
or U476 (N_476,In_532,In_887);
and U477 (N_477,In_1459,N_211);
and U478 (N_478,N_280,In_557);
nor U479 (N_479,N_114,N_182);
nand U480 (N_480,In_571,In_1509);
nor U481 (N_481,In_1131,N_312);
or U482 (N_482,In_220,N_348);
and U483 (N_483,In_1426,N_167);
and U484 (N_484,In_580,In_1364);
xor U485 (N_485,In_1533,In_1916);
xnor U486 (N_486,In_831,N_307);
nand U487 (N_487,In_1272,N_209);
or U488 (N_488,In_1589,In_419);
or U489 (N_489,In_265,In_263);
nor U490 (N_490,In_1660,N_193);
and U491 (N_491,N_338,In_1880);
nor U492 (N_492,In_270,In_1497);
xor U493 (N_493,In_1652,N_33);
or U494 (N_494,In_768,In_702);
or U495 (N_495,In_211,N_35);
nor U496 (N_496,N_402,N_241);
nand U497 (N_497,In_1633,N_275);
and U498 (N_498,N_180,In_1485);
nor U499 (N_499,In_1836,In_750);
nand U500 (N_500,In_687,In_215);
and U501 (N_501,In_1462,In_783);
and U502 (N_502,In_610,In_526);
and U503 (N_503,In_1276,In_613);
or U504 (N_504,N_18,In_1196);
and U505 (N_505,In_752,In_1010);
and U506 (N_506,In_1831,In_1938);
and U507 (N_507,N_90,N_454);
nand U508 (N_508,In_1798,In_1969);
and U509 (N_509,In_1562,In_1148);
nand U510 (N_510,In_1246,In_524);
nor U511 (N_511,N_261,In_1647);
and U512 (N_512,N_223,In_280);
xor U513 (N_513,N_2,In_45);
xnor U514 (N_514,In_1865,In_1329);
nor U515 (N_515,In_78,N_472);
nor U516 (N_516,In_921,In_392);
or U517 (N_517,In_43,In_1270);
and U518 (N_518,In_1103,In_1873);
nand U519 (N_519,In_429,In_1409);
or U520 (N_520,In_1926,In_1138);
nand U521 (N_521,In_965,In_723);
and U522 (N_522,In_1167,In_1205);
and U523 (N_523,N_285,N_321);
nor U524 (N_524,In_1905,In_1452);
and U525 (N_525,In_151,N_368);
xor U526 (N_526,N_77,In_498);
and U527 (N_527,In_510,In_1369);
or U528 (N_528,N_289,In_1871);
or U529 (N_529,In_278,In_782);
nor U530 (N_530,In_202,In_1569);
or U531 (N_531,In_1136,In_791);
nor U532 (N_532,In_1532,In_788);
xor U533 (N_533,In_1389,In_1841);
xnor U534 (N_534,In_1097,In_876);
nand U535 (N_535,N_208,N_385);
or U536 (N_536,N_17,In_1581);
and U537 (N_537,N_374,In_912);
and U538 (N_538,In_1584,In_1190);
and U539 (N_539,N_259,In_1465);
or U540 (N_540,In_352,N_464);
or U541 (N_541,In_946,In_922);
or U542 (N_542,N_161,In_1939);
and U543 (N_543,In_1126,In_1083);
xor U544 (N_544,N_311,In_404);
xor U545 (N_545,In_1667,In_93);
and U546 (N_546,N_471,In_1338);
or U547 (N_547,N_270,In_200);
and U548 (N_548,In_1074,In_1165);
and U549 (N_549,N_49,N_24);
nor U550 (N_550,N_46,In_165);
xnor U551 (N_551,In_1955,In_1412);
nor U552 (N_552,In_1666,In_206);
xor U553 (N_553,In_221,N_478);
nand U554 (N_554,N_111,In_1807);
nor U555 (N_555,In_636,In_1358);
or U556 (N_556,In_997,N_394);
and U557 (N_557,In_383,N_107);
and U558 (N_558,In_1017,N_34);
nand U559 (N_559,N_430,In_680);
nor U560 (N_560,In_1529,In_925);
nand U561 (N_561,In_1984,In_1787);
and U562 (N_562,In_194,In_1234);
or U563 (N_563,N_150,In_1944);
nor U564 (N_564,N_134,In_394);
nor U565 (N_565,In_1472,In_1245);
or U566 (N_566,N_191,In_666);
nor U567 (N_567,In_325,In_623);
nor U568 (N_568,In_1071,In_525);
or U569 (N_569,In_1751,In_1204);
and U570 (N_570,In_1840,In_1528);
nor U571 (N_571,In_277,In_1508);
nand U572 (N_572,In_927,In_796);
and U573 (N_573,In_1240,In_869);
and U574 (N_574,In_1631,In_490);
nor U575 (N_575,In_763,In_348);
nor U576 (N_576,N_449,In_1636);
or U577 (N_577,In_1671,In_701);
and U578 (N_578,In_877,N_88);
or U579 (N_579,In_516,N_371);
nor U580 (N_580,In_232,In_879);
nand U581 (N_581,N_398,In_1812);
nor U582 (N_582,In_1324,In_1510);
nand U583 (N_583,In_799,In_967);
nor U584 (N_584,N_328,In_811);
and U585 (N_585,In_1056,N_8);
nand U586 (N_586,In_1669,N_362);
or U587 (N_587,N_228,In_122);
nand U588 (N_588,In_519,In_1924);
nor U589 (N_589,In_915,In_993);
and U590 (N_590,In_1540,In_361);
nor U591 (N_591,In_305,In_1493);
or U592 (N_592,In_23,In_1286);
xor U593 (N_593,In_464,In_179);
xnor U594 (N_594,In_615,In_1575);
nand U595 (N_595,In_149,In_972);
and U596 (N_596,In_1577,In_1160);
nor U597 (N_597,In_1118,In_770);
and U598 (N_598,In_239,N_412);
and U599 (N_599,In_637,In_51);
and U600 (N_600,In_718,In_412);
or U601 (N_601,In_1576,N_441);
nor U602 (N_602,In_1656,In_1383);
nor U603 (N_603,In_1527,In_503);
nand U604 (N_604,N_403,In_403);
nand U605 (N_605,In_445,In_271);
nor U606 (N_606,In_1549,In_1028);
or U607 (N_607,N_147,In_1009);
or U608 (N_608,In_1145,In_1834);
nand U609 (N_609,In_1963,In_955);
nor U610 (N_610,In_1019,In_656);
nand U611 (N_611,N_376,In_1551);
and U612 (N_612,In_1496,In_1744);
nand U613 (N_613,In_1727,In_1263);
and U614 (N_614,N_141,N_126);
or U615 (N_615,N_372,In_427);
nor U616 (N_616,N_375,In_1375);
nor U617 (N_617,In_1777,In_337);
and U618 (N_618,In_1249,In_986);
and U619 (N_619,N_249,In_250);
and U620 (N_620,In_1335,In_1269);
nand U621 (N_621,In_1282,In_389);
or U622 (N_622,In_1482,In_1818);
nand U623 (N_623,In_1974,In_307);
nand U624 (N_624,N_220,In_1302);
nor U625 (N_625,N_177,In_1814);
nor U626 (N_626,In_1896,In_1756);
nor U627 (N_627,In_899,N_354);
or U628 (N_628,In_171,N_226);
or U629 (N_629,In_691,N_373);
or U630 (N_630,In_709,In_387);
and U631 (N_631,N_198,In_1909);
and U632 (N_632,N_465,N_51);
and U633 (N_633,In_183,In_1535);
or U634 (N_634,In_130,In_1044);
nor U635 (N_635,In_794,In_286);
nor U636 (N_636,In_2,In_1564);
xnor U637 (N_637,In_452,N_287);
or U638 (N_638,N_105,In_137);
or U639 (N_639,In_1424,In_1014);
nand U640 (N_640,N_605,In_1431);
xor U641 (N_641,In_494,N_57);
nor U642 (N_642,In_367,N_240);
and U643 (N_643,In_628,N_639);
nand U644 (N_644,In_276,In_870);
nor U645 (N_645,N_543,N_120);
and U646 (N_646,In_1106,N_501);
nand U647 (N_647,N_625,In_95);
xor U648 (N_648,In_188,N_576);
or U649 (N_649,In_1817,N_561);
or U650 (N_650,In_1184,In_1013);
nor U651 (N_651,N_317,In_708);
nand U652 (N_652,In_1121,In_1253);
and U653 (N_653,N_266,N_526);
and U654 (N_654,In_598,N_621);
and U655 (N_655,In_1390,In_1275);
or U656 (N_656,In_746,In_1897);
or U657 (N_657,In_777,N_582);
and U658 (N_658,N_411,N_383);
nand U659 (N_659,In_803,N_230);
and U660 (N_660,N_350,N_583);
nor U661 (N_661,N_595,N_565);
and U662 (N_662,In_868,In_142);
nand U663 (N_663,In_1423,In_397);
nand U664 (N_664,In_1162,N_397);
and U665 (N_665,N_190,In_1407);
and U666 (N_666,In_386,N_222);
nor U667 (N_667,In_1657,In_1128);
and U668 (N_668,In_883,In_1473);
nand U669 (N_669,In_778,N_377);
nand U670 (N_670,In_1117,In_247);
nand U671 (N_671,In_981,In_744);
nor U672 (N_672,In_947,In_1612);
and U673 (N_673,In_1682,In_1466);
or U674 (N_674,In_201,In_147);
nand U675 (N_675,In_1864,N_163);
nand U676 (N_676,In_773,N_212);
nand U677 (N_677,In_1042,In_1699);
nor U678 (N_678,N_437,In_1687);
nand U679 (N_679,In_1451,In_1749);
and U680 (N_680,In_1618,In_509);
xnor U681 (N_681,N_518,In_1507);
nor U682 (N_682,In_850,In_1936);
or U683 (N_683,N_529,In_714);
nand U684 (N_684,N_213,N_181);
or U685 (N_685,N_562,N_300);
nand U686 (N_686,In_706,In_235);
or U687 (N_687,In_456,N_254);
nand U688 (N_688,In_1988,N_299);
or U689 (N_689,In_1313,N_560);
and U690 (N_690,In_1561,N_158);
and U691 (N_691,In_565,N_355);
nor U692 (N_692,In_400,In_1273);
or U693 (N_693,In_35,In_48);
and U694 (N_694,In_1480,In_1867);
or U695 (N_695,N_325,N_622);
nor U696 (N_696,N_499,In_479);
or U697 (N_697,In_1586,In_155);
or U698 (N_698,N_305,N_507);
and U699 (N_699,N_564,N_400);
or U700 (N_700,In_1590,In_1374);
nand U701 (N_701,N_210,In_730);
nor U702 (N_702,N_159,In_1487);
and U703 (N_703,In_451,In_1953);
nand U704 (N_704,In_1290,In_913);
and U705 (N_705,N_52,In_1900);
or U706 (N_706,N_614,In_582);
and U707 (N_707,In_33,N_255);
nor U708 (N_708,N_12,N_440);
nand U709 (N_709,In_1020,N_620);
xnor U710 (N_710,In_716,N_341);
nand U711 (N_711,N_497,In_242);
nand U712 (N_712,N_290,In_1129);
and U713 (N_713,In_1645,In_1729);
nand U714 (N_714,N_108,In_1892);
and U715 (N_715,N_532,In_1399);
xnor U716 (N_716,In_1922,In_1008);
or U717 (N_717,N_94,In_1765);
and U718 (N_718,In_1567,N_123);
nand U719 (N_719,N_585,In_39);
xnor U720 (N_720,N_366,In_225);
nor U721 (N_721,N_1,N_382);
nand U722 (N_722,In_1770,In_1844);
or U723 (N_723,N_340,In_518);
and U724 (N_724,In_1402,In_476);
nor U725 (N_725,N_601,N_50);
or U726 (N_726,N_466,In_343);
nor U727 (N_727,In_1824,In_855);
and U728 (N_728,N_429,In_1021);
nand U729 (N_729,In_1889,N_293);
or U730 (N_730,In_1262,In_1684);
and U731 (N_731,In_836,In_1404);
nand U732 (N_732,In_724,In_1946);
nand U733 (N_733,N_483,In_523);
and U734 (N_734,N_422,N_333);
and U735 (N_735,In_1241,In_1100);
or U736 (N_736,In_1680,In_619);
nor U737 (N_737,N_129,In_1503);
and U738 (N_738,N_479,In_1692);
nor U739 (N_739,In_902,In_1725);
or U740 (N_740,In_481,In_1084);
or U741 (N_741,N_396,In_1259);
and U742 (N_742,In_1846,N_579);
nor U743 (N_743,In_1601,N_42);
or U744 (N_744,In_682,In_3);
or U745 (N_745,In_805,N_474);
or U746 (N_746,In_573,In_1672);
or U747 (N_747,In_363,In_1632);
and U748 (N_748,N_263,N_152);
xor U749 (N_749,N_30,In_1717);
nor U750 (N_750,N_467,In_41);
and U751 (N_751,In_145,In_1971);
nor U752 (N_752,In_620,In_1808);
and U753 (N_753,In_1792,N_353);
xor U754 (N_754,N_633,N_179);
or U755 (N_755,In_1928,In_1619);
nand U756 (N_756,N_557,In_954);
nor U757 (N_757,N_205,N_14);
nor U758 (N_758,N_184,In_1769);
nor U759 (N_759,N_343,In_694);
xnor U760 (N_760,N_406,N_100);
and U761 (N_761,In_1210,In_1432);
or U762 (N_762,In_1096,In_1149);
nand U763 (N_763,In_324,In_784);
nor U764 (N_764,In_58,In_1498);
or U765 (N_765,In_74,In_283);
nand U766 (N_766,In_536,In_1236);
nor U767 (N_767,In_408,N_154);
nand U768 (N_768,In_1790,N_476);
nand U769 (N_769,In_1353,N_535);
and U770 (N_770,In_1810,N_283);
nor U771 (N_771,N_623,N_433);
xor U772 (N_772,In_1248,N_272);
and U773 (N_773,N_460,In_1467);
and U774 (N_774,N_435,In_670);
or U775 (N_775,In_444,In_629);
or U776 (N_776,In_538,In_710);
nor U777 (N_777,N_214,N_445);
and U778 (N_778,In_1235,In_1091);
nor U779 (N_779,N_591,In_1733);
and U780 (N_780,N_618,N_569);
xnor U781 (N_781,In_822,N_575);
xor U782 (N_782,In_1740,N_132);
or U783 (N_783,N_568,In_1888);
xnor U784 (N_784,N_473,In_1525);
or U785 (N_785,In_754,N_314);
nand U786 (N_786,N_175,In_1414);
nor U787 (N_787,In_269,N_143);
or U788 (N_788,N_502,In_1045);
and U789 (N_789,In_713,N_48);
or U790 (N_790,N_188,In_496);
and U791 (N_791,In_1311,N_248);
and U792 (N_792,In_1077,In_1116);
and U793 (N_793,In_353,In_722);
or U794 (N_794,N_401,In_1036);
and U795 (N_795,In_885,In_460);
or U796 (N_796,In_631,In_1280);
nor U797 (N_797,N_523,N_584);
nand U798 (N_798,In_69,N_25);
nor U799 (N_799,N_596,N_468);
or U800 (N_800,In_1421,In_1317);
or U801 (N_801,In_564,In_1959);
xor U802 (N_802,N_566,N_588);
nand U803 (N_803,N_799,In_181);
nor U804 (N_804,In_1538,In_1070);
and U805 (N_805,N_166,In_705);
or U806 (N_806,In_1224,In_1861);
or U807 (N_807,In_1209,In_28);
nand U808 (N_808,In_1300,In_357);
or U809 (N_809,In_1862,N_85);
and U810 (N_810,In_1977,N_237);
or U811 (N_811,N_357,N_688);
nand U812 (N_812,In_1,In_409);
and U813 (N_813,In_1688,N_630);
nor U814 (N_814,In_168,N_653);
nor U815 (N_815,N_701,N_784);
nand U816 (N_816,N_626,N_793);
xnor U817 (N_817,N_219,N_386);
nand U818 (N_818,N_603,In_124);
or U819 (N_819,In_1232,In_1881);
or U820 (N_820,In_12,N_110);
nor U821 (N_821,In_366,In_1665);
nand U822 (N_822,In_1919,N_390);
or U823 (N_823,N_480,N_344);
nand U824 (N_824,In_742,In_1661);
and U825 (N_825,N_511,In_16);
nor U826 (N_826,In_550,In_1380);
nor U827 (N_827,In_648,In_1182);
or U828 (N_828,In_1016,In_1155);
and U829 (N_829,In_939,N_475);
and U830 (N_830,N_482,In_1966);
and U831 (N_831,In_475,N_678);
or U832 (N_832,In_858,N_727);
nand U833 (N_833,N_587,In_1172);
or U834 (N_834,In_378,N_418);
nor U835 (N_835,N_556,N_231);
or U836 (N_836,In_227,N_524);
and U837 (N_837,In_787,N_29);
and U838 (N_838,In_1394,N_734);
or U839 (N_839,In_446,In_1537);
or U840 (N_840,In_196,N_365);
and U841 (N_841,N_494,In_815);
and U842 (N_842,In_1227,In_938);
nor U843 (N_843,In_83,N_144);
or U844 (N_844,In_948,N_766);
nand U845 (N_845,N_187,In_1908);
nand U846 (N_846,In_253,In_1463);
and U847 (N_847,In_973,In_304);
nand U848 (N_848,In_651,In_1761);
nor U849 (N_849,In_934,In_554);
nor U850 (N_850,In_38,In_1141);
nand U851 (N_851,In_1199,In_461);
and U852 (N_852,N_666,In_1022);
nand U853 (N_853,In_1332,N_615);
or U854 (N_854,In_1762,N_790);
xnor U855 (N_855,In_1479,In_1161);
nor U856 (N_856,In_103,In_988);
or U857 (N_857,In_1845,In_1449);
nor U858 (N_858,N_651,N_11);
nand U859 (N_859,N_707,In_989);
and U860 (N_860,In_732,In_1743);
nor U861 (N_861,In_262,In_761);
and U862 (N_862,In_268,In_37);
and U863 (N_863,In_1250,In_1040);
or U864 (N_864,In_1349,N_173);
xor U865 (N_865,In_1883,In_851);
nor U866 (N_866,In_1360,In_1004);
or U867 (N_867,N_745,In_1526);
nor U868 (N_868,In_1572,In_872);
nor U869 (N_869,In_1132,N_541);
nand U870 (N_870,In_1268,In_298);
xnor U871 (N_871,In_1058,N_760);
nand U872 (N_872,In_719,In_1352);
xor U873 (N_873,In_1685,N_703);
or U874 (N_874,In_842,N_586);
nand U875 (N_875,In_535,N_257);
nor U876 (N_876,N_747,In_184);
and U877 (N_877,In_1038,N_367);
nor U878 (N_878,In_246,N_489);
and U879 (N_879,In_703,N_643);
nand U880 (N_880,In_1637,In_1755);
or U881 (N_881,In_120,In_1580);
xor U882 (N_882,In_739,N_294);
or U883 (N_883,In_1003,In_1566);
or U884 (N_884,In_1809,In_64);
nand U885 (N_885,In_1827,In_1968);
xnor U886 (N_886,N_641,N_544);
nor U887 (N_887,N_631,In_1681);
xnor U888 (N_888,N_698,In_529);
nor U889 (N_889,N_298,N_432);
or U890 (N_890,N_540,N_525);
or U891 (N_891,In_994,N_74);
nor U892 (N_892,N_97,N_306);
nor U893 (N_893,In_852,N_722);
nor U894 (N_894,In_728,In_26);
or U895 (N_895,N_604,In_528);
or U896 (N_896,In_695,N_654);
and U897 (N_897,In_1330,N_670);
and U898 (N_898,N_642,N_347);
and U899 (N_899,In_407,N_735);
nand U900 (N_900,In_1663,N_6);
or U901 (N_901,N_81,In_743);
and U902 (N_902,N_660,In_172);
nor U903 (N_903,In_1464,N_73);
or U904 (N_904,In_1791,In_25);
nor U905 (N_905,N_530,In_910);
and U906 (N_906,N_260,In_567);
and U907 (N_907,In_1430,N_415);
nor U908 (N_908,In_1133,N_172);
and U909 (N_909,In_664,In_1385);
and U910 (N_910,N_117,In_1295);
nand U911 (N_911,In_1626,N_610);
nand U912 (N_912,In_1746,N_130);
xnor U913 (N_913,In_1243,In_1994);
and U914 (N_914,In_1444,In_231);
nor U915 (N_915,N_777,In_1368);
nand U916 (N_916,N_748,In_1705);
and U917 (N_917,N_469,In_1341);
nor U918 (N_918,N_554,N_577);
and U919 (N_919,N_322,In_841);
nor U920 (N_920,In_466,In_1030);
and U921 (N_921,In_1438,In_1031);
and U922 (N_922,In_1719,In_907);
nor U923 (N_923,N_450,N_736);
xnor U924 (N_924,N_613,N_28);
nor U925 (N_925,In_860,N_627);
or U926 (N_926,In_951,N_488);
nor U927 (N_927,N_508,In_1261);
xnor U928 (N_928,N_427,In_375);
and U929 (N_929,In_91,In_881);
and U930 (N_930,In_1795,In_371);
nor U931 (N_931,In_1076,N_318);
nand U932 (N_932,N_550,In_1450);
and U933 (N_933,In_449,In_1195);
xnor U934 (N_934,In_190,N_455);
nand U935 (N_935,In_1958,In_1174);
nor U936 (N_936,In_484,N_65);
nor U937 (N_937,In_1760,In_563);
and U938 (N_938,N_764,In_653);
nand U939 (N_939,In_107,In_1942);
or U940 (N_940,N_714,N_59);
nor U941 (N_941,N_416,In_222);
and U942 (N_942,In_595,In_1779);
nor U943 (N_943,N_379,In_1895);
nand U944 (N_944,In_150,N_717);
and U945 (N_945,In_1228,N_165);
or U946 (N_946,N_345,In_1256);
and U947 (N_947,N_99,N_19);
xor U948 (N_948,In_561,In_1910);
nor U949 (N_949,In_1811,In_176);
nor U950 (N_950,In_161,In_440);
and U951 (N_951,In_1568,In_635);
and U952 (N_952,In_1439,N_552);
nor U953 (N_953,N_531,N_4);
nor U954 (N_954,N_536,N_407);
nand U955 (N_955,N_751,In_1156);
xnor U956 (N_956,N_176,N_742);
or U957 (N_957,In_1143,N_235);
and U958 (N_958,N_710,N_506);
nor U959 (N_959,In_652,N_315);
nor U960 (N_960,In_71,N_833);
nand U961 (N_961,In_105,In_1991);
nand U962 (N_962,N_514,N_133);
and U963 (N_963,In_1033,In_665);
and U964 (N_964,N_935,In_602);
or U965 (N_965,N_534,N_324);
nor U966 (N_966,In_1221,N_186);
and U967 (N_967,In_1455,N_854);
nor U968 (N_968,In_1403,In_284);
nor U969 (N_969,N_689,N_949);
and U970 (N_970,In_6,In_1709);
nor U971 (N_971,N_239,N_923);
nand U972 (N_972,In_1797,In_1638);
or U973 (N_973,N_805,N_957);
nand U974 (N_974,In_678,N_925);
nand U975 (N_975,In_1171,In_1734);
nand U976 (N_976,N_932,N_477);
nor U977 (N_977,N_456,In_820);
or U978 (N_978,N_504,N_517);
xor U979 (N_979,N_646,In_894);
or U980 (N_980,In_587,In_941);
xnor U981 (N_981,N_856,N_725);
nand U982 (N_982,In_1950,In_1759);
and U983 (N_983,In_256,In_1642);
nand U984 (N_984,In_59,N_859);
nand U985 (N_985,N_726,In_1050);
and U986 (N_986,In_923,In_1731);
nand U987 (N_987,In_1934,N_792);
nand U988 (N_988,In_1754,N_787);
xor U989 (N_989,In_544,In_1492);
nand U990 (N_990,N_697,N_951);
nor U991 (N_991,In_1707,In_643);
nor U992 (N_992,In_658,In_167);
nor U993 (N_993,In_182,In_1411);
nand U994 (N_994,In_1981,In_1605);
nand U995 (N_995,In_1327,N_817);
nor U996 (N_996,In_1109,N_911);
or U997 (N_997,In_1386,In_10);
nand U998 (N_998,N_944,N_66);
and U999 (N_999,In_1478,N_204);
and U1000 (N_1000,In_79,N_720);
nand U1001 (N_1001,In_1635,N_264);
nor U1002 (N_1002,N_816,In_144);
nor U1003 (N_1003,N_426,N_442);
nand U1004 (N_1004,N_796,N_772);
and U1005 (N_1005,N_738,N_888);
and U1006 (N_1006,N_858,N_485);
and U1007 (N_1007,N_910,N_749);
nand U1008 (N_1008,N_895,N_548);
nand U1009 (N_1009,N_800,In_1826);
nor U1010 (N_1010,N_882,In_1776);
nor U1011 (N_1011,In_1344,N_744);
nor U1012 (N_1012,In_1556,In_1337);
nor U1013 (N_1013,In_684,N_673);
or U1014 (N_1014,In_248,In_1401);
and U1015 (N_1015,In_1630,N_723);
nor U1016 (N_1016,N_349,N_786);
nand U1017 (N_1017,N_127,In_495);
and U1018 (N_1018,In_624,In_1105);
and U1019 (N_1019,N_952,In_372);
nand U1020 (N_1020,N_644,N_574);
nor U1021 (N_1021,In_1088,N_959);
nor U1022 (N_1022,In_186,In_942);
xor U1023 (N_1023,In_1935,N_828);
nand U1024 (N_1024,In_1396,N_758);
and U1025 (N_1025,In_1715,In_1063);
nor U1026 (N_1026,In_1346,N_715);
nor U1027 (N_1027,In_1505,N_808);
nand U1028 (N_1028,N_754,In_1154);
nand U1029 (N_1029,In_1728,N_571);
or U1030 (N_1030,N_537,N_258);
or U1031 (N_1031,In_1320,In_226);
xor U1032 (N_1032,In_1410,N_706);
nand U1033 (N_1033,N_206,In_1391);
nand U1034 (N_1034,In_1223,N_15);
nand U1035 (N_1035,N_484,In_1370);
or U1036 (N_1036,N_936,In_1127);
and U1037 (N_1037,N_592,N_342);
or U1038 (N_1038,N_136,N_361);
and U1039 (N_1039,N_875,N_788);
and U1040 (N_1040,N_71,N_39);
or U1041 (N_1041,In_1893,In_1326);
and U1042 (N_1042,In_212,N_578);
or U1043 (N_1043,In_1361,N_505);
and U1044 (N_1044,In_1843,N_281);
xnor U1045 (N_1045,N_451,In_1220);
and U1046 (N_1046,In_1768,In_1877);
nand U1047 (N_1047,N_555,In_1319);
or U1048 (N_1048,N_680,N_795);
and U1049 (N_1049,N_761,In_143);
nor U1050 (N_1050,In_1354,N_813);
or U1051 (N_1051,In_297,N_252);
nor U1052 (N_1052,N_674,In_1345);
and U1053 (N_1053,In_729,In_421);
nand U1054 (N_1054,N_203,N_243);
or U1055 (N_1055,In_174,In_734);
nand U1056 (N_1056,N_515,N_337);
nand U1057 (N_1057,In_721,In_1940);
nand U1058 (N_1058,N_837,N_619);
nor U1059 (N_1059,In_1730,In_667);
nor U1060 (N_1060,N_528,N_291);
or U1061 (N_1061,In_205,In_1962);
and U1062 (N_1062,N_174,N_712);
nor U1063 (N_1063,In_1388,N_496);
nand U1064 (N_1064,In_621,In_1703);
nand U1065 (N_1065,In_627,In_971);
or U1066 (N_1066,In_511,In_195);
or U1067 (N_1067,In_306,N_826);
nand U1068 (N_1068,In_699,N_391);
nor U1069 (N_1069,In_472,N_750);
nand U1070 (N_1070,In_1102,In_329);
or U1071 (N_1071,N_329,In_1995);
nor U1072 (N_1072,In_1229,N_955);
nand U1073 (N_1073,N_693,In_219);
nor U1074 (N_1074,In_1448,In_1736);
nor U1075 (N_1075,N_247,In_1460);
or U1076 (N_1076,In_592,In_810);
and U1077 (N_1077,N_879,N_943);
nand U1078 (N_1078,N_510,In_545);
and U1079 (N_1079,N_323,N_765);
nor U1080 (N_1080,N_731,N_956);
and U1081 (N_1081,N_559,In_1957);
xnor U1082 (N_1082,In_1454,N_16);
or U1083 (N_1083,N_954,N_945);
or U1084 (N_1084,In_1679,N_53);
and U1085 (N_1085,In_1169,N_938);
xnor U1086 (N_1086,N_794,N_138);
or U1087 (N_1087,N_388,N_851);
nor U1088 (N_1088,N_599,N_863);
nand U1089 (N_1089,In_1784,N_444);
nor U1090 (N_1090,In_558,N_803);
xor U1091 (N_1091,N_847,In_625);
nand U1092 (N_1092,In_5,In_1945);
nand U1093 (N_1093,N_327,In_180);
and U1094 (N_1094,In_1144,N_807);
nand U1095 (N_1095,N_831,In_482);
or U1096 (N_1096,N_774,N_481);
and U1097 (N_1097,In_809,N_447);
and U1098 (N_1098,N_195,N_267);
and U1099 (N_1099,In_101,N_866);
xor U1100 (N_1100,N_677,N_171);
and U1101 (N_1101,In_261,N_647);
nor U1102 (N_1102,In_349,In_230);
nor U1103 (N_1103,In_164,In_1980);
or U1104 (N_1104,N_937,N_487);
nand U1105 (N_1105,N_870,N_358);
nand U1106 (N_1106,N_768,N_843);
and U1107 (N_1107,N_913,N_590);
or U1108 (N_1108,In_1627,In_360);
nand U1109 (N_1109,In_47,N_44);
and U1110 (N_1110,In_825,N_309);
and U1111 (N_1111,N_459,In_1854);
nor U1112 (N_1112,In_1458,In_96);
nor U1113 (N_1113,In_208,N_869);
xor U1114 (N_1114,N_687,In_1218);
nor U1115 (N_1115,In_506,N_23);
nor U1116 (N_1116,N_785,In_1428);
and U1117 (N_1117,N_75,In_808);
nor U1118 (N_1118,In_880,In_916);
nor U1119 (N_1119,N_145,N_370);
nand U1120 (N_1120,N_522,In_432);
nor U1121 (N_1121,In_756,N_533);
or U1122 (N_1122,N_907,N_589);
and U1123 (N_1123,In_15,N_874);
or U1124 (N_1124,N_91,In_1365);
nand U1125 (N_1125,N_122,N_116);
nor U1126 (N_1126,In_80,In_1547);
and U1127 (N_1127,N_278,N_563);
or U1128 (N_1128,N_164,N_527);
nor U1129 (N_1129,N_699,In_441);
nor U1130 (N_1130,In_1625,In_332);
and U1131 (N_1131,N_279,N_72);
nand U1132 (N_1132,In_974,N_989);
and U1133 (N_1133,N_739,In_594);
xnor U1134 (N_1134,In_639,In_1194);
and U1135 (N_1135,N_378,N_1066);
nand U1136 (N_1136,N_896,N_431);
nor U1137 (N_1137,N_802,N_832);
or U1138 (N_1138,N_775,In_861);
and U1139 (N_1139,N_351,N_183);
or U1140 (N_1140,N_704,N_873);
xnor U1141 (N_1141,N_446,N_1096);
xnor U1142 (N_1142,N_1057,In_1907);
nor U1143 (N_1143,N_381,N_1111);
nor U1144 (N_1144,N_232,In_1607);
nand U1145 (N_1145,N_1069,N_773);
and U1146 (N_1146,N_70,N_492);
nor U1147 (N_1147,In_1956,In_313);
or U1148 (N_1148,In_1646,N_887);
xor U1149 (N_1149,N_716,N_393);
nand U1150 (N_1150,N_405,N_1090);
nor U1151 (N_1151,In_459,N_1002);
or U1152 (N_1152,N_1028,In_1381);
nand U1153 (N_1153,In_1238,N_634);
nor U1154 (N_1154,N_966,N_919);
and U1155 (N_1155,N_894,N_1050);
or U1156 (N_1156,In_933,N_558);
or U1157 (N_1157,In_1442,In_780);
and U1158 (N_1158,N_356,In_1334);
xnor U1159 (N_1159,N_658,N_994);
nand U1160 (N_1160,In_1932,In_823);
xnor U1161 (N_1161,N_684,In_1816);
or U1162 (N_1162,In_1213,N_834);
nand U1163 (N_1163,N_339,N_899);
xnor U1164 (N_1164,In_1325,N_980);
or U1165 (N_1165,In_689,N_931);
or U1166 (N_1166,N_812,N_520);
or U1167 (N_1167,In_483,In_675);
or U1168 (N_1168,In_154,In_1005);
or U1169 (N_1169,In_574,N_974);
nor U1170 (N_1170,In_463,N_617);
nand U1171 (N_1171,In_673,In_1837);
nand U1172 (N_1172,N_1047,In_1674);
and U1173 (N_1173,N_7,N_410);
and U1174 (N_1174,In_749,In_390);
xnor U1175 (N_1175,In_1882,N_972);
nand U1176 (N_1176,In_81,N_753);
nor U1177 (N_1177,N_713,In_191);
and U1178 (N_1178,N_162,N_995);
or U1179 (N_1179,N_922,In_1047);
nor U1180 (N_1180,N_814,N_86);
nor U1181 (N_1181,N_927,In_1265);
or U1182 (N_1182,N_1080,N_809);
nor U1183 (N_1183,N_655,N_637);
and U1184 (N_1184,N_934,N_436);
xnor U1185 (N_1185,N_690,N_336);
nand U1186 (N_1186,In_1523,In_234);
nor U1187 (N_1187,In_1554,N_852);
and U1188 (N_1188,N_101,N_964);
xnor U1189 (N_1189,N_421,In_1735);
and U1190 (N_1190,N_609,N_1013);
nor U1191 (N_1191,N_741,N_728);
or U1192 (N_1192,In_736,In_949);
nor U1193 (N_1193,N_594,In_1522);
xor U1194 (N_1194,N_906,N_877);
nand U1195 (N_1195,N_389,In_1961);
nor U1196 (N_1196,In_1474,In_1315);
or U1197 (N_1197,In_1855,In_1701);
or U1198 (N_1198,N_878,N_822);
nor U1199 (N_1199,N_657,In_1574);
nor U1200 (N_1200,In_1073,N_256);
or U1201 (N_1201,N_649,N_1074);
and U1202 (N_1202,In_1373,N_1075);
or U1203 (N_1203,In_1054,N_908);
xor U1204 (N_1204,In_606,N_286);
or U1205 (N_1205,N_1063,In_504);
nor U1206 (N_1206,N_903,In_859);
and U1207 (N_1207,N_1046,N_352);
nand U1208 (N_1208,N_463,N_1067);
nor U1209 (N_1209,N_63,N_920);
or U1210 (N_1210,In_1284,N_233);
and U1211 (N_1211,N_705,N_917);
nand U1212 (N_1212,N_409,N_1044);
nor U1213 (N_1213,N_201,N_438);
and U1214 (N_1214,In_632,N_200);
nor U1215 (N_1215,N_770,N_5);
or U1216 (N_1216,N_1081,In_549);
and U1217 (N_1217,In_382,N_763);
nand U1218 (N_1218,In_1085,N_304);
nor U1219 (N_1219,N_985,In_54);
and U1220 (N_1220,N_271,In_758);
or U1221 (N_1221,N_663,In_320);
xnor U1222 (N_1222,N_549,N_1024);
or U1223 (N_1223,N_1003,N_1103);
nand U1224 (N_1224,In_1898,N_334);
or U1225 (N_1225,N_380,N_776);
nor U1226 (N_1226,N_1100,N_930);
nor U1227 (N_1227,N_992,N_310);
nor U1228 (N_1228,N_1018,N_302);
and U1229 (N_1229,N_572,N_640);
nand U1230 (N_1230,N_880,N_645);
nand U1231 (N_1231,In_901,N_918);
nor U1232 (N_1232,N_1079,In_502);
nor U1233 (N_1233,N_21,N_929);
nor U1234 (N_1234,N_743,N_709);
nand U1235 (N_1235,In_1997,In_806);
and U1236 (N_1236,N_1084,In_56);
and U1237 (N_1237,In_1739,In_1461);
and U1238 (N_1238,N_538,N_947);
and U1239 (N_1239,In_1713,N_789);
or U1240 (N_1240,N_1006,N_60);
or U1241 (N_1241,In_1230,N_940);
or U1242 (N_1242,N_846,N_1020);
and U1243 (N_1243,In_1534,N_1027);
and U1244 (N_1244,N_733,In_458);
and U1245 (N_1245,In_1333,In_1279);
nor U1246 (N_1246,N_1012,N_282);
or U1247 (N_1247,N_901,N_982);
or U1248 (N_1248,In_1949,N_1026);
or U1249 (N_1249,In_829,N_976);
nor U1250 (N_1250,N_909,N_681);
and U1251 (N_1251,N_1043,In_1704);
nor U1252 (N_1252,In_65,In_1722);
nand U1253 (N_1253,N_667,In_1079);
and U1254 (N_1254,N_1015,N_971);
nor U1255 (N_1255,N_636,In_640);
nand U1256 (N_1256,N_824,N_1061);
or U1257 (N_1257,N_841,In_82);
or U1258 (N_1258,N_276,In_192);
and U1259 (N_1259,N_1098,N_1091);
and U1260 (N_1260,N_915,In_527);
and U1261 (N_1261,N_185,In_584);
and U1262 (N_1262,N_1059,N_652);
nor U1263 (N_1263,In_1555,N_1110);
and U1264 (N_1264,N_914,In_311);
nand U1265 (N_1265,In_1998,N_360);
nor U1266 (N_1266,In_679,In_1975);
xnor U1267 (N_1267,In_1293,N_509);
and U1268 (N_1268,N_1105,In_1960);
or U1269 (N_1269,In_125,N_197);
and U1270 (N_1270,N_1102,N_251);
or U1271 (N_1271,In_1648,N_926);
nor U1272 (N_1272,In_1059,N_928);
and U1273 (N_1273,N_1113,N_1001);
xor U1274 (N_1274,In_889,In_890);
and U1275 (N_1275,N_990,N_897);
nand U1276 (N_1276,In_1815,In_1766);
nand U1277 (N_1277,In_335,In_1545);
nand U1278 (N_1278,In_257,In_351);
xnor U1279 (N_1279,In_1550,N_1094);
xor U1280 (N_1280,N_1266,N_387);
nand U1281 (N_1281,N_933,N_1171);
or U1282 (N_1282,In_1973,N_580);
nand U1283 (N_1283,In_50,N_1041);
or U1284 (N_1284,N_892,N_984);
nor U1285 (N_1285,N_791,In_1025);
nor U1286 (N_1286,N_93,N_1154);
nor U1287 (N_1287,N_1141,N_612);
nor U1288 (N_1288,N_978,N_486);
and U1289 (N_1289,N_898,In_274);
or U1290 (N_1290,N_194,N_1125);
and U1291 (N_1291,In_801,N_1172);
and U1292 (N_1292,N_1180,N_332);
and U1293 (N_1293,N_1274,In_100);
or U1294 (N_1294,N_1149,N_1209);
nand U1295 (N_1295,N_1119,N_711);
and U1296 (N_1296,N_1232,N_845);
and U1297 (N_1297,N_835,N_836);
nor U1298 (N_1298,N_1186,N_662);
and U1299 (N_1299,N_865,N_207);
or U1300 (N_1300,In_1951,N_273);
or U1301 (N_1301,N_1261,In_738);
nand U1302 (N_1302,N_810,N_1144);
xnor U1303 (N_1303,In_1233,In_1520);
nor U1304 (N_1304,In_1135,N_820);
and U1305 (N_1305,N_384,N_665);
and U1306 (N_1306,N_363,N_1129);
and U1307 (N_1307,N_1014,N_1056);
or U1308 (N_1308,In_488,N_1210);
or U1309 (N_1309,N_1181,N_392);
xor U1310 (N_1310,N_448,In_1499);
nand U1311 (N_1311,N_885,In_1115);
and U1312 (N_1312,N_47,In_1125);
nand U1313 (N_1313,In_272,In_448);
and U1314 (N_1314,N_1121,N_884);
nand U1315 (N_1315,N_238,In_77);
nor U1316 (N_1316,In_1585,N_1055);
or U1317 (N_1317,In_1427,N_399);
or U1318 (N_1318,N_1189,In_1543);
and U1319 (N_1319,N_246,N_1243);
or U1320 (N_1320,In_1696,N_551);
nand U1321 (N_1321,N_692,In_583);
nand U1322 (N_1322,In_1114,N_1065);
nor U1323 (N_1323,In_943,N_490);
nor U1324 (N_1324,N_1218,N_498);
or U1325 (N_1325,In_1417,N_960);
or U1326 (N_1326,N_125,N_1138);
or U1327 (N_1327,In_84,N_1163);
or U1328 (N_1328,In_1392,N_1086);
xnor U1329 (N_1329,N_82,N_1022);
nand U1330 (N_1330,In_1215,N_262);
nand U1331 (N_1331,In_932,In_60);
nor U1332 (N_1332,N_1053,N_916);
nor U1333 (N_1333,N_675,In_846);
nand U1334 (N_1334,N_1007,In_1675);
nor U1335 (N_1335,N_628,In_49);
nand U1336 (N_1336,N_861,N_519);
nor U1337 (N_1337,In_1789,N_1245);
nor U1338 (N_1338,N_1216,In_462);
or U1339 (N_1339,N_724,N_1145);
nand U1340 (N_1340,In_1378,In_1578);
xnor U1341 (N_1341,N_900,In_1763);
nand U1342 (N_1342,N_844,N_1253);
nor U1343 (N_1343,N_702,N_1165);
and U1344 (N_1344,N_1252,N_1068);
nand U1345 (N_1345,N_1264,N_1040);
nand U1346 (N_1346,N_1244,In_671);
nor U1347 (N_1347,N_616,N_1267);
nor U1348 (N_1348,N_778,In_1264);
and U1349 (N_1349,N_1011,N_848);
nor U1350 (N_1350,N_924,In_1152);
or U1351 (N_1351,N_1156,In_88);
or U1352 (N_1352,N_1249,N_912);
nand U1353 (N_1353,N_1064,In_1678);
nand U1354 (N_1354,N_1124,N_503);
nand U1355 (N_1355,N_691,N_602);
and U1356 (N_1356,In_769,In_340);
or U1357 (N_1357,N_849,N_1197);
xor U1358 (N_1358,N_864,N_783);
or U1359 (N_1359,In_1041,In_87);
and U1360 (N_1360,N_1221,N_570);
nor U1361 (N_1361,N_1045,N_977);
or U1362 (N_1362,N_521,N_798);
and U1363 (N_1363,N_1048,N_1260);
nor U1364 (N_1364,N_853,N_404);
nor U1365 (N_1365,N_1153,N_452);
and U1366 (N_1366,In_213,N_56);
or U1367 (N_1367,N_825,N_632);
or U1368 (N_1368,N_1269,In_1092);
nor U1369 (N_1369,N_815,N_694);
and U1370 (N_1370,In_1764,In_886);
nor U1371 (N_1371,In_854,In_1911);
and U1372 (N_1372,In_1806,N_811);
and U1373 (N_1373,N_1220,N_1025);
and U1374 (N_1374,N_1195,N_823);
nor U1375 (N_1375,N_1060,N_890);
nand U1376 (N_1376,In_604,N_1147);
or U1377 (N_1377,N_1214,N_970);
nor U1378 (N_1378,N_326,N_1211);
and U1379 (N_1379,N_1175,N_779);
nand U1380 (N_1380,N_1095,N_9);
and U1381 (N_1381,N_759,N_1134);
nor U1382 (N_1382,N_1193,N_1250);
and U1383 (N_1383,In_1299,N_1148);
xnor U1384 (N_1384,N_1265,N_567);
nand U1385 (N_1385,N_1092,N_650);
xnor U1386 (N_1386,N_1161,N_1035);
nand U1387 (N_1387,N_1179,N_1031);
nor U1388 (N_1388,N_1234,In_20);
xnor U1389 (N_1389,N_320,In_659);
nor U1390 (N_1390,N_413,N_419);
or U1391 (N_1391,N_245,N_1029);
xor U1392 (N_1392,N_1030,In_579);
nand U1393 (N_1393,N_965,In_1089);
xor U1394 (N_1394,N_661,N_1054);
nand U1395 (N_1395,N_729,N_629);
and U1396 (N_1396,N_967,N_757);
and U1397 (N_1397,N_671,In_418);
and U1398 (N_1398,N_1206,N_1176);
xor U1399 (N_1399,N_1240,N_719);
and U1400 (N_1400,N_461,N_905);
xor U1401 (N_1401,N_1268,N_1089);
nand U1402 (N_1402,N_1192,N_1164);
or U1403 (N_1403,N_553,N_335);
nor U1404 (N_1404,N_1017,N_1231);
or U1405 (N_1405,N_242,In_1277);
or U1406 (N_1406,N_762,In_468);
and U1407 (N_1407,In_1653,N_581);
xor U1408 (N_1408,N_1213,N_1135);
nor U1409 (N_1409,N_999,N_1005);
and U1410 (N_1410,N_1202,N_423);
and U1411 (N_1411,N_1076,N_839);
and U1412 (N_1412,N_1257,N_1248);
or U1413 (N_1413,N_1010,N_1137);
nor U1414 (N_1414,N_996,N_986);
nand U1415 (N_1415,N_491,In_1297);
or U1416 (N_1416,N_128,N_1070);
or U1417 (N_1417,N_1215,N_648);
or U1418 (N_1418,In_267,N_600);
nand U1419 (N_1419,N_797,N_983);
nor U1420 (N_1420,N_963,In_251);
and U1421 (N_1421,In_1923,N_1049);
and U1422 (N_1422,In_952,N_225);
or U1423 (N_1423,N_1198,N_1132);
nor U1424 (N_1424,N_1205,N_1093);
xor U1425 (N_1425,In_223,In_826);
and U1426 (N_1426,N_838,N_740);
nor U1427 (N_1427,N_1109,In_1894);
nor U1428 (N_1428,N_434,N_668);
nand U1429 (N_1429,N_1118,N_1225);
nor U1430 (N_1430,N_1151,N_346);
or U1431 (N_1431,In_1773,N_1016);
nor U1432 (N_1432,N_1127,In_776);
and U1433 (N_1433,In_1514,In_1885);
nand U1434 (N_1434,In_681,In_741);
nand U1435 (N_1435,N_767,In_1948);
and U1436 (N_1436,N_1062,N_547);
and U1437 (N_1437,In_1979,N_1019);
and U1438 (N_1438,N_598,N_608);
and U1439 (N_1439,In_1741,In_551);
and U1440 (N_1440,N_1276,N_1254);
nor U1441 (N_1441,In_725,In_1941);
nand U1442 (N_1442,In_61,N_1273);
nand U1443 (N_1443,N_1332,N_1411);
nand U1444 (N_1444,N_1255,N_1229);
and U1445 (N_1445,N_1037,N_1396);
and U1446 (N_1446,In_373,N_883);
and U1447 (N_1447,N_1152,In_1904);
nand U1448 (N_1448,In_1622,N_1190);
and U1449 (N_1449,In_1065,N_1344);
nand U1450 (N_1450,N_862,In_1359);
and U1451 (N_1451,N_1359,N_827);
or U1452 (N_1452,In_288,In_1673);
xnor U1453 (N_1453,N_1427,N_1364);
nand U1454 (N_1454,N_1130,In_1303);
nand U1455 (N_1455,In_560,N_801);
or U1456 (N_1456,N_1373,N_142);
or U1457 (N_1457,N_102,N_939);
and U1458 (N_1458,N_1328,N_804);
and U1459 (N_1459,In_1217,In_177);
or U1460 (N_1460,In_1440,In_960);
nor U1461 (N_1461,N_1389,N_1296);
nor U1462 (N_1462,N_752,N_1348);
and U1463 (N_1463,N_1227,N_1042);
xor U1464 (N_1464,N_1302,In_996);
or U1465 (N_1465,N_546,N_1128);
and U1466 (N_1466,In_1828,N_1428);
and U1467 (N_1467,N_941,N_1307);
nor U1468 (N_1468,N_993,In_1495);
or U1469 (N_1469,N_1375,N_1319);
or U1470 (N_1470,N_1365,N_1325);
xnor U1471 (N_1471,N_539,N_1291);
xor U1472 (N_1472,N_1160,N_1204);
nand U1473 (N_1473,N_1287,In_1376);
and U1474 (N_1474,N_1350,N_1351);
nor U1475 (N_1475,N_683,N_1330);
nor U1476 (N_1476,N_676,N_948);
and U1477 (N_1477,N_170,N_953);
or U1478 (N_1478,N_470,N_316);
or U1479 (N_1479,N_1278,N_462);
nor U1480 (N_1480,N_1309,N_1342);
xnor U1481 (N_1481,N_1208,N_593);
and U1482 (N_1482,N_369,N_1136);
nor U1483 (N_1483,N_821,In_354);
nand U1484 (N_1484,N_1406,N_359);
and U1485 (N_1485,In_14,In_918);
nand U1486 (N_1486,N_458,N_1073);
xor U1487 (N_1487,N_1106,In_1312);
nand U1488 (N_1488,N_1349,N_1432);
or U1489 (N_1489,N_1275,N_1413);
nor U1490 (N_1490,In_1168,In_1347);
and U1491 (N_1491,N_1104,In_603);
nor U1492 (N_1492,N_139,N_857);
and U1493 (N_1493,N_1420,N_1140);
nand U1494 (N_1494,N_1353,N_1292);
nor U1495 (N_1495,N_958,N_1391);
nand U1496 (N_1496,N_1230,N_516);
nand U1497 (N_1497,N_1417,N_1334);
nor U1498 (N_1498,N_1023,In_1200);
nand U1499 (N_1499,N_904,In_1634);
nor U1500 (N_1500,N_1158,N_1116);
nor U1501 (N_1501,N_1223,N_1314);
and U1502 (N_1502,In_426,N_780);
nand U1503 (N_1503,In_937,N_573);
and U1504 (N_1504,In_57,N_607);
xnor U1505 (N_1505,N_1117,N_1036);
or U1506 (N_1506,N_1199,N_1366);
and U1507 (N_1507,N_1434,In_487);
nor U1508 (N_1508,In_1591,N_1228);
nor U1509 (N_1509,N_1439,In_751);
and U1510 (N_1510,N_1078,N_1184);
or U1511 (N_1511,N_1357,N_1277);
nand U1512 (N_1512,N_1303,In_1258);
and U1513 (N_1513,N_942,N_746);
nand U1514 (N_1514,N_1239,In_1868);
nand U1515 (N_1515,N_1360,In_135);
nand U1516 (N_1516,In_1173,In_711);
nor U1517 (N_1517,In_513,N_1320);
nor U1518 (N_1518,N_1323,In_160);
nand U1519 (N_1519,N_1281,N_1279);
or U1520 (N_1520,N_1377,N_1183);
or U1521 (N_1521,N_1347,N_1107);
nor U1522 (N_1522,N_1301,In_1801);
xnor U1523 (N_1523,N_1177,In_1595);
nor U1524 (N_1524,N_950,N_439);
nand U1525 (N_1525,N_217,In_1435);
or U1526 (N_1526,N_1139,N_1341);
and U1527 (N_1527,N_417,In_1015);
nand U1528 (N_1528,In_1583,In_1506);
xnor U1529 (N_1529,N_1423,N_756);
nor U1530 (N_1530,In_650,N_1072);
or U1531 (N_1531,N_1311,N_1437);
or U1532 (N_1532,N_1399,N_998);
nor U1533 (N_1533,N_1408,N_1306);
nor U1534 (N_1534,N_975,N_1237);
nor U1535 (N_1535,N_1431,N_829);
or U1536 (N_1536,N_1162,In_1075);
and U1537 (N_1537,N_1238,N_20);
and U1538 (N_1538,N_1415,In_388);
nor U1539 (N_1539,N_1304,N_443);
nor U1540 (N_1540,N_414,In_279);
nand U1541 (N_1541,N_1159,N_493);
nor U1542 (N_1542,N_1372,N_1414);
and U1543 (N_1543,N_886,N_1187);
nand U1544 (N_1544,N_1133,N_1430);
xnor U1545 (N_1545,N_1122,N_1368);
and U1546 (N_1546,N_1433,N_295);
nand U1547 (N_1547,N_1339,N_1370);
nand U1548 (N_1548,N_696,N_1283);
nor U1549 (N_1549,N_1416,N_1395);
nor U1550 (N_1550,N_1295,N_781);
or U1551 (N_1551,N_682,N_868);
and U1552 (N_1552,N_973,N_1108);
or U1553 (N_1553,N_1087,N_1188);
or U1554 (N_1554,N_1410,N_1400);
and U1555 (N_1555,In_1051,N_819);
nor U1556 (N_1556,N_695,N_638);
nand U1557 (N_1557,N_1009,N_1101);
xor U1558 (N_1558,In_112,N_1272);
or U1559 (N_1559,In_816,N_1308);
or U1560 (N_1560,N_1298,N_1352);
nor U1561 (N_1561,N_1219,N_1185);
nor U1562 (N_1562,N_1371,N_1297);
nor U1563 (N_1563,In_1481,N_1426);
nor U1564 (N_1564,N_301,N_1358);
or U1565 (N_1565,N_224,In_1714);
nor U1566 (N_1566,N_686,N_1321);
and U1567 (N_1567,N_1422,N_1051);
or U1568 (N_1568,N_1436,N_1355);
and U1569 (N_1569,In_1061,N_1157);
nand U1570 (N_1570,N_876,In_425);
or U1571 (N_1571,In_1965,N_1246);
nor U1572 (N_1572,N_1097,In_255);
nor U1573 (N_1573,In_607,N_1284);
nor U1574 (N_1574,N_331,N_1285);
or U1575 (N_1575,N_1217,N_453);
or U1576 (N_1576,In_668,In_501);
and U1577 (N_1577,N_1082,In_1803);
or U1578 (N_1578,N_1385,N_1182);
or U1579 (N_1579,N_700,N_1242);
and U1580 (N_1580,N_1174,N_1343);
nand U1581 (N_1581,N_730,N_1404);
or U1582 (N_1582,N_1305,N_1392);
nand U1583 (N_1583,N_1315,N_1407);
nor U1584 (N_1584,In_760,N_1169);
nand U1585 (N_1585,N_234,In_1027);
xnor U1586 (N_1586,N_755,N_1376);
or U1587 (N_1587,In_688,N_597);
nor U1588 (N_1588,N_1280,N_1077);
and U1589 (N_1589,N_871,N_718);
or U1590 (N_1590,N_1438,N_1114);
nand U1591 (N_1591,N_330,N_1387);
xor U1592 (N_1592,N_988,N_1126);
or U1593 (N_1593,N_1258,N_1324);
and U1594 (N_1594,N_1329,N_1052);
nor U1595 (N_1595,N_1004,N_1289);
or U1596 (N_1596,In_929,N_1259);
xor U1597 (N_1597,N_420,In_396);
nand U1598 (N_1598,N_1099,N_1008);
nand U1599 (N_1599,N_1032,N_881);
or U1600 (N_1600,N_1492,N_1535);
and U1601 (N_1601,N_1544,In_237);
xnor U1602 (N_1602,N_1568,N_1585);
or U1603 (N_1603,N_1386,N_1313);
nor U1604 (N_1604,N_1299,N_842);
nand U1605 (N_1605,N_1450,N_1142);
xor U1606 (N_1606,N_1083,N_1596);
nor U1607 (N_1607,In_415,In_1285);
nand U1608 (N_1608,N_1226,N_1482);
nor U1609 (N_1609,N_840,In_436);
or U1610 (N_1610,N_89,N_1576);
or U1611 (N_1611,N_424,N_1191);
and U1612 (N_1612,N_495,N_1300);
or U1613 (N_1613,N_1572,N_1233);
and U1614 (N_1614,N_1405,N_1346);
and U1615 (N_1615,N_1469,N_1516);
nor U1616 (N_1616,N_1333,N_1501);
nor U1617 (N_1617,N_1345,N_1200);
xor U1618 (N_1618,In_919,N_1262);
nor U1619 (N_1619,N_1123,In_1308);
and U1620 (N_1620,N_1316,N_1598);
nand U1621 (N_1621,N_1574,N_1379);
or U1622 (N_1622,In_530,N_1336);
nand U1623 (N_1623,N_1021,N_1578);
and U1624 (N_1624,N_1514,N_1488);
or U1625 (N_1625,N_1588,N_1456);
and U1626 (N_1626,N_408,N_721);
or U1627 (N_1627,In_676,In_1400);
nand U1628 (N_1628,N_1463,In_310);
xor U1629 (N_1629,N_818,In_73);
and U1630 (N_1630,N_1458,N_1593);
and U1631 (N_1631,N_850,N_1378);
nand U1632 (N_1632,N_1337,N_1455);
or U1633 (N_1633,N_1533,N_1486);
nor U1634 (N_1634,N_997,In_119);
nor U1635 (N_1635,N_1338,N_1527);
and U1636 (N_1636,N_1468,In_1976);
and U1637 (N_1637,N_1120,N_1497);
nor U1638 (N_1638,N_606,N_769);
and U1639 (N_1639,N_1471,N_1442);
and U1640 (N_1640,N_1380,N_1537);
or U1641 (N_1641,N_893,N_1548);
and U1642 (N_1642,N_545,N_867);
xnor U1643 (N_1643,N_1584,N_782);
or U1644 (N_1644,N_1440,In_677);
nand U1645 (N_1645,N_611,In_961);
and U1646 (N_1646,N_991,N_1494);
or U1647 (N_1647,In_1930,N_1581);
nor U1648 (N_1648,N_1058,In_1180);
and U1649 (N_1649,N_1312,In_1099);
nand U1650 (N_1650,In_1137,In_94);
nor U1651 (N_1651,N_1470,N_1212);
nor U1652 (N_1652,N_1327,N_962);
or U1653 (N_1653,N_1173,N_679);
nor U1654 (N_1654,N_1224,N_891);
or U1655 (N_1655,In_128,N_1491);
xnor U1656 (N_1656,N_1201,N_1393);
or U1657 (N_1657,N_1167,In_1608);
and U1658 (N_1658,In_1305,N_1429);
xnor U1659 (N_1659,N_1143,N_1503);
nor U1660 (N_1660,N_1331,N_656);
xnor U1661 (N_1661,N_1088,N_1477);
xor U1662 (N_1662,N_624,N_1508);
or U1663 (N_1663,In_1906,N_1445);
nor U1664 (N_1664,N_1554,N_1384);
and U1665 (N_1665,In_273,In_541);
nor U1666 (N_1666,N_981,N_1466);
and U1667 (N_1667,N_1131,N_1170);
and U1668 (N_1668,N_1443,N_1461);
xnor U1669 (N_1669,N_1525,In_1802);
nand U1670 (N_1670,In_1443,N_1462);
and U1671 (N_1671,N_1447,N_1326);
or U1672 (N_1672,N_1479,N_1480);
or U1673 (N_1673,N_708,N_1565);
nand U1674 (N_1674,N_1115,N_1564);
nand U1675 (N_1675,N_500,N_1577);
nand U1676 (N_1676,N_1452,In_44);
or U1677 (N_1677,In_1912,N_1178);
nand U1678 (N_1678,N_1039,N_1381);
nand U1679 (N_1679,In_1644,N_1536);
nand U1680 (N_1680,In_962,N_1340);
and U1681 (N_1681,N_1506,N_1496);
nand U1682 (N_1682,N_512,In_1429);
or U1683 (N_1683,N_1522,N_1474);
nor U1684 (N_1684,N_1459,N_1546);
nor U1685 (N_1685,N_1529,N_1421);
nand U1686 (N_1686,N_1476,N_1561);
and U1687 (N_1687,N_1322,N_1369);
or U1688 (N_1688,In_669,N_987);
or U1689 (N_1689,N_1481,N_1435);
xor U1690 (N_1690,N_1361,N_1263);
xor U1691 (N_1691,N_1580,N_1553);
or U1692 (N_1692,N_1388,In_727);
nor U1693 (N_1693,N_1518,N_969);
xnor U1694 (N_1694,N_664,N_1085);
or U1695 (N_1695,N_1545,N_1256);
nor U1696 (N_1696,N_244,N_860);
nor U1697 (N_1697,N_1586,N_1394);
nor U1698 (N_1698,In_477,N_1532);
or U1699 (N_1699,N_1567,N_672);
and U1700 (N_1700,N_1454,N_1499);
and U1701 (N_1701,N_1196,N_1583);
and U1702 (N_1702,N_1446,N_457);
or U1703 (N_1703,N_1318,N_1402);
nor U1704 (N_1704,N_1540,N_1150);
nor U1705 (N_1705,N_1505,N_1478);
nand U1706 (N_1706,N_425,N_1517);
xor U1707 (N_1707,N_946,N_1472);
nor U1708 (N_1708,N_1597,N_1409);
nand U1709 (N_1709,In_346,N_1509);
nor U1710 (N_1710,N_236,N_979);
or U1711 (N_1711,N_1484,In_1055);
and U1712 (N_1712,N_296,N_1549);
nor U1713 (N_1713,N_889,N_1485);
nor U1714 (N_1714,In_1080,N_1551);
or U1715 (N_1715,N_1552,In_1593);
and U1716 (N_1716,N_1566,N_685);
nand U1717 (N_1717,N_1523,In_1614);
or U1718 (N_1718,N_1362,N_1556);
nand U1719 (N_1719,In_1553,N_1579);
xor U1720 (N_1720,In_1231,N_1390);
and U1721 (N_1721,In_356,N_1569);
xnor U1722 (N_1722,In_696,N_1573);
nor U1723 (N_1723,N_1530,N_1487);
xnor U1724 (N_1724,N_1591,N_1425);
nand U1725 (N_1725,N_1403,N_1534);
and U1726 (N_1726,In_374,N_1207);
or U1727 (N_1727,N_1475,N_1542);
and U1728 (N_1728,N_1335,N_1465);
and U1729 (N_1729,N_1511,N_1033);
or U1730 (N_1730,N_1570,N_1441);
nor U1731 (N_1731,N_1571,In_156);
and U1732 (N_1732,N_1034,N_1449);
xor U1733 (N_1733,N_732,N_1367);
or U1734 (N_1734,N_921,In_1616);
and U1735 (N_1735,N_1550,N_1317);
xnor U1736 (N_1736,In_1433,N_1236);
nor U1737 (N_1737,N_1398,N_1356);
or U1738 (N_1738,N_1166,N_1270);
or U1739 (N_1739,In_891,N_513);
nor U1740 (N_1740,N_1293,N_1557);
xor U1741 (N_1741,In_1989,N_855);
nand U1742 (N_1742,In_336,N_1524);
and U1743 (N_1743,N_1521,N_1194);
xnor U1744 (N_1744,N_1587,N_1203);
nor U1745 (N_1745,N_1397,N_1541);
nor U1746 (N_1746,N_635,N_771);
nor U1747 (N_1747,In_1512,N_1288);
or U1748 (N_1748,N_1271,N_830);
or U1749 (N_1749,N_1513,N_1495);
and U1750 (N_1750,N_1555,N_1363);
nand U1751 (N_1751,N_1473,N_1000);
nor U1752 (N_1752,N_1168,In_1251);
or U1753 (N_1753,N_1560,N_395);
nor U1754 (N_1754,N_1594,N_1507);
or U1755 (N_1755,N_1247,N_1515);
or U1756 (N_1756,N_1448,N_1595);
or U1757 (N_1757,N_1592,N_1382);
nor U1758 (N_1758,N_1222,N_806);
xnor U1759 (N_1759,N_1582,N_13);
and U1760 (N_1760,N_1604,N_1653);
or U1761 (N_1761,N_1662,N_1636);
and U1762 (N_1762,N_1654,N_1562);
and U1763 (N_1763,N_1631,N_1661);
and U1764 (N_1764,N_1759,N_1746);
nand U1765 (N_1765,N_1698,N_1722);
nand U1766 (N_1766,N_1689,N_1672);
nor U1767 (N_1767,N_961,N_669);
nor U1768 (N_1768,N_1688,N_1690);
and U1769 (N_1769,N_1629,In_608);
nand U1770 (N_1770,N_1374,N_1756);
or U1771 (N_1771,N_1643,N_1575);
and U1772 (N_1772,N_1614,N_659);
and U1773 (N_1773,N_1493,N_1589);
nor U1774 (N_1774,N_1618,N_1613);
nor U1775 (N_1775,N_1251,N_1282);
nand U1776 (N_1776,N_1630,N_1711);
nand U1777 (N_1777,N_1504,N_1687);
or U1778 (N_1778,N_1729,N_1723);
nor U1779 (N_1779,N_1616,N_1676);
nand U1780 (N_1780,N_1502,N_1747);
xnor U1781 (N_1781,N_1650,N_1451);
and U1782 (N_1782,In_904,N_1453);
nand U1783 (N_1783,N_1743,N_1651);
xor U1784 (N_1784,N_1692,N_1641);
nand U1785 (N_1785,N_1728,N_1725);
or U1786 (N_1786,N_1235,N_1685);
xnor U1787 (N_1787,In_1328,N_1647);
nor U1788 (N_1788,N_428,N_1640);
or U1789 (N_1789,N_1623,N_1701);
nor U1790 (N_1790,N_542,N_968);
or U1791 (N_1791,N_1538,N_1599);
or U1792 (N_1792,N_1286,In_491);
nor U1793 (N_1793,N_1620,N_1691);
and U1794 (N_1794,N_1412,N_1483);
nor U1795 (N_1795,N_1038,N_1707);
xnor U1796 (N_1796,N_1658,N_1700);
nor U1797 (N_1797,N_1294,N_1727);
or U1798 (N_1798,N_1730,N_1609);
and U1799 (N_1799,N_1611,N_1600);
nand U1800 (N_1800,N_1753,N_1750);
nand U1801 (N_1801,N_1622,N_1667);
xor U1802 (N_1802,N_1705,N_1693);
nand U1803 (N_1803,N_1617,N_1602);
nand U1804 (N_1804,N_1719,N_1558);
or U1805 (N_1805,N_1696,N_1563);
and U1806 (N_1806,N_1526,N_1637);
and U1807 (N_1807,N_1539,N_1758);
nand U1808 (N_1808,N_1752,N_1713);
xnor U1809 (N_1809,N_1659,N_1714);
and U1810 (N_1810,N_1755,N_1754);
and U1811 (N_1811,N_1290,N_1241);
and U1812 (N_1812,N_1632,N_1737);
nor U1813 (N_1813,N_1657,In_52);
or U1814 (N_1814,N_1642,N_1627);
xor U1815 (N_1815,N_1146,N_1424);
nand U1816 (N_1816,N_1419,N_1697);
nor U1817 (N_1817,In_292,N_1740);
xor U1818 (N_1818,N_1528,N_1634);
and U1819 (N_1819,N_1715,N_1071);
nand U1820 (N_1820,N_1619,N_1669);
or U1821 (N_1821,N_1678,N_1628);
nand U1822 (N_1822,N_1490,N_1738);
nor U1823 (N_1823,N_1652,N_1418);
nand U1824 (N_1824,N_1656,N_1649);
and U1825 (N_1825,N_1663,N_1666);
nor U1826 (N_1826,N_1734,N_1610);
or U1827 (N_1827,N_1735,N_1626);
nand U1828 (N_1828,N_1703,N_1531);
nor U1829 (N_1829,N_1720,N_1721);
xnor U1830 (N_1830,N_1621,N_1668);
nand U1831 (N_1831,N_1559,N_1547);
nor U1832 (N_1832,N_1489,N_1670);
or U1833 (N_1833,N_1708,In_416);
or U1834 (N_1834,N_1683,N_1702);
nor U1835 (N_1835,N_1675,In_1943);
nand U1836 (N_1836,N_1681,N_1660);
nand U1837 (N_1837,N_1615,N_1682);
nand U1838 (N_1838,N_1709,In_735);
and U1839 (N_1839,N_1638,N_1710);
nand U1840 (N_1840,N_1695,N_1716);
or U1841 (N_1841,N_1590,N_1457);
and U1842 (N_1842,N_1686,N_1633);
or U1843 (N_1843,N_1444,N_364);
nor U1844 (N_1844,N_1665,N_1510);
or U1845 (N_1845,N_1704,N_1724);
and U1846 (N_1846,N_1603,N_1625);
nor U1847 (N_1847,N_1748,N_1742);
or U1848 (N_1848,N_1354,N_1112);
xor U1849 (N_1849,N_1673,N_1717);
nand U1850 (N_1850,N_1757,N_1645);
and U1851 (N_1851,N_1731,In_1571);
nor U1852 (N_1852,N_1155,In_1307);
and U1853 (N_1853,N_1601,N_872);
nor U1854 (N_1854,N_1644,N_1684);
nor U1855 (N_1855,N_1745,N_1607);
nor U1856 (N_1856,N_1718,N_1677);
nor U1857 (N_1857,N_1460,N_1543);
and U1858 (N_1858,In_936,N_1612);
nand U1859 (N_1859,N_1467,N_1706);
or U1860 (N_1860,N_1680,N_1606);
nor U1861 (N_1861,In_393,N_1608);
and U1862 (N_1862,In_618,N_1664);
nand U1863 (N_1863,N_1726,N_1741);
and U1864 (N_1864,N_1733,N_1310);
or U1865 (N_1865,N_1635,N_1464);
and U1866 (N_1866,N_1519,N_1744);
nor U1867 (N_1867,N_1500,In_473);
nand U1868 (N_1868,N_1512,N_1498);
nor U1869 (N_1869,N_1749,N_1679);
nand U1870 (N_1870,N_1732,N_1383);
or U1871 (N_1871,N_1694,N_737);
nor U1872 (N_1872,N_902,N_1736);
and U1873 (N_1873,N_1624,N_1712);
and U1874 (N_1874,N_1648,N_1520);
and U1875 (N_1875,N_1401,N_1699);
or U1876 (N_1876,N_1655,N_1639);
nand U1877 (N_1877,N_1646,N_1605);
and U1878 (N_1878,N_1751,N_1739);
nand U1879 (N_1879,N_1671,N_1674);
and U1880 (N_1880,In_618,N_1623);
and U1881 (N_1881,N_1282,N_1607);
nand U1882 (N_1882,N_1732,N_1733);
nor U1883 (N_1883,N_1453,N_1631);
or U1884 (N_1884,N_1563,N_1241);
or U1885 (N_1885,N_1653,N_1710);
and U1886 (N_1886,N_1660,N_1617);
nor U1887 (N_1887,N_1615,N_1681);
nor U1888 (N_1888,N_902,N_1467);
and U1889 (N_1889,N_1647,N_1620);
xor U1890 (N_1890,N_1749,N_1724);
and U1891 (N_1891,N_1752,N_1707);
nor U1892 (N_1892,N_1647,In_52);
xnor U1893 (N_1893,N_1500,N_1686);
nor U1894 (N_1894,N_1658,N_1736);
or U1895 (N_1895,N_1653,In_416);
and U1896 (N_1896,N_1294,N_1412);
nor U1897 (N_1897,N_872,N_1667);
and U1898 (N_1898,N_1743,N_1735);
and U1899 (N_1899,N_1644,N_1647);
and U1900 (N_1900,N_1698,In_608);
and U1901 (N_1901,N_1667,N_1662);
or U1902 (N_1902,N_1235,N_1626);
nand U1903 (N_1903,N_1628,N_1633);
nand U1904 (N_1904,N_1729,N_1603);
xor U1905 (N_1905,N_1617,In_936);
nand U1906 (N_1906,N_1684,N_1673);
or U1907 (N_1907,N_737,N_1728);
nor U1908 (N_1908,N_1611,N_1748);
nor U1909 (N_1909,N_1526,N_1666);
nor U1910 (N_1910,N_1616,N_1383);
and U1911 (N_1911,N_1457,N_1539);
nand U1912 (N_1912,In_904,N_1624);
and U1913 (N_1913,N_1717,N_1676);
nor U1914 (N_1914,N_1710,N_1632);
and U1915 (N_1915,N_1493,N_1614);
nor U1916 (N_1916,N_1669,N_1724);
nand U1917 (N_1917,N_1751,N_1490);
and U1918 (N_1918,N_1520,N_1726);
nor U1919 (N_1919,N_1698,N_1716);
or U1920 (N_1920,N_1862,N_1870);
and U1921 (N_1921,N_1802,N_1864);
nor U1922 (N_1922,N_1835,N_1914);
and U1923 (N_1923,N_1800,N_1825);
and U1924 (N_1924,N_1878,N_1805);
nor U1925 (N_1925,N_1777,N_1771);
or U1926 (N_1926,N_1868,N_1902);
nand U1927 (N_1927,N_1837,N_1772);
and U1928 (N_1928,N_1827,N_1764);
or U1929 (N_1929,N_1904,N_1819);
nor U1930 (N_1930,N_1816,N_1801);
and U1931 (N_1931,N_1849,N_1797);
nand U1932 (N_1932,N_1910,N_1790);
nand U1933 (N_1933,N_1883,N_1915);
nand U1934 (N_1934,N_1907,N_1793);
nand U1935 (N_1935,N_1832,N_1887);
and U1936 (N_1936,N_1774,N_1873);
xnor U1937 (N_1937,N_1833,N_1893);
xor U1938 (N_1938,N_1905,N_1789);
nand U1939 (N_1939,N_1831,N_1810);
or U1940 (N_1940,N_1840,N_1820);
or U1941 (N_1941,N_1913,N_1898);
nor U1942 (N_1942,N_1881,N_1906);
nand U1943 (N_1943,N_1763,N_1779);
and U1944 (N_1944,N_1776,N_1806);
and U1945 (N_1945,N_1808,N_1916);
nand U1946 (N_1946,N_1788,N_1885);
and U1947 (N_1947,N_1894,N_1791);
and U1948 (N_1948,N_1886,N_1795);
or U1949 (N_1949,N_1850,N_1858);
nor U1950 (N_1950,N_1855,N_1880);
nor U1951 (N_1951,N_1857,N_1804);
and U1952 (N_1952,N_1859,N_1863);
or U1953 (N_1953,N_1854,N_1796);
nand U1954 (N_1954,N_1828,N_1872);
nor U1955 (N_1955,N_1908,N_1818);
or U1956 (N_1956,N_1856,N_1861);
and U1957 (N_1957,N_1794,N_1778);
or U1958 (N_1958,N_1853,N_1845);
and U1959 (N_1959,N_1900,N_1811);
nand U1960 (N_1960,N_1775,N_1839);
or U1961 (N_1961,N_1798,N_1918);
and U1962 (N_1962,N_1890,N_1836);
or U1963 (N_1963,N_1892,N_1899);
xor U1964 (N_1964,N_1879,N_1760);
and U1965 (N_1965,N_1768,N_1851);
or U1966 (N_1966,N_1889,N_1787);
nand U1967 (N_1967,N_1912,N_1766);
nand U1968 (N_1968,N_1792,N_1903);
nand U1969 (N_1969,N_1875,N_1829);
nor U1970 (N_1970,N_1844,N_1848);
and U1971 (N_1971,N_1767,N_1869);
or U1972 (N_1972,N_1895,N_1891);
and U1973 (N_1973,N_1838,N_1799);
and U1974 (N_1974,N_1784,N_1762);
xnor U1975 (N_1975,N_1877,N_1901);
xnor U1976 (N_1976,N_1782,N_1765);
or U1977 (N_1977,N_1841,N_1817);
nand U1978 (N_1978,N_1824,N_1847);
or U1979 (N_1979,N_1761,N_1871);
and U1980 (N_1980,N_1812,N_1919);
nor U1981 (N_1981,N_1781,N_1846);
or U1982 (N_1982,N_1843,N_1897);
and U1983 (N_1983,N_1867,N_1842);
nand U1984 (N_1984,N_1896,N_1865);
nor U1985 (N_1985,N_1780,N_1884);
and U1986 (N_1986,N_1770,N_1783);
nor U1987 (N_1987,N_1814,N_1882);
nor U1988 (N_1988,N_1822,N_1911);
and U1989 (N_1989,N_1786,N_1909);
nor U1990 (N_1990,N_1866,N_1803);
nor U1991 (N_1991,N_1834,N_1773);
nand U1992 (N_1992,N_1874,N_1821);
nor U1993 (N_1993,N_1917,N_1807);
nor U1994 (N_1994,N_1815,N_1826);
nand U1995 (N_1995,N_1888,N_1860);
nor U1996 (N_1996,N_1813,N_1809);
or U1997 (N_1997,N_1876,N_1823);
and U1998 (N_1998,N_1852,N_1785);
or U1999 (N_1999,N_1769,N_1830);
nor U2000 (N_2000,N_1834,N_1792);
and U2001 (N_2001,N_1806,N_1801);
and U2002 (N_2002,N_1845,N_1842);
and U2003 (N_2003,N_1803,N_1766);
or U2004 (N_2004,N_1802,N_1818);
nand U2005 (N_2005,N_1847,N_1879);
nor U2006 (N_2006,N_1774,N_1814);
nand U2007 (N_2007,N_1891,N_1903);
nor U2008 (N_2008,N_1784,N_1825);
nor U2009 (N_2009,N_1825,N_1846);
nor U2010 (N_2010,N_1828,N_1844);
or U2011 (N_2011,N_1915,N_1893);
and U2012 (N_2012,N_1905,N_1781);
nand U2013 (N_2013,N_1845,N_1779);
or U2014 (N_2014,N_1821,N_1790);
or U2015 (N_2015,N_1782,N_1914);
and U2016 (N_2016,N_1761,N_1860);
xor U2017 (N_2017,N_1862,N_1841);
nor U2018 (N_2018,N_1815,N_1834);
nor U2019 (N_2019,N_1830,N_1833);
and U2020 (N_2020,N_1854,N_1762);
nor U2021 (N_2021,N_1905,N_1783);
nand U2022 (N_2022,N_1798,N_1842);
or U2023 (N_2023,N_1903,N_1854);
or U2024 (N_2024,N_1851,N_1862);
and U2025 (N_2025,N_1791,N_1875);
nor U2026 (N_2026,N_1814,N_1825);
and U2027 (N_2027,N_1837,N_1907);
and U2028 (N_2028,N_1763,N_1894);
and U2029 (N_2029,N_1913,N_1832);
and U2030 (N_2030,N_1813,N_1908);
and U2031 (N_2031,N_1905,N_1851);
or U2032 (N_2032,N_1788,N_1882);
nor U2033 (N_2033,N_1795,N_1893);
xor U2034 (N_2034,N_1796,N_1833);
or U2035 (N_2035,N_1874,N_1849);
nor U2036 (N_2036,N_1901,N_1832);
xor U2037 (N_2037,N_1821,N_1863);
or U2038 (N_2038,N_1830,N_1907);
and U2039 (N_2039,N_1778,N_1834);
and U2040 (N_2040,N_1882,N_1851);
xnor U2041 (N_2041,N_1867,N_1781);
and U2042 (N_2042,N_1768,N_1778);
nand U2043 (N_2043,N_1885,N_1778);
nor U2044 (N_2044,N_1828,N_1864);
and U2045 (N_2045,N_1849,N_1900);
and U2046 (N_2046,N_1871,N_1815);
or U2047 (N_2047,N_1786,N_1783);
nor U2048 (N_2048,N_1840,N_1876);
xnor U2049 (N_2049,N_1857,N_1917);
and U2050 (N_2050,N_1869,N_1788);
or U2051 (N_2051,N_1900,N_1763);
nor U2052 (N_2052,N_1882,N_1846);
and U2053 (N_2053,N_1899,N_1830);
nand U2054 (N_2054,N_1860,N_1842);
or U2055 (N_2055,N_1821,N_1889);
and U2056 (N_2056,N_1838,N_1829);
nand U2057 (N_2057,N_1843,N_1833);
and U2058 (N_2058,N_1777,N_1897);
nor U2059 (N_2059,N_1808,N_1809);
and U2060 (N_2060,N_1896,N_1776);
nand U2061 (N_2061,N_1895,N_1793);
nor U2062 (N_2062,N_1795,N_1798);
or U2063 (N_2063,N_1760,N_1829);
and U2064 (N_2064,N_1873,N_1763);
and U2065 (N_2065,N_1908,N_1857);
and U2066 (N_2066,N_1898,N_1804);
or U2067 (N_2067,N_1913,N_1874);
nor U2068 (N_2068,N_1902,N_1882);
nor U2069 (N_2069,N_1882,N_1792);
and U2070 (N_2070,N_1879,N_1792);
or U2071 (N_2071,N_1812,N_1872);
and U2072 (N_2072,N_1798,N_1814);
and U2073 (N_2073,N_1918,N_1807);
or U2074 (N_2074,N_1912,N_1896);
nand U2075 (N_2075,N_1826,N_1879);
or U2076 (N_2076,N_1780,N_1864);
nor U2077 (N_2077,N_1818,N_1851);
or U2078 (N_2078,N_1813,N_1808);
or U2079 (N_2079,N_1831,N_1827);
and U2080 (N_2080,N_1933,N_1994);
nand U2081 (N_2081,N_1993,N_1990);
or U2082 (N_2082,N_1948,N_1980);
nand U2083 (N_2083,N_2029,N_2070);
or U2084 (N_2084,N_2005,N_1930);
nor U2085 (N_2085,N_1972,N_1949);
nor U2086 (N_2086,N_1969,N_2009);
nand U2087 (N_2087,N_1952,N_1977);
nand U2088 (N_2088,N_2022,N_2078);
nor U2089 (N_2089,N_1934,N_1976);
xor U2090 (N_2090,N_1921,N_2025);
and U2091 (N_2091,N_2054,N_2055);
or U2092 (N_2092,N_1957,N_2047);
nand U2093 (N_2093,N_2019,N_2057);
nand U2094 (N_2094,N_1932,N_1959);
xnor U2095 (N_2095,N_2033,N_1936);
and U2096 (N_2096,N_1923,N_1926);
nand U2097 (N_2097,N_1996,N_2059);
or U2098 (N_2098,N_2043,N_1940);
nand U2099 (N_2099,N_1991,N_2063);
nor U2100 (N_2100,N_1985,N_1965);
nor U2101 (N_2101,N_1924,N_1978);
xnor U2102 (N_2102,N_1928,N_2026);
xnor U2103 (N_2103,N_1925,N_1951);
or U2104 (N_2104,N_1955,N_2064);
and U2105 (N_2105,N_2069,N_2011);
xnor U2106 (N_2106,N_1938,N_2040);
or U2107 (N_2107,N_1979,N_2030);
nor U2108 (N_2108,N_2032,N_2062);
or U2109 (N_2109,N_2001,N_2035);
nor U2110 (N_2110,N_1997,N_2060);
and U2111 (N_2111,N_2034,N_1966);
or U2112 (N_2112,N_2044,N_2020);
nand U2113 (N_2113,N_1931,N_1929);
nand U2114 (N_2114,N_1981,N_2016);
nand U2115 (N_2115,N_1992,N_1974);
nand U2116 (N_2116,N_1935,N_2000);
nand U2117 (N_2117,N_1941,N_2008);
nand U2118 (N_2118,N_1958,N_1964);
nand U2119 (N_2119,N_2021,N_2066);
nand U2120 (N_2120,N_2028,N_2015);
or U2121 (N_2121,N_2071,N_2077);
and U2122 (N_2122,N_1982,N_2068);
nor U2123 (N_2123,N_2017,N_2010);
or U2124 (N_2124,N_2024,N_2051);
or U2125 (N_2125,N_1927,N_2036);
nor U2126 (N_2126,N_1939,N_1989);
or U2127 (N_2127,N_1937,N_1999);
nor U2128 (N_2128,N_2061,N_2076);
nor U2129 (N_2129,N_1962,N_1943);
or U2130 (N_2130,N_1967,N_2048);
nand U2131 (N_2131,N_2052,N_1968);
nand U2132 (N_2132,N_1998,N_1970);
nor U2133 (N_2133,N_1971,N_2013);
and U2134 (N_2134,N_1946,N_2067);
and U2135 (N_2135,N_1975,N_2075);
and U2136 (N_2136,N_2056,N_2049);
or U2137 (N_2137,N_1944,N_2074);
and U2138 (N_2138,N_1960,N_2018);
or U2139 (N_2139,N_2014,N_1987);
nor U2140 (N_2140,N_1956,N_2073);
xor U2141 (N_2141,N_2072,N_1953);
nand U2142 (N_2142,N_2079,N_1950);
and U2143 (N_2143,N_1947,N_1942);
and U2144 (N_2144,N_2041,N_2004);
or U2145 (N_2145,N_1984,N_2058);
and U2146 (N_2146,N_2007,N_2023);
or U2147 (N_2147,N_1922,N_1988);
xor U2148 (N_2148,N_2003,N_2045);
nand U2149 (N_2149,N_2053,N_1983);
nor U2150 (N_2150,N_1961,N_2042);
nor U2151 (N_2151,N_2006,N_1995);
xor U2152 (N_2152,N_1954,N_1945);
nand U2153 (N_2153,N_1920,N_2050);
and U2154 (N_2154,N_1973,N_1963);
or U2155 (N_2155,N_2039,N_2065);
and U2156 (N_2156,N_2027,N_2002);
nand U2157 (N_2157,N_2031,N_1986);
nor U2158 (N_2158,N_2037,N_2012);
nor U2159 (N_2159,N_2038,N_2046);
and U2160 (N_2160,N_1951,N_1984);
xor U2161 (N_2161,N_1944,N_2008);
nor U2162 (N_2162,N_2058,N_1932);
nand U2163 (N_2163,N_2073,N_2006);
and U2164 (N_2164,N_2009,N_2020);
xnor U2165 (N_2165,N_2006,N_1957);
or U2166 (N_2166,N_2038,N_2068);
or U2167 (N_2167,N_2020,N_1949);
nor U2168 (N_2168,N_2025,N_1943);
or U2169 (N_2169,N_2038,N_2069);
nor U2170 (N_2170,N_2001,N_2040);
nand U2171 (N_2171,N_2040,N_2048);
or U2172 (N_2172,N_1931,N_2053);
xnor U2173 (N_2173,N_2020,N_1933);
or U2174 (N_2174,N_2008,N_2063);
nand U2175 (N_2175,N_1991,N_1950);
and U2176 (N_2176,N_2046,N_2068);
or U2177 (N_2177,N_2000,N_1968);
nand U2178 (N_2178,N_1990,N_2026);
and U2179 (N_2179,N_1970,N_1964);
nor U2180 (N_2180,N_1955,N_1967);
and U2181 (N_2181,N_2004,N_1928);
or U2182 (N_2182,N_1936,N_1934);
and U2183 (N_2183,N_2050,N_2035);
and U2184 (N_2184,N_2009,N_2022);
nor U2185 (N_2185,N_1961,N_1934);
or U2186 (N_2186,N_2041,N_1951);
and U2187 (N_2187,N_2020,N_1942);
or U2188 (N_2188,N_1940,N_2059);
nor U2189 (N_2189,N_1920,N_2053);
or U2190 (N_2190,N_1931,N_1952);
or U2191 (N_2191,N_2055,N_2043);
nand U2192 (N_2192,N_1942,N_1984);
and U2193 (N_2193,N_2008,N_2045);
and U2194 (N_2194,N_1987,N_1990);
and U2195 (N_2195,N_1964,N_2049);
nor U2196 (N_2196,N_1975,N_1959);
or U2197 (N_2197,N_2035,N_2044);
and U2198 (N_2198,N_1928,N_1983);
nor U2199 (N_2199,N_2023,N_1937);
and U2200 (N_2200,N_1965,N_1931);
or U2201 (N_2201,N_2018,N_1994);
and U2202 (N_2202,N_1944,N_1930);
and U2203 (N_2203,N_2003,N_1934);
nand U2204 (N_2204,N_2019,N_2041);
or U2205 (N_2205,N_2040,N_2027);
nor U2206 (N_2206,N_1945,N_2053);
nor U2207 (N_2207,N_1965,N_2058);
and U2208 (N_2208,N_2056,N_1931);
nand U2209 (N_2209,N_2036,N_1947);
nand U2210 (N_2210,N_2045,N_1946);
nor U2211 (N_2211,N_1958,N_1979);
nand U2212 (N_2212,N_1988,N_2038);
nor U2213 (N_2213,N_2061,N_1977);
and U2214 (N_2214,N_1997,N_2014);
and U2215 (N_2215,N_1943,N_2063);
and U2216 (N_2216,N_2066,N_2042);
nand U2217 (N_2217,N_2048,N_2036);
or U2218 (N_2218,N_2013,N_1928);
or U2219 (N_2219,N_1929,N_1968);
nor U2220 (N_2220,N_2062,N_1945);
nand U2221 (N_2221,N_2046,N_2051);
or U2222 (N_2222,N_1938,N_1929);
nor U2223 (N_2223,N_1984,N_1966);
nand U2224 (N_2224,N_1937,N_1929);
nor U2225 (N_2225,N_2072,N_2045);
nand U2226 (N_2226,N_2073,N_1924);
or U2227 (N_2227,N_1971,N_1938);
and U2228 (N_2228,N_2001,N_2078);
xnor U2229 (N_2229,N_2026,N_2042);
and U2230 (N_2230,N_1989,N_1995);
nand U2231 (N_2231,N_1973,N_1964);
and U2232 (N_2232,N_2051,N_2006);
nand U2233 (N_2233,N_2021,N_1996);
nand U2234 (N_2234,N_1933,N_2044);
and U2235 (N_2235,N_2010,N_1921);
and U2236 (N_2236,N_1986,N_1972);
nand U2237 (N_2237,N_2012,N_1961);
nor U2238 (N_2238,N_1993,N_2027);
nand U2239 (N_2239,N_2043,N_1979);
or U2240 (N_2240,N_2126,N_2211);
nor U2241 (N_2241,N_2165,N_2162);
or U2242 (N_2242,N_2125,N_2127);
nand U2243 (N_2243,N_2218,N_2195);
or U2244 (N_2244,N_2095,N_2215);
nor U2245 (N_2245,N_2205,N_2140);
and U2246 (N_2246,N_2239,N_2201);
nand U2247 (N_2247,N_2204,N_2132);
or U2248 (N_2248,N_2129,N_2128);
nand U2249 (N_2249,N_2091,N_2133);
nand U2250 (N_2250,N_2191,N_2123);
nand U2251 (N_2251,N_2089,N_2170);
nor U2252 (N_2252,N_2176,N_2206);
and U2253 (N_2253,N_2082,N_2097);
nand U2254 (N_2254,N_2157,N_2137);
or U2255 (N_2255,N_2146,N_2136);
nor U2256 (N_2256,N_2203,N_2160);
and U2257 (N_2257,N_2214,N_2186);
and U2258 (N_2258,N_2210,N_2138);
nand U2259 (N_2259,N_2233,N_2238);
and U2260 (N_2260,N_2083,N_2142);
nor U2261 (N_2261,N_2149,N_2171);
xnor U2262 (N_2262,N_2164,N_2086);
or U2263 (N_2263,N_2225,N_2209);
nand U2264 (N_2264,N_2122,N_2084);
and U2265 (N_2265,N_2236,N_2096);
or U2266 (N_2266,N_2158,N_2234);
and U2267 (N_2267,N_2085,N_2114);
and U2268 (N_2268,N_2151,N_2183);
nor U2269 (N_2269,N_2194,N_2202);
and U2270 (N_2270,N_2232,N_2155);
nor U2271 (N_2271,N_2168,N_2144);
nand U2272 (N_2272,N_2116,N_2150);
nand U2273 (N_2273,N_2222,N_2227);
nand U2274 (N_2274,N_2098,N_2111);
and U2275 (N_2275,N_2216,N_2212);
and U2276 (N_2276,N_2231,N_2094);
and U2277 (N_2277,N_2099,N_2179);
nor U2278 (N_2278,N_2115,N_2147);
nor U2279 (N_2279,N_2235,N_2121);
and U2280 (N_2280,N_2088,N_2185);
or U2281 (N_2281,N_2229,N_2112);
nand U2282 (N_2282,N_2220,N_2101);
or U2283 (N_2283,N_2224,N_2159);
nor U2284 (N_2284,N_2230,N_2187);
nor U2285 (N_2285,N_2174,N_2197);
or U2286 (N_2286,N_2169,N_2184);
and U2287 (N_2287,N_2134,N_2108);
or U2288 (N_2288,N_2166,N_2196);
nor U2289 (N_2289,N_2213,N_2104);
or U2290 (N_2290,N_2120,N_2207);
xor U2291 (N_2291,N_2188,N_2105);
nand U2292 (N_2292,N_2237,N_2154);
nand U2293 (N_2293,N_2118,N_2182);
or U2294 (N_2294,N_2192,N_2223);
nand U2295 (N_2295,N_2080,N_2102);
nand U2296 (N_2296,N_2180,N_2130);
nor U2297 (N_2297,N_2228,N_2163);
nand U2298 (N_2298,N_2106,N_2139);
nor U2299 (N_2299,N_2109,N_2081);
nand U2300 (N_2300,N_2193,N_2093);
nor U2301 (N_2301,N_2148,N_2103);
xnor U2302 (N_2302,N_2208,N_2152);
nand U2303 (N_2303,N_2189,N_2221);
and U2304 (N_2304,N_2219,N_2145);
nor U2305 (N_2305,N_2178,N_2087);
and U2306 (N_2306,N_2199,N_2173);
nor U2307 (N_2307,N_2190,N_2124);
nand U2308 (N_2308,N_2107,N_2167);
nor U2309 (N_2309,N_2110,N_2175);
and U2310 (N_2310,N_2141,N_2156);
or U2311 (N_2311,N_2177,N_2100);
or U2312 (N_2312,N_2135,N_2143);
and U2313 (N_2313,N_2131,N_2217);
and U2314 (N_2314,N_2172,N_2090);
and U2315 (N_2315,N_2226,N_2092);
xnor U2316 (N_2316,N_2181,N_2198);
nor U2317 (N_2317,N_2153,N_2113);
or U2318 (N_2318,N_2119,N_2117);
nand U2319 (N_2319,N_2161,N_2200);
and U2320 (N_2320,N_2213,N_2157);
or U2321 (N_2321,N_2182,N_2202);
nor U2322 (N_2322,N_2154,N_2234);
xor U2323 (N_2323,N_2226,N_2087);
nor U2324 (N_2324,N_2116,N_2139);
xnor U2325 (N_2325,N_2178,N_2229);
nand U2326 (N_2326,N_2104,N_2181);
nand U2327 (N_2327,N_2104,N_2237);
and U2328 (N_2328,N_2122,N_2150);
nor U2329 (N_2329,N_2164,N_2157);
xnor U2330 (N_2330,N_2099,N_2096);
and U2331 (N_2331,N_2206,N_2167);
xor U2332 (N_2332,N_2198,N_2132);
or U2333 (N_2333,N_2181,N_2134);
or U2334 (N_2334,N_2170,N_2126);
xnor U2335 (N_2335,N_2087,N_2192);
nand U2336 (N_2336,N_2222,N_2108);
or U2337 (N_2337,N_2210,N_2170);
and U2338 (N_2338,N_2097,N_2093);
nor U2339 (N_2339,N_2111,N_2182);
xnor U2340 (N_2340,N_2220,N_2237);
nor U2341 (N_2341,N_2108,N_2213);
xnor U2342 (N_2342,N_2182,N_2166);
nand U2343 (N_2343,N_2165,N_2125);
or U2344 (N_2344,N_2164,N_2169);
and U2345 (N_2345,N_2154,N_2110);
xnor U2346 (N_2346,N_2100,N_2168);
or U2347 (N_2347,N_2096,N_2224);
nand U2348 (N_2348,N_2095,N_2105);
or U2349 (N_2349,N_2089,N_2169);
and U2350 (N_2350,N_2219,N_2196);
nor U2351 (N_2351,N_2112,N_2088);
and U2352 (N_2352,N_2201,N_2165);
or U2353 (N_2353,N_2160,N_2127);
nor U2354 (N_2354,N_2155,N_2096);
and U2355 (N_2355,N_2141,N_2209);
or U2356 (N_2356,N_2119,N_2110);
xor U2357 (N_2357,N_2161,N_2159);
or U2358 (N_2358,N_2239,N_2144);
or U2359 (N_2359,N_2180,N_2157);
nor U2360 (N_2360,N_2203,N_2201);
nand U2361 (N_2361,N_2160,N_2181);
nand U2362 (N_2362,N_2165,N_2129);
or U2363 (N_2363,N_2117,N_2139);
nand U2364 (N_2364,N_2128,N_2117);
and U2365 (N_2365,N_2184,N_2166);
xnor U2366 (N_2366,N_2171,N_2124);
or U2367 (N_2367,N_2111,N_2200);
and U2368 (N_2368,N_2177,N_2142);
nand U2369 (N_2369,N_2167,N_2237);
nand U2370 (N_2370,N_2084,N_2189);
nor U2371 (N_2371,N_2221,N_2122);
xor U2372 (N_2372,N_2080,N_2112);
or U2373 (N_2373,N_2112,N_2110);
and U2374 (N_2374,N_2085,N_2199);
nand U2375 (N_2375,N_2123,N_2154);
or U2376 (N_2376,N_2224,N_2091);
or U2377 (N_2377,N_2123,N_2157);
and U2378 (N_2378,N_2104,N_2190);
or U2379 (N_2379,N_2132,N_2084);
or U2380 (N_2380,N_2115,N_2186);
and U2381 (N_2381,N_2225,N_2197);
nand U2382 (N_2382,N_2189,N_2147);
nand U2383 (N_2383,N_2105,N_2120);
nand U2384 (N_2384,N_2181,N_2081);
nor U2385 (N_2385,N_2081,N_2197);
and U2386 (N_2386,N_2230,N_2156);
and U2387 (N_2387,N_2183,N_2095);
and U2388 (N_2388,N_2221,N_2179);
nor U2389 (N_2389,N_2081,N_2099);
and U2390 (N_2390,N_2159,N_2207);
or U2391 (N_2391,N_2204,N_2179);
and U2392 (N_2392,N_2090,N_2216);
and U2393 (N_2393,N_2117,N_2105);
nand U2394 (N_2394,N_2158,N_2161);
nor U2395 (N_2395,N_2134,N_2147);
and U2396 (N_2396,N_2145,N_2163);
nor U2397 (N_2397,N_2105,N_2106);
or U2398 (N_2398,N_2147,N_2195);
nor U2399 (N_2399,N_2203,N_2149);
nor U2400 (N_2400,N_2351,N_2280);
nor U2401 (N_2401,N_2380,N_2307);
nand U2402 (N_2402,N_2350,N_2265);
nand U2403 (N_2403,N_2397,N_2311);
and U2404 (N_2404,N_2282,N_2346);
or U2405 (N_2405,N_2301,N_2304);
and U2406 (N_2406,N_2343,N_2240);
xnor U2407 (N_2407,N_2257,N_2322);
nand U2408 (N_2408,N_2308,N_2283);
nor U2409 (N_2409,N_2394,N_2362);
and U2410 (N_2410,N_2375,N_2312);
or U2411 (N_2411,N_2399,N_2297);
nand U2412 (N_2412,N_2390,N_2363);
and U2413 (N_2413,N_2245,N_2371);
nor U2414 (N_2414,N_2319,N_2263);
and U2415 (N_2415,N_2339,N_2258);
or U2416 (N_2416,N_2378,N_2298);
and U2417 (N_2417,N_2340,N_2335);
nor U2418 (N_2418,N_2296,N_2243);
nand U2419 (N_2419,N_2344,N_2281);
or U2420 (N_2420,N_2347,N_2295);
nand U2421 (N_2421,N_2269,N_2328);
or U2422 (N_2422,N_2255,N_2361);
nand U2423 (N_2423,N_2373,N_2294);
or U2424 (N_2424,N_2355,N_2264);
nand U2425 (N_2425,N_2268,N_2267);
or U2426 (N_2426,N_2254,N_2248);
or U2427 (N_2427,N_2377,N_2315);
nand U2428 (N_2428,N_2324,N_2366);
or U2429 (N_2429,N_2381,N_2259);
nor U2430 (N_2430,N_2293,N_2342);
or U2431 (N_2431,N_2289,N_2285);
and U2432 (N_2432,N_2320,N_2246);
or U2433 (N_2433,N_2274,N_2360);
nand U2434 (N_2434,N_2327,N_2241);
and U2435 (N_2435,N_2253,N_2306);
and U2436 (N_2436,N_2310,N_2333);
or U2437 (N_2437,N_2290,N_2341);
nor U2438 (N_2438,N_2331,N_2266);
and U2439 (N_2439,N_2299,N_2396);
nor U2440 (N_2440,N_2352,N_2385);
or U2441 (N_2441,N_2279,N_2348);
or U2442 (N_2442,N_2389,N_2330);
or U2443 (N_2443,N_2372,N_2383);
and U2444 (N_2444,N_2286,N_2261);
or U2445 (N_2445,N_2345,N_2247);
nand U2446 (N_2446,N_2278,N_2323);
nor U2447 (N_2447,N_2272,N_2317);
or U2448 (N_2448,N_2384,N_2250);
xnor U2449 (N_2449,N_2398,N_2357);
nor U2450 (N_2450,N_2338,N_2392);
and U2451 (N_2451,N_2356,N_2277);
nor U2452 (N_2452,N_2291,N_2354);
and U2453 (N_2453,N_2364,N_2332);
and U2454 (N_2454,N_2386,N_2292);
nor U2455 (N_2455,N_2242,N_2359);
nor U2456 (N_2456,N_2334,N_2321);
and U2457 (N_2457,N_2368,N_2275);
nor U2458 (N_2458,N_2244,N_2284);
and U2459 (N_2459,N_2270,N_2318);
nor U2460 (N_2460,N_2382,N_2326);
nand U2461 (N_2461,N_2251,N_2369);
or U2462 (N_2462,N_2329,N_2276);
and U2463 (N_2463,N_2393,N_2262);
or U2464 (N_2464,N_2353,N_2271);
nor U2465 (N_2465,N_2358,N_2388);
or U2466 (N_2466,N_2387,N_2370);
or U2467 (N_2467,N_2309,N_2305);
nor U2468 (N_2468,N_2256,N_2336);
nand U2469 (N_2469,N_2273,N_2365);
nand U2470 (N_2470,N_2288,N_2325);
nand U2471 (N_2471,N_2300,N_2303);
and U2472 (N_2472,N_2349,N_2379);
and U2473 (N_2473,N_2376,N_2314);
or U2474 (N_2474,N_2395,N_2367);
nand U2475 (N_2475,N_2287,N_2252);
nand U2476 (N_2476,N_2260,N_2337);
nand U2477 (N_2477,N_2302,N_2316);
and U2478 (N_2478,N_2391,N_2313);
or U2479 (N_2479,N_2374,N_2249);
nor U2480 (N_2480,N_2275,N_2293);
nand U2481 (N_2481,N_2286,N_2322);
and U2482 (N_2482,N_2288,N_2369);
or U2483 (N_2483,N_2286,N_2383);
and U2484 (N_2484,N_2290,N_2396);
nand U2485 (N_2485,N_2302,N_2362);
and U2486 (N_2486,N_2323,N_2306);
and U2487 (N_2487,N_2379,N_2351);
and U2488 (N_2488,N_2307,N_2247);
and U2489 (N_2489,N_2264,N_2244);
and U2490 (N_2490,N_2381,N_2258);
nor U2491 (N_2491,N_2245,N_2344);
nand U2492 (N_2492,N_2323,N_2365);
nand U2493 (N_2493,N_2370,N_2350);
nor U2494 (N_2494,N_2361,N_2396);
xnor U2495 (N_2495,N_2356,N_2350);
nor U2496 (N_2496,N_2285,N_2342);
or U2497 (N_2497,N_2377,N_2297);
and U2498 (N_2498,N_2328,N_2302);
nor U2499 (N_2499,N_2288,N_2267);
nand U2500 (N_2500,N_2252,N_2340);
nor U2501 (N_2501,N_2385,N_2376);
nand U2502 (N_2502,N_2397,N_2355);
nor U2503 (N_2503,N_2352,N_2390);
or U2504 (N_2504,N_2311,N_2299);
nand U2505 (N_2505,N_2241,N_2272);
nand U2506 (N_2506,N_2312,N_2319);
nor U2507 (N_2507,N_2341,N_2312);
nor U2508 (N_2508,N_2261,N_2289);
and U2509 (N_2509,N_2253,N_2369);
and U2510 (N_2510,N_2286,N_2254);
xnor U2511 (N_2511,N_2304,N_2367);
nor U2512 (N_2512,N_2240,N_2276);
nor U2513 (N_2513,N_2397,N_2259);
nor U2514 (N_2514,N_2347,N_2308);
nor U2515 (N_2515,N_2252,N_2306);
and U2516 (N_2516,N_2388,N_2257);
nand U2517 (N_2517,N_2314,N_2267);
or U2518 (N_2518,N_2349,N_2337);
nand U2519 (N_2519,N_2266,N_2315);
nand U2520 (N_2520,N_2295,N_2385);
or U2521 (N_2521,N_2378,N_2307);
nor U2522 (N_2522,N_2246,N_2262);
xnor U2523 (N_2523,N_2396,N_2253);
or U2524 (N_2524,N_2302,N_2275);
or U2525 (N_2525,N_2256,N_2352);
and U2526 (N_2526,N_2253,N_2387);
or U2527 (N_2527,N_2252,N_2250);
nor U2528 (N_2528,N_2245,N_2243);
nand U2529 (N_2529,N_2275,N_2391);
nor U2530 (N_2530,N_2329,N_2396);
or U2531 (N_2531,N_2379,N_2281);
nand U2532 (N_2532,N_2291,N_2269);
nand U2533 (N_2533,N_2365,N_2397);
nor U2534 (N_2534,N_2293,N_2366);
and U2535 (N_2535,N_2269,N_2388);
nor U2536 (N_2536,N_2280,N_2240);
nor U2537 (N_2537,N_2393,N_2268);
nor U2538 (N_2538,N_2373,N_2338);
or U2539 (N_2539,N_2355,N_2268);
and U2540 (N_2540,N_2261,N_2242);
and U2541 (N_2541,N_2288,N_2313);
xnor U2542 (N_2542,N_2264,N_2248);
or U2543 (N_2543,N_2300,N_2371);
nor U2544 (N_2544,N_2284,N_2323);
or U2545 (N_2545,N_2323,N_2352);
and U2546 (N_2546,N_2305,N_2310);
xnor U2547 (N_2547,N_2292,N_2299);
and U2548 (N_2548,N_2320,N_2270);
nand U2549 (N_2549,N_2241,N_2357);
nor U2550 (N_2550,N_2299,N_2253);
nand U2551 (N_2551,N_2348,N_2304);
nand U2552 (N_2552,N_2344,N_2283);
or U2553 (N_2553,N_2349,N_2290);
and U2554 (N_2554,N_2304,N_2262);
xnor U2555 (N_2555,N_2277,N_2359);
nor U2556 (N_2556,N_2240,N_2328);
nor U2557 (N_2557,N_2356,N_2389);
nand U2558 (N_2558,N_2349,N_2399);
or U2559 (N_2559,N_2343,N_2381);
nand U2560 (N_2560,N_2502,N_2465);
nor U2561 (N_2561,N_2546,N_2483);
and U2562 (N_2562,N_2550,N_2409);
and U2563 (N_2563,N_2410,N_2541);
nand U2564 (N_2564,N_2453,N_2457);
nand U2565 (N_2565,N_2493,N_2537);
nor U2566 (N_2566,N_2495,N_2479);
nor U2567 (N_2567,N_2451,N_2532);
nand U2568 (N_2568,N_2531,N_2452);
or U2569 (N_2569,N_2519,N_2400);
nand U2570 (N_2570,N_2506,N_2503);
and U2571 (N_2571,N_2413,N_2428);
and U2572 (N_2572,N_2497,N_2415);
xnor U2573 (N_2573,N_2478,N_2548);
or U2574 (N_2574,N_2458,N_2491);
and U2575 (N_2575,N_2402,N_2484);
nor U2576 (N_2576,N_2448,N_2508);
and U2577 (N_2577,N_2481,N_2547);
nor U2578 (N_2578,N_2456,N_2439);
nand U2579 (N_2579,N_2486,N_2435);
and U2580 (N_2580,N_2433,N_2529);
or U2581 (N_2581,N_2553,N_2445);
or U2582 (N_2582,N_2404,N_2545);
or U2583 (N_2583,N_2462,N_2432);
and U2584 (N_2584,N_2510,N_2450);
nand U2585 (N_2585,N_2437,N_2496);
and U2586 (N_2586,N_2468,N_2549);
nand U2587 (N_2587,N_2438,N_2431);
nand U2588 (N_2588,N_2473,N_2408);
nand U2589 (N_2589,N_2426,N_2518);
and U2590 (N_2590,N_2471,N_2512);
and U2591 (N_2591,N_2405,N_2418);
nor U2592 (N_2592,N_2469,N_2425);
and U2593 (N_2593,N_2513,N_2515);
nor U2594 (N_2594,N_2476,N_2434);
xor U2595 (N_2595,N_2521,N_2422);
nor U2596 (N_2596,N_2470,N_2558);
nand U2597 (N_2597,N_2464,N_2528);
nand U2598 (N_2598,N_2534,N_2460);
or U2599 (N_2599,N_2505,N_2429);
and U2600 (N_2600,N_2416,N_2504);
and U2601 (N_2601,N_2480,N_2485);
and U2602 (N_2602,N_2459,N_2419);
nand U2603 (N_2603,N_2556,N_2430);
nand U2604 (N_2604,N_2499,N_2444);
or U2605 (N_2605,N_2492,N_2551);
xnor U2606 (N_2606,N_2509,N_2488);
nand U2607 (N_2607,N_2441,N_2542);
nand U2608 (N_2608,N_2474,N_2522);
nand U2609 (N_2609,N_2498,N_2477);
nand U2610 (N_2610,N_2423,N_2552);
and U2611 (N_2611,N_2555,N_2427);
and U2612 (N_2612,N_2501,N_2455);
xor U2613 (N_2613,N_2401,N_2412);
nor U2614 (N_2614,N_2511,N_2533);
nand U2615 (N_2615,N_2527,N_2543);
xnor U2616 (N_2616,N_2446,N_2475);
nor U2617 (N_2617,N_2466,N_2539);
or U2618 (N_2618,N_2524,N_2514);
nor U2619 (N_2619,N_2517,N_2443);
and U2620 (N_2620,N_2406,N_2490);
nand U2621 (N_2621,N_2461,N_2411);
nor U2622 (N_2622,N_2424,N_2540);
or U2623 (N_2623,N_2544,N_2507);
and U2624 (N_2624,N_2414,N_2447);
or U2625 (N_2625,N_2538,N_2554);
and U2626 (N_2626,N_2525,N_2472);
and U2627 (N_2627,N_2516,N_2440);
nand U2628 (N_2628,N_2436,N_2535);
or U2629 (N_2629,N_2526,N_2417);
and U2630 (N_2630,N_2421,N_2520);
nor U2631 (N_2631,N_2463,N_2454);
xor U2632 (N_2632,N_2500,N_2442);
xor U2633 (N_2633,N_2536,N_2557);
xnor U2634 (N_2634,N_2482,N_2523);
nor U2635 (N_2635,N_2494,N_2420);
or U2636 (N_2636,N_2487,N_2489);
or U2637 (N_2637,N_2403,N_2559);
nor U2638 (N_2638,N_2467,N_2530);
nor U2639 (N_2639,N_2407,N_2449);
nor U2640 (N_2640,N_2550,N_2417);
nand U2641 (N_2641,N_2484,N_2540);
nand U2642 (N_2642,N_2442,N_2514);
or U2643 (N_2643,N_2426,N_2414);
nor U2644 (N_2644,N_2558,N_2530);
nand U2645 (N_2645,N_2541,N_2418);
or U2646 (N_2646,N_2514,N_2431);
nand U2647 (N_2647,N_2559,N_2480);
nor U2648 (N_2648,N_2514,N_2434);
and U2649 (N_2649,N_2530,N_2485);
xnor U2650 (N_2650,N_2438,N_2493);
nor U2651 (N_2651,N_2413,N_2494);
or U2652 (N_2652,N_2511,N_2460);
nor U2653 (N_2653,N_2519,N_2504);
xor U2654 (N_2654,N_2487,N_2417);
nand U2655 (N_2655,N_2481,N_2416);
xor U2656 (N_2656,N_2535,N_2472);
nor U2657 (N_2657,N_2511,N_2518);
xnor U2658 (N_2658,N_2474,N_2521);
nor U2659 (N_2659,N_2509,N_2500);
nand U2660 (N_2660,N_2505,N_2453);
and U2661 (N_2661,N_2524,N_2490);
nand U2662 (N_2662,N_2451,N_2429);
nand U2663 (N_2663,N_2418,N_2501);
or U2664 (N_2664,N_2448,N_2454);
and U2665 (N_2665,N_2403,N_2483);
and U2666 (N_2666,N_2498,N_2511);
and U2667 (N_2667,N_2422,N_2424);
nor U2668 (N_2668,N_2481,N_2444);
and U2669 (N_2669,N_2509,N_2408);
and U2670 (N_2670,N_2445,N_2403);
nor U2671 (N_2671,N_2525,N_2489);
or U2672 (N_2672,N_2545,N_2554);
nor U2673 (N_2673,N_2535,N_2483);
xor U2674 (N_2674,N_2422,N_2455);
nor U2675 (N_2675,N_2451,N_2434);
or U2676 (N_2676,N_2502,N_2531);
or U2677 (N_2677,N_2485,N_2522);
nand U2678 (N_2678,N_2495,N_2501);
and U2679 (N_2679,N_2527,N_2403);
and U2680 (N_2680,N_2476,N_2540);
xor U2681 (N_2681,N_2553,N_2556);
xnor U2682 (N_2682,N_2475,N_2408);
and U2683 (N_2683,N_2523,N_2530);
or U2684 (N_2684,N_2472,N_2501);
and U2685 (N_2685,N_2530,N_2539);
or U2686 (N_2686,N_2527,N_2469);
nor U2687 (N_2687,N_2493,N_2514);
nor U2688 (N_2688,N_2489,N_2411);
and U2689 (N_2689,N_2483,N_2412);
nand U2690 (N_2690,N_2419,N_2410);
and U2691 (N_2691,N_2468,N_2489);
nand U2692 (N_2692,N_2425,N_2522);
and U2693 (N_2693,N_2430,N_2513);
nor U2694 (N_2694,N_2507,N_2470);
or U2695 (N_2695,N_2503,N_2417);
and U2696 (N_2696,N_2542,N_2471);
nand U2697 (N_2697,N_2511,N_2420);
or U2698 (N_2698,N_2479,N_2530);
nor U2699 (N_2699,N_2508,N_2422);
nor U2700 (N_2700,N_2424,N_2544);
nand U2701 (N_2701,N_2471,N_2406);
and U2702 (N_2702,N_2492,N_2508);
or U2703 (N_2703,N_2480,N_2434);
or U2704 (N_2704,N_2498,N_2425);
xor U2705 (N_2705,N_2426,N_2409);
or U2706 (N_2706,N_2413,N_2400);
xor U2707 (N_2707,N_2535,N_2424);
xnor U2708 (N_2708,N_2543,N_2513);
nand U2709 (N_2709,N_2461,N_2547);
nor U2710 (N_2710,N_2477,N_2439);
and U2711 (N_2711,N_2469,N_2511);
nor U2712 (N_2712,N_2443,N_2400);
and U2713 (N_2713,N_2536,N_2544);
nand U2714 (N_2714,N_2472,N_2556);
and U2715 (N_2715,N_2462,N_2426);
nor U2716 (N_2716,N_2480,N_2410);
xnor U2717 (N_2717,N_2401,N_2450);
or U2718 (N_2718,N_2549,N_2548);
or U2719 (N_2719,N_2460,N_2537);
or U2720 (N_2720,N_2606,N_2624);
and U2721 (N_2721,N_2594,N_2694);
and U2722 (N_2722,N_2658,N_2649);
and U2723 (N_2723,N_2561,N_2697);
xnor U2724 (N_2724,N_2705,N_2693);
or U2725 (N_2725,N_2566,N_2619);
and U2726 (N_2726,N_2716,N_2709);
and U2727 (N_2727,N_2632,N_2615);
nor U2728 (N_2728,N_2569,N_2698);
and U2729 (N_2729,N_2590,N_2682);
nand U2730 (N_2730,N_2580,N_2562);
nand U2731 (N_2731,N_2611,N_2651);
nand U2732 (N_2732,N_2687,N_2644);
nor U2733 (N_2733,N_2599,N_2655);
or U2734 (N_2734,N_2598,N_2672);
nor U2735 (N_2735,N_2674,N_2690);
and U2736 (N_2736,N_2581,N_2616);
and U2737 (N_2737,N_2684,N_2662);
or U2738 (N_2738,N_2686,N_2717);
nand U2739 (N_2739,N_2592,N_2669);
nor U2740 (N_2740,N_2646,N_2608);
nor U2741 (N_2741,N_2579,N_2623);
nor U2742 (N_2742,N_2691,N_2703);
nand U2743 (N_2743,N_2650,N_2663);
and U2744 (N_2744,N_2702,N_2696);
nor U2745 (N_2745,N_2596,N_2588);
and U2746 (N_2746,N_2645,N_2701);
nand U2747 (N_2747,N_2583,N_2635);
xor U2748 (N_2748,N_2637,N_2638);
and U2749 (N_2749,N_2677,N_2710);
xor U2750 (N_2750,N_2571,N_2620);
or U2751 (N_2751,N_2667,N_2671);
xnor U2752 (N_2752,N_2679,N_2714);
nand U2753 (N_2753,N_2614,N_2613);
nand U2754 (N_2754,N_2653,N_2657);
xor U2755 (N_2755,N_2586,N_2633);
and U2756 (N_2756,N_2692,N_2640);
nand U2757 (N_2757,N_2708,N_2678);
xor U2758 (N_2758,N_2576,N_2618);
and U2759 (N_2759,N_2680,N_2584);
xnor U2760 (N_2760,N_2572,N_2719);
nor U2761 (N_2761,N_2565,N_2564);
nor U2762 (N_2762,N_2683,N_2612);
nand U2763 (N_2763,N_2641,N_2603);
xnor U2764 (N_2764,N_2634,N_2595);
or U2765 (N_2765,N_2666,N_2673);
nand U2766 (N_2766,N_2648,N_2605);
xor U2767 (N_2767,N_2715,N_2688);
or U2768 (N_2768,N_2695,N_2570);
and U2769 (N_2769,N_2706,N_2601);
or U2770 (N_2770,N_2676,N_2610);
nor U2771 (N_2771,N_2628,N_2699);
nor U2772 (N_2772,N_2626,N_2607);
xnor U2773 (N_2773,N_2681,N_2589);
and U2774 (N_2774,N_2578,N_2660);
and U2775 (N_2775,N_2631,N_2656);
nor U2776 (N_2776,N_2560,N_2668);
xor U2777 (N_2777,N_2568,N_2670);
or U2778 (N_2778,N_2689,N_2629);
or U2779 (N_2779,N_2707,N_2713);
xor U2780 (N_2780,N_2712,N_2573);
and U2781 (N_2781,N_2621,N_2630);
or U2782 (N_2782,N_2643,N_2652);
and U2783 (N_2783,N_2582,N_2685);
nand U2784 (N_2784,N_2622,N_2577);
nor U2785 (N_2785,N_2675,N_2704);
nand U2786 (N_2786,N_2659,N_2639);
or U2787 (N_2787,N_2711,N_2563);
and U2788 (N_2788,N_2600,N_2585);
and U2789 (N_2789,N_2627,N_2597);
nand U2790 (N_2790,N_2593,N_2642);
nor U2791 (N_2791,N_2617,N_2587);
or U2792 (N_2792,N_2661,N_2604);
nand U2793 (N_2793,N_2718,N_2567);
nor U2794 (N_2794,N_2636,N_2647);
nand U2795 (N_2795,N_2574,N_2700);
and U2796 (N_2796,N_2654,N_2591);
nor U2797 (N_2797,N_2665,N_2625);
and U2798 (N_2798,N_2575,N_2602);
nand U2799 (N_2799,N_2609,N_2664);
xor U2800 (N_2800,N_2613,N_2611);
nand U2801 (N_2801,N_2709,N_2622);
xnor U2802 (N_2802,N_2680,N_2695);
nor U2803 (N_2803,N_2598,N_2710);
and U2804 (N_2804,N_2641,N_2567);
and U2805 (N_2805,N_2573,N_2671);
nor U2806 (N_2806,N_2625,N_2590);
xor U2807 (N_2807,N_2652,N_2694);
or U2808 (N_2808,N_2630,N_2692);
and U2809 (N_2809,N_2576,N_2710);
nor U2810 (N_2810,N_2609,N_2638);
or U2811 (N_2811,N_2668,N_2680);
nand U2812 (N_2812,N_2579,N_2642);
nand U2813 (N_2813,N_2643,N_2635);
nor U2814 (N_2814,N_2619,N_2620);
or U2815 (N_2815,N_2566,N_2653);
or U2816 (N_2816,N_2608,N_2585);
nand U2817 (N_2817,N_2597,N_2578);
nand U2818 (N_2818,N_2655,N_2699);
nand U2819 (N_2819,N_2694,N_2710);
nor U2820 (N_2820,N_2654,N_2561);
nand U2821 (N_2821,N_2717,N_2708);
or U2822 (N_2822,N_2624,N_2663);
nor U2823 (N_2823,N_2679,N_2637);
and U2824 (N_2824,N_2578,N_2695);
nor U2825 (N_2825,N_2654,N_2600);
nor U2826 (N_2826,N_2587,N_2657);
and U2827 (N_2827,N_2635,N_2692);
nand U2828 (N_2828,N_2640,N_2672);
nor U2829 (N_2829,N_2603,N_2655);
nor U2830 (N_2830,N_2663,N_2614);
or U2831 (N_2831,N_2583,N_2622);
and U2832 (N_2832,N_2604,N_2639);
nor U2833 (N_2833,N_2626,N_2582);
and U2834 (N_2834,N_2628,N_2598);
xor U2835 (N_2835,N_2711,N_2675);
and U2836 (N_2836,N_2655,N_2578);
and U2837 (N_2837,N_2606,N_2615);
or U2838 (N_2838,N_2666,N_2683);
nor U2839 (N_2839,N_2653,N_2594);
nand U2840 (N_2840,N_2645,N_2638);
nor U2841 (N_2841,N_2570,N_2702);
or U2842 (N_2842,N_2575,N_2652);
nor U2843 (N_2843,N_2660,N_2692);
and U2844 (N_2844,N_2668,N_2683);
nand U2845 (N_2845,N_2583,N_2666);
nor U2846 (N_2846,N_2702,N_2710);
nand U2847 (N_2847,N_2593,N_2569);
nor U2848 (N_2848,N_2578,N_2642);
and U2849 (N_2849,N_2687,N_2641);
or U2850 (N_2850,N_2658,N_2597);
nor U2851 (N_2851,N_2644,N_2594);
nand U2852 (N_2852,N_2635,N_2578);
nand U2853 (N_2853,N_2674,N_2705);
nand U2854 (N_2854,N_2695,N_2568);
or U2855 (N_2855,N_2595,N_2636);
nand U2856 (N_2856,N_2698,N_2587);
nand U2857 (N_2857,N_2605,N_2562);
nand U2858 (N_2858,N_2642,N_2679);
nand U2859 (N_2859,N_2607,N_2622);
nor U2860 (N_2860,N_2617,N_2585);
nand U2861 (N_2861,N_2639,N_2698);
nand U2862 (N_2862,N_2604,N_2574);
nand U2863 (N_2863,N_2635,N_2653);
nor U2864 (N_2864,N_2596,N_2686);
nor U2865 (N_2865,N_2715,N_2680);
and U2866 (N_2866,N_2589,N_2610);
or U2867 (N_2867,N_2651,N_2591);
nand U2868 (N_2868,N_2716,N_2620);
and U2869 (N_2869,N_2639,N_2705);
nor U2870 (N_2870,N_2656,N_2616);
nand U2871 (N_2871,N_2626,N_2597);
and U2872 (N_2872,N_2604,N_2692);
and U2873 (N_2873,N_2591,N_2626);
and U2874 (N_2874,N_2707,N_2681);
nor U2875 (N_2875,N_2708,N_2663);
nor U2876 (N_2876,N_2694,N_2627);
nor U2877 (N_2877,N_2590,N_2701);
or U2878 (N_2878,N_2568,N_2586);
and U2879 (N_2879,N_2656,N_2697);
nor U2880 (N_2880,N_2825,N_2810);
xnor U2881 (N_2881,N_2814,N_2729);
or U2882 (N_2882,N_2796,N_2851);
nand U2883 (N_2883,N_2778,N_2877);
nand U2884 (N_2884,N_2783,N_2732);
xor U2885 (N_2885,N_2782,N_2779);
and U2886 (N_2886,N_2835,N_2840);
and U2887 (N_2887,N_2820,N_2739);
nor U2888 (N_2888,N_2817,N_2836);
or U2889 (N_2889,N_2876,N_2807);
and U2890 (N_2890,N_2758,N_2741);
nor U2891 (N_2891,N_2873,N_2768);
and U2892 (N_2892,N_2766,N_2855);
xnor U2893 (N_2893,N_2770,N_2867);
or U2894 (N_2894,N_2781,N_2813);
and U2895 (N_2895,N_2842,N_2748);
nand U2896 (N_2896,N_2856,N_2799);
and U2897 (N_2897,N_2833,N_2795);
or U2898 (N_2898,N_2720,N_2790);
or U2899 (N_2899,N_2776,N_2747);
and U2900 (N_2900,N_2750,N_2734);
nand U2901 (N_2901,N_2870,N_2763);
nor U2902 (N_2902,N_2859,N_2727);
xor U2903 (N_2903,N_2845,N_2721);
and U2904 (N_2904,N_2846,N_2854);
nor U2905 (N_2905,N_2723,N_2743);
nor U2906 (N_2906,N_2849,N_2733);
or U2907 (N_2907,N_2744,N_2843);
and U2908 (N_2908,N_2822,N_2777);
nand U2909 (N_2909,N_2831,N_2760);
or U2910 (N_2910,N_2737,N_2740);
and U2911 (N_2911,N_2738,N_2751);
nand U2912 (N_2912,N_2728,N_2761);
nor U2913 (N_2913,N_2784,N_2844);
nand U2914 (N_2914,N_2722,N_2756);
nor U2915 (N_2915,N_2786,N_2874);
nor U2916 (N_2916,N_2753,N_2823);
nor U2917 (N_2917,N_2757,N_2818);
or U2918 (N_2918,N_2811,N_2785);
and U2919 (N_2919,N_2746,N_2724);
nor U2920 (N_2920,N_2827,N_2752);
or U2921 (N_2921,N_2839,N_2801);
nand U2922 (N_2922,N_2791,N_2793);
xor U2923 (N_2923,N_2850,N_2774);
nor U2924 (N_2924,N_2787,N_2804);
and U2925 (N_2925,N_2780,N_2730);
nand U2926 (N_2926,N_2860,N_2819);
or U2927 (N_2927,N_2755,N_2834);
xor U2928 (N_2928,N_2794,N_2745);
xnor U2929 (N_2929,N_2731,N_2764);
nor U2930 (N_2930,N_2762,N_2853);
and U2931 (N_2931,N_2830,N_2769);
xor U2932 (N_2932,N_2868,N_2865);
nor U2933 (N_2933,N_2806,N_2771);
nor U2934 (N_2934,N_2879,N_2871);
nand U2935 (N_2935,N_2725,N_2858);
nor U2936 (N_2936,N_2861,N_2841);
and U2937 (N_2937,N_2726,N_2821);
nand U2938 (N_2938,N_2788,N_2828);
or U2939 (N_2939,N_2792,N_2852);
nor U2940 (N_2940,N_2797,N_2829);
or U2941 (N_2941,N_2869,N_2866);
nand U2942 (N_2942,N_2863,N_2803);
nor U2943 (N_2943,N_2800,N_2759);
and U2944 (N_2944,N_2816,N_2805);
or U2945 (N_2945,N_2847,N_2789);
or U2946 (N_2946,N_2767,N_2826);
nand U2947 (N_2947,N_2812,N_2878);
and U2948 (N_2948,N_2862,N_2742);
and U2949 (N_2949,N_2838,N_2837);
nor U2950 (N_2950,N_2875,N_2775);
nor U2951 (N_2951,N_2864,N_2802);
and U2952 (N_2952,N_2832,N_2809);
and U2953 (N_2953,N_2808,N_2824);
nand U2954 (N_2954,N_2773,N_2872);
nand U2955 (N_2955,N_2798,N_2765);
and U2956 (N_2956,N_2749,N_2848);
or U2957 (N_2957,N_2754,N_2857);
xor U2958 (N_2958,N_2735,N_2815);
xor U2959 (N_2959,N_2772,N_2736);
nor U2960 (N_2960,N_2804,N_2808);
nand U2961 (N_2961,N_2744,N_2754);
nor U2962 (N_2962,N_2859,N_2799);
nand U2963 (N_2963,N_2752,N_2878);
nor U2964 (N_2964,N_2760,N_2736);
nand U2965 (N_2965,N_2787,N_2843);
nor U2966 (N_2966,N_2871,N_2797);
xnor U2967 (N_2967,N_2873,N_2764);
nand U2968 (N_2968,N_2728,N_2865);
and U2969 (N_2969,N_2754,N_2810);
and U2970 (N_2970,N_2857,N_2759);
nand U2971 (N_2971,N_2861,N_2734);
or U2972 (N_2972,N_2782,N_2760);
nor U2973 (N_2973,N_2727,N_2732);
or U2974 (N_2974,N_2770,N_2748);
nor U2975 (N_2975,N_2740,N_2776);
nand U2976 (N_2976,N_2876,N_2858);
nand U2977 (N_2977,N_2809,N_2783);
and U2978 (N_2978,N_2850,N_2723);
nor U2979 (N_2979,N_2841,N_2797);
and U2980 (N_2980,N_2766,N_2834);
nor U2981 (N_2981,N_2724,N_2854);
nand U2982 (N_2982,N_2867,N_2782);
nand U2983 (N_2983,N_2747,N_2731);
and U2984 (N_2984,N_2721,N_2822);
or U2985 (N_2985,N_2833,N_2799);
nand U2986 (N_2986,N_2803,N_2763);
or U2987 (N_2987,N_2736,N_2818);
and U2988 (N_2988,N_2741,N_2770);
nor U2989 (N_2989,N_2744,N_2784);
and U2990 (N_2990,N_2731,N_2862);
nor U2991 (N_2991,N_2790,N_2853);
xnor U2992 (N_2992,N_2780,N_2764);
or U2993 (N_2993,N_2879,N_2770);
or U2994 (N_2994,N_2838,N_2755);
nand U2995 (N_2995,N_2738,N_2796);
nand U2996 (N_2996,N_2750,N_2794);
and U2997 (N_2997,N_2811,N_2875);
nand U2998 (N_2998,N_2734,N_2774);
and U2999 (N_2999,N_2784,N_2827);
nor U3000 (N_3000,N_2748,N_2747);
and U3001 (N_3001,N_2808,N_2793);
nand U3002 (N_3002,N_2804,N_2814);
xor U3003 (N_3003,N_2826,N_2875);
nand U3004 (N_3004,N_2861,N_2876);
or U3005 (N_3005,N_2748,N_2829);
and U3006 (N_3006,N_2834,N_2797);
nor U3007 (N_3007,N_2872,N_2820);
and U3008 (N_3008,N_2755,N_2720);
nor U3009 (N_3009,N_2731,N_2773);
xnor U3010 (N_3010,N_2865,N_2869);
and U3011 (N_3011,N_2879,N_2865);
or U3012 (N_3012,N_2820,N_2759);
nor U3013 (N_3013,N_2824,N_2790);
nor U3014 (N_3014,N_2873,N_2829);
nand U3015 (N_3015,N_2772,N_2874);
nor U3016 (N_3016,N_2725,N_2769);
nor U3017 (N_3017,N_2727,N_2786);
nor U3018 (N_3018,N_2721,N_2761);
nand U3019 (N_3019,N_2726,N_2860);
or U3020 (N_3020,N_2722,N_2868);
and U3021 (N_3021,N_2853,N_2851);
and U3022 (N_3022,N_2810,N_2791);
nand U3023 (N_3023,N_2814,N_2859);
nand U3024 (N_3024,N_2874,N_2736);
and U3025 (N_3025,N_2742,N_2820);
nand U3026 (N_3026,N_2864,N_2748);
and U3027 (N_3027,N_2800,N_2818);
nor U3028 (N_3028,N_2801,N_2835);
nor U3029 (N_3029,N_2805,N_2758);
xor U3030 (N_3030,N_2723,N_2751);
xor U3031 (N_3031,N_2799,N_2851);
xor U3032 (N_3032,N_2823,N_2865);
xnor U3033 (N_3033,N_2858,N_2724);
or U3034 (N_3034,N_2729,N_2763);
xor U3035 (N_3035,N_2745,N_2779);
xnor U3036 (N_3036,N_2877,N_2759);
or U3037 (N_3037,N_2834,N_2865);
nand U3038 (N_3038,N_2830,N_2760);
and U3039 (N_3039,N_2730,N_2751);
nor U3040 (N_3040,N_3033,N_3032);
nand U3041 (N_3041,N_2971,N_3014);
nand U3042 (N_3042,N_2914,N_3022);
and U3043 (N_3043,N_2918,N_2958);
nor U3044 (N_3044,N_2932,N_2935);
nand U3045 (N_3045,N_2946,N_2906);
and U3046 (N_3046,N_2908,N_2982);
nor U3047 (N_3047,N_2942,N_2917);
and U3048 (N_3048,N_2987,N_2997);
or U3049 (N_3049,N_2944,N_2952);
nor U3050 (N_3050,N_3036,N_2937);
or U3051 (N_3051,N_2950,N_2986);
nor U3052 (N_3052,N_2895,N_2940);
and U3053 (N_3053,N_2976,N_2911);
and U3054 (N_3054,N_2977,N_2913);
xnor U3055 (N_3055,N_3008,N_3028);
nand U3056 (N_3056,N_3039,N_2883);
or U3057 (N_3057,N_2961,N_2890);
nand U3058 (N_3058,N_3005,N_3030);
nand U3059 (N_3059,N_2999,N_3038);
nor U3060 (N_3060,N_2991,N_2909);
xnor U3061 (N_3061,N_2980,N_2985);
xor U3062 (N_3062,N_2931,N_2926);
or U3063 (N_3063,N_2885,N_2934);
or U3064 (N_3064,N_2981,N_2922);
or U3065 (N_3065,N_2953,N_3037);
nor U3066 (N_3066,N_2897,N_3001);
and U3067 (N_3067,N_2910,N_2888);
nand U3068 (N_3068,N_3009,N_2967);
nor U3069 (N_3069,N_3017,N_2916);
nor U3070 (N_3070,N_2886,N_3007);
nand U3071 (N_3071,N_2929,N_3029);
xnor U3072 (N_3072,N_2983,N_2954);
nand U3073 (N_3073,N_2905,N_2904);
and U3074 (N_3074,N_2969,N_2960);
nor U3075 (N_3075,N_2891,N_3011);
and U3076 (N_3076,N_2898,N_2992);
xnor U3077 (N_3077,N_2941,N_2893);
or U3078 (N_3078,N_3023,N_2968);
nand U3079 (N_3079,N_2892,N_2993);
nor U3080 (N_3080,N_3025,N_3027);
or U3081 (N_3081,N_2887,N_2956);
or U3082 (N_3082,N_3013,N_2963);
nand U3083 (N_3083,N_2882,N_3021);
nor U3084 (N_3084,N_2945,N_2990);
nand U3085 (N_3085,N_2951,N_2974);
and U3086 (N_3086,N_2949,N_2881);
nand U3087 (N_3087,N_2925,N_3031);
nand U3088 (N_3088,N_3034,N_2903);
nor U3089 (N_3089,N_2948,N_2919);
nand U3090 (N_3090,N_2975,N_2936);
or U3091 (N_3091,N_2884,N_2964);
nand U3092 (N_3092,N_2907,N_3020);
or U3093 (N_3093,N_3010,N_2984);
nor U3094 (N_3094,N_2965,N_3003);
and U3095 (N_3095,N_2880,N_3035);
nor U3096 (N_3096,N_2902,N_2994);
and U3097 (N_3097,N_3016,N_2923);
or U3098 (N_3098,N_2912,N_2973);
nand U3099 (N_3099,N_2955,N_2998);
xor U3100 (N_3100,N_2947,N_2900);
and U3101 (N_3101,N_2943,N_3006);
or U3102 (N_3102,N_2988,N_2896);
or U3103 (N_3103,N_3019,N_3000);
and U3104 (N_3104,N_3002,N_2978);
xor U3105 (N_3105,N_2989,N_3024);
nand U3106 (N_3106,N_2939,N_2938);
nand U3107 (N_3107,N_2927,N_2959);
nor U3108 (N_3108,N_2966,N_2901);
nor U3109 (N_3109,N_2915,N_2899);
and U3110 (N_3110,N_2928,N_2889);
and U3111 (N_3111,N_2972,N_2962);
nor U3112 (N_3112,N_2924,N_2957);
nor U3113 (N_3113,N_3004,N_2894);
or U3114 (N_3114,N_2920,N_3018);
nand U3115 (N_3115,N_2995,N_3012);
and U3116 (N_3116,N_2921,N_2979);
or U3117 (N_3117,N_2930,N_2933);
xnor U3118 (N_3118,N_3026,N_2996);
nand U3119 (N_3119,N_2970,N_3015);
xor U3120 (N_3120,N_2954,N_2921);
and U3121 (N_3121,N_2987,N_3000);
and U3122 (N_3122,N_2940,N_2917);
and U3123 (N_3123,N_3025,N_3003);
nor U3124 (N_3124,N_2963,N_3012);
or U3125 (N_3125,N_2982,N_2925);
nor U3126 (N_3126,N_2899,N_2979);
nor U3127 (N_3127,N_2935,N_2964);
xor U3128 (N_3128,N_2931,N_2954);
and U3129 (N_3129,N_2952,N_3010);
or U3130 (N_3130,N_3030,N_2998);
or U3131 (N_3131,N_2991,N_2988);
nand U3132 (N_3132,N_2930,N_2881);
nor U3133 (N_3133,N_2950,N_2992);
xnor U3134 (N_3134,N_2920,N_2918);
nor U3135 (N_3135,N_2943,N_2973);
nand U3136 (N_3136,N_2987,N_2995);
and U3137 (N_3137,N_2952,N_2890);
or U3138 (N_3138,N_2983,N_2995);
nor U3139 (N_3139,N_2971,N_2951);
nand U3140 (N_3140,N_2897,N_2956);
and U3141 (N_3141,N_3007,N_2992);
or U3142 (N_3142,N_2979,N_2897);
and U3143 (N_3143,N_3000,N_2997);
nand U3144 (N_3144,N_2918,N_3036);
nand U3145 (N_3145,N_2897,N_3024);
and U3146 (N_3146,N_3023,N_2973);
nor U3147 (N_3147,N_3028,N_2990);
and U3148 (N_3148,N_2995,N_2957);
xnor U3149 (N_3149,N_2955,N_2898);
nor U3150 (N_3150,N_3021,N_2893);
xnor U3151 (N_3151,N_2975,N_2989);
nand U3152 (N_3152,N_2914,N_2917);
nor U3153 (N_3153,N_2898,N_3035);
nand U3154 (N_3154,N_3012,N_3015);
nor U3155 (N_3155,N_2902,N_2991);
nand U3156 (N_3156,N_3000,N_2937);
or U3157 (N_3157,N_2887,N_2901);
and U3158 (N_3158,N_2945,N_2971);
and U3159 (N_3159,N_3003,N_2999);
and U3160 (N_3160,N_3011,N_3005);
xnor U3161 (N_3161,N_2965,N_2966);
nand U3162 (N_3162,N_2994,N_3003);
nor U3163 (N_3163,N_3007,N_3036);
xnor U3164 (N_3164,N_2957,N_2947);
nor U3165 (N_3165,N_2922,N_3012);
xnor U3166 (N_3166,N_2971,N_2887);
nor U3167 (N_3167,N_2958,N_2899);
nor U3168 (N_3168,N_2969,N_2899);
nor U3169 (N_3169,N_2950,N_2956);
or U3170 (N_3170,N_3003,N_2972);
xor U3171 (N_3171,N_2973,N_2963);
nand U3172 (N_3172,N_2992,N_3033);
or U3173 (N_3173,N_3022,N_2969);
nand U3174 (N_3174,N_2935,N_3029);
nand U3175 (N_3175,N_2990,N_2984);
nor U3176 (N_3176,N_2976,N_2915);
nor U3177 (N_3177,N_2935,N_2908);
nor U3178 (N_3178,N_3005,N_3016);
nor U3179 (N_3179,N_2977,N_2981);
and U3180 (N_3180,N_3033,N_2883);
and U3181 (N_3181,N_3025,N_2890);
nand U3182 (N_3182,N_2905,N_2992);
nor U3183 (N_3183,N_2902,N_3002);
or U3184 (N_3184,N_2890,N_2975);
nor U3185 (N_3185,N_2918,N_2896);
nand U3186 (N_3186,N_2914,N_2908);
or U3187 (N_3187,N_2896,N_3022);
nand U3188 (N_3188,N_2976,N_2972);
or U3189 (N_3189,N_3003,N_2946);
or U3190 (N_3190,N_2959,N_2964);
xnor U3191 (N_3191,N_2993,N_2955);
or U3192 (N_3192,N_3035,N_3026);
or U3193 (N_3193,N_2934,N_2954);
nor U3194 (N_3194,N_2948,N_3007);
or U3195 (N_3195,N_3016,N_3013);
nand U3196 (N_3196,N_2891,N_2886);
nor U3197 (N_3197,N_2900,N_2898);
or U3198 (N_3198,N_3002,N_2885);
or U3199 (N_3199,N_3004,N_3030);
nor U3200 (N_3200,N_3123,N_3098);
xnor U3201 (N_3201,N_3050,N_3074);
and U3202 (N_3202,N_3063,N_3177);
nand U3203 (N_3203,N_3110,N_3122);
and U3204 (N_3204,N_3188,N_3145);
or U3205 (N_3205,N_3092,N_3130);
or U3206 (N_3206,N_3153,N_3192);
xor U3207 (N_3207,N_3101,N_3171);
nor U3208 (N_3208,N_3072,N_3167);
nor U3209 (N_3209,N_3165,N_3174);
and U3210 (N_3210,N_3133,N_3156);
nand U3211 (N_3211,N_3089,N_3047);
and U3212 (N_3212,N_3056,N_3132);
and U3213 (N_3213,N_3182,N_3191);
and U3214 (N_3214,N_3057,N_3172);
and U3215 (N_3215,N_3138,N_3065);
and U3216 (N_3216,N_3094,N_3180);
nor U3217 (N_3217,N_3189,N_3155);
or U3218 (N_3218,N_3120,N_3114);
and U3219 (N_3219,N_3135,N_3176);
nand U3220 (N_3220,N_3186,N_3137);
nor U3221 (N_3221,N_3149,N_3051);
and U3222 (N_3222,N_3157,N_3069);
or U3223 (N_3223,N_3161,N_3158);
nor U3224 (N_3224,N_3040,N_3127);
nand U3225 (N_3225,N_3068,N_3093);
nand U3226 (N_3226,N_3151,N_3116);
nor U3227 (N_3227,N_3199,N_3077);
nor U3228 (N_3228,N_3170,N_3196);
xnor U3229 (N_3229,N_3087,N_3198);
or U3230 (N_3230,N_3108,N_3136);
xnor U3231 (N_3231,N_3084,N_3194);
or U3232 (N_3232,N_3042,N_3091);
nor U3233 (N_3233,N_3066,N_3140);
or U3234 (N_3234,N_3195,N_3046);
or U3235 (N_3235,N_3081,N_3179);
or U3236 (N_3236,N_3141,N_3187);
nand U3237 (N_3237,N_3090,N_3160);
nand U3238 (N_3238,N_3146,N_3163);
and U3239 (N_3239,N_3162,N_3178);
or U3240 (N_3240,N_3104,N_3111);
and U3241 (N_3241,N_3044,N_3097);
nor U3242 (N_3242,N_3070,N_3049);
nand U3243 (N_3243,N_3197,N_3166);
and U3244 (N_3244,N_3175,N_3059);
and U3245 (N_3245,N_3129,N_3086);
or U3246 (N_3246,N_3142,N_3054);
or U3247 (N_3247,N_3121,N_3060);
or U3248 (N_3248,N_3168,N_3144);
xor U3249 (N_3249,N_3190,N_3100);
nand U3250 (N_3250,N_3043,N_3152);
nor U3251 (N_3251,N_3126,N_3107);
and U3252 (N_3252,N_3109,N_3125);
nand U3253 (N_3253,N_3164,N_3143);
or U3254 (N_3254,N_3115,N_3173);
or U3255 (N_3255,N_3147,N_3064);
and U3256 (N_3256,N_3193,N_3124);
or U3257 (N_3257,N_3071,N_3103);
or U3258 (N_3258,N_3183,N_3169);
or U3259 (N_3259,N_3075,N_3088);
and U3260 (N_3260,N_3099,N_3150);
nor U3261 (N_3261,N_3117,N_3052);
nand U3262 (N_3262,N_3106,N_3184);
xor U3263 (N_3263,N_3139,N_3113);
nand U3264 (N_3264,N_3048,N_3067);
nand U3265 (N_3265,N_3083,N_3062);
or U3266 (N_3266,N_3045,N_3080);
nand U3267 (N_3267,N_3061,N_3159);
xnor U3268 (N_3268,N_3128,N_3181);
and U3269 (N_3269,N_3148,N_3102);
or U3270 (N_3270,N_3095,N_3131);
and U3271 (N_3271,N_3185,N_3053);
and U3272 (N_3272,N_3105,N_3058);
and U3273 (N_3273,N_3076,N_3078);
and U3274 (N_3274,N_3073,N_3119);
xor U3275 (N_3275,N_3112,N_3154);
xnor U3276 (N_3276,N_3079,N_3055);
nor U3277 (N_3277,N_3085,N_3041);
nand U3278 (N_3278,N_3096,N_3082);
xor U3279 (N_3279,N_3134,N_3118);
nor U3280 (N_3280,N_3180,N_3195);
nand U3281 (N_3281,N_3190,N_3111);
nand U3282 (N_3282,N_3136,N_3120);
nor U3283 (N_3283,N_3183,N_3054);
and U3284 (N_3284,N_3053,N_3090);
nand U3285 (N_3285,N_3048,N_3112);
nor U3286 (N_3286,N_3123,N_3125);
and U3287 (N_3287,N_3154,N_3087);
nand U3288 (N_3288,N_3082,N_3097);
or U3289 (N_3289,N_3128,N_3044);
nand U3290 (N_3290,N_3158,N_3168);
nand U3291 (N_3291,N_3086,N_3110);
nor U3292 (N_3292,N_3092,N_3091);
xor U3293 (N_3293,N_3166,N_3097);
nand U3294 (N_3294,N_3061,N_3158);
nand U3295 (N_3295,N_3131,N_3072);
or U3296 (N_3296,N_3046,N_3135);
and U3297 (N_3297,N_3169,N_3188);
xor U3298 (N_3298,N_3078,N_3093);
nor U3299 (N_3299,N_3126,N_3134);
nor U3300 (N_3300,N_3120,N_3142);
nand U3301 (N_3301,N_3169,N_3098);
nand U3302 (N_3302,N_3138,N_3061);
and U3303 (N_3303,N_3052,N_3194);
and U3304 (N_3304,N_3187,N_3156);
nor U3305 (N_3305,N_3180,N_3156);
and U3306 (N_3306,N_3158,N_3114);
and U3307 (N_3307,N_3136,N_3183);
nor U3308 (N_3308,N_3064,N_3041);
nor U3309 (N_3309,N_3121,N_3050);
nand U3310 (N_3310,N_3079,N_3197);
xnor U3311 (N_3311,N_3061,N_3095);
and U3312 (N_3312,N_3111,N_3169);
nand U3313 (N_3313,N_3185,N_3170);
and U3314 (N_3314,N_3157,N_3066);
nor U3315 (N_3315,N_3165,N_3064);
nand U3316 (N_3316,N_3165,N_3196);
nand U3317 (N_3317,N_3132,N_3051);
nand U3318 (N_3318,N_3098,N_3181);
nand U3319 (N_3319,N_3081,N_3113);
nand U3320 (N_3320,N_3157,N_3172);
or U3321 (N_3321,N_3152,N_3040);
and U3322 (N_3322,N_3111,N_3087);
and U3323 (N_3323,N_3187,N_3193);
and U3324 (N_3324,N_3136,N_3186);
and U3325 (N_3325,N_3185,N_3174);
and U3326 (N_3326,N_3049,N_3173);
or U3327 (N_3327,N_3153,N_3166);
nand U3328 (N_3328,N_3188,N_3053);
and U3329 (N_3329,N_3123,N_3147);
nor U3330 (N_3330,N_3124,N_3122);
and U3331 (N_3331,N_3113,N_3103);
xnor U3332 (N_3332,N_3089,N_3194);
and U3333 (N_3333,N_3146,N_3116);
xnor U3334 (N_3334,N_3104,N_3170);
nand U3335 (N_3335,N_3198,N_3139);
or U3336 (N_3336,N_3189,N_3069);
nor U3337 (N_3337,N_3123,N_3111);
or U3338 (N_3338,N_3110,N_3178);
nand U3339 (N_3339,N_3071,N_3060);
and U3340 (N_3340,N_3056,N_3049);
nor U3341 (N_3341,N_3159,N_3142);
or U3342 (N_3342,N_3160,N_3158);
nand U3343 (N_3343,N_3148,N_3185);
xnor U3344 (N_3344,N_3054,N_3082);
xnor U3345 (N_3345,N_3096,N_3155);
nand U3346 (N_3346,N_3094,N_3192);
nand U3347 (N_3347,N_3078,N_3147);
xor U3348 (N_3348,N_3167,N_3146);
nor U3349 (N_3349,N_3147,N_3079);
nor U3350 (N_3350,N_3137,N_3049);
nand U3351 (N_3351,N_3122,N_3146);
and U3352 (N_3352,N_3196,N_3144);
or U3353 (N_3353,N_3134,N_3059);
and U3354 (N_3354,N_3145,N_3051);
nand U3355 (N_3355,N_3175,N_3159);
and U3356 (N_3356,N_3160,N_3199);
nand U3357 (N_3357,N_3062,N_3109);
or U3358 (N_3358,N_3155,N_3162);
or U3359 (N_3359,N_3042,N_3065);
nor U3360 (N_3360,N_3204,N_3254);
or U3361 (N_3361,N_3274,N_3332);
or U3362 (N_3362,N_3306,N_3327);
nand U3363 (N_3363,N_3307,N_3252);
nor U3364 (N_3364,N_3203,N_3334);
and U3365 (N_3365,N_3270,N_3271);
nor U3366 (N_3366,N_3237,N_3328);
nor U3367 (N_3367,N_3224,N_3305);
and U3368 (N_3368,N_3300,N_3341);
nand U3369 (N_3369,N_3358,N_3253);
xor U3370 (N_3370,N_3338,N_3344);
or U3371 (N_3371,N_3275,N_3264);
nor U3372 (N_3372,N_3310,N_3346);
and U3373 (N_3373,N_3220,N_3209);
nor U3374 (N_3374,N_3352,N_3284);
or U3375 (N_3375,N_3208,N_3298);
and U3376 (N_3376,N_3315,N_3256);
or U3377 (N_3377,N_3299,N_3247);
nand U3378 (N_3378,N_3329,N_3309);
or U3379 (N_3379,N_3226,N_3211);
or U3380 (N_3380,N_3359,N_3322);
or U3381 (N_3381,N_3317,N_3339);
or U3382 (N_3382,N_3357,N_3356);
nor U3383 (N_3383,N_3304,N_3236);
nand U3384 (N_3384,N_3207,N_3290);
or U3385 (N_3385,N_3292,N_3244);
nand U3386 (N_3386,N_3326,N_3325);
or U3387 (N_3387,N_3276,N_3295);
and U3388 (N_3388,N_3333,N_3240);
and U3389 (N_3389,N_3319,N_3234);
nor U3390 (N_3390,N_3301,N_3331);
nor U3391 (N_3391,N_3206,N_3350);
nand U3392 (N_3392,N_3221,N_3243);
nand U3393 (N_3393,N_3296,N_3251);
or U3394 (N_3394,N_3213,N_3235);
nand U3395 (N_3395,N_3250,N_3216);
nor U3396 (N_3396,N_3308,N_3278);
nand U3397 (N_3397,N_3230,N_3205);
or U3398 (N_3398,N_3242,N_3316);
or U3399 (N_3399,N_3225,N_3268);
and U3400 (N_3400,N_3342,N_3215);
or U3401 (N_3401,N_3210,N_3238);
and U3402 (N_3402,N_3287,N_3291);
and U3403 (N_3403,N_3200,N_3265);
or U3404 (N_3404,N_3289,N_3281);
nor U3405 (N_3405,N_3202,N_3349);
nor U3406 (N_3406,N_3228,N_3262);
nor U3407 (N_3407,N_3285,N_3241);
nand U3408 (N_3408,N_3353,N_3320);
or U3409 (N_3409,N_3219,N_3231);
nor U3410 (N_3410,N_3201,N_3288);
and U3411 (N_3411,N_3269,N_3212);
nand U3412 (N_3412,N_3222,N_3233);
nand U3413 (N_3413,N_3214,N_3312);
nor U3414 (N_3414,N_3227,N_3283);
and U3415 (N_3415,N_3260,N_3245);
nor U3416 (N_3416,N_3330,N_3255);
or U3417 (N_3417,N_3335,N_3282);
or U3418 (N_3418,N_3248,N_3311);
nand U3419 (N_3419,N_3277,N_3223);
and U3420 (N_3420,N_3232,N_3318);
nand U3421 (N_3421,N_3286,N_3217);
nor U3422 (N_3422,N_3354,N_3259);
or U3423 (N_3423,N_3343,N_3261);
nor U3424 (N_3424,N_3258,N_3337);
and U3425 (N_3425,N_3249,N_3239);
or U3426 (N_3426,N_3340,N_3229);
or U3427 (N_3427,N_3355,N_3280);
or U3428 (N_3428,N_3345,N_3351);
or U3429 (N_3429,N_3321,N_3279);
nand U3430 (N_3430,N_3266,N_3257);
nand U3431 (N_3431,N_3348,N_3323);
and U3432 (N_3432,N_3263,N_3336);
and U3433 (N_3433,N_3218,N_3324);
nor U3434 (N_3434,N_3246,N_3303);
or U3435 (N_3435,N_3267,N_3302);
or U3436 (N_3436,N_3272,N_3273);
or U3437 (N_3437,N_3297,N_3293);
nand U3438 (N_3438,N_3313,N_3347);
nor U3439 (N_3439,N_3294,N_3314);
or U3440 (N_3440,N_3318,N_3252);
nor U3441 (N_3441,N_3312,N_3333);
nor U3442 (N_3442,N_3268,N_3284);
and U3443 (N_3443,N_3264,N_3287);
or U3444 (N_3444,N_3219,N_3319);
and U3445 (N_3445,N_3316,N_3275);
and U3446 (N_3446,N_3245,N_3331);
nor U3447 (N_3447,N_3257,N_3325);
and U3448 (N_3448,N_3306,N_3219);
or U3449 (N_3449,N_3241,N_3245);
or U3450 (N_3450,N_3315,N_3235);
xnor U3451 (N_3451,N_3336,N_3223);
or U3452 (N_3452,N_3357,N_3326);
nand U3453 (N_3453,N_3211,N_3252);
or U3454 (N_3454,N_3305,N_3233);
nor U3455 (N_3455,N_3343,N_3348);
and U3456 (N_3456,N_3271,N_3346);
nand U3457 (N_3457,N_3238,N_3258);
nor U3458 (N_3458,N_3228,N_3206);
nor U3459 (N_3459,N_3285,N_3354);
or U3460 (N_3460,N_3358,N_3279);
and U3461 (N_3461,N_3351,N_3320);
nor U3462 (N_3462,N_3300,N_3272);
and U3463 (N_3463,N_3344,N_3275);
nor U3464 (N_3464,N_3357,N_3253);
nor U3465 (N_3465,N_3246,N_3263);
and U3466 (N_3466,N_3231,N_3204);
nor U3467 (N_3467,N_3217,N_3220);
nor U3468 (N_3468,N_3316,N_3215);
or U3469 (N_3469,N_3215,N_3210);
nor U3470 (N_3470,N_3221,N_3230);
or U3471 (N_3471,N_3285,N_3263);
nand U3472 (N_3472,N_3229,N_3302);
nand U3473 (N_3473,N_3233,N_3272);
or U3474 (N_3474,N_3238,N_3242);
xor U3475 (N_3475,N_3248,N_3323);
nand U3476 (N_3476,N_3272,N_3248);
nor U3477 (N_3477,N_3279,N_3353);
and U3478 (N_3478,N_3286,N_3288);
and U3479 (N_3479,N_3349,N_3297);
nor U3480 (N_3480,N_3243,N_3323);
nor U3481 (N_3481,N_3300,N_3240);
and U3482 (N_3482,N_3307,N_3280);
nor U3483 (N_3483,N_3274,N_3333);
and U3484 (N_3484,N_3353,N_3357);
or U3485 (N_3485,N_3252,N_3228);
nor U3486 (N_3486,N_3215,N_3208);
xor U3487 (N_3487,N_3243,N_3319);
or U3488 (N_3488,N_3216,N_3315);
or U3489 (N_3489,N_3240,N_3202);
nor U3490 (N_3490,N_3217,N_3282);
and U3491 (N_3491,N_3323,N_3324);
nor U3492 (N_3492,N_3234,N_3353);
nor U3493 (N_3493,N_3318,N_3225);
or U3494 (N_3494,N_3290,N_3299);
nand U3495 (N_3495,N_3232,N_3297);
nor U3496 (N_3496,N_3308,N_3336);
and U3497 (N_3497,N_3357,N_3206);
nand U3498 (N_3498,N_3356,N_3231);
or U3499 (N_3499,N_3250,N_3264);
nor U3500 (N_3500,N_3226,N_3204);
nor U3501 (N_3501,N_3304,N_3311);
or U3502 (N_3502,N_3246,N_3220);
or U3503 (N_3503,N_3263,N_3226);
nor U3504 (N_3504,N_3218,N_3242);
xnor U3505 (N_3505,N_3336,N_3283);
or U3506 (N_3506,N_3283,N_3331);
or U3507 (N_3507,N_3256,N_3300);
nand U3508 (N_3508,N_3236,N_3273);
nor U3509 (N_3509,N_3305,N_3202);
nand U3510 (N_3510,N_3216,N_3203);
and U3511 (N_3511,N_3204,N_3217);
nor U3512 (N_3512,N_3228,N_3328);
nand U3513 (N_3513,N_3300,N_3235);
xnor U3514 (N_3514,N_3205,N_3268);
nor U3515 (N_3515,N_3265,N_3269);
xnor U3516 (N_3516,N_3224,N_3310);
nor U3517 (N_3517,N_3241,N_3350);
or U3518 (N_3518,N_3352,N_3323);
and U3519 (N_3519,N_3343,N_3245);
xnor U3520 (N_3520,N_3366,N_3468);
xnor U3521 (N_3521,N_3439,N_3399);
nor U3522 (N_3522,N_3404,N_3370);
xnor U3523 (N_3523,N_3482,N_3460);
nand U3524 (N_3524,N_3487,N_3475);
and U3525 (N_3525,N_3499,N_3381);
and U3526 (N_3526,N_3365,N_3422);
nand U3527 (N_3527,N_3377,N_3513);
or U3528 (N_3528,N_3379,N_3409);
or U3529 (N_3529,N_3497,N_3383);
nor U3530 (N_3530,N_3433,N_3481);
or U3531 (N_3531,N_3362,N_3466);
xor U3532 (N_3532,N_3503,N_3430);
and U3533 (N_3533,N_3413,N_3392);
and U3534 (N_3534,N_3411,N_3457);
and U3535 (N_3535,N_3375,N_3420);
and U3536 (N_3536,N_3469,N_3372);
nand U3537 (N_3537,N_3376,N_3495);
xnor U3538 (N_3538,N_3510,N_3516);
nor U3539 (N_3539,N_3398,N_3455);
nand U3540 (N_3540,N_3461,N_3435);
and U3541 (N_3541,N_3458,N_3502);
nand U3542 (N_3542,N_3432,N_3456);
or U3543 (N_3543,N_3416,N_3448);
and U3544 (N_3544,N_3427,N_3385);
nand U3545 (N_3545,N_3408,N_3401);
nor U3546 (N_3546,N_3443,N_3382);
and U3547 (N_3547,N_3489,N_3415);
and U3548 (N_3548,N_3424,N_3515);
nor U3549 (N_3549,N_3491,N_3445);
nor U3550 (N_3550,N_3373,N_3480);
nor U3551 (N_3551,N_3403,N_3467);
nor U3552 (N_3552,N_3418,N_3444);
or U3553 (N_3553,N_3454,N_3386);
nand U3554 (N_3554,N_3485,N_3407);
and U3555 (N_3555,N_3374,N_3384);
and U3556 (N_3556,N_3506,N_3395);
and U3557 (N_3557,N_3494,N_3446);
nor U3558 (N_3558,N_3423,N_3472);
nor U3559 (N_3559,N_3429,N_3517);
nor U3560 (N_3560,N_3447,N_3389);
nor U3561 (N_3561,N_3470,N_3406);
and U3562 (N_3562,N_3465,N_3371);
nand U3563 (N_3563,N_3512,N_3378);
nand U3564 (N_3564,N_3473,N_3390);
nand U3565 (N_3565,N_3361,N_3436);
or U3566 (N_3566,N_3471,N_3396);
and U3567 (N_3567,N_3501,N_3462);
or U3568 (N_3568,N_3486,N_3388);
nor U3569 (N_3569,N_3508,N_3360);
and U3570 (N_3570,N_3511,N_3449);
xor U3571 (N_3571,N_3414,N_3412);
or U3572 (N_3572,N_3405,N_3363);
nand U3573 (N_3573,N_3498,N_3410);
and U3574 (N_3574,N_3474,N_3477);
or U3575 (N_3575,N_3492,N_3391);
or U3576 (N_3576,N_3369,N_3426);
nand U3577 (N_3577,N_3507,N_3438);
or U3578 (N_3578,N_3402,N_3451);
or U3579 (N_3579,N_3514,N_3459);
and U3580 (N_3580,N_3478,N_3479);
nand U3581 (N_3581,N_3500,N_3450);
or U3582 (N_3582,N_3425,N_3434);
or U3583 (N_3583,N_3380,N_3476);
nor U3584 (N_3584,N_3397,N_3368);
nor U3585 (N_3585,N_3417,N_3463);
or U3586 (N_3586,N_3442,N_3483);
and U3587 (N_3587,N_3387,N_3519);
nand U3588 (N_3588,N_3509,N_3490);
xnor U3589 (N_3589,N_3504,N_3393);
xnor U3590 (N_3590,N_3394,N_3518);
nor U3591 (N_3591,N_3452,N_3428);
nand U3592 (N_3592,N_3367,N_3488);
or U3593 (N_3593,N_3421,N_3484);
nand U3594 (N_3594,N_3437,N_3419);
or U3595 (N_3595,N_3496,N_3505);
nand U3596 (N_3596,N_3364,N_3440);
or U3597 (N_3597,N_3400,N_3431);
and U3598 (N_3598,N_3493,N_3453);
nand U3599 (N_3599,N_3441,N_3464);
nand U3600 (N_3600,N_3409,N_3514);
nor U3601 (N_3601,N_3419,N_3447);
nand U3602 (N_3602,N_3467,N_3425);
and U3603 (N_3603,N_3407,N_3382);
or U3604 (N_3604,N_3379,N_3497);
nand U3605 (N_3605,N_3472,N_3463);
or U3606 (N_3606,N_3472,N_3467);
nand U3607 (N_3607,N_3468,N_3433);
nand U3608 (N_3608,N_3430,N_3373);
nor U3609 (N_3609,N_3447,N_3443);
or U3610 (N_3610,N_3372,N_3446);
nor U3611 (N_3611,N_3497,N_3470);
xor U3612 (N_3612,N_3403,N_3517);
nand U3613 (N_3613,N_3488,N_3364);
and U3614 (N_3614,N_3409,N_3495);
nor U3615 (N_3615,N_3368,N_3454);
or U3616 (N_3616,N_3386,N_3489);
and U3617 (N_3617,N_3500,N_3519);
nor U3618 (N_3618,N_3419,N_3441);
or U3619 (N_3619,N_3429,N_3421);
and U3620 (N_3620,N_3484,N_3496);
or U3621 (N_3621,N_3414,N_3381);
nor U3622 (N_3622,N_3504,N_3466);
nand U3623 (N_3623,N_3474,N_3368);
and U3624 (N_3624,N_3483,N_3439);
and U3625 (N_3625,N_3364,N_3490);
nand U3626 (N_3626,N_3406,N_3380);
nand U3627 (N_3627,N_3438,N_3479);
nor U3628 (N_3628,N_3479,N_3492);
nand U3629 (N_3629,N_3395,N_3364);
xor U3630 (N_3630,N_3517,N_3438);
or U3631 (N_3631,N_3371,N_3446);
nor U3632 (N_3632,N_3419,N_3507);
or U3633 (N_3633,N_3430,N_3511);
xnor U3634 (N_3634,N_3509,N_3371);
nor U3635 (N_3635,N_3488,N_3411);
and U3636 (N_3636,N_3436,N_3444);
or U3637 (N_3637,N_3384,N_3388);
and U3638 (N_3638,N_3451,N_3441);
or U3639 (N_3639,N_3446,N_3515);
nor U3640 (N_3640,N_3361,N_3386);
and U3641 (N_3641,N_3449,N_3484);
nor U3642 (N_3642,N_3443,N_3426);
and U3643 (N_3643,N_3503,N_3392);
nor U3644 (N_3644,N_3415,N_3446);
or U3645 (N_3645,N_3478,N_3510);
nand U3646 (N_3646,N_3388,N_3475);
xnor U3647 (N_3647,N_3403,N_3445);
nor U3648 (N_3648,N_3449,N_3442);
nor U3649 (N_3649,N_3368,N_3380);
and U3650 (N_3650,N_3407,N_3412);
xnor U3651 (N_3651,N_3370,N_3376);
or U3652 (N_3652,N_3391,N_3464);
and U3653 (N_3653,N_3429,N_3456);
or U3654 (N_3654,N_3421,N_3373);
and U3655 (N_3655,N_3396,N_3494);
or U3656 (N_3656,N_3441,N_3484);
and U3657 (N_3657,N_3436,N_3501);
nor U3658 (N_3658,N_3428,N_3369);
nand U3659 (N_3659,N_3480,N_3369);
or U3660 (N_3660,N_3509,N_3415);
or U3661 (N_3661,N_3501,N_3497);
and U3662 (N_3662,N_3473,N_3410);
nor U3663 (N_3663,N_3398,N_3364);
nor U3664 (N_3664,N_3396,N_3371);
nand U3665 (N_3665,N_3424,N_3361);
nor U3666 (N_3666,N_3448,N_3462);
or U3667 (N_3667,N_3461,N_3502);
and U3668 (N_3668,N_3462,N_3450);
nand U3669 (N_3669,N_3451,N_3480);
nand U3670 (N_3670,N_3446,N_3470);
or U3671 (N_3671,N_3487,N_3518);
nand U3672 (N_3672,N_3407,N_3370);
and U3673 (N_3673,N_3492,N_3503);
nand U3674 (N_3674,N_3427,N_3390);
nor U3675 (N_3675,N_3456,N_3464);
nand U3676 (N_3676,N_3415,N_3419);
nor U3677 (N_3677,N_3369,N_3401);
nor U3678 (N_3678,N_3437,N_3510);
nor U3679 (N_3679,N_3488,N_3368);
and U3680 (N_3680,N_3628,N_3551);
nor U3681 (N_3681,N_3544,N_3569);
or U3682 (N_3682,N_3658,N_3643);
and U3683 (N_3683,N_3588,N_3530);
and U3684 (N_3684,N_3629,N_3572);
or U3685 (N_3685,N_3574,N_3578);
or U3686 (N_3686,N_3669,N_3621);
nor U3687 (N_3687,N_3618,N_3631);
and U3688 (N_3688,N_3556,N_3600);
or U3689 (N_3689,N_3651,N_3577);
and U3690 (N_3690,N_3653,N_3533);
nor U3691 (N_3691,N_3585,N_3625);
xor U3692 (N_3692,N_3624,N_3555);
or U3693 (N_3693,N_3620,N_3584);
nand U3694 (N_3694,N_3564,N_3614);
xnor U3695 (N_3695,N_3520,N_3675);
nand U3696 (N_3696,N_3527,N_3666);
or U3697 (N_3697,N_3526,N_3659);
or U3698 (N_3698,N_3672,N_3667);
or U3699 (N_3699,N_3630,N_3525);
nor U3700 (N_3700,N_3674,N_3576);
nand U3701 (N_3701,N_3673,N_3586);
nand U3702 (N_3702,N_3655,N_3647);
xnor U3703 (N_3703,N_3677,N_3635);
nor U3704 (N_3704,N_3639,N_3590);
and U3705 (N_3705,N_3605,N_3622);
and U3706 (N_3706,N_3531,N_3549);
or U3707 (N_3707,N_3565,N_3594);
or U3708 (N_3708,N_3599,N_3552);
or U3709 (N_3709,N_3603,N_3521);
nor U3710 (N_3710,N_3613,N_3561);
nand U3711 (N_3711,N_3595,N_3636);
or U3712 (N_3712,N_3633,N_3676);
nor U3713 (N_3713,N_3529,N_3632);
nor U3714 (N_3714,N_3665,N_3601);
or U3715 (N_3715,N_3640,N_3654);
and U3716 (N_3716,N_3575,N_3604);
xnor U3717 (N_3717,N_3612,N_3587);
and U3718 (N_3718,N_3543,N_3634);
nand U3719 (N_3719,N_3656,N_3522);
nand U3720 (N_3720,N_3542,N_3583);
nand U3721 (N_3721,N_3679,N_3609);
nand U3722 (N_3722,N_3582,N_3663);
and U3723 (N_3723,N_3598,N_3539);
nand U3724 (N_3724,N_3596,N_3589);
and U3725 (N_3725,N_3626,N_3593);
nand U3726 (N_3726,N_3540,N_3608);
and U3727 (N_3727,N_3546,N_3617);
nand U3728 (N_3728,N_3645,N_3562);
or U3729 (N_3729,N_3662,N_3550);
nand U3730 (N_3730,N_3547,N_3528);
or U3731 (N_3731,N_3650,N_3568);
nor U3732 (N_3732,N_3623,N_3537);
nor U3733 (N_3733,N_3559,N_3670);
and U3734 (N_3734,N_3668,N_3616);
and U3735 (N_3735,N_3566,N_3592);
or U3736 (N_3736,N_3548,N_3638);
nor U3737 (N_3737,N_3597,N_3541);
nor U3738 (N_3738,N_3657,N_3567);
and U3739 (N_3739,N_3615,N_3563);
nand U3740 (N_3740,N_3602,N_3571);
nand U3741 (N_3741,N_3523,N_3660);
nand U3742 (N_3742,N_3606,N_3580);
xor U3743 (N_3743,N_3535,N_3536);
nor U3744 (N_3744,N_3553,N_3671);
or U3745 (N_3745,N_3644,N_3532);
nor U3746 (N_3746,N_3678,N_3664);
nand U3747 (N_3747,N_3641,N_3538);
nand U3748 (N_3748,N_3579,N_3649);
xnor U3749 (N_3749,N_3619,N_3557);
and U3750 (N_3750,N_3610,N_3534);
xnor U3751 (N_3751,N_3570,N_3607);
or U3752 (N_3752,N_3646,N_3611);
or U3753 (N_3753,N_3554,N_3573);
xor U3754 (N_3754,N_3524,N_3642);
or U3755 (N_3755,N_3545,N_3652);
and U3756 (N_3756,N_3627,N_3581);
or U3757 (N_3757,N_3637,N_3560);
nand U3758 (N_3758,N_3591,N_3648);
and U3759 (N_3759,N_3661,N_3558);
or U3760 (N_3760,N_3549,N_3554);
nor U3761 (N_3761,N_3612,N_3557);
and U3762 (N_3762,N_3587,N_3647);
xnor U3763 (N_3763,N_3536,N_3582);
and U3764 (N_3764,N_3679,N_3600);
and U3765 (N_3765,N_3550,N_3577);
or U3766 (N_3766,N_3628,N_3670);
nand U3767 (N_3767,N_3529,N_3588);
nand U3768 (N_3768,N_3565,N_3577);
or U3769 (N_3769,N_3641,N_3622);
nand U3770 (N_3770,N_3577,N_3618);
and U3771 (N_3771,N_3634,N_3597);
nand U3772 (N_3772,N_3659,N_3523);
xor U3773 (N_3773,N_3569,N_3597);
and U3774 (N_3774,N_3652,N_3618);
nor U3775 (N_3775,N_3544,N_3639);
and U3776 (N_3776,N_3558,N_3621);
and U3777 (N_3777,N_3639,N_3670);
nand U3778 (N_3778,N_3612,N_3558);
nand U3779 (N_3779,N_3637,N_3613);
nand U3780 (N_3780,N_3614,N_3678);
or U3781 (N_3781,N_3552,N_3656);
and U3782 (N_3782,N_3547,N_3668);
or U3783 (N_3783,N_3564,N_3583);
nand U3784 (N_3784,N_3569,N_3537);
and U3785 (N_3785,N_3574,N_3615);
xnor U3786 (N_3786,N_3663,N_3579);
nor U3787 (N_3787,N_3624,N_3549);
nand U3788 (N_3788,N_3615,N_3677);
and U3789 (N_3789,N_3520,N_3525);
nor U3790 (N_3790,N_3565,N_3656);
nand U3791 (N_3791,N_3647,N_3546);
nor U3792 (N_3792,N_3560,N_3617);
nand U3793 (N_3793,N_3592,N_3651);
or U3794 (N_3794,N_3673,N_3601);
nor U3795 (N_3795,N_3590,N_3592);
nor U3796 (N_3796,N_3551,N_3605);
and U3797 (N_3797,N_3634,N_3568);
or U3798 (N_3798,N_3674,N_3540);
nor U3799 (N_3799,N_3643,N_3674);
and U3800 (N_3800,N_3648,N_3629);
nor U3801 (N_3801,N_3659,N_3576);
nand U3802 (N_3802,N_3665,N_3630);
nor U3803 (N_3803,N_3580,N_3609);
or U3804 (N_3804,N_3619,N_3520);
or U3805 (N_3805,N_3573,N_3612);
or U3806 (N_3806,N_3614,N_3578);
and U3807 (N_3807,N_3661,N_3601);
or U3808 (N_3808,N_3627,N_3666);
or U3809 (N_3809,N_3670,N_3658);
nand U3810 (N_3810,N_3558,N_3576);
nand U3811 (N_3811,N_3554,N_3634);
or U3812 (N_3812,N_3561,N_3586);
or U3813 (N_3813,N_3632,N_3586);
nand U3814 (N_3814,N_3582,N_3524);
nor U3815 (N_3815,N_3656,N_3661);
or U3816 (N_3816,N_3566,N_3602);
xor U3817 (N_3817,N_3663,N_3608);
nor U3818 (N_3818,N_3614,N_3532);
nor U3819 (N_3819,N_3540,N_3631);
nand U3820 (N_3820,N_3539,N_3571);
nand U3821 (N_3821,N_3582,N_3629);
and U3822 (N_3822,N_3642,N_3567);
and U3823 (N_3823,N_3656,N_3531);
and U3824 (N_3824,N_3603,N_3677);
nor U3825 (N_3825,N_3672,N_3552);
or U3826 (N_3826,N_3648,N_3524);
nand U3827 (N_3827,N_3528,N_3623);
nand U3828 (N_3828,N_3642,N_3544);
xor U3829 (N_3829,N_3615,N_3592);
and U3830 (N_3830,N_3667,N_3550);
or U3831 (N_3831,N_3656,N_3629);
and U3832 (N_3832,N_3536,N_3576);
nor U3833 (N_3833,N_3641,N_3596);
nor U3834 (N_3834,N_3552,N_3579);
nor U3835 (N_3835,N_3591,N_3601);
xnor U3836 (N_3836,N_3548,N_3602);
or U3837 (N_3837,N_3550,N_3554);
and U3838 (N_3838,N_3544,N_3529);
nand U3839 (N_3839,N_3614,N_3548);
or U3840 (N_3840,N_3749,N_3702);
or U3841 (N_3841,N_3698,N_3808);
and U3842 (N_3842,N_3828,N_3807);
or U3843 (N_3843,N_3786,N_3696);
nor U3844 (N_3844,N_3690,N_3779);
or U3845 (N_3845,N_3689,N_3726);
nand U3846 (N_3846,N_3734,N_3716);
nor U3847 (N_3847,N_3760,N_3789);
or U3848 (N_3848,N_3816,N_3839);
or U3849 (N_3849,N_3705,N_3692);
or U3850 (N_3850,N_3806,N_3835);
nor U3851 (N_3851,N_3811,N_3742);
or U3852 (N_3852,N_3833,N_3803);
or U3853 (N_3853,N_3836,N_3761);
nand U3854 (N_3854,N_3715,N_3737);
xor U3855 (N_3855,N_3682,N_3691);
or U3856 (N_3856,N_3683,N_3824);
or U3857 (N_3857,N_3809,N_3699);
nand U3858 (N_3858,N_3798,N_3838);
and U3859 (N_3859,N_3722,N_3815);
nor U3860 (N_3860,N_3713,N_3754);
or U3861 (N_3861,N_3810,N_3800);
xnor U3862 (N_3862,N_3762,N_3746);
nand U3863 (N_3863,N_3733,N_3738);
nand U3864 (N_3864,N_3687,N_3684);
or U3865 (N_3865,N_3729,N_3744);
nand U3866 (N_3866,N_3755,N_3708);
nor U3867 (N_3867,N_3688,N_3748);
or U3868 (N_3868,N_3701,N_3757);
nand U3869 (N_3869,N_3785,N_3750);
nand U3870 (N_3870,N_3720,N_3730);
or U3871 (N_3871,N_3700,N_3751);
nor U3872 (N_3872,N_3685,N_3743);
nand U3873 (N_3873,N_3718,N_3818);
nor U3874 (N_3874,N_3741,N_3707);
nand U3875 (N_3875,N_3790,N_3776);
and U3876 (N_3876,N_3782,N_3686);
nor U3877 (N_3877,N_3728,N_3739);
nor U3878 (N_3878,N_3765,N_3788);
xor U3879 (N_3879,N_3825,N_3680);
and U3880 (N_3880,N_3768,N_3723);
and U3881 (N_3881,N_3781,N_3740);
nand U3882 (N_3882,N_3832,N_3759);
nand U3883 (N_3883,N_3766,N_3802);
or U3884 (N_3884,N_3819,N_3717);
nand U3885 (N_3885,N_3693,N_3732);
nand U3886 (N_3886,N_3709,N_3780);
and U3887 (N_3887,N_3787,N_3719);
and U3888 (N_3888,N_3796,N_3783);
nor U3889 (N_3889,N_3771,N_3710);
xnor U3890 (N_3890,N_3794,N_3764);
nor U3891 (N_3891,N_3821,N_3801);
and U3892 (N_3892,N_3727,N_3822);
xnor U3893 (N_3893,N_3704,N_3777);
nand U3894 (N_3894,N_3797,N_3736);
or U3895 (N_3895,N_3775,N_3712);
or U3896 (N_3896,N_3770,N_3745);
nor U3897 (N_3897,N_3804,N_3694);
nand U3898 (N_3898,N_3747,N_3817);
or U3899 (N_3899,N_3697,N_3774);
and U3900 (N_3900,N_3826,N_3725);
and U3901 (N_3901,N_3731,N_3772);
xnor U3902 (N_3902,N_3756,N_3778);
or U3903 (N_3903,N_3753,N_3711);
nand U3904 (N_3904,N_3831,N_3805);
nor U3905 (N_3905,N_3829,N_3791);
or U3906 (N_3906,N_3763,N_3767);
nand U3907 (N_3907,N_3758,N_3752);
and U3908 (N_3908,N_3834,N_3721);
nor U3909 (N_3909,N_3820,N_3814);
or U3910 (N_3910,N_3681,N_3795);
and U3911 (N_3911,N_3724,N_3837);
or U3912 (N_3912,N_3703,N_3784);
and U3913 (N_3913,N_3827,N_3714);
or U3914 (N_3914,N_3773,N_3793);
and U3915 (N_3915,N_3823,N_3706);
xor U3916 (N_3916,N_3695,N_3813);
and U3917 (N_3917,N_3799,N_3812);
nand U3918 (N_3918,N_3830,N_3792);
nor U3919 (N_3919,N_3769,N_3735);
or U3920 (N_3920,N_3804,N_3749);
nor U3921 (N_3921,N_3759,N_3779);
nand U3922 (N_3922,N_3799,N_3803);
nor U3923 (N_3923,N_3777,N_3710);
nor U3924 (N_3924,N_3759,N_3801);
or U3925 (N_3925,N_3753,N_3757);
nand U3926 (N_3926,N_3697,N_3732);
nor U3927 (N_3927,N_3789,N_3764);
nor U3928 (N_3928,N_3811,N_3683);
nand U3929 (N_3929,N_3753,N_3803);
nor U3930 (N_3930,N_3733,N_3705);
or U3931 (N_3931,N_3778,N_3774);
and U3932 (N_3932,N_3801,N_3707);
or U3933 (N_3933,N_3832,N_3806);
nor U3934 (N_3934,N_3786,N_3699);
nor U3935 (N_3935,N_3831,N_3685);
nor U3936 (N_3936,N_3706,N_3824);
nor U3937 (N_3937,N_3796,N_3682);
nor U3938 (N_3938,N_3709,N_3830);
or U3939 (N_3939,N_3773,N_3806);
or U3940 (N_3940,N_3723,N_3721);
nand U3941 (N_3941,N_3792,N_3816);
and U3942 (N_3942,N_3769,N_3767);
and U3943 (N_3943,N_3816,N_3743);
nor U3944 (N_3944,N_3806,N_3767);
nor U3945 (N_3945,N_3821,N_3720);
nor U3946 (N_3946,N_3779,N_3793);
or U3947 (N_3947,N_3753,N_3696);
or U3948 (N_3948,N_3692,N_3814);
nor U3949 (N_3949,N_3764,N_3791);
xnor U3950 (N_3950,N_3730,N_3700);
nor U3951 (N_3951,N_3818,N_3782);
and U3952 (N_3952,N_3737,N_3780);
and U3953 (N_3953,N_3817,N_3728);
xor U3954 (N_3954,N_3778,N_3808);
nor U3955 (N_3955,N_3762,N_3788);
and U3956 (N_3956,N_3812,N_3736);
or U3957 (N_3957,N_3805,N_3694);
and U3958 (N_3958,N_3752,N_3708);
or U3959 (N_3959,N_3732,N_3775);
or U3960 (N_3960,N_3812,N_3711);
nor U3961 (N_3961,N_3783,N_3738);
or U3962 (N_3962,N_3687,N_3809);
nor U3963 (N_3963,N_3682,N_3760);
and U3964 (N_3964,N_3686,N_3803);
nor U3965 (N_3965,N_3777,N_3828);
and U3966 (N_3966,N_3685,N_3748);
or U3967 (N_3967,N_3704,N_3727);
and U3968 (N_3968,N_3833,N_3784);
xor U3969 (N_3969,N_3809,N_3765);
nand U3970 (N_3970,N_3757,N_3702);
nand U3971 (N_3971,N_3801,N_3766);
and U3972 (N_3972,N_3785,N_3691);
or U3973 (N_3973,N_3768,N_3698);
nor U3974 (N_3974,N_3803,N_3781);
and U3975 (N_3975,N_3712,N_3694);
nand U3976 (N_3976,N_3790,N_3732);
nand U3977 (N_3977,N_3728,N_3787);
nand U3978 (N_3978,N_3724,N_3801);
nand U3979 (N_3979,N_3780,N_3770);
or U3980 (N_3980,N_3778,N_3760);
nor U3981 (N_3981,N_3743,N_3692);
and U3982 (N_3982,N_3695,N_3772);
or U3983 (N_3983,N_3809,N_3744);
nand U3984 (N_3984,N_3745,N_3787);
and U3985 (N_3985,N_3829,N_3777);
nand U3986 (N_3986,N_3819,N_3714);
xor U3987 (N_3987,N_3829,N_3794);
and U3988 (N_3988,N_3819,N_3716);
or U3989 (N_3989,N_3819,N_3793);
nand U3990 (N_3990,N_3797,N_3809);
or U3991 (N_3991,N_3835,N_3802);
and U3992 (N_3992,N_3765,N_3818);
xor U3993 (N_3993,N_3797,N_3830);
nand U3994 (N_3994,N_3693,N_3703);
xor U3995 (N_3995,N_3792,N_3798);
nand U3996 (N_3996,N_3767,N_3832);
and U3997 (N_3997,N_3717,N_3708);
and U3998 (N_3998,N_3767,N_3745);
and U3999 (N_3999,N_3701,N_3792);
and U4000 (N_4000,N_3902,N_3864);
nor U4001 (N_4001,N_3844,N_3867);
nor U4002 (N_4002,N_3956,N_3976);
xnor U4003 (N_4003,N_3905,N_3887);
xnor U4004 (N_4004,N_3999,N_3873);
and U4005 (N_4005,N_3960,N_3889);
or U4006 (N_4006,N_3950,N_3896);
or U4007 (N_4007,N_3935,N_3962);
nor U4008 (N_4008,N_3880,N_3953);
nor U4009 (N_4009,N_3847,N_3933);
nor U4010 (N_4010,N_3906,N_3983);
xor U4011 (N_4011,N_3884,N_3897);
nor U4012 (N_4012,N_3938,N_3927);
or U4013 (N_4013,N_3920,N_3946);
xor U4014 (N_4014,N_3911,N_3908);
nor U4015 (N_4015,N_3975,N_3947);
nor U4016 (N_4016,N_3865,N_3972);
and U4017 (N_4017,N_3890,N_3858);
nand U4018 (N_4018,N_3932,N_3915);
nor U4019 (N_4019,N_3845,N_3919);
and U4020 (N_4020,N_3878,N_3941);
and U4021 (N_4021,N_3944,N_3912);
or U4022 (N_4022,N_3883,N_3863);
and U4023 (N_4023,N_3969,N_3978);
and U4024 (N_4024,N_3990,N_3886);
and U4025 (N_4025,N_3917,N_3965);
nor U4026 (N_4026,N_3988,N_3846);
and U4027 (N_4027,N_3954,N_3955);
nor U4028 (N_4028,N_3870,N_3854);
and U4029 (N_4029,N_3925,N_3931);
nand U4030 (N_4030,N_3849,N_3980);
or U4031 (N_4031,N_3848,N_3952);
or U4032 (N_4032,N_3986,N_3868);
and U4033 (N_4033,N_3945,N_3852);
and U4034 (N_4034,N_3910,N_3898);
or U4035 (N_4035,N_3872,N_3977);
nor U4036 (N_4036,N_3966,N_3918);
nand U4037 (N_4037,N_3979,N_3851);
nor U4038 (N_4038,N_3984,N_3885);
nand U4039 (N_4039,N_3940,N_3923);
nand U4040 (N_4040,N_3840,N_3951);
or U4041 (N_4041,N_3894,N_3996);
nand U4042 (N_4042,N_3866,N_3862);
or U4043 (N_4043,N_3929,N_3892);
or U4044 (N_4044,N_3998,N_3921);
nor U4045 (N_4045,N_3963,N_3850);
nor U4046 (N_4046,N_3959,N_3971);
or U4047 (N_4047,N_3991,N_3958);
and U4048 (N_4048,N_3900,N_3993);
and U4049 (N_4049,N_3857,N_3895);
nand U4050 (N_4050,N_3877,N_3882);
nor U4051 (N_4051,N_3869,N_3974);
or U4052 (N_4052,N_3874,N_3871);
nand U4053 (N_4053,N_3994,N_3859);
nor U4054 (N_4054,N_3914,N_3891);
nand U4055 (N_4055,N_3843,N_3893);
nor U4056 (N_4056,N_3875,N_3888);
or U4057 (N_4057,N_3937,N_3841);
nand U4058 (N_4058,N_3997,N_3970);
and U4059 (N_4059,N_3899,N_3936);
and U4060 (N_4060,N_3992,N_3855);
nor U4061 (N_4061,N_3995,N_3907);
or U4062 (N_4062,N_3973,N_3982);
and U4063 (N_4063,N_3948,N_3987);
or U4064 (N_4064,N_3957,N_3881);
or U4065 (N_4065,N_3903,N_3961);
and U4066 (N_4066,N_3964,N_3860);
nor U4067 (N_4067,N_3876,N_3926);
nor U4068 (N_4068,N_3942,N_3981);
and U4069 (N_4069,N_3913,N_3904);
nor U4070 (N_4070,N_3901,N_3967);
or U4071 (N_4071,N_3924,N_3856);
and U4072 (N_4072,N_3943,N_3879);
or U4073 (N_4073,N_3842,N_3909);
nor U4074 (N_4074,N_3939,N_3985);
and U4075 (N_4075,N_3916,N_3861);
nand U4076 (N_4076,N_3928,N_3989);
xor U4077 (N_4077,N_3853,N_3968);
and U4078 (N_4078,N_3949,N_3930);
nand U4079 (N_4079,N_3922,N_3934);
nand U4080 (N_4080,N_3928,N_3869);
or U4081 (N_4081,N_3921,N_3915);
nand U4082 (N_4082,N_3940,N_3902);
xnor U4083 (N_4083,N_3977,N_3940);
nor U4084 (N_4084,N_3869,N_3921);
and U4085 (N_4085,N_3884,N_3996);
nor U4086 (N_4086,N_3863,N_3874);
or U4087 (N_4087,N_3848,N_3999);
nand U4088 (N_4088,N_3982,N_3862);
or U4089 (N_4089,N_3891,N_3937);
and U4090 (N_4090,N_3913,N_3978);
and U4091 (N_4091,N_3881,N_3899);
xor U4092 (N_4092,N_3940,N_3945);
nand U4093 (N_4093,N_3969,N_3872);
nor U4094 (N_4094,N_3923,N_3884);
nor U4095 (N_4095,N_3980,N_3982);
nand U4096 (N_4096,N_3923,N_3967);
and U4097 (N_4097,N_3972,N_3869);
or U4098 (N_4098,N_3907,N_3872);
xor U4099 (N_4099,N_3924,N_3889);
and U4100 (N_4100,N_3914,N_3893);
and U4101 (N_4101,N_3902,N_3974);
or U4102 (N_4102,N_3996,N_3842);
or U4103 (N_4103,N_3887,N_3912);
xor U4104 (N_4104,N_3920,N_3919);
nor U4105 (N_4105,N_3853,N_3925);
and U4106 (N_4106,N_3967,N_3915);
nor U4107 (N_4107,N_3893,N_3989);
nand U4108 (N_4108,N_3964,N_3864);
and U4109 (N_4109,N_3898,N_3872);
xnor U4110 (N_4110,N_3886,N_3927);
and U4111 (N_4111,N_3883,N_3912);
nor U4112 (N_4112,N_3964,N_3859);
and U4113 (N_4113,N_3872,N_3928);
or U4114 (N_4114,N_3936,N_3883);
xnor U4115 (N_4115,N_3909,N_3902);
or U4116 (N_4116,N_3930,N_3887);
and U4117 (N_4117,N_3977,N_3996);
and U4118 (N_4118,N_3907,N_3876);
nand U4119 (N_4119,N_3939,N_3872);
or U4120 (N_4120,N_3884,N_3911);
nand U4121 (N_4121,N_3993,N_3947);
and U4122 (N_4122,N_3871,N_3990);
xnor U4123 (N_4123,N_3910,N_3925);
or U4124 (N_4124,N_3844,N_3866);
nor U4125 (N_4125,N_3969,N_3995);
nand U4126 (N_4126,N_3982,N_3875);
nand U4127 (N_4127,N_3911,N_3936);
nand U4128 (N_4128,N_3894,N_3955);
xor U4129 (N_4129,N_3948,N_3933);
nand U4130 (N_4130,N_3852,N_3966);
or U4131 (N_4131,N_3898,N_3926);
nand U4132 (N_4132,N_3863,N_3992);
nor U4133 (N_4133,N_3910,N_3878);
nand U4134 (N_4134,N_3964,N_3900);
xor U4135 (N_4135,N_3878,N_3942);
or U4136 (N_4136,N_3913,N_3950);
or U4137 (N_4137,N_3920,N_3943);
and U4138 (N_4138,N_3914,N_3850);
and U4139 (N_4139,N_3872,N_3998);
and U4140 (N_4140,N_3961,N_3925);
nand U4141 (N_4141,N_3906,N_3878);
and U4142 (N_4142,N_3987,N_3978);
nor U4143 (N_4143,N_3943,N_3923);
and U4144 (N_4144,N_3867,N_3862);
and U4145 (N_4145,N_3916,N_3889);
or U4146 (N_4146,N_3989,N_3977);
or U4147 (N_4147,N_3918,N_3950);
xnor U4148 (N_4148,N_3887,N_3894);
xnor U4149 (N_4149,N_3940,N_3850);
or U4150 (N_4150,N_3911,N_3938);
nand U4151 (N_4151,N_3859,N_3904);
nor U4152 (N_4152,N_3984,N_3895);
nor U4153 (N_4153,N_3942,N_3921);
and U4154 (N_4154,N_3982,N_3848);
and U4155 (N_4155,N_3971,N_3872);
nor U4156 (N_4156,N_3841,N_3973);
nor U4157 (N_4157,N_3897,N_3860);
or U4158 (N_4158,N_3916,N_3994);
nand U4159 (N_4159,N_3952,N_3898);
and U4160 (N_4160,N_4008,N_4122);
nor U4161 (N_4161,N_4010,N_4106);
xor U4162 (N_4162,N_4094,N_4139);
or U4163 (N_4163,N_4079,N_4136);
and U4164 (N_4164,N_4001,N_4054);
xor U4165 (N_4165,N_4044,N_4086);
or U4166 (N_4166,N_4115,N_4154);
nor U4167 (N_4167,N_4032,N_4016);
or U4168 (N_4168,N_4133,N_4064);
or U4169 (N_4169,N_4142,N_4149);
nor U4170 (N_4170,N_4029,N_4098);
or U4171 (N_4171,N_4150,N_4063);
nand U4172 (N_4172,N_4125,N_4124);
or U4173 (N_4173,N_4073,N_4112);
and U4174 (N_4174,N_4104,N_4030);
or U4175 (N_4175,N_4121,N_4126);
and U4176 (N_4176,N_4083,N_4041);
nor U4177 (N_4177,N_4092,N_4002);
and U4178 (N_4178,N_4039,N_4075);
and U4179 (N_4179,N_4143,N_4036);
or U4180 (N_4180,N_4009,N_4020);
and U4181 (N_4181,N_4153,N_4105);
nor U4182 (N_4182,N_4060,N_4110);
or U4183 (N_4183,N_4082,N_4091);
nor U4184 (N_4184,N_4006,N_4151);
nand U4185 (N_4185,N_4021,N_4061);
nor U4186 (N_4186,N_4102,N_4103);
and U4187 (N_4187,N_4088,N_4107);
or U4188 (N_4188,N_4037,N_4113);
nand U4189 (N_4189,N_4156,N_4062);
xor U4190 (N_4190,N_4051,N_4146);
or U4191 (N_4191,N_4065,N_4159);
xor U4192 (N_4192,N_4132,N_4134);
nand U4193 (N_4193,N_4117,N_4093);
or U4194 (N_4194,N_4024,N_4127);
nor U4195 (N_4195,N_4089,N_4128);
xnor U4196 (N_4196,N_4074,N_4042);
or U4197 (N_4197,N_4111,N_4097);
nand U4198 (N_4198,N_4071,N_4043);
xnor U4199 (N_4199,N_4022,N_4019);
xor U4200 (N_4200,N_4057,N_4116);
or U4201 (N_4201,N_4095,N_4040);
and U4202 (N_4202,N_4090,N_4144);
or U4203 (N_4203,N_4080,N_4109);
nor U4204 (N_4204,N_4017,N_4048);
or U4205 (N_4205,N_4026,N_4081);
nor U4206 (N_4206,N_4015,N_4027);
nand U4207 (N_4207,N_4101,N_4078);
or U4208 (N_4208,N_4119,N_4035);
and U4209 (N_4209,N_4011,N_4049);
xnor U4210 (N_4210,N_4157,N_4077);
xnor U4211 (N_4211,N_4158,N_4047);
xor U4212 (N_4212,N_4031,N_4155);
nand U4213 (N_4213,N_4003,N_4145);
and U4214 (N_4214,N_4123,N_4033);
nor U4215 (N_4215,N_4038,N_4005);
xnor U4216 (N_4216,N_4058,N_4137);
nor U4217 (N_4217,N_4076,N_4135);
and U4218 (N_4218,N_4100,N_4068);
or U4219 (N_4219,N_4007,N_4000);
or U4220 (N_4220,N_4152,N_4053);
nor U4221 (N_4221,N_4072,N_4023);
nand U4222 (N_4222,N_4070,N_4130);
nand U4223 (N_4223,N_4014,N_4056);
and U4224 (N_4224,N_4025,N_4087);
or U4225 (N_4225,N_4069,N_4066);
xor U4226 (N_4226,N_4129,N_4059);
nand U4227 (N_4227,N_4084,N_4138);
or U4228 (N_4228,N_4114,N_4067);
and U4229 (N_4229,N_4096,N_4028);
and U4230 (N_4230,N_4131,N_4050);
nor U4231 (N_4231,N_4141,N_4120);
and U4232 (N_4232,N_4140,N_4055);
nand U4233 (N_4233,N_4118,N_4148);
nand U4234 (N_4234,N_4099,N_4034);
xor U4235 (N_4235,N_4004,N_4052);
nand U4236 (N_4236,N_4012,N_4085);
and U4237 (N_4237,N_4045,N_4108);
and U4238 (N_4238,N_4018,N_4147);
nand U4239 (N_4239,N_4046,N_4013);
nor U4240 (N_4240,N_4096,N_4072);
or U4241 (N_4241,N_4010,N_4144);
nor U4242 (N_4242,N_4124,N_4153);
and U4243 (N_4243,N_4121,N_4065);
and U4244 (N_4244,N_4103,N_4001);
nor U4245 (N_4245,N_4139,N_4061);
or U4246 (N_4246,N_4077,N_4158);
or U4247 (N_4247,N_4117,N_4054);
and U4248 (N_4248,N_4059,N_4134);
nand U4249 (N_4249,N_4094,N_4136);
nor U4250 (N_4250,N_4033,N_4109);
nor U4251 (N_4251,N_4126,N_4020);
and U4252 (N_4252,N_4148,N_4123);
and U4253 (N_4253,N_4028,N_4112);
nand U4254 (N_4254,N_4045,N_4003);
or U4255 (N_4255,N_4013,N_4132);
nand U4256 (N_4256,N_4028,N_4023);
and U4257 (N_4257,N_4100,N_4039);
nor U4258 (N_4258,N_4004,N_4159);
nand U4259 (N_4259,N_4014,N_4002);
nand U4260 (N_4260,N_4148,N_4018);
and U4261 (N_4261,N_4102,N_4138);
nor U4262 (N_4262,N_4063,N_4018);
and U4263 (N_4263,N_4157,N_4112);
and U4264 (N_4264,N_4070,N_4107);
or U4265 (N_4265,N_4057,N_4003);
or U4266 (N_4266,N_4081,N_4052);
xnor U4267 (N_4267,N_4037,N_4007);
or U4268 (N_4268,N_4076,N_4019);
and U4269 (N_4269,N_4034,N_4070);
and U4270 (N_4270,N_4157,N_4151);
nor U4271 (N_4271,N_4073,N_4096);
nor U4272 (N_4272,N_4043,N_4047);
xor U4273 (N_4273,N_4106,N_4003);
nand U4274 (N_4274,N_4098,N_4009);
nand U4275 (N_4275,N_4062,N_4113);
nand U4276 (N_4276,N_4089,N_4131);
nand U4277 (N_4277,N_4053,N_4069);
nand U4278 (N_4278,N_4096,N_4131);
and U4279 (N_4279,N_4035,N_4021);
or U4280 (N_4280,N_4058,N_4136);
nor U4281 (N_4281,N_4082,N_4019);
nand U4282 (N_4282,N_4015,N_4053);
nor U4283 (N_4283,N_4026,N_4157);
nand U4284 (N_4284,N_4071,N_4045);
nand U4285 (N_4285,N_4037,N_4060);
and U4286 (N_4286,N_4116,N_4110);
nand U4287 (N_4287,N_4140,N_4013);
nand U4288 (N_4288,N_4158,N_4003);
nand U4289 (N_4289,N_4022,N_4066);
and U4290 (N_4290,N_4062,N_4080);
nor U4291 (N_4291,N_4027,N_4066);
nor U4292 (N_4292,N_4085,N_4013);
or U4293 (N_4293,N_4108,N_4031);
and U4294 (N_4294,N_4077,N_4054);
nor U4295 (N_4295,N_4027,N_4070);
nand U4296 (N_4296,N_4006,N_4114);
or U4297 (N_4297,N_4119,N_4112);
and U4298 (N_4298,N_4059,N_4067);
or U4299 (N_4299,N_4062,N_4142);
and U4300 (N_4300,N_4082,N_4065);
and U4301 (N_4301,N_4026,N_4086);
nor U4302 (N_4302,N_4096,N_4141);
nor U4303 (N_4303,N_4115,N_4152);
nand U4304 (N_4304,N_4013,N_4122);
nor U4305 (N_4305,N_4037,N_4140);
nor U4306 (N_4306,N_4140,N_4002);
and U4307 (N_4307,N_4149,N_4020);
nand U4308 (N_4308,N_4015,N_4119);
nor U4309 (N_4309,N_4056,N_4127);
xnor U4310 (N_4310,N_4074,N_4113);
and U4311 (N_4311,N_4010,N_4035);
and U4312 (N_4312,N_4127,N_4081);
or U4313 (N_4313,N_4153,N_4051);
nor U4314 (N_4314,N_4077,N_4022);
and U4315 (N_4315,N_4003,N_4026);
nor U4316 (N_4316,N_4051,N_4052);
nand U4317 (N_4317,N_4029,N_4000);
or U4318 (N_4318,N_4092,N_4143);
and U4319 (N_4319,N_4080,N_4145);
and U4320 (N_4320,N_4299,N_4208);
or U4321 (N_4321,N_4249,N_4238);
and U4322 (N_4322,N_4293,N_4167);
nor U4323 (N_4323,N_4224,N_4211);
or U4324 (N_4324,N_4185,N_4162);
or U4325 (N_4325,N_4285,N_4172);
or U4326 (N_4326,N_4188,N_4281);
nor U4327 (N_4327,N_4182,N_4246);
and U4328 (N_4328,N_4264,N_4221);
nand U4329 (N_4329,N_4222,N_4244);
nand U4330 (N_4330,N_4260,N_4165);
or U4331 (N_4331,N_4181,N_4289);
nand U4332 (N_4332,N_4287,N_4234);
or U4333 (N_4333,N_4207,N_4252);
nand U4334 (N_4334,N_4161,N_4272);
or U4335 (N_4335,N_4312,N_4227);
nor U4336 (N_4336,N_4197,N_4242);
xnor U4337 (N_4337,N_4219,N_4191);
nor U4338 (N_4338,N_4163,N_4291);
or U4339 (N_4339,N_4267,N_4300);
nor U4340 (N_4340,N_4269,N_4239);
and U4341 (N_4341,N_4253,N_4236);
or U4342 (N_4342,N_4228,N_4195);
or U4343 (N_4343,N_4308,N_4218);
nor U4344 (N_4344,N_4261,N_4307);
nor U4345 (N_4345,N_4213,N_4317);
nand U4346 (N_4346,N_4266,N_4316);
and U4347 (N_4347,N_4235,N_4212);
nand U4348 (N_4348,N_4231,N_4202);
nor U4349 (N_4349,N_4171,N_4262);
or U4350 (N_4350,N_4205,N_4256);
and U4351 (N_4351,N_4318,N_4278);
or U4352 (N_4352,N_4210,N_4192);
or U4353 (N_4353,N_4174,N_4319);
or U4354 (N_4354,N_4232,N_4241);
and U4355 (N_4355,N_4288,N_4305);
nand U4356 (N_4356,N_4180,N_4279);
xor U4357 (N_4357,N_4311,N_4255);
or U4358 (N_4358,N_4226,N_4200);
nor U4359 (N_4359,N_4290,N_4280);
and U4360 (N_4360,N_4247,N_4284);
nor U4361 (N_4361,N_4168,N_4215);
nand U4362 (N_4362,N_4304,N_4250);
xor U4363 (N_4363,N_4303,N_4230);
or U4364 (N_4364,N_4190,N_4177);
or U4365 (N_4365,N_4240,N_4298);
and U4366 (N_4366,N_4187,N_4251);
nor U4367 (N_4367,N_4173,N_4265);
nand U4368 (N_4368,N_4229,N_4223);
and U4369 (N_4369,N_4274,N_4237);
nor U4370 (N_4370,N_4166,N_4292);
or U4371 (N_4371,N_4286,N_4270);
nand U4372 (N_4372,N_4282,N_4214);
nor U4373 (N_4373,N_4216,N_4271);
xor U4374 (N_4374,N_4301,N_4259);
or U4375 (N_4375,N_4263,N_4254);
and U4376 (N_4376,N_4201,N_4170);
nand U4377 (N_4377,N_4194,N_4283);
or U4378 (N_4378,N_4186,N_4203);
and U4379 (N_4379,N_4225,N_4245);
and U4380 (N_4380,N_4209,N_4313);
nor U4381 (N_4381,N_4196,N_4248);
nand U4382 (N_4382,N_4176,N_4184);
and U4383 (N_4383,N_4268,N_4178);
nand U4384 (N_4384,N_4310,N_4277);
or U4385 (N_4385,N_4179,N_4199);
and U4386 (N_4386,N_4217,N_4294);
nor U4387 (N_4387,N_4314,N_4295);
nor U4388 (N_4388,N_4183,N_4315);
nor U4389 (N_4389,N_4276,N_4257);
or U4390 (N_4390,N_4175,N_4189);
and U4391 (N_4391,N_4297,N_4306);
and U4392 (N_4392,N_4275,N_4233);
nor U4393 (N_4393,N_4243,N_4198);
xnor U4394 (N_4394,N_4220,N_4160);
nand U4395 (N_4395,N_4302,N_4204);
and U4396 (N_4396,N_4164,N_4309);
and U4397 (N_4397,N_4296,N_4258);
and U4398 (N_4398,N_4273,N_4169);
and U4399 (N_4399,N_4206,N_4193);
or U4400 (N_4400,N_4165,N_4282);
nand U4401 (N_4401,N_4206,N_4268);
or U4402 (N_4402,N_4212,N_4211);
and U4403 (N_4403,N_4287,N_4270);
or U4404 (N_4404,N_4224,N_4307);
nor U4405 (N_4405,N_4257,N_4218);
or U4406 (N_4406,N_4253,N_4178);
nor U4407 (N_4407,N_4164,N_4272);
nand U4408 (N_4408,N_4189,N_4252);
nor U4409 (N_4409,N_4282,N_4190);
nand U4410 (N_4410,N_4293,N_4296);
nand U4411 (N_4411,N_4296,N_4173);
nor U4412 (N_4412,N_4178,N_4311);
and U4413 (N_4413,N_4247,N_4212);
nor U4414 (N_4414,N_4296,N_4241);
nor U4415 (N_4415,N_4244,N_4218);
nor U4416 (N_4416,N_4203,N_4174);
nor U4417 (N_4417,N_4291,N_4238);
nand U4418 (N_4418,N_4199,N_4210);
nor U4419 (N_4419,N_4301,N_4176);
or U4420 (N_4420,N_4319,N_4314);
nand U4421 (N_4421,N_4182,N_4240);
and U4422 (N_4422,N_4299,N_4241);
and U4423 (N_4423,N_4200,N_4314);
nand U4424 (N_4424,N_4192,N_4167);
nand U4425 (N_4425,N_4252,N_4190);
xnor U4426 (N_4426,N_4210,N_4303);
or U4427 (N_4427,N_4206,N_4272);
nand U4428 (N_4428,N_4257,N_4169);
or U4429 (N_4429,N_4239,N_4247);
and U4430 (N_4430,N_4299,N_4237);
and U4431 (N_4431,N_4266,N_4196);
nand U4432 (N_4432,N_4177,N_4202);
or U4433 (N_4433,N_4228,N_4245);
or U4434 (N_4434,N_4255,N_4278);
or U4435 (N_4435,N_4201,N_4212);
nand U4436 (N_4436,N_4207,N_4273);
and U4437 (N_4437,N_4185,N_4240);
nand U4438 (N_4438,N_4272,N_4254);
nand U4439 (N_4439,N_4317,N_4204);
nor U4440 (N_4440,N_4315,N_4200);
and U4441 (N_4441,N_4192,N_4253);
nand U4442 (N_4442,N_4197,N_4272);
nor U4443 (N_4443,N_4289,N_4163);
and U4444 (N_4444,N_4274,N_4278);
nand U4445 (N_4445,N_4160,N_4289);
nor U4446 (N_4446,N_4318,N_4264);
xor U4447 (N_4447,N_4258,N_4248);
nor U4448 (N_4448,N_4192,N_4231);
nand U4449 (N_4449,N_4291,N_4311);
nor U4450 (N_4450,N_4216,N_4275);
nand U4451 (N_4451,N_4293,N_4210);
nor U4452 (N_4452,N_4247,N_4303);
or U4453 (N_4453,N_4314,N_4210);
or U4454 (N_4454,N_4234,N_4175);
nor U4455 (N_4455,N_4265,N_4243);
nand U4456 (N_4456,N_4291,N_4254);
nor U4457 (N_4457,N_4174,N_4285);
nor U4458 (N_4458,N_4273,N_4223);
and U4459 (N_4459,N_4204,N_4269);
and U4460 (N_4460,N_4303,N_4206);
nor U4461 (N_4461,N_4308,N_4161);
nor U4462 (N_4462,N_4319,N_4167);
xor U4463 (N_4463,N_4313,N_4255);
nor U4464 (N_4464,N_4202,N_4225);
nor U4465 (N_4465,N_4255,N_4177);
or U4466 (N_4466,N_4184,N_4198);
and U4467 (N_4467,N_4286,N_4217);
xor U4468 (N_4468,N_4202,N_4163);
xor U4469 (N_4469,N_4310,N_4319);
and U4470 (N_4470,N_4182,N_4193);
nand U4471 (N_4471,N_4263,N_4221);
or U4472 (N_4472,N_4315,N_4252);
and U4473 (N_4473,N_4267,N_4191);
or U4474 (N_4474,N_4215,N_4197);
or U4475 (N_4475,N_4299,N_4183);
nand U4476 (N_4476,N_4177,N_4242);
or U4477 (N_4477,N_4312,N_4309);
xnor U4478 (N_4478,N_4247,N_4171);
nor U4479 (N_4479,N_4219,N_4167);
nor U4480 (N_4480,N_4465,N_4410);
and U4481 (N_4481,N_4332,N_4380);
or U4482 (N_4482,N_4468,N_4397);
nand U4483 (N_4483,N_4422,N_4405);
nand U4484 (N_4484,N_4473,N_4447);
or U4485 (N_4485,N_4442,N_4418);
nor U4486 (N_4486,N_4324,N_4430);
or U4487 (N_4487,N_4376,N_4429);
nor U4488 (N_4488,N_4359,N_4350);
nand U4489 (N_4489,N_4362,N_4372);
or U4490 (N_4490,N_4354,N_4394);
xor U4491 (N_4491,N_4441,N_4340);
nand U4492 (N_4492,N_4407,N_4339);
and U4493 (N_4493,N_4426,N_4444);
xor U4494 (N_4494,N_4401,N_4369);
nand U4495 (N_4495,N_4478,N_4445);
and U4496 (N_4496,N_4328,N_4446);
and U4497 (N_4497,N_4406,N_4335);
xnor U4498 (N_4498,N_4425,N_4462);
nand U4499 (N_4499,N_4474,N_4355);
nor U4500 (N_4500,N_4463,N_4333);
and U4501 (N_4501,N_4388,N_4379);
and U4502 (N_4502,N_4464,N_4365);
or U4503 (N_4503,N_4423,N_4360);
nand U4504 (N_4504,N_4338,N_4368);
nand U4505 (N_4505,N_4460,N_4427);
nor U4506 (N_4506,N_4386,N_4448);
nand U4507 (N_4507,N_4436,N_4443);
nand U4508 (N_4508,N_4342,N_4449);
nor U4509 (N_4509,N_4403,N_4402);
xor U4510 (N_4510,N_4475,N_4373);
nand U4511 (N_4511,N_4472,N_4346);
and U4512 (N_4512,N_4323,N_4451);
nor U4513 (N_4513,N_4466,N_4391);
nand U4514 (N_4514,N_4452,N_4456);
nand U4515 (N_4515,N_4420,N_4404);
or U4516 (N_4516,N_4467,N_4428);
and U4517 (N_4517,N_4434,N_4400);
nor U4518 (N_4518,N_4352,N_4432);
nor U4519 (N_4519,N_4392,N_4437);
nand U4520 (N_4520,N_4381,N_4471);
nor U4521 (N_4521,N_4382,N_4399);
or U4522 (N_4522,N_4469,N_4455);
nand U4523 (N_4523,N_4383,N_4348);
nand U4524 (N_4524,N_4454,N_4396);
nand U4525 (N_4525,N_4377,N_4385);
nand U4526 (N_4526,N_4470,N_4357);
nand U4527 (N_4527,N_4337,N_4457);
or U4528 (N_4528,N_4364,N_4413);
nor U4529 (N_4529,N_4343,N_4440);
nand U4530 (N_4530,N_4330,N_4344);
nand U4531 (N_4531,N_4320,N_4458);
nand U4532 (N_4532,N_4353,N_4439);
nand U4533 (N_4533,N_4433,N_4479);
nand U4534 (N_4534,N_4363,N_4378);
xor U4535 (N_4535,N_4329,N_4389);
nor U4536 (N_4536,N_4412,N_4367);
nor U4537 (N_4537,N_4345,N_4358);
and U4538 (N_4538,N_4370,N_4390);
nor U4539 (N_4539,N_4417,N_4419);
nor U4540 (N_4540,N_4374,N_4476);
or U4541 (N_4541,N_4327,N_4325);
xor U4542 (N_4542,N_4411,N_4331);
nor U4543 (N_4543,N_4322,N_4450);
or U4544 (N_4544,N_4347,N_4349);
nor U4545 (N_4545,N_4409,N_4366);
nand U4546 (N_4546,N_4398,N_4477);
nor U4547 (N_4547,N_4414,N_4356);
nand U4548 (N_4548,N_4408,N_4461);
nor U4549 (N_4549,N_4424,N_4351);
and U4550 (N_4550,N_4375,N_4393);
nor U4551 (N_4551,N_4431,N_4321);
nor U4552 (N_4552,N_4341,N_4421);
and U4553 (N_4553,N_4453,N_4438);
or U4554 (N_4554,N_4415,N_4361);
nand U4555 (N_4555,N_4435,N_4371);
nor U4556 (N_4556,N_4334,N_4416);
or U4557 (N_4557,N_4336,N_4384);
nand U4558 (N_4558,N_4459,N_4326);
and U4559 (N_4559,N_4387,N_4395);
nor U4560 (N_4560,N_4448,N_4369);
nand U4561 (N_4561,N_4452,N_4447);
nand U4562 (N_4562,N_4422,N_4432);
or U4563 (N_4563,N_4446,N_4325);
nor U4564 (N_4564,N_4425,N_4389);
xnor U4565 (N_4565,N_4324,N_4352);
nand U4566 (N_4566,N_4322,N_4386);
nand U4567 (N_4567,N_4360,N_4467);
nand U4568 (N_4568,N_4451,N_4423);
xnor U4569 (N_4569,N_4475,N_4338);
xor U4570 (N_4570,N_4435,N_4345);
or U4571 (N_4571,N_4382,N_4384);
nand U4572 (N_4572,N_4473,N_4427);
or U4573 (N_4573,N_4446,N_4408);
and U4574 (N_4574,N_4367,N_4441);
or U4575 (N_4575,N_4470,N_4437);
or U4576 (N_4576,N_4424,N_4394);
and U4577 (N_4577,N_4400,N_4350);
or U4578 (N_4578,N_4350,N_4478);
nor U4579 (N_4579,N_4398,N_4359);
nor U4580 (N_4580,N_4384,N_4440);
nand U4581 (N_4581,N_4343,N_4410);
and U4582 (N_4582,N_4389,N_4373);
nand U4583 (N_4583,N_4415,N_4443);
nor U4584 (N_4584,N_4464,N_4470);
or U4585 (N_4585,N_4353,N_4367);
xnor U4586 (N_4586,N_4360,N_4381);
nand U4587 (N_4587,N_4327,N_4341);
and U4588 (N_4588,N_4391,N_4333);
or U4589 (N_4589,N_4362,N_4333);
nor U4590 (N_4590,N_4425,N_4375);
nand U4591 (N_4591,N_4389,N_4327);
nor U4592 (N_4592,N_4370,N_4417);
nand U4593 (N_4593,N_4326,N_4388);
or U4594 (N_4594,N_4415,N_4369);
nand U4595 (N_4595,N_4380,N_4357);
nor U4596 (N_4596,N_4370,N_4438);
xnor U4597 (N_4597,N_4477,N_4440);
and U4598 (N_4598,N_4461,N_4352);
or U4599 (N_4599,N_4449,N_4320);
nand U4600 (N_4600,N_4463,N_4421);
or U4601 (N_4601,N_4419,N_4479);
nand U4602 (N_4602,N_4450,N_4391);
or U4603 (N_4603,N_4432,N_4345);
nor U4604 (N_4604,N_4425,N_4377);
nand U4605 (N_4605,N_4401,N_4337);
nor U4606 (N_4606,N_4337,N_4431);
nand U4607 (N_4607,N_4442,N_4386);
nor U4608 (N_4608,N_4400,N_4432);
nor U4609 (N_4609,N_4341,N_4423);
nor U4610 (N_4610,N_4382,N_4347);
or U4611 (N_4611,N_4320,N_4350);
xor U4612 (N_4612,N_4327,N_4411);
nand U4613 (N_4613,N_4338,N_4346);
nor U4614 (N_4614,N_4367,N_4430);
or U4615 (N_4615,N_4346,N_4422);
or U4616 (N_4616,N_4389,N_4340);
nor U4617 (N_4617,N_4455,N_4457);
and U4618 (N_4618,N_4378,N_4452);
xor U4619 (N_4619,N_4431,N_4356);
xor U4620 (N_4620,N_4461,N_4452);
and U4621 (N_4621,N_4404,N_4367);
nand U4622 (N_4622,N_4475,N_4387);
and U4623 (N_4623,N_4439,N_4430);
nor U4624 (N_4624,N_4321,N_4345);
nand U4625 (N_4625,N_4400,N_4435);
nand U4626 (N_4626,N_4433,N_4389);
nand U4627 (N_4627,N_4391,N_4331);
and U4628 (N_4628,N_4325,N_4462);
nor U4629 (N_4629,N_4474,N_4475);
xnor U4630 (N_4630,N_4373,N_4383);
nor U4631 (N_4631,N_4460,N_4433);
or U4632 (N_4632,N_4462,N_4448);
and U4633 (N_4633,N_4345,N_4371);
xnor U4634 (N_4634,N_4428,N_4448);
nor U4635 (N_4635,N_4437,N_4352);
and U4636 (N_4636,N_4320,N_4419);
nand U4637 (N_4637,N_4376,N_4403);
nand U4638 (N_4638,N_4367,N_4341);
nand U4639 (N_4639,N_4375,N_4402);
nor U4640 (N_4640,N_4529,N_4600);
and U4641 (N_4641,N_4517,N_4493);
or U4642 (N_4642,N_4545,N_4515);
and U4643 (N_4643,N_4575,N_4584);
nor U4644 (N_4644,N_4582,N_4592);
and U4645 (N_4645,N_4542,N_4534);
nand U4646 (N_4646,N_4590,N_4622);
nor U4647 (N_4647,N_4553,N_4580);
or U4648 (N_4648,N_4574,N_4508);
nand U4649 (N_4649,N_4609,N_4480);
nand U4650 (N_4650,N_4626,N_4629);
or U4651 (N_4651,N_4633,N_4623);
nand U4652 (N_4652,N_4569,N_4585);
nor U4653 (N_4653,N_4516,N_4612);
nor U4654 (N_4654,N_4631,N_4496);
and U4655 (N_4655,N_4625,N_4531);
or U4656 (N_4656,N_4573,N_4521);
and U4657 (N_4657,N_4602,N_4618);
and U4658 (N_4658,N_4539,N_4558);
nand U4659 (N_4659,N_4607,N_4616);
nand U4660 (N_4660,N_4639,N_4490);
or U4661 (N_4661,N_4559,N_4549);
xnor U4662 (N_4662,N_4621,N_4610);
or U4663 (N_4663,N_4624,N_4540);
xnor U4664 (N_4664,N_4550,N_4567);
or U4665 (N_4665,N_4500,N_4520);
nand U4666 (N_4666,N_4620,N_4595);
and U4667 (N_4667,N_4587,N_4510);
nand U4668 (N_4668,N_4617,N_4525);
nand U4669 (N_4669,N_4572,N_4603);
nor U4670 (N_4670,N_4576,N_4494);
nand U4671 (N_4671,N_4591,N_4605);
nor U4672 (N_4672,N_4489,N_4638);
or U4673 (N_4673,N_4483,N_4537);
nor U4674 (N_4674,N_4548,N_4527);
and U4675 (N_4675,N_4634,N_4583);
or U4676 (N_4676,N_4506,N_4613);
and U4677 (N_4677,N_4492,N_4488);
or U4678 (N_4678,N_4557,N_4594);
or U4679 (N_4679,N_4555,N_4499);
or U4680 (N_4680,N_4530,N_4561);
or U4681 (N_4681,N_4546,N_4505);
or U4682 (N_4682,N_4522,N_4611);
nor U4683 (N_4683,N_4596,N_4556);
nor U4684 (N_4684,N_4528,N_4619);
nor U4685 (N_4685,N_4599,N_4563);
nand U4686 (N_4686,N_4571,N_4485);
nand U4687 (N_4687,N_4635,N_4511);
or U4688 (N_4688,N_4501,N_4509);
and U4689 (N_4689,N_4562,N_4589);
or U4690 (N_4690,N_4568,N_4484);
nand U4691 (N_4691,N_4487,N_4523);
and U4692 (N_4692,N_4627,N_4514);
and U4693 (N_4693,N_4614,N_4497);
and U4694 (N_4694,N_4536,N_4544);
nand U4695 (N_4695,N_4601,N_4486);
or U4696 (N_4696,N_4637,N_4504);
and U4697 (N_4697,N_4565,N_4547);
xnor U4698 (N_4698,N_4554,N_4566);
nor U4699 (N_4699,N_4526,N_4535);
xor U4700 (N_4700,N_4579,N_4564);
and U4701 (N_4701,N_4578,N_4482);
nor U4702 (N_4702,N_4495,N_4541);
and U4703 (N_4703,N_4593,N_4491);
nor U4704 (N_4704,N_4551,N_4586);
or U4705 (N_4705,N_4606,N_4502);
or U4706 (N_4706,N_4513,N_4503);
nor U4707 (N_4707,N_4533,N_4498);
or U4708 (N_4708,N_4581,N_4588);
xor U4709 (N_4709,N_4628,N_4552);
and U4710 (N_4710,N_4512,N_4630);
nand U4711 (N_4711,N_4577,N_4570);
or U4712 (N_4712,N_4507,N_4604);
nor U4713 (N_4713,N_4560,N_4615);
and U4714 (N_4714,N_4608,N_4538);
and U4715 (N_4715,N_4632,N_4636);
nand U4716 (N_4716,N_4597,N_4543);
nand U4717 (N_4717,N_4518,N_4524);
nor U4718 (N_4718,N_4481,N_4519);
or U4719 (N_4719,N_4532,N_4598);
nand U4720 (N_4720,N_4557,N_4556);
nor U4721 (N_4721,N_4624,N_4572);
and U4722 (N_4722,N_4527,N_4579);
or U4723 (N_4723,N_4493,N_4535);
or U4724 (N_4724,N_4517,N_4482);
or U4725 (N_4725,N_4621,N_4519);
or U4726 (N_4726,N_4576,N_4579);
nor U4727 (N_4727,N_4546,N_4535);
nor U4728 (N_4728,N_4591,N_4621);
nand U4729 (N_4729,N_4577,N_4571);
nor U4730 (N_4730,N_4614,N_4543);
and U4731 (N_4731,N_4521,N_4566);
and U4732 (N_4732,N_4498,N_4532);
nand U4733 (N_4733,N_4539,N_4532);
or U4734 (N_4734,N_4564,N_4638);
and U4735 (N_4735,N_4549,N_4501);
and U4736 (N_4736,N_4577,N_4540);
or U4737 (N_4737,N_4560,N_4627);
xor U4738 (N_4738,N_4497,N_4552);
and U4739 (N_4739,N_4625,N_4544);
nor U4740 (N_4740,N_4482,N_4541);
or U4741 (N_4741,N_4607,N_4522);
xor U4742 (N_4742,N_4494,N_4516);
or U4743 (N_4743,N_4627,N_4523);
and U4744 (N_4744,N_4486,N_4520);
and U4745 (N_4745,N_4576,N_4595);
nand U4746 (N_4746,N_4545,N_4574);
or U4747 (N_4747,N_4585,N_4486);
or U4748 (N_4748,N_4506,N_4536);
nor U4749 (N_4749,N_4483,N_4562);
or U4750 (N_4750,N_4583,N_4498);
or U4751 (N_4751,N_4578,N_4565);
or U4752 (N_4752,N_4570,N_4612);
nand U4753 (N_4753,N_4516,N_4532);
or U4754 (N_4754,N_4532,N_4543);
nand U4755 (N_4755,N_4495,N_4499);
or U4756 (N_4756,N_4510,N_4505);
and U4757 (N_4757,N_4529,N_4548);
or U4758 (N_4758,N_4508,N_4588);
or U4759 (N_4759,N_4553,N_4620);
or U4760 (N_4760,N_4522,N_4613);
and U4761 (N_4761,N_4506,N_4584);
and U4762 (N_4762,N_4600,N_4525);
nand U4763 (N_4763,N_4574,N_4488);
nand U4764 (N_4764,N_4480,N_4544);
nor U4765 (N_4765,N_4484,N_4511);
xor U4766 (N_4766,N_4538,N_4619);
or U4767 (N_4767,N_4601,N_4611);
and U4768 (N_4768,N_4582,N_4512);
or U4769 (N_4769,N_4480,N_4559);
or U4770 (N_4770,N_4594,N_4511);
and U4771 (N_4771,N_4482,N_4619);
and U4772 (N_4772,N_4637,N_4621);
nor U4773 (N_4773,N_4617,N_4543);
xnor U4774 (N_4774,N_4607,N_4556);
or U4775 (N_4775,N_4606,N_4527);
nor U4776 (N_4776,N_4604,N_4572);
nor U4777 (N_4777,N_4632,N_4526);
and U4778 (N_4778,N_4597,N_4515);
xnor U4779 (N_4779,N_4536,N_4494);
or U4780 (N_4780,N_4485,N_4491);
xnor U4781 (N_4781,N_4602,N_4518);
nand U4782 (N_4782,N_4639,N_4532);
xnor U4783 (N_4783,N_4601,N_4607);
nor U4784 (N_4784,N_4508,N_4505);
nand U4785 (N_4785,N_4506,N_4616);
nand U4786 (N_4786,N_4514,N_4525);
nor U4787 (N_4787,N_4598,N_4523);
or U4788 (N_4788,N_4514,N_4491);
or U4789 (N_4789,N_4531,N_4494);
and U4790 (N_4790,N_4639,N_4591);
or U4791 (N_4791,N_4566,N_4513);
nor U4792 (N_4792,N_4625,N_4497);
or U4793 (N_4793,N_4637,N_4531);
and U4794 (N_4794,N_4488,N_4568);
or U4795 (N_4795,N_4578,N_4562);
and U4796 (N_4796,N_4620,N_4509);
and U4797 (N_4797,N_4565,N_4592);
nor U4798 (N_4798,N_4490,N_4575);
and U4799 (N_4799,N_4572,N_4522);
nand U4800 (N_4800,N_4752,N_4664);
xor U4801 (N_4801,N_4799,N_4713);
nand U4802 (N_4802,N_4659,N_4797);
or U4803 (N_4803,N_4743,N_4795);
or U4804 (N_4804,N_4739,N_4787);
or U4805 (N_4805,N_4709,N_4723);
nor U4806 (N_4806,N_4661,N_4668);
nand U4807 (N_4807,N_4715,N_4658);
nand U4808 (N_4808,N_4790,N_4655);
or U4809 (N_4809,N_4733,N_4747);
or U4810 (N_4810,N_4749,N_4679);
and U4811 (N_4811,N_4643,N_4786);
nor U4812 (N_4812,N_4788,N_4699);
nor U4813 (N_4813,N_4707,N_4703);
nor U4814 (N_4814,N_4704,N_4684);
or U4815 (N_4815,N_4690,N_4735);
or U4816 (N_4816,N_4774,N_4717);
nand U4817 (N_4817,N_4745,N_4666);
or U4818 (N_4818,N_4662,N_4779);
and U4819 (N_4819,N_4646,N_4705);
xnor U4820 (N_4820,N_4706,N_4680);
and U4821 (N_4821,N_4697,N_4711);
nor U4822 (N_4822,N_4692,N_4759);
nand U4823 (N_4823,N_4769,N_4792);
nor U4824 (N_4824,N_4742,N_4781);
and U4825 (N_4825,N_4721,N_4689);
nor U4826 (N_4826,N_4675,N_4731);
and U4827 (N_4827,N_4798,N_4716);
and U4828 (N_4828,N_4762,N_4714);
nor U4829 (N_4829,N_4738,N_4640);
or U4830 (N_4830,N_4728,N_4729);
nand U4831 (N_4831,N_4732,N_4663);
nor U4832 (N_4832,N_4794,N_4754);
or U4833 (N_4833,N_4796,N_4771);
nor U4834 (N_4834,N_4667,N_4722);
and U4835 (N_4835,N_4688,N_4652);
and U4836 (N_4836,N_4693,N_4702);
nor U4837 (N_4837,N_4683,N_4757);
or U4838 (N_4838,N_4657,N_4671);
nor U4839 (N_4839,N_4691,N_4753);
nand U4840 (N_4840,N_4763,N_4764);
and U4841 (N_4841,N_4686,N_4783);
and U4842 (N_4842,N_4712,N_4653);
nand U4843 (N_4843,N_4674,N_4672);
and U4844 (N_4844,N_4645,N_4758);
nor U4845 (N_4845,N_4708,N_4760);
nand U4846 (N_4846,N_4726,N_4656);
xor U4847 (N_4847,N_4694,N_4685);
nor U4848 (N_4848,N_4701,N_4718);
nand U4849 (N_4849,N_4682,N_4698);
and U4850 (N_4850,N_4782,N_4642);
or U4851 (N_4851,N_4725,N_4681);
nand U4852 (N_4852,N_4750,N_4644);
and U4853 (N_4853,N_4737,N_4647);
or U4854 (N_4854,N_4670,N_4751);
nor U4855 (N_4855,N_4687,N_4660);
nand U4856 (N_4856,N_4665,N_4734);
and U4857 (N_4857,N_4767,N_4746);
or U4858 (N_4858,N_4677,N_4776);
and U4859 (N_4859,N_4676,N_4777);
or U4860 (N_4860,N_4785,N_4789);
nand U4861 (N_4861,N_4766,N_4756);
nand U4862 (N_4862,N_4695,N_4793);
and U4863 (N_4863,N_4654,N_4770);
nor U4864 (N_4864,N_4678,N_4650);
xnor U4865 (N_4865,N_4773,N_4780);
nor U4866 (N_4866,N_4768,N_4710);
or U4867 (N_4867,N_4772,N_4791);
or U4868 (N_4868,N_4736,N_4719);
or U4869 (N_4869,N_4727,N_4648);
and U4870 (N_4870,N_4741,N_4649);
or U4871 (N_4871,N_4740,N_4730);
nand U4872 (N_4872,N_4669,N_4775);
nor U4873 (N_4873,N_4673,N_4651);
nand U4874 (N_4874,N_4696,N_4761);
or U4875 (N_4875,N_4755,N_4778);
and U4876 (N_4876,N_4748,N_4641);
or U4877 (N_4877,N_4744,N_4724);
nand U4878 (N_4878,N_4765,N_4700);
and U4879 (N_4879,N_4784,N_4720);
and U4880 (N_4880,N_4788,N_4774);
nor U4881 (N_4881,N_4728,N_4699);
nor U4882 (N_4882,N_4651,N_4768);
nor U4883 (N_4883,N_4791,N_4738);
nor U4884 (N_4884,N_4667,N_4766);
nand U4885 (N_4885,N_4687,N_4778);
or U4886 (N_4886,N_4708,N_4721);
xnor U4887 (N_4887,N_4704,N_4655);
nor U4888 (N_4888,N_4765,N_4789);
nand U4889 (N_4889,N_4695,N_4795);
nand U4890 (N_4890,N_4749,N_4700);
nand U4891 (N_4891,N_4687,N_4738);
nor U4892 (N_4892,N_4771,N_4785);
xnor U4893 (N_4893,N_4776,N_4692);
nand U4894 (N_4894,N_4781,N_4762);
nor U4895 (N_4895,N_4715,N_4785);
or U4896 (N_4896,N_4654,N_4718);
or U4897 (N_4897,N_4741,N_4712);
nand U4898 (N_4898,N_4723,N_4674);
nor U4899 (N_4899,N_4780,N_4760);
or U4900 (N_4900,N_4690,N_4665);
nand U4901 (N_4901,N_4744,N_4716);
nand U4902 (N_4902,N_4646,N_4699);
xor U4903 (N_4903,N_4794,N_4772);
and U4904 (N_4904,N_4650,N_4656);
and U4905 (N_4905,N_4796,N_4698);
or U4906 (N_4906,N_4747,N_4791);
and U4907 (N_4907,N_4729,N_4737);
nand U4908 (N_4908,N_4770,N_4773);
and U4909 (N_4909,N_4710,N_4748);
nor U4910 (N_4910,N_4647,N_4793);
and U4911 (N_4911,N_4719,N_4645);
nor U4912 (N_4912,N_4659,N_4767);
and U4913 (N_4913,N_4717,N_4722);
and U4914 (N_4914,N_4681,N_4660);
xnor U4915 (N_4915,N_4664,N_4716);
xor U4916 (N_4916,N_4778,N_4662);
or U4917 (N_4917,N_4659,N_4652);
or U4918 (N_4918,N_4791,N_4663);
nor U4919 (N_4919,N_4649,N_4693);
nand U4920 (N_4920,N_4654,N_4773);
nor U4921 (N_4921,N_4713,N_4736);
nor U4922 (N_4922,N_4726,N_4716);
or U4923 (N_4923,N_4710,N_4654);
nand U4924 (N_4924,N_4796,N_4648);
xnor U4925 (N_4925,N_4768,N_4798);
or U4926 (N_4926,N_4670,N_4782);
nor U4927 (N_4927,N_4768,N_4762);
or U4928 (N_4928,N_4743,N_4647);
nor U4929 (N_4929,N_4781,N_4641);
nor U4930 (N_4930,N_4748,N_4701);
and U4931 (N_4931,N_4723,N_4685);
nand U4932 (N_4932,N_4687,N_4790);
nand U4933 (N_4933,N_4777,N_4669);
or U4934 (N_4934,N_4711,N_4755);
and U4935 (N_4935,N_4721,N_4666);
nor U4936 (N_4936,N_4780,N_4745);
xnor U4937 (N_4937,N_4680,N_4789);
nor U4938 (N_4938,N_4657,N_4760);
nand U4939 (N_4939,N_4681,N_4721);
nand U4940 (N_4940,N_4740,N_4775);
nor U4941 (N_4941,N_4669,N_4728);
nand U4942 (N_4942,N_4771,N_4656);
or U4943 (N_4943,N_4708,N_4644);
nand U4944 (N_4944,N_4665,N_4700);
or U4945 (N_4945,N_4659,N_4754);
xor U4946 (N_4946,N_4701,N_4647);
or U4947 (N_4947,N_4681,N_4762);
nand U4948 (N_4948,N_4717,N_4698);
or U4949 (N_4949,N_4728,N_4722);
and U4950 (N_4950,N_4731,N_4713);
nand U4951 (N_4951,N_4647,N_4677);
xor U4952 (N_4952,N_4711,N_4783);
or U4953 (N_4953,N_4641,N_4659);
and U4954 (N_4954,N_4661,N_4786);
and U4955 (N_4955,N_4698,N_4667);
nand U4956 (N_4956,N_4676,N_4682);
and U4957 (N_4957,N_4649,N_4681);
and U4958 (N_4958,N_4745,N_4682);
nand U4959 (N_4959,N_4643,N_4706);
or U4960 (N_4960,N_4925,N_4895);
nor U4961 (N_4961,N_4952,N_4873);
nor U4962 (N_4962,N_4905,N_4838);
nand U4963 (N_4963,N_4906,N_4854);
and U4964 (N_4964,N_4823,N_4856);
or U4965 (N_4965,N_4821,N_4872);
nand U4966 (N_4966,N_4939,N_4914);
and U4967 (N_4967,N_4836,N_4936);
xor U4968 (N_4968,N_4849,N_4817);
nand U4969 (N_4969,N_4917,N_4860);
nor U4970 (N_4970,N_4948,N_4950);
or U4971 (N_4971,N_4807,N_4841);
or U4972 (N_4972,N_4846,N_4889);
nand U4973 (N_4973,N_4848,N_4913);
nand U4974 (N_4974,N_4837,N_4899);
and U4975 (N_4975,N_4953,N_4883);
and U4976 (N_4976,N_4813,N_4942);
or U4977 (N_4977,N_4903,N_4945);
or U4978 (N_4978,N_4874,N_4835);
or U4979 (N_4979,N_4830,N_4800);
or U4980 (N_4980,N_4891,N_4922);
nand U4981 (N_4981,N_4926,N_4845);
nor U4982 (N_4982,N_4944,N_4943);
or U4983 (N_4983,N_4855,N_4858);
nand U4984 (N_4984,N_4904,N_4894);
nand U4985 (N_4985,N_4920,N_4892);
nor U4986 (N_4986,N_4957,N_4912);
nor U4987 (N_4987,N_4818,N_4842);
or U4988 (N_4988,N_4941,N_4916);
xnor U4989 (N_4989,N_4870,N_4859);
or U4990 (N_4990,N_4875,N_4863);
and U4991 (N_4991,N_4816,N_4820);
nand U4992 (N_4992,N_4814,N_4831);
nor U4993 (N_4993,N_4958,N_4919);
nand U4994 (N_4994,N_4898,N_4839);
nor U4995 (N_4995,N_4824,N_4804);
nor U4996 (N_4996,N_4907,N_4929);
nand U4997 (N_4997,N_4949,N_4956);
nor U4998 (N_4998,N_4933,N_4880);
and U4999 (N_4999,N_4828,N_4827);
xor U5000 (N_5000,N_4868,N_4815);
nand U5001 (N_5001,N_4927,N_4843);
nand U5002 (N_5002,N_4822,N_4896);
nand U5003 (N_5003,N_4946,N_4881);
and U5004 (N_5004,N_4951,N_4887);
or U5005 (N_5005,N_4923,N_4885);
nor U5006 (N_5006,N_4853,N_4834);
nor U5007 (N_5007,N_4900,N_4832);
xor U5008 (N_5008,N_4850,N_4862);
and U5009 (N_5009,N_4861,N_4811);
and U5010 (N_5010,N_4866,N_4921);
nor U5011 (N_5011,N_4871,N_4930);
nand U5012 (N_5012,N_4959,N_4908);
nor U5013 (N_5013,N_4864,N_4893);
xnor U5014 (N_5014,N_4826,N_4954);
nand U5015 (N_5015,N_4915,N_4809);
nand U5016 (N_5016,N_4851,N_4934);
and U5017 (N_5017,N_4847,N_4947);
nand U5018 (N_5018,N_4829,N_4810);
or U5019 (N_5019,N_4888,N_4901);
and U5020 (N_5020,N_4897,N_4879);
nand U5021 (N_5021,N_4928,N_4819);
xor U5022 (N_5022,N_4955,N_4877);
and U5023 (N_5023,N_4911,N_4884);
or U5024 (N_5024,N_4932,N_4886);
or U5025 (N_5025,N_4902,N_4909);
nor U5026 (N_5026,N_4910,N_4924);
or U5027 (N_5027,N_4938,N_4940);
and U5028 (N_5028,N_4833,N_4844);
and U5029 (N_5029,N_4878,N_4805);
xnor U5030 (N_5030,N_4808,N_4852);
or U5031 (N_5031,N_4801,N_4857);
nor U5032 (N_5032,N_4803,N_4890);
nand U5033 (N_5033,N_4825,N_4840);
nand U5034 (N_5034,N_4935,N_4937);
or U5035 (N_5035,N_4876,N_4869);
nor U5036 (N_5036,N_4865,N_4931);
nand U5037 (N_5037,N_4802,N_4812);
nand U5038 (N_5038,N_4806,N_4882);
nor U5039 (N_5039,N_4867,N_4918);
or U5040 (N_5040,N_4877,N_4811);
nand U5041 (N_5041,N_4909,N_4821);
or U5042 (N_5042,N_4835,N_4849);
nand U5043 (N_5043,N_4818,N_4836);
and U5044 (N_5044,N_4875,N_4911);
or U5045 (N_5045,N_4928,N_4903);
and U5046 (N_5046,N_4903,N_4867);
nor U5047 (N_5047,N_4857,N_4864);
nand U5048 (N_5048,N_4849,N_4873);
and U5049 (N_5049,N_4862,N_4918);
nand U5050 (N_5050,N_4878,N_4924);
or U5051 (N_5051,N_4875,N_4937);
nor U5052 (N_5052,N_4824,N_4915);
nor U5053 (N_5053,N_4907,N_4866);
or U5054 (N_5054,N_4868,N_4938);
nand U5055 (N_5055,N_4937,N_4850);
and U5056 (N_5056,N_4938,N_4934);
and U5057 (N_5057,N_4877,N_4914);
and U5058 (N_5058,N_4818,N_4835);
or U5059 (N_5059,N_4944,N_4955);
and U5060 (N_5060,N_4921,N_4824);
and U5061 (N_5061,N_4858,N_4893);
xor U5062 (N_5062,N_4825,N_4822);
and U5063 (N_5063,N_4915,N_4902);
or U5064 (N_5064,N_4868,N_4901);
nand U5065 (N_5065,N_4826,N_4935);
and U5066 (N_5066,N_4874,N_4864);
nand U5067 (N_5067,N_4939,N_4826);
nand U5068 (N_5068,N_4886,N_4891);
and U5069 (N_5069,N_4957,N_4817);
or U5070 (N_5070,N_4922,N_4884);
nor U5071 (N_5071,N_4817,N_4870);
nor U5072 (N_5072,N_4941,N_4959);
nor U5073 (N_5073,N_4914,N_4944);
or U5074 (N_5074,N_4924,N_4913);
nor U5075 (N_5075,N_4868,N_4867);
nand U5076 (N_5076,N_4875,N_4871);
nor U5077 (N_5077,N_4895,N_4955);
and U5078 (N_5078,N_4854,N_4869);
nor U5079 (N_5079,N_4883,N_4827);
nor U5080 (N_5080,N_4873,N_4856);
or U5081 (N_5081,N_4893,N_4914);
and U5082 (N_5082,N_4943,N_4827);
and U5083 (N_5083,N_4802,N_4952);
nand U5084 (N_5084,N_4953,N_4894);
nor U5085 (N_5085,N_4925,N_4951);
and U5086 (N_5086,N_4887,N_4867);
nand U5087 (N_5087,N_4930,N_4822);
nand U5088 (N_5088,N_4906,N_4843);
or U5089 (N_5089,N_4934,N_4917);
or U5090 (N_5090,N_4839,N_4831);
nor U5091 (N_5091,N_4824,N_4882);
xnor U5092 (N_5092,N_4826,N_4810);
or U5093 (N_5093,N_4843,N_4944);
nor U5094 (N_5094,N_4855,N_4847);
xor U5095 (N_5095,N_4807,N_4934);
nand U5096 (N_5096,N_4873,N_4874);
or U5097 (N_5097,N_4940,N_4953);
nor U5098 (N_5098,N_4938,N_4957);
and U5099 (N_5099,N_4840,N_4950);
and U5100 (N_5100,N_4955,N_4881);
and U5101 (N_5101,N_4920,N_4915);
and U5102 (N_5102,N_4807,N_4951);
and U5103 (N_5103,N_4954,N_4914);
nand U5104 (N_5104,N_4814,N_4878);
xnor U5105 (N_5105,N_4922,N_4880);
and U5106 (N_5106,N_4922,N_4804);
nor U5107 (N_5107,N_4828,N_4908);
nor U5108 (N_5108,N_4847,N_4954);
nand U5109 (N_5109,N_4870,N_4872);
nor U5110 (N_5110,N_4906,N_4916);
and U5111 (N_5111,N_4856,N_4936);
nand U5112 (N_5112,N_4879,N_4855);
nand U5113 (N_5113,N_4826,N_4853);
nand U5114 (N_5114,N_4819,N_4943);
nand U5115 (N_5115,N_4835,N_4801);
nor U5116 (N_5116,N_4925,N_4918);
xor U5117 (N_5117,N_4829,N_4854);
nor U5118 (N_5118,N_4894,N_4938);
nor U5119 (N_5119,N_4816,N_4956);
nand U5120 (N_5120,N_4967,N_5042);
or U5121 (N_5121,N_4995,N_4989);
nand U5122 (N_5122,N_5096,N_5077);
or U5123 (N_5123,N_5114,N_4977);
nand U5124 (N_5124,N_5036,N_5101);
nand U5125 (N_5125,N_5002,N_5035);
nor U5126 (N_5126,N_5005,N_5078);
nand U5127 (N_5127,N_5093,N_5022);
or U5128 (N_5128,N_4976,N_5061);
nor U5129 (N_5129,N_5046,N_4984);
or U5130 (N_5130,N_4971,N_5050);
nand U5131 (N_5131,N_5118,N_5068);
nor U5132 (N_5132,N_5014,N_5003);
nor U5133 (N_5133,N_5010,N_4970);
or U5134 (N_5134,N_5065,N_4965);
and U5135 (N_5135,N_5079,N_5094);
nor U5136 (N_5136,N_5012,N_4960);
nor U5137 (N_5137,N_5004,N_5099);
nand U5138 (N_5138,N_5116,N_4997);
nor U5139 (N_5139,N_5080,N_5029);
and U5140 (N_5140,N_5030,N_4974);
nand U5141 (N_5141,N_5084,N_5064);
and U5142 (N_5142,N_5097,N_5016);
nor U5143 (N_5143,N_5054,N_5088);
and U5144 (N_5144,N_5000,N_5060);
nor U5145 (N_5145,N_4979,N_5047);
nor U5146 (N_5146,N_4964,N_5011);
nor U5147 (N_5147,N_5020,N_5015);
and U5148 (N_5148,N_5034,N_5053);
nand U5149 (N_5149,N_5063,N_5082);
xnor U5150 (N_5150,N_5040,N_5106);
nand U5151 (N_5151,N_4975,N_5073);
nand U5152 (N_5152,N_4982,N_5028);
nand U5153 (N_5153,N_5115,N_5025);
and U5154 (N_5154,N_5087,N_5108);
and U5155 (N_5155,N_5008,N_4990);
nand U5156 (N_5156,N_5049,N_5103);
nor U5157 (N_5157,N_5039,N_5074);
or U5158 (N_5158,N_4999,N_5062);
or U5159 (N_5159,N_5081,N_5095);
and U5160 (N_5160,N_5102,N_4962);
or U5161 (N_5161,N_5091,N_5056);
nand U5162 (N_5162,N_5021,N_4994);
and U5163 (N_5163,N_5086,N_5006);
nor U5164 (N_5164,N_5019,N_5009);
or U5165 (N_5165,N_5032,N_5109);
nor U5166 (N_5166,N_4981,N_5098);
nand U5167 (N_5167,N_5018,N_4998);
nand U5168 (N_5168,N_5037,N_4961);
nand U5169 (N_5169,N_5001,N_5043);
nor U5170 (N_5170,N_5044,N_4972);
and U5171 (N_5171,N_5026,N_4968);
and U5172 (N_5172,N_5083,N_5075);
nand U5173 (N_5173,N_5112,N_5066);
and U5174 (N_5174,N_5113,N_5072);
nand U5175 (N_5175,N_4996,N_4985);
and U5176 (N_5176,N_5023,N_5089);
or U5177 (N_5177,N_5117,N_5071);
and U5178 (N_5178,N_5104,N_5110);
nor U5179 (N_5179,N_5059,N_5051);
or U5180 (N_5180,N_4987,N_5092);
xnor U5181 (N_5181,N_5085,N_5055);
xnor U5182 (N_5182,N_5119,N_4978);
or U5183 (N_5183,N_5031,N_5090);
or U5184 (N_5184,N_4983,N_5045);
nor U5185 (N_5185,N_4988,N_5067);
and U5186 (N_5186,N_5107,N_5033);
nand U5187 (N_5187,N_4973,N_5007);
nand U5188 (N_5188,N_5111,N_5017);
nor U5189 (N_5189,N_5013,N_4991);
nor U5190 (N_5190,N_5057,N_4980);
nand U5191 (N_5191,N_5041,N_5100);
or U5192 (N_5192,N_5105,N_4986);
or U5193 (N_5193,N_5069,N_5076);
or U5194 (N_5194,N_5027,N_5058);
nand U5195 (N_5195,N_4966,N_5052);
nor U5196 (N_5196,N_5038,N_4993);
nor U5197 (N_5197,N_5070,N_5048);
nand U5198 (N_5198,N_5024,N_4969);
nand U5199 (N_5199,N_4992,N_4963);
and U5200 (N_5200,N_5117,N_5064);
nand U5201 (N_5201,N_5038,N_5083);
xnor U5202 (N_5202,N_5089,N_5051);
or U5203 (N_5203,N_5109,N_5064);
nand U5204 (N_5204,N_5028,N_5008);
and U5205 (N_5205,N_5117,N_5034);
or U5206 (N_5206,N_4970,N_5082);
or U5207 (N_5207,N_5109,N_5053);
and U5208 (N_5208,N_5103,N_5045);
xor U5209 (N_5209,N_5056,N_5000);
and U5210 (N_5210,N_4966,N_5086);
xor U5211 (N_5211,N_5055,N_5001);
or U5212 (N_5212,N_4962,N_4997);
and U5213 (N_5213,N_5107,N_5036);
or U5214 (N_5214,N_4988,N_5052);
xor U5215 (N_5215,N_4970,N_5098);
and U5216 (N_5216,N_5074,N_5064);
and U5217 (N_5217,N_5116,N_5014);
nor U5218 (N_5218,N_5087,N_4965);
and U5219 (N_5219,N_4968,N_4974);
nand U5220 (N_5220,N_5007,N_4978);
nand U5221 (N_5221,N_5089,N_5018);
nor U5222 (N_5222,N_5010,N_5109);
nor U5223 (N_5223,N_4965,N_4977);
or U5224 (N_5224,N_5049,N_4986);
nor U5225 (N_5225,N_5002,N_5098);
xor U5226 (N_5226,N_5008,N_5043);
nand U5227 (N_5227,N_5020,N_5074);
nand U5228 (N_5228,N_4979,N_5090);
and U5229 (N_5229,N_5077,N_5088);
nor U5230 (N_5230,N_4963,N_5028);
xnor U5231 (N_5231,N_5068,N_5043);
nor U5232 (N_5232,N_5048,N_5051);
or U5233 (N_5233,N_5075,N_4965);
or U5234 (N_5234,N_5050,N_5055);
and U5235 (N_5235,N_5039,N_5057);
xor U5236 (N_5236,N_5069,N_5094);
nand U5237 (N_5237,N_4987,N_4996);
and U5238 (N_5238,N_5084,N_5085);
nor U5239 (N_5239,N_4968,N_5109);
nor U5240 (N_5240,N_5076,N_5048);
nand U5241 (N_5241,N_5094,N_5043);
nor U5242 (N_5242,N_5015,N_5115);
xor U5243 (N_5243,N_5072,N_5030);
and U5244 (N_5244,N_4984,N_4972);
nand U5245 (N_5245,N_5097,N_4968);
nand U5246 (N_5246,N_5112,N_5068);
xnor U5247 (N_5247,N_5093,N_5095);
or U5248 (N_5248,N_5065,N_5047);
xnor U5249 (N_5249,N_4965,N_5048);
and U5250 (N_5250,N_5111,N_5082);
nand U5251 (N_5251,N_5004,N_4974);
nand U5252 (N_5252,N_5073,N_5062);
nor U5253 (N_5253,N_5006,N_5010);
and U5254 (N_5254,N_4986,N_5070);
or U5255 (N_5255,N_5025,N_4980);
nand U5256 (N_5256,N_4964,N_5052);
nand U5257 (N_5257,N_5054,N_5017);
nor U5258 (N_5258,N_5104,N_5008);
or U5259 (N_5259,N_4988,N_4968);
and U5260 (N_5260,N_5059,N_4996);
and U5261 (N_5261,N_5073,N_5019);
and U5262 (N_5262,N_5011,N_5082);
and U5263 (N_5263,N_5008,N_5059);
or U5264 (N_5264,N_4986,N_5106);
nand U5265 (N_5265,N_5099,N_5015);
nor U5266 (N_5266,N_5004,N_5045);
nor U5267 (N_5267,N_5103,N_5108);
nor U5268 (N_5268,N_5075,N_5055);
and U5269 (N_5269,N_5072,N_5062);
nor U5270 (N_5270,N_4988,N_4977);
nand U5271 (N_5271,N_5067,N_5042);
and U5272 (N_5272,N_5104,N_5090);
nand U5273 (N_5273,N_5091,N_4988);
nand U5274 (N_5274,N_5084,N_5070);
nor U5275 (N_5275,N_5040,N_5029);
nor U5276 (N_5276,N_5066,N_4978);
and U5277 (N_5277,N_5040,N_5063);
nand U5278 (N_5278,N_5011,N_5040);
or U5279 (N_5279,N_5021,N_5085);
xor U5280 (N_5280,N_5268,N_5223);
nor U5281 (N_5281,N_5200,N_5187);
and U5282 (N_5282,N_5147,N_5219);
nor U5283 (N_5283,N_5228,N_5172);
and U5284 (N_5284,N_5243,N_5148);
nand U5285 (N_5285,N_5146,N_5255);
nor U5286 (N_5286,N_5231,N_5238);
and U5287 (N_5287,N_5161,N_5263);
nor U5288 (N_5288,N_5171,N_5135);
nand U5289 (N_5289,N_5168,N_5261);
xor U5290 (N_5290,N_5217,N_5136);
and U5291 (N_5291,N_5155,N_5203);
and U5292 (N_5292,N_5209,N_5273);
nand U5293 (N_5293,N_5252,N_5153);
nor U5294 (N_5294,N_5242,N_5165);
nand U5295 (N_5295,N_5218,N_5193);
and U5296 (N_5296,N_5144,N_5139);
nand U5297 (N_5297,N_5237,N_5207);
xnor U5298 (N_5298,N_5227,N_5258);
or U5299 (N_5299,N_5244,N_5234);
nand U5300 (N_5300,N_5213,N_5142);
and U5301 (N_5301,N_5190,N_5210);
nor U5302 (N_5302,N_5152,N_5271);
and U5303 (N_5303,N_5145,N_5253);
or U5304 (N_5304,N_5245,N_5141);
nand U5305 (N_5305,N_5236,N_5275);
and U5306 (N_5306,N_5195,N_5225);
or U5307 (N_5307,N_5143,N_5140);
nand U5308 (N_5308,N_5177,N_5166);
nor U5309 (N_5309,N_5270,N_5160);
nor U5310 (N_5310,N_5204,N_5254);
nand U5311 (N_5311,N_5189,N_5150);
xnor U5312 (N_5312,N_5251,N_5176);
xnor U5313 (N_5313,N_5182,N_5274);
nand U5314 (N_5314,N_5130,N_5260);
or U5315 (N_5315,N_5157,N_5239);
or U5316 (N_5316,N_5235,N_5196);
nor U5317 (N_5317,N_5259,N_5159);
and U5318 (N_5318,N_5170,N_5128);
and U5319 (N_5319,N_5137,N_5269);
nand U5320 (N_5320,N_5198,N_5241);
or U5321 (N_5321,N_5246,N_5191);
nand U5322 (N_5322,N_5192,N_5179);
xor U5323 (N_5323,N_5158,N_5233);
nor U5324 (N_5324,N_5277,N_5216);
nand U5325 (N_5325,N_5131,N_5124);
nor U5326 (N_5326,N_5224,N_5262);
nand U5327 (N_5327,N_5247,N_5126);
or U5328 (N_5328,N_5167,N_5202);
and U5329 (N_5329,N_5123,N_5178);
and U5330 (N_5330,N_5154,N_5221);
and U5331 (N_5331,N_5220,N_5215);
nand U5332 (N_5332,N_5149,N_5240);
or U5333 (N_5333,N_5120,N_5183);
nor U5334 (N_5334,N_5276,N_5164);
or U5335 (N_5335,N_5249,N_5197);
xor U5336 (N_5336,N_5162,N_5278);
nand U5337 (N_5337,N_5129,N_5229);
or U5338 (N_5338,N_5186,N_5169);
or U5339 (N_5339,N_5180,N_5151);
nor U5340 (N_5340,N_5173,N_5256);
nor U5341 (N_5341,N_5125,N_5199);
xnor U5342 (N_5342,N_5133,N_5266);
or U5343 (N_5343,N_5279,N_5127);
nand U5344 (N_5344,N_5122,N_5184);
and U5345 (N_5345,N_5257,N_5185);
nor U5346 (N_5346,N_5265,N_5134);
and U5347 (N_5347,N_5163,N_5267);
nand U5348 (N_5348,N_5181,N_5121);
xnor U5349 (N_5349,N_5208,N_5188);
nor U5350 (N_5350,N_5230,N_5264);
nor U5351 (N_5351,N_5232,N_5212);
nor U5352 (N_5352,N_5250,N_5205);
or U5353 (N_5353,N_5222,N_5156);
nor U5354 (N_5354,N_5194,N_5201);
or U5355 (N_5355,N_5226,N_5211);
or U5356 (N_5356,N_5175,N_5272);
xnor U5357 (N_5357,N_5214,N_5248);
or U5358 (N_5358,N_5132,N_5206);
or U5359 (N_5359,N_5138,N_5174);
nor U5360 (N_5360,N_5228,N_5210);
or U5361 (N_5361,N_5169,N_5132);
and U5362 (N_5362,N_5208,N_5235);
nor U5363 (N_5363,N_5272,N_5191);
nor U5364 (N_5364,N_5214,N_5275);
xnor U5365 (N_5365,N_5145,N_5255);
and U5366 (N_5366,N_5228,N_5175);
nand U5367 (N_5367,N_5167,N_5219);
nor U5368 (N_5368,N_5276,N_5194);
nand U5369 (N_5369,N_5232,N_5261);
nor U5370 (N_5370,N_5191,N_5216);
nor U5371 (N_5371,N_5163,N_5258);
or U5372 (N_5372,N_5222,N_5254);
or U5373 (N_5373,N_5161,N_5127);
nand U5374 (N_5374,N_5235,N_5147);
nor U5375 (N_5375,N_5124,N_5272);
nor U5376 (N_5376,N_5217,N_5259);
nor U5377 (N_5377,N_5194,N_5157);
nand U5378 (N_5378,N_5233,N_5178);
nor U5379 (N_5379,N_5240,N_5157);
and U5380 (N_5380,N_5248,N_5255);
or U5381 (N_5381,N_5160,N_5250);
or U5382 (N_5382,N_5125,N_5168);
or U5383 (N_5383,N_5210,N_5267);
nor U5384 (N_5384,N_5265,N_5260);
nor U5385 (N_5385,N_5269,N_5133);
nor U5386 (N_5386,N_5221,N_5127);
and U5387 (N_5387,N_5183,N_5273);
and U5388 (N_5388,N_5203,N_5258);
nand U5389 (N_5389,N_5262,N_5185);
and U5390 (N_5390,N_5254,N_5245);
and U5391 (N_5391,N_5256,N_5192);
and U5392 (N_5392,N_5174,N_5120);
nand U5393 (N_5393,N_5217,N_5233);
and U5394 (N_5394,N_5207,N_5185);
or U5395 (N_5395,N_5197,N_5260);
and U5396 (N_5396,N_5245,N_5164);
nand U5397 (N_5397,N_5262,N_5279);
and U5398 (N_5398,N_5137,N_5233);
and U5399 (N_5399,N_5175,N_5186);
and U5400 (N_5400,N_5244,N_5180);
or U5401 (N_5401,N_5277,N_5273);
nand U5402 (N_5402,N_5252,N_5242);
xnor U5403 (N_5403,N_5179,N_5210);
nor U5404 (N_5404,N_5260,N_5156);
or U5405 (N_5405,N_5144,N_5128);
nor U5406 (N_5406,N_5123,N_5208);
or U5407 (N_5407,N_5181,N_5127);
nor U5408 (N_5408,N_5248,N_5171);
nand U5409 (N_5409,N_5240,N_5205);
nand U5410 (N_5410,N_5186,N_5131);
nor U5411 (N_5411,N_5264,N_5199);
or U5412 (N_5412,N_5236,N_5217);
nand U5413 (N_5413,N_5237,N_5264);
or U5414 (N_5414,N_5227,N_5230);
and U5415 (N_5415,N_5228,N_5278);
or U5416 (N_5416,N_5189,N_5242);
or U5417 (N_5417,N_5278,N_5141);
xor U5418 (N_5418,N_5191,N_5219);
nand U5419 (N_5419,N_5141,N_5212);
nand U5420 (N_5420,N_5236,N_5240);
nor U5421 (N_5421,N_5241,N_5133);
or U5422 (N_5422,N_5166,N_5241);
nand U5423 (N_5423,N_5240,N_5156);
nand U5424 (N_5424,N_5213,N_5277);
and U5425 (N_5425,N_5149,N_5166);
nand U5426 (N_5426,N_5193,N_5234);
and U5427 (N_5427,N_5249,N_5183);
nand U5428 (N_5428,N_5218,N_5260);
or U5429 (N_5429,N_5137,N_5213);
xnor U5430 (N_5430,N_5221,N_5153);
and U5431 (N_5431,N_5223,N_5190);
nand U5432 (N_5432,N_5137,N_5165);
or U5433 (N_5433,N_5123,N_5197);
and U5434 (N_5434,N_5245,N_5183);
or U5435 (N_5435,N_5232,N_5213);
nand U5436 (N_5436,N_5185,N_5271);
or U5437 (N_5437,N_5196,N_5274);
and U5438 (N_5438,N_5200,N_5141);
or U5439 (N_5439,N_5266,N_5144);
or U5440 (N_5440,N_5343,N_5386);
and U5441 (N_5441,N_5307,N_5344);
nor U5442 (N_5442,N_5366,N_5355);
nor U5443 (N_5443,N_5282,N_5364);
nor U5444 (N_5444,N_5384,N_5432);
nand U5445 (N_5445,N_5362,N_5318);
nor U5446 (N_5446,N_5357,N_5289);
nor U5447 (N_5447,N_5306,N_5377);
or U5448 (N_5448,N_5397,N_5321);
nor U5449 (N_5449,N_5437,N_5418);
and U5450 (N_5450,N_5330,N_5436);
xor U5451 (N_5451,N_5373,N_5303);
nor U5452 (N_5452,N_5298,N_5398);
or U5453 (N_5453,N_5425,N_5319);
xor U5454 (N_5454,N_5288,N_5300);
and U5455 (N_5455,N_5421,N_5414);
nor U5456 (N_5456,N_5299,N_5308);
nand U5457 (N_5457,N_5345,N_5360);
and U5458 (N_5458,N_5416,N_5412);
nand U5459 (N_5459,N_5424,N_5348);
nor U5460 (N_5460,N_5375,N_5405);
nor U5461 (N_5461,N_5406,N_5356);
nor U5462 (N_5462,N_5342,N_5296);
or U5463 (N_5463,N_5391,N_5431);
nor U5464 (N_5464,N_5317,N_5326);
nand U5465 (N_5465,N_5428,N_5379);
or U5466 (N_5466,N_5291,N_5280);
and U5467 (N_5467,N_5388,N_5395);
or U5468 (N_5468,N_5337,N_5334);
and U5469 (N_5469,N_5434,N_5385);
and U5470 (N_5470,N_5336,N_5404);
or U5471 (N_5471,N_5320,N_5417);
nor U5472 (N_5472,N_5340,N_5295);
nor U5473 (N_5473,N_5323,N_5426);
or U5474 (N_5474,N_5292,N_5304);
and U5475 (N_5475,N_5314,N_5411);
nor U5476 (N_5476,N_5286,N_5420);
nor U5477 (N_5477,N_5281,N_5410);
nor U5478 (N_5478,N_5394,N_5338);
nand U5479 (N_5479,N_5302,N_5396);
and U5480 (N_5480,N_5407,N_5438);
nor U5481 (N_5481,N_5341,N_5381);
and U5482 (N_5482,N_5358,N_5389);
and U5483 (N_5483,N_5370,N_5301);
or U5484 (N_5484,N_5413,N_5402);
nor U5485 (N_5485,N_5339,N_5439);
xnor U5486 (N_5486,N_5419,N_5376);
or U5487 (N_5487,N_5369,N_5392);
nand U5488 (N_5488,N_5283,N_5287);
and U5489 (N_5489,N_5316,N_5315);
nor U5490 (N_5490,N_5427,N_5387);
nor U5491 (N_5491,N_5350,N_5312);
nor U5492 (N_5492,N_5285,N_5329);
and U5493 (N_5493,N_5313,N_5325);
and U5494 (N_5494,N_5346,N_5429);
or U5495 (N_5495,N_5328,N_5327);
nand U5496 (N_5496,N_5294,N_5349);
nand U5497 (N_5497,N_5331,N_5354);
nand U5498 (N_5498,N_5374,N_5367);
and U5499 (N_5499,N_5322,N_5290);
and U5500 (N_5500,N_5433,N_5324);
and U5501 (N_5501,N_5430,N_5365);
nand U5502 (N_5502,N_5380,N_5409);
and U5503 (N_5503,N_5305,N_5332);
xor U5504 (N_5504,N_5382,N_5353);
and U5505 (N_5505,N_5422,N_5423);
and U5506 (N_5506,N_5390,N_5371);
nand U5507 (N_5507,N_5347,N_5351);
or U5508 (N_5508,N_5372,N_5352);
xnor U5509 (N_5509,N_5399,N_5383);
nand U5510 (N_5510,N_5363,N_5393);
and U5511 (N_5511,N_5368,N_5435);
and U5512 (N_5512,N_5310,N_5361);
xnor U5513 (N_5513,N_5335,N_5284);
and U5514 (N_5514,N_5309,N_5415);
and U5515 (N_5515,N_5403,N_5401);
xor U5516 (N_5516,N_5408,N_5400);
nand U5517 (N_5517,N_5293,N_5297);
or U5518 (N_5518,N_5311,N_5333);
and U5519 (N_5519,N_5359,N_5378);
and U5520 (N_5520,N_5345,N_5379);
or U5521 (N_5521,N_5420,N_5426);
or U5522 (N_5522,N_5381,N_5407);
nor U5523 (N_5523,N_5386,N_5362);
and U5524 (N_5524,N_5303,N_5361);
and U5525 (N_5525,N_5361,N_5333);
nor U5526 (N_5526,N_5344,N_5424);
nor U5527 (N_5527,N_5358,N_5418);
and U5528 (N_5528,N_5307,N_5430);
nand U5529 (N_5529,N_5426,N_5331);
nor U5530 (N_5530,N_5333,N_5404);
nor U5531 (N_5531,N_5313,N_5353);
xor U5532 (N_5532,N_5308,N_5354);
nand U5533 (N_5533,N_5306,N_5353);
and U5534 (N_5534,N_5424,N_5357);
nor U5535 (N_5535,N_5383,N_5280);
nand U5536 (N_5536,N_5421,N_5409);
and U5537 (N_5537,N_5428,N_5411);
nand U5538 (N_5538,N_5349,N_5348);
and U5539 (N_5539,N_5397,N_5349);
and U5540 (N_5540,N_5284,N_5400);
nand U5541 (N_5541,N_5345,N_5438);
xnor U5542 (N_5542,N_5325,N_5315);
nor U5543 (N_5543,N_5288,N_5283);
and U5544 (N_5544,N_5421,N_5423);
nor U5545 (N_5545,N_5282,N_5289);
or U5546 (N_5546,N_5420,N_5357);
or U5547 (N_5547,N_5298,N_5350);
or U5548 (N_5548,N_5301,N_5309);
xor U5549 (N_5549,N_5287,N_5433);
or U5550 (N_5550,N_5298,N_5397);
nand U5551 (N_5551,N_5340,N_5404);
and U5552 (N_5552,N_5353,N_5303);
and U5553 (N_5553,N_5433,N_5434);
or U5554 (N_5554,N_5436,N_5375);
and U5555 (N_5555,N_5334,N_5411);
xnor U5556 (N_5556,N_5349,N_5306);
or U5557 (N_5557,N_5328,N_5289);
nor U5558 (N_5558,N_5409,N_5437);
nand U5559 (N_5559,N_5354,N_5300);
nor U5560 (N_5560,N_5366,N_5427);
nor U5561 (N_5561,N_5415,N_5298);
and U5562 (N_5562,N_5303,N_5405);
nor U5563 (N_5563,N_5301,N_5358);
and U5564 (N_5564,N_5314,N_5356);
and U5565 (N_5565,N_5367,N_5433);
and U5566 (N_5566,N_5420,N_5292);
and U5567 (N_5567,N_5336,N_5322);
or U5568 (N_5568,N_5336,N_5302);
nand U5569 (N_5569,N_5385,N_5340);
and U5570 (N_5570,N_5372,N_5428);
nor U5571 (N_5571,N_5288,N_5358);
and U5572 (N_5572,N_5299,N_5302);
nand U5573 (N_5573,N_5412,N_5433);
nand U5574 (N_5574,N_5427,N_5300);
nand U5575 (N_5575,N_5385,N_5343);
and U5576 (N_5576,N_5406,N_5368);
nand U5577 (N_5577,N_5285,N_5316);
or U5578 (N_5578,N_5358,N_5365);
nand U5579 (N_5579,N_5424,N_5342);
or U5580 (N_5580,N_5382,N_5306);
xor U5581 (N_5581,N_5296,N_5421);
and U5582 (N_5582,N_5306,N_5433);
and U5583 (N_5583,N_5312,N_5369);
and U5584 (N_5584,N_5370,N_5407);
nand U5585 (N_5585,N_5353,N_5370);
xor U5586 (N_5586,N_5298,N_5369);
xor U5587 (N_5587,N_5330,N_5331);
nand U5588 (N_5588,N_5287,N_5409);
or U5589 (N_5589,N_5409,N_5391);
nor U5590 (N_5590,N_5309,N_5284);
and U5591 (N_5591,N_5291,N_5337);
and U5592 (N_5592,N_5290,N_5287);
or U5593 (N_5593,N_5356,N_5288);
xor U5594 (N_5594,N_5423,N_5290);
or U5595 (N_5595,N_5340,N_5383);
nand U5596 (N_5596,N_5331,N_5365);
nor U5597 (N_5597,N_5329,N_5426);
and U5598 (N_5598,N_5375,N_5430);
nand U5599 (N_5599,N_5335,N_5321);
nor U5600 (N_5600,N_5578,N_5511);
and U5601 (N_5601,N_5461,N_5531);
and U5602 (N_5602,N_5469,N_5554);
nor U5603 (N_5603,N_5575,N_5577);
and U5604 (N_5604,N_5488,N_5523);
nor U5605 (N_5605,N_5486,N_5593);
or U5606 (N_5606,N_5499,N_5572);
nand U5607 (N_5607,N_5563,N_5579);
or U5608 (N_5608,N_5559,N_5529);
and U5609 (N_5609,N_5582,N_5494);
nor U5610 (N_5610,N_5503,N_5589);
nor U5611 (N_5611,N_5440,N_5476);
or U5612 (N_5612,N_5552,N_5448);
nor U5613 (N_5613,N_5567,N_5497);
nor U5614 (N_5614,N_5468,N_5587);
nor U5615 (N_5615,N_5447,N_5450);
nand U5616 (N_5616,N_5510,N_5576);
or U5617 (N_5617,N_5473,N_5539);
nor U5618 (N_5618,N_5547,N_5596);
nor U5619 (N_5619,N_5472,N_5508);
or U5620 (N_5620,N_5457,N_5487);
xor U5621 (N_5621,N_5588,N_5498);
or U5622 (N_5622,N_5561,N_5528);
nor U5623 (N_5623,N_5483,N_5555);
nor U5624 (N_5624,N_5568,N_5550);
or U5625 (N_5625,N_5543,N_5493);
or U5626 (N_5626,N_5479,N_5553);
xnor U5627 (N_5627,N_5522,N_5532);
nand U5628 (N_5628,N_5462,N_5548);
nor U5629 (N_5629,N_5557,N_5474);
or U5630 (N_5630,N_5592,N_5594);
nor U5631 (N_5631,N_5585,N_5590);
and U5632 (N_5632,N_5513,N_5442);
and U5633 (N_5633,N_5441,N_5455);
xnor U5634 (N_5634,N_5534,N_5507);
nand U5635 (N_5635,N_5466,N_5558);
nand U5636 (N_5636,N_5595,N_5445);
nor U5637 (N_5637,N_5453,N_5512);
or U5638 (N_5638,N_5495,N_5591);
nand U5639 (N_5639,N_5599,N_5500);
or U5640 (N_5640,N_5506,N_5485);
nand U5641 (N_5641,N_5451,N_5549);
and U5642 (N_5642,N_5516,N_5519);
nor U5643 (N_5643,N_5551,N_5533);
nor U5644 (N_5644,N_5537,N_5484);
and U5645 (N_5645,N_5454,N_5481);
nand U5646 (N_5646,N_5446,N_5584);
nand U5647 (N_5647,N_5560,N_5444);
and U5648 (N_5648,N_5460,N_5598);
xnor U5649 (N_5649,N_5489,N_5477);
nand U5650 (N_5650,N_5501,N_5562);
nor U5651 (N_5651,N_5443,N_5470);
nand U5652 (N_5652,N_5541,N_5544);
nor U5653 (N_5653,N_5574,N_5491);
xnor U5654 (N_5654,N_5545,N_5458);
or U5655 (N_5655,N_5509,N_5530);
nor U5656 (N_5656,N_5540,N_5490);
nor U5657 (N_5657,N_5535,N_5475);
nand U5658 (N_5658,N_5467,N_5526);
or U5659 (N_5659,N_5478,N_5449);
or U5660 (N_5660,N_5456,N_5465);
or U5661 (N_5661,N_5517,N_5536);
xnor U5662 (N_5662,N_5482,N_5505);
nor U5663 (N_5663,N_5542,N_5464);
nand U5664 (N_5664,N_5581,N_5471);
or U5665 (N_5665,N_5459,N_5515);
or U5666 (N_5666,N_5527,N_5463);
or U5667 (N_5667,N_5521,N_5583);
nand U5668 (N_5668,N_5586,N_5571);
nor U5669 (N_5669,N_5502,N_5538);
and U5670 (N_5670,N_5564,N_5452);
xor U5671 (N_5671,N_5580,N_5520);
or U5672 (N_5672,N_5504,N_5569);
nand U5673 (N_5673,N_5597,N_5525);
nand U5674 (N_5674,N_5546,N_5565);
and U5675 (N_5675,N_5480,N_5570);
nor U5676 (N_5676,N_5556,N_5573);
xnor U5677 (N_5677,N_5524,N_5496);
and U5678 (N_5678,N_5514,N_5518);
nand U5679 (N_5679,N_5566,N_5492);
xnor U5680 (N_5680,N_5523,N_5494);
or U5681 (N_5681,N_5519,N_5596);
and U5682 (N_5682,N_5543,N_5465);
xor U5683 (N_5683,N_5527,N_5547);
nor U5684 (N_5684,N_5519,N_5575);
or U5685 (N_5685,N_5472,N_5588);
and U5686 (N_5686,N_5575,N_5472);
nor U5687 (N_5687,N_5444,N_5593);
and U5688 (N_5688,N_5472,N_5517);
or U5689 (N_5689,N_5440,N_5586);
nand U5690 (N_5690,N_5478,N_5474);
and U5691 (N_5691,N_5487,N_5568);
or U5692 (N_5692,N_5548,N_5536);
nand U5693 (N_5693,N_5596,N_5570);
nand U5694 (N_5694,N_5528,N_5488);
nand U5695 (N_5695,N_5562,N_5535);
nand U5696 (N_5696,N_5453,N_5477);
and U5697 (N_5697,N_5589,N_5532);
nand U5698 (N_5698,N_5508,N_5468);
nand U5699 (N_5699,N_5470,N_5594);
or U5700 (N_5700,N_5540,N_5474);
and U5701 (N_5701,N_5507,N_5539);
or U5702 (N_5702,N_5597,N_5581);
and U5703 (N_5703,N_5569,N_5483);
nand U5704 (N_5704,N_5569,N_5502);
or U5705 (N_5705,N_5527,N_5452);
nand U5706 (N_5706,N_5448,N_5510);
or U5707 (N_5707,N_5592,N_5557);
or U5708 (N_5708,N_5489,N_5590);
nand U5709 (N_5709,N_5445,N_5527);
or U5710 (N_5710,N_5526,N_5557);
nor U5711 (N_5711,N_5549,N_5525);
nor U5712 (N_5712,N_5540,N_5536);
nor U5713 (N_5713,N_5463,N_5524);
nand U5714 (N_5714,N_5532,N_5491);
nor U5715 (N_5715,N_5518,N_5599);
nor U5716 (N_5716,N_5532,N_5573);
or U5717 (N_5717,N_5453,N_5571);
nor U5718 (N_5718,N_5531,N_5568);
nor U5719 (N_5719,N_5591,N_5571);
nor U5720 (N_5720,N_5524,N_5505);
and U5721 (N_5721,N_5523,N_5493);
or U5722 (N_5722,N_5463,N_5482);
nand U5723 (N_5723,N_5511,N_5576);
nor U5724 (N_5724,N_5462,N_5487);
or U5725 (N_5725,N_5483,N_5528);
and U5726 (N_5726,N_5525,N_5440);
nor U5727 (N_5727,N_5541,N_5526);
nand U5728 (N_5728,N_5530,N_5536);
and U5729 (N_5729,N_5531,N_5578);
nor U5730 (N_5730,N_5482,N_5480);
and U5731 (N_5731,N_5505,N_5558);
nor U5732 (N_5732,N_5550,N_5462);
xor U5733 (N_5733,N_5519,N_5504);
nor U5734 (N_5734,N_5514,N_5502);
or U5735 (N_5735,N_5512,N_5546);
and U5736 (N_5736,N_5574,N_5581);
and U5737 (N_5737,N_5588,N_5540);
and U5738 (N_5738,N_5576,N_5541);
or U5739 (N_5739,N_5549,N_5567);
and U5740 (N_5740,N_5589,N_5593);
or U5741 (N_5741,N_5513,N_5583);
and U5742 (N_5742,N_5573,N_5518);
nand U5743 (N_5743,N_5582,N_5599);
xnor U5744 (N_5744,N_5468,N_5478);
and U5745 (N_5745,N_5479,N_5511);
and U5746 (N_5746,N_5561,N_5487);
or U5747 (N_5747,N_5451,N_5582);
xor U5748 (N_5748,N_5557,N_5514);
nor U5749 (N_5749,N_5495,N_5520);
and U5750 (N_5750,N_5441,N_5515);
and U5751 (N_5751,N_5477,N_5599);
nand U5752 (N_5752,N_5453,N_5580);
or U5753 (N_5753,N_5598,N_5471);
nand U5754 (N_5754,N_5521,N_5447);
and U5755 (N_5755,N_5520,N_5509);
xnor U5756 (N_5756,N_5490,N_5469);
nor U5757 (N_5757,N_5527,N_5553);
or U5758 (N_5758,N_5530,N_5443);
xnor U5759 (N_5759,N_5556,N_5550);
nor U5760 (N_5760,N_5713,N_5670);
nand U5761 (N_5761,N_5619,N_5671);
nor U5762 (N_5762,N_5627,N_5641);
and U5763 (N_5763,N_5733,N_5697);
nand U5764 (N_5764,N_5633,N_5726);
nand U5765 (N_5765,N_5658,N_5661);
or U5766 (N_5766,N_5637,N_5605);
and U5767 (N_5767,N_5604,N_5652);
xor U5768 (N_5768,N_5752,N_5701);
or U5769 (N_5769,N_5738,N_5756);
nand U5770 (N_5770,N_5629,N_5741);
or U5771 (N_5771,N_5727,N_5721);
nor U5772 (N_5772,N_5609,N_5690);
and U5773 (N_5773,N_5606,N_5612);
xor U5774 (N_5774,N_5646,N_5755);
or U5775 (N_5775,N_5618,N_5615);
nor U5776 (N_5776,N_5685,N_5695);
or U5777 (N_5777,N_5630,N_5711);
nand U5778 (N_5778,N_5736,N_5636);
and U5779 (N_5779,N_5718,N_5719);
xor U5780 (N_5780,N_5600,N_5623);
and U5781 (N_5781,N_5684,N_5621);
nor U5782 (N_5782,N_5696,N_5674);
nand U5783 (N_5783,N_5745,N_5643);
or U5784 (N_5784,N_5626,N_5645);
nor U5785 (N_5785,N_5679,N_5642);
or U5786 (N_5786,N_5707,N_5632);
nand U5787 (N_5787,N_5634,N_5617);
or U5788 (N_5788,N_5704,N_5700);
and U5789 (N_5789,N_5675,N_5740);
or U5790 (N_5790,N_5725,N_5724);
xor U5791 (N_5791,N_5625,N_5759);
nand U5792 (N_5792,N_5687,N_5706);
and U5793 (N_5793,N_5691,N_5620);
xor U5794 (N_5794,N_5639,N_5729);
nor U5795 (N_5795,N_5657,N_5667);
xor U5796 (N_5796,N_5666,N_5716);
nand U5797 (N_5797,N_5688,N_5659);
nor U5798 (N_5798,N_5715,N_5672);
and U5799 (N_5799,N_5747,N_5673);
nor U5800 (N_5800,N_5603,N_5647);
nand U5801 (N_5801,N_5631,N_5744);
nand U5802 (N_5802,N_5693,N_5757);
or U5803 (N_5803,N_5677,N_5710);
and U5804 (N_5804,N_5720,N_5653);
nor U5805 (N_5805,N_5692,N_5709);
and U5806 (N_5806,N_5686,N_5601);
or U5807 (N_5807,N_5610,N_5616);
nor U5808 (N_5808,N_5699,N_5735);
or U5809 (N_5809,N_5739,N_5654);
xnor U5810 (N_5810,N_5742,N_5705);
and U5811 (N_5811,N_5614,N_5669);
and U5812 (N_5812,N_5743,N_5753);
or U5813 (N_5813,N_5608,N_5731);
nor U5814 (N_5814,N_5655,N_5728);
and U5815 (N_5815,N_5613,N_5681);
or U5816 (N_5816,N_5751,N_5648);
or U5817 (N_5817,N_5664,N_5734);
nor U5818 (N_5818,N_5611,N_5624);
or U5819 (N_5819,N_5678,N_5732);
and U5820 (N_5820,N_5662,N_5714);
nor U5821 (N_5821,N_5665,N_5656);
and U5822 (N_5822,N_5622,N_5676);
nor U5823 (N_5823,N_5628,N_5703);
or U5824 (N_5824,N_5723,N_5694);
or U5825 (N_5825,N_5644,N_5660);
xnor U5826 (N_5826,N_5649,N_5638);
or U5827 (N_5827,N_5640,N_5749);
and U5828 (N_5828,N_5746,N_5712);
nor U5829 (N_5829,N_5750,N_5722);
nor U5830 (N_5830,N_5635,N_5682);
nor U5831 (N_5831,N_5754,N_5698);
nor U5832 (N_5832,N_5737,N_5602);
nand U5833 (N_5833,N_5708,N_5717);
or U5834 (N_5834,N_5663,N_5651);
nand U5835 (N_5835,N_5683,N_5748);
nor U5836 (N_5836,N_5702,N_5680);
nand U5837 (N_5837,N_5607,N_5689);
or U5838 (N_5838,N_5758,N_5650);
nand U5839 (N_5839,N_5668,N_5730);
nand U5840 (N_5840,N_5621,N_5630);
nor U5841 (N_5841,N_5690,N_5711);
and U5842 (N_5842,N_5739,N_5683);
nor U5843 (N_5843,N_5639,N_5691);
xnor U5844 (N_5844,N_5734,N_5603);
nor U5845 (N_5845,N_5749,N_5642);
and U5846 (N_5846,N_5716,N_5695);
or U5847 (N_5847,N_5699,N_5672);
nor U5848 (N_5848,N_5740,N_5642);
xnor U5849 (N_5849,N_5619,N_5700);
or U5850 (N_5850,N_5690,N_5640);
nor U5851 (N_5851,N_5698,N_5666);
nand U5852 (N_5852,N_5651,N_5664);
nor U5853 (N_5853,N_5659,N_5626);
nor U5854 (N_5854,N_5731,N_5698);
or U5855 (N_5855,N_5670,N_5717);
or U5856 (N_5856,N_5656,N_5623);
and U5857 (N_5857,N_5601,N_5711);
nor U5858 (N_5858,N_5647,N_5666);
nand U5859 (N_5859,N_5742,N_5737);
nand U5860 (N_5860,N_5611,N_5614);
or U5861 (N_5861,N_5750,N_5635);
and U5862 (N_5862,N_5637,N_5604);
and U5863 (N_5863,N_5678,N_5759);
or U5864 (N_5864,N_5737,N_5608);
nand U5865 (N_5865,N_5704,N_5746);
nand U5866 (N_5866,N_5672,N_5704);
and U5867 (N_5867,N_5627,N_5728);
or U5868 (N_5868,N_5640,N_5604);
or U5869 (N_5869,N_5626,N_5729);
nand U5870 (N_5870,N_5752,N_5622);
nor U5871 (N_5871,N_5646,N_5718);
and U5872 (N_5872,N_5718,N_5602);
nand U5873 (N_5873,N_5692,N_5734);
and U5874 (N_5874,N_5668,N_5646);
and U5875 (N_5875,N_5742,N_5664);
nand U5876 (N_5876,N_5756,N_5658);
or U5877 (N_5877,N_5680,N_5673);
and U5878 (N_5878,N_5653,N_5648);
or U5879 (N_5879,N_5756,N_5612);
xnor U5880 (N_5880,N_5718,N_5723);
or U5881 (N_5881,N_5689,N_5636);
and U5882 (N_5882,N_5699,N_5642);
nor U5883 (N_5883,N_5747,N_5663);
xor U5884 (N_5884,N_5708,N_5753);
nand U5885 (N_5885,N_5739,N_5691);
nand U5886 (N_5886,N_5613,N_5724);
nand U5887 (N_5887,N_5630,N_5633);
nor U5888 (N_5888,N_5613,N_5635);
and U5889 (N_5889,N_5634,N_5743);
nor U5890 (N_5890,N_5735,N_5747);
nor U5891 (N_5891,N_5632,N_5619);
xnor U5892 (N_5892,N_5671,N_5720);
nand U5893 (N_5893,N_5681,N_5733);
or U5894 (N_5894,N_5626,N_5711);
or U5895 (N_5895,N_5721,N_5623);
or U5896 (N_5896,N_5745,N_5612);
nand U5897 (N_5897,N_5698,N_5719);
or U5898 (N_5898,N_5712,N_5753);
and U5899 (N_5899,N_5678,N_5610);
and U5900 (N_5900,N_5656,N_5644);
and U5901 (N_5901,N_5736,N_5713);
nor U5902 (N_5902,N_5626,N_5735);
or U5903 (N_5903,N_5731,N_5695);
and U5904 (N_5904,N_5623,N_5750);
and U5905 (N_5905,N_5658,N_5643);
and U5906 (N_5906,N_5709,N_5636);
xor U5907 (N_5907,N_5601,N_5640);
or U5908 (N_5908,N_5657,N_5741);
xor U5909 (N_5909,N_5663,N_5646);
and U5910 (N_5910,N_5666,N_5686);
or U5911 (N_5911,N_5665,N_5600);
xor U5912 (N_5912,N_5669,N_5689);
xor U5913 (N_5913,N_5708,N_5694);
nor U5914 (N_5914,N_5732,N_5623);
nor U5915 (N_5915,N_5674,N_5650);
and U5916 (N_5916,N_5727,N_5616);
and U5917 (N_5917,N_5677,N_5631);
and U5918 (N_5918,N_5678,N_5641);
and U5919 (N_5919,N_5680,N_5723);
nand U5920 (N_5920,N_5819,N_5873);
or U5921 (N_5921,N_5863,N_5768);
xnor U5922 (N_5922,N_5868,N_5916);
or U5923 (N_5923,N_5856,N_5893);
or U5924 (N_5924,N_5816,N_5882);
and U5925 (N_5925,N_5844,N_5903);
nor U5926 (N_5926,N_5912,N_5778);
nor U5927 (N_5927,N_5799,N_5794);
or U5928 (N_5928,N_5765,N_5811);
nor U5929 (N_5929,N_5793,N_5814);
or U5930 (N_5930,N_5866,N_5766);
xnor U5931 (N_5931,N_5853,N_5786);
nor U5932 (N_5932,N_5895,N_5802);
or U5933 (N_5933,N_5810,N_5909);
nand U5934 (N_5934,N_5854,N_5845);
nor U5935 (N_5935,N_5847,N_5874);
or U5936 (N_5936,N_5869,N_5776);
or U5937 (N_5937,N_5795,N_5907);
and U5938 (N_5938,N_5889,N_5911);
and U5939 (N_5939,N_5910,N_5904);
nor U5940 (N_5940,N_5838,N_5783);
and U5941 (N_5941,N_5823,N_5867);
nand U5942 (N_5942,N_5846,N_5803);
and U5943 (N_5943,N_5821,N_5900);
or U5944 (N_5944,N_5851,N_5773);
or U5945 (N_5945,N_5862,N_5859);
nor U5946 (N_5946,N_5858,N_5800);
nor U5947 (N_5947,N_5809,N_5798);
nor U5948 (N_5948,N_5788,N_5840);
nor U5949 (N_5949,N_5781,N_5843);
and U5950 (N_5950,N_5870,N_5899);
nor U5951 (N_5951,N_5782,N_5892);
nor U5952 (N_5952,N_5855,N_5864);
nand U5953 (N_5953,N_5876,N_5825);
or U5954 (N_5954,N_5877,N_5852);
nand U5955 (N_5955,N_5771,N_5784);
nor U5956 (N_5956,N_5818,N_5914);
nand U5957 (N_5957,N_5774,N_5761);
nor U5958 (N_5958,N_5913,N_5790);
nand U5959 (N_5959,N_5762,N_5850);
and U5960 (N_5960,N_5832,N_5906);
or U5961 (N_5961,N_5772,N_5836);
nor U5962 (N_5962,N_5769,N_5839);
or U5963 (N_5963,N_5806,N_5861);
nor U5964 (N_5964,N_5901,N_5787);
and U5965 (N_5965,N_5808,N_5890);
nand U5966 (N_5966,N_5883,N_5831);
nand U5967 (N_5967,N_5849,N_5815);
nand U5968 (N_5968,N_5807,N_5887);
or U5969 (N_5969,N_5865,N_5841);
or U5970 (N_5970,N_5860,N_5898);
nor U5971 (N_5971,N_5760,N_5896);
or U5972 (N_5972,N_5777,N_5881);
nand U5973 (N_5973,N_5791,N_5875);
nor U5974 (N_5974,N_5812,N_5779);
nand U5975 (N_5975,N_5908,N_5894);
nand U5976 (N_5976,N_5820,N_5785);
xor U5977 (N_5977,N_5872,N_5822);
and U5978 (N_5978,N_5780,N_5888);
nand U5979 (N_5979,N_5834,N_5789);
or U5980 (N_5980,N_5770,N_5792);
nor U5981 (N_5981,N_5767,N_5835);
nand U5982 (N_5982,N_5830,N_5897);
nor U5983 (N_5983,N_5902,N_5891);
nand U5984 (N_5984,N_5824,N_5917);
or U5985 (N_5985,N_5918,N_5884);
or U5986 (N_5986,N_5919,N_5905);
xor U5987 (N_5987,N_5796,N_5817);
and U5988 (N_5988,N_5842,N_5885);
or U5989 (N_5989,N_5880,N_5837);
xor U5990 (N_5990,N_5813,N_5915);
nor U5991 (N_5991,N_5763,N_5805);
nand U5992 (N_5992,N_5797,N_5886);
nand U5993 (N_5993,N_5826,N_5857);
nand U5994 (N_5994,N_5828,N_5833);
and U5995 (N_5995,N_5871,N_5801);
nor U5996 (N_5996,N_5764,N_5879);
or U5997 (N_5997,N_5775,N_5829);
and U5998 (N_5998,N_5848,N_5804);
and U5999 (N_5999,N_5878,N_5827);
nor U6000 (N_6000,N_5916,N_5827);
nand U6001 (N_6001,N_5827,N_5773);
or U6002 (N_6002,N_5814,N_5889);
and U6003 (N_6003,N_5831,N_5916);
and U6004 (N_6004,N_5891,N_5918);
and U6005 (N_6005,N_5890,N_5868);
nor U6006 (N_6006,N_5765,N_5884);
xnor U6007 (N_6007,N_5842,N_5769);
nor U6008 (N_6008,N_5892,N_5875);
nand U6009 (N_6009,N_5799,N_5782);
and U6010 (N_6010,N_5774,N_5855);
nand U6011 (N_6011,N_5869,N_5840);
and U6012 (N_6012,N_5868,N_5766);
or U6013 (N_6013,N_5793,N_5903);
xnor U6014 (N_6014,N_5810,N_5854);
nor U6015 (N_6015,N_5825,N_5820);
or U6016 (N_6016,N_5860,N_5801);
nand U6017 (N_6017,N_5877,N_5831);
and U6018 (N_6018,N_5838,N_5842);
nand U6019 (N_6019,N_5885,N_5847);
or U6020 (N_6020,N_5876,N_5834);
nor U6021 (N_6021,N_5866,N_5896);
or U6022 (N_6022,N_5770,N_5911);
nor U6023 (N_6023,N_5791,N_5877);
xnor U6024 (N_6024,N_5796,N_5861);
or U6025 (N_6025,N_5875,N_5804);
and U6026 (N_6026,N_5827,N_5808);
or U6027 (N_6027,N_5764,N_5914);
and U6028 (N_6028,N_5868,N_5850);
nand U6029 (N_6029,N_5864,N_5868);
or U6030 (N_6030,N_5874,N_5767);
nand U6031 (N_6031,N_5828,N_5805);
nand U6032 (N_6032,N_5907,N_5893);
or U6033 (N_6033,N_5836,N_5840);
and U6034 (N_6034,N_5870,N_5874);
nor U6035 (N_6035,N_5778,N_5891);
and U6036 (N_6036,N_5915,N_5857);
or U6037 (N_6037,N_5905,N_5867);
nor U6038 (N_6038,N_5827,N_5919);
or U6039 (N_6039,N_5867,N_5860);
or U6040 (N_6040,N_5909,N_5798);
and U6041 (N_6041,N_5783,N_5814);
or U6042 (N_6042,N_5878,N_5803);
or U6043 (N_6043,N_5777,N_5837);
nor U6044 (N_6044,N_5815,N_5844);
nor U6045 (N_6045,N_5919,N_5810);
and U6046 (N_6046,N_5776,N_5899);
and U6047 (N_6047,N_5860,N_5834);
nor U6048 (N_6048,N_5836,N_5841);
nor U6049 (N_6049,N_5869,N_5811);
nor U6050 (N_6050,N_5867,N_5802);
nor U6051 (N_6051,N_5847,N_5852);
and U6052 (N_6052,N_5869,N_5822);
nand U6053 (N_6053,N_5888,N_5893);
or U6054 (N_6054,N_5915,N_5850);
nor U6055 (N_6055,N_5801,N_5838);
nand U6056 (N_6056,N_5813,N_5822);
nand U6057 (N_6057,N_5906,N_5836);
or U6058 (N_6058,N_5832,N_5786);
and U6059 (N_6059,N_5841,N_5906);
or U6060 (N_6060,N_5776,N_5875);
nand U6061 (N_6061,N_5853,N_5825);
nor U6062 (N_6062,N_5833,N_5902);
and U6063 (N_6063,N_5822,N_5792);
or U6064 (N_6064,N_5794,N_5893);
nand U6065 (N_6065,N_5829,N_5785);
nand U6066 (N_6066,N_5815,N_5863);
nand U6067 (N_6067,N_5915,N_5836);
nand U6068 (N_6068,N_5799,N_5858);
nor U6069 (N_6069,N_5799,N_5797);
and U6070 (N_6070,N_5829,N_5772);
xnor U6071 (N_6071,N_5831,N_5858);
or U6072 (N_6072,N_5795,N_5772);
or U6073 (N_6073,N_5779,N_5789);
and U6074 (N_6074,N_5860,N_5905);
nand U6075 (N_6075,N_5892,N_5761);
nand U6076 (N_6076,N_5912,N_5858);
nand U6077 (N_6077,N_5767,N_5794);
and U6078 (N_6078,N_5836,N_5852);
or U6079 (N_6079,N_5868,N_5829);
nand U6080 (N_6080,N_5936,N_5968);
nor U6081 (N_6081,N_5971,N_6032);
or U6082 (N_6082,N_6070,N_6048);
xnor U6083 (N_6083,N_5935,N_6064);
and U6084 (N_6084,N_6075,N_6046);
nand U6085 (N_6085,N_6050,N_5977);
xnor U6086 (N_6086,N_6010,N_6066);
or U6087 (N_6087,N_5993,N_5982);
and U6088 (N_6088,N_5948,N_5926);
nor U6089 (N_6089,N_5942,N_6056);
and U6090 (N_6090,N_6001,N_5974);
nor U6091 (N_6091,N_6041,N_5945);
nand U6092 (N_6092,N_6038,N_5985);
and U6093 (N_6093,N_5959,N_6042);
nand U6094 (N_6094,N_5949,N_5998);
nand U6095 (N_6095,N_6055,N_6009);
and U6096 (N_6096,N_6030,N_6003);
nand U6097 (N_6097,N_6018,N_5995);
or U6098 (N_6098,N_5920,N_6026);
nand U6099 (N_6099,N_5962,N_6019);
nand U6100 (N_6100,N_6051,N_6044);
or U6101 (N_6101,N_6035,N_6036);
and U6102 (N_6102,N_5930,N_6023);
nor U6103 (N_6103,N_5996,N_6014);
xor U6104 (N_6104,N_6021,N_5992);
nand U6105 (N_6105,N_5956,N_6079);
nand U6106 (N_6106,N_6060,N_5939);
and U6107 (N_6107,N_5955,N_6063);
nand U6108 (N_6108,N_6008,N_5989);
nand U6109 (N_6109,N_6004,N_6013);
nand U6110 (N_6110,N_5951,N_5938);
nand U6111 (N_6111,N_5966,N_6022);
nand U6112 (N_6112,N_5922,N_5929);
and U6113 (N_6113,N_5967,N_5983);
or U6114 (N_6114,N_5970,N_5927);
and U6115 (N_6115,N_5941,N_5997);
or U6116 (N_6116,N_6054,N_5944);
or U6117 (N_6117,N_5924,N_5961);
xor U6118 (N_6118,N_6061,N_5990);
xnor U6119 (N_6119,N_5972,N_6011);
nand U6120 (N_6120,N_6074,N_6033);
or U6121 (N_6121,N_5925,N_5931);
nand U6122 (N_6122,N_6073,N_5973);
nor U6123 (N_6123,N_6062,N_6024);
nor U6124 (N_6124,N_5940,N_5932);
nand U6125 (N_6125,N_5947,N_5980);
nand U6126 (N_6126,N_6067,N_6005);
nand U6127 (N_6127,N_6012,N_6031);
nand U6128 (N_6128,N_5960,N_5987);
or U6129 (N_6129,N_6006,N_6000);
or U6130 (N_6130,N_5937,N_6049);
or U6131 (N_6131,N_6039,N_6007);
and U6132 (N_6132,N_6052,N_6034);
nor U6133 (N_6133,N_5984,N_6077);
and U6134 (N_6134,N_5957,N_5965);
and U6135 (N_6135,N_6043,N_5988);
nor U6136 (N_6136,N_6025,N_6078);
or U6137 (N_6137,N_5933,N_6068);
or U6138 (N_6138,N_5975,N_5928);
or U6139 (N_6139,N_5986,N_5923);
nand U6140 (N_6140,N_6027,N_5921);
and U6141 (N_6141,N_6059,N_5976);
nand U6142 (N_6142,N_5950,N_6037);
xnor U6143 (N_6143,N_6058,N_5946);
nand U6144 (N_6144,N_6002,N_6071);
and U6145 (N_6145,N_6015,N_5979);
nand U6146 (N_6146,N_5994,N_5954);
nor U6147 (N_6147,N_6045,N_5981);
and U6148 (N_6148,N_6029,N_5964);
and U6149 (N_6149,N_5991,N_6017);
nand U6150 (N_6150,N_6076,N_6020);
nand U6151 (N_6151,N_5958,N_6047);
nand U6152 (N_6152,N_5953,N_5943);
nor U6153 (N_6153,N_5978,N_6016);
nand U6154 (N_6154,N_6072,N_5969);
nor U6155 (N_6155,N_6069,N_6028);
nand U6156 (N_6156,N_6053,N_6057);
xnor U6157 (N_6157,N_5952,N_6040);
nor U6158 (N_6158,N_6065,N_5934);
or U6159 (N_6159,N_5999,N_5963);
or U6160 (N_6160,N_5949,N_6037);
and U6161 (N_6161,N_6005,N_6034);
nor U6162 (N_6162,N_6003,N_5959);
or U6163 (N_6163,N_6047,N_6043);
nand U6164 (N_6164,N_6021,N_5950);
nor U6165 (N_6165,N_5965,N_5942);
xnor U6166 (N_6166,N_5975,N_6050);
nand U6167 (N_6167,N_5991,N_5937);
nor U6168 (N_6168,N_6028,N_5955);
xnor U6169 (N_6169,N_6066,N_6068);
nor U6170 (N_6170,N_5976,N_5923);
nor U6171 (N_6171,N_6042,N_6016);
and U6172 (N_6172,N_5971,N_6042);
nor U6173 (N_6173,N_5946,N_6070);
nand U6174 (N_6174,N_6018,N_6024);
nand U6175 (N_6175,N_6049,N_6011);
xnor U6176 (N_6176,N_5952,N_6073);
and U6177 (N_6177,N_6052,N_6006);
nand U6178 (N_6178,N_5998,N_5920);
xor U6179 (N_6179,N_5989,N_5944);
nand U6180 (N_6180,N_5965,N_6007);
nand U6181 (N_6181,N_5956,N_5948);
and U6182 (N_6182,N_5978,N_6049);
or U6183 (N_6183,N_5991,N_6007);
xor U6184 (N_6184,N_6026,N_6046);
nor U6185 (N_6185,N_6066,N_6078);
xor U6186 (N_6186,N_5932,N_5969);
and U6187 (N_6187,N_6063,N_5973);
xor U6188 (N_6188,N_5954,N_5941);
nor U6189 (N_6189,N_5973,N_6067);
or U6190 (N_6190,N_6072,N_6008);
nor U6191 (N_6191,N_5984,N_5978);
nor U6192 (N_6192,N_6041,N_5965);
nor U6193 (N_6193,N_5976,N_5965);
xnor U6194 (N_6194,N_5939,N_6042);
or U6195 (N_6195,N_6021,N_6014);
or U6196 (N_6196,N_6025,N_5962);
xor U6197 (N_6197,N_5999,N_5950);
and U6198 (N_6198,N_5953,N_6023);
nor U6199 (N_6199,N_5925,N_5999);
nor U6200 (N_6200,N_6050,N_5994);
or U6201 (N_6201,N_5959,N_5932);
nor U6202 (N_6202,N_5974,N_6060);
and U6203 (N_6203,N_5959,N_6026);
nand U6204 (N_6204,N_6051,N_5970);
or U6205 (N_6205,N_5950,N_5956);
and U6206 (N_6206,N_5955,N_5940);
xnor U6207 (N_6207,N_6065,N_5960);
nand U6208 (N_6208,N_6020,N_5962);
and U6209 (N_6209,N_6060,N_6032);
nand U6210 (N_6210,N_5943,N_5942);
xor U6211 (N_6211,N_5958,N_6020);
or U6212 (N_6212,N_6070,N_6006);
or U6213 (N_6213,N_5938,N_5987);
nor U6214 (N_6214,N_6053,N_5923);
xor U6215 (N_6215,N_6067,N_5948);
and U6216 (N_6216,N_5921,N_6008);
and U6217 (N_6217,N_5942,N_5921);
or U6218 (N_6218,N_5930,N_6061);
or U6219 (N_6219,N_6059,N_5968);
or U6220 (N_6220,N_6018,N_5977);
or U6221 (N_6221,N_5943,N_5947);
xor U6222 (N_6222,N_5997,N_6079);
and U6223 (N_6223,N_5923,N_5947);
nand U6224 (N_6224,N_5966,N_6066);
and U6225 (N_6225,N_5938,N_6032);
and U6226 (N_6226,N_6078,N_6048);
xor U6227 (N_6227,N_6071,N_6025);
nand U6228 (N_6228,N_6034,N_6047);
nor U6229 (N_6229,N_5948,N_5975);
nor U6230 (N_6230,N_6008,N_5926);
nand U6231 (N_6231,N_5928,N_5966);
nand U6232 (N_6232,N_5996,N_5922);
or U6233 (N_6233,N_6017,N_6032);
nand U6234 (N_6234,N_6023,N_5941);
nor U6235 (N_6235,N_6035,N_5942);
nand U6236 (N_6236,N_6035,N_6071);
xnor U6237 (N_6237,N_6011,N_5923);
and U6238 (N_6238,N_5974,N_6026);
and U6239 (N_6239,N_6020,N_5979);
nor U6240 (N_6240,N_6156,N_6148);
nand U6241 (N_6241,N_6161,N_6147);
nand U6242 (N_6242,N_6230,N_6192);
nand U6243 (N_6243,N_6091,N_6179);
or U6244 (N_6244,N_6218,N_6126);
and U6245 (N_6245,N_6206,N_6116);
nand U6246 (N_6246,N_6088,N_6202);
and U6247 (N_6247,N_6210,N_6085);
or U6248 (N_6248,N_6146,N_6086);
or U6249 (N_6249,N_6190,N_6196);
nand U6250 (N_6250,N_6193,N_6205);
nand U6251 (N_6251,N_6168,N_6159);
or U6252 (N_6252,N_6098,N_6106);
nor U6253 (N_6253,N_6092,N_6133);
and U6254 (N_6254,N_6233,N_6109);
nand U6255 (N_6255,N_6110,N_6171);
or U6256 (N_6256,N_6203,N_6219);
or U6257 (N_6257,N_6238,N_6103);
or U6258 (N_6258,N_6199,N_6142);
nor U6259 (N_6259,N_6151,N_6144);
nor U6260 (N_6260,N_6130,N_6225);
nand U6261 (N_6261,N_6181,N_6084);
nor U6262 (N_6262,N_6154,N_6224);
and U6263 (N_6263,N_6176,N_6235);
nand U6264 (N_6264,N_6215,N_6163);
xnor U6265 (N_6265,N_6239,N_6195);
or U6266 (N_6266,N_6090,N_6152);
and U6267 (N_6267,N_6119,N_6102);
nand U6268 (N_6268,N_6115,N_6214);
nand U6269 (N_6269,N_6234,N_6172);
or U6270 (N_6270,N_6112,N_6157);
and U6271 (N_6271,N_6138,N_6182);
or U6272 (N_6272,N_6140,N_6134);
nor U6273 (N_6273,N_6155,N_6213);
or U6274 (N_6274,N_6178,N_6167);
and U6275 (N_6275,N_6096,N_6204);
nor U6276 (N_6276,N_6137,N_6093);
xor U6277 (N_6277,N_6217,N_6207);
nor U6278 (N_6278,N_6097,N_6122);
or U6279 (N_6279,N_6127,N_6183);
nor U6280 (N_6280,N_6114,N_6211);
nor U6281 (N_6281,N_6132,N_6177);
nand U6282 (N_6282,N_6105,N_6180);
or U6283 (N_6283,N_6185,N_6222);
xnor U6284 (N_6284,N_6221,N_6123);
nand U6285 (N_6285,N_6162,N_6125);
nor U6286 (N_6286,N_6186,N_6153);
xor U6287 (N_6287,N_6216,N_6191);
nand U6288 (N_6288,N_6173,N_6107);
and U6289 (N_6289,N_6184,N_6111);
and U6290 (N_6290,N_6228,N_6081);
and U6291 (N_6291,N_6229,N_6220);
nand U6292 (N_6292,N_6200,N_6170);
and U6293 (N_6293,N_6139,N_6095);
xnor U6294 (N_6294,N_6201,N_6209);
nand U6295 (N_6295,N_6121,N_6197);
nor U6296 (N_6296,N_6141,N_6124);
and U6297 (N_6297,N_6194,N_6113);
nand U6298 (N_6298,N_6231,N_6188);
or U6299 (N_6299,N_6120,N_6117);
xnor U6300 (N_6300,N_6237,N_6087);
nor U6301 (N_6301,N_6083,N_6080);
xnor U6302 (N_6302,N_6135,N_6128);
and U6303 (N_6303,N_6089,N_6212);
nand U6304 (N_6304,N_6198,N_6108);
or U6305 (N_6305,N_6169,N_6104);
and U6306 (N_6306,N_6165,N_6149);
and U6307 (N_6307,N_6129,N_6164);
or U6308 (N_6308,N_6158,N_6160);
or U6309 (N_6309,N_6227,N_6166);
and U6310 (N_6310,N_6208,N_6187);
and U6311 (N_6311,N_6150,N_6145);
and U6312 (N_6312,N_6236,N_6099);
nand U6313 (N_6313,N_6189,N_6223);
or U6314 (N_6314,N_6118,N_6136);
xnor U6315 (N_6315,N_6101,N_6175);
nand U6316 (N_6316,N_6226,N_6232);
nor U6317 (N_6317,N_6131,N_6143);
xnor U6318 (N_6318,N_6082,N_6100);
or U6319 (N_6319,N_6174,N_6094);
and U6320 (N_6320,N_6195,N_6085);
nor U6321 (N_6321,N_6177,N_6123);
nor U6322 (N_6322,N_6169,N_6140);
and U6323 (N_6323,N_6163,N_6091);
nand U6324 (N_6324,N_6153,N_6204);
xnor U6325 (N_6325,N_6106,N_6229);
and U6326 (N_6326,N_6118,N_6153);
and U6327 (N_6327,N_6091,N_6111);
nand U6328 (N_6328,N_6171,N_6218);
xnor U6329 (N_6329,N_6152,N_6092);
and U6330 (N_6330,N_6167,N_6194);
or U6331 (N_6331,N_6166,N_6211);
nand U6332 (N_6332,N_6211,N_6208);
nand U6333 (N_6333,N_6180,N_6191);
or U6334 (N_6334,N_6205,N_6190);
xnor U6335 (N_6335,N_6097,N_6123);
or U6336 (N_6336,N_6190,N_6212);
nor U6337 (N_6337,N_6098,N_6172);
nor U6338 (N_6338,N_6211,N_6127);
nand U6339 (N_6339,N_6197,N_6231);
and U6340 (N_6340,N_6110,N_6142);
or U6341 (N_6341,N_6178,N_6150);
and U6342 (N_6342,N_6229,N_6230);
nand U6343 (N_6343,N_6232,N_6089);
or U6344 (N_6344,N_6189,N_6202);
and U6345 (N_6345,N_6216,N_6217);
nor U6346 (N_6346,N_6123,N_6083);
xor U6347 (N_6347,N_6183,N_6202);
or U6348 (N_6348,N_6082,N_6123);
nor U6349 (N_6349,N_6182,N_6152);
nor U6350 (N_6350,N_6174,N_6226);
or U6351 (N_6351,N_6143,N_6118);
nand U6352 (N_6352,N_6099,N_6172);
nand U6353 (N_6353,N_6137,N_6156);
or U6354 (N_6354,N_6177,N_6197);
xor U6355 (N_6355,N_6218,N_6203);
and U6356 (N_6356,N_6124,N_6162);
nand U6357 (N_6357,N_6095,N_6104);
nor U6358 (N_6358,N_6221,N_6169);
and U6359 (N_6359,N_6182,N_6160);
or U6360 (N_6360,N_6127,N_6153);
nor U6361 (N_6361,N_6214,N_6143);
nor U6362 (N_6362,N_6092,N_6225);
or U6363 (N_6363,N_6103,N_6115);
and U6364 (N_6364,N_6173,N_6227);
xnor U6365 (N_6365,N_6185,N_6197);
and U6366 (N_6366,N_6221,N_6100);
nand U6367 (N_6367,N_6162,N_6100);
nor U6368 (N_6368,N_6215,N_6089);
nand U6369 (N_6369,N_6234,N_6216);
or U6370 (N_6370,N_6200,N_6142);
nor U6371 (N_6371,N_6080,N_6118);
and U6372 (N_6372,N_6142,N_6083);
or U6373 (N_6373,N_6163,N_6231);
nand U6374 (N_6374,N_6192,N_6111);
nand U6375 (N_6375,N_6222,N_6111);
nor U6376 (N_6376,N_6124,N_6136);
and U6377 (N_6377,N_6109,N_6127);
nor U6378 (N_6378,N_6125,N_6168);
nand U6379 (N_6379,N_6236,N_6133);
or U6380 (N_6380,N_6113,N_6115);
nand U6381 (N_6381,N_6163,N_6094);
nor U6382 (N_6382,N_6081,N_6225);
nor U6383 (N_6383,N_6118,N_6130);
and U6384 (N_6384,N_6082,N_6210);
and U6385 (N_6385,N_6185,N_6228);
nor U6386 (N_6386,N_6239,N_6127);
and U6387 (N_6387,N_6202,N_6106);
and U6388 (N_6388,N_6120,N_6105);
nor U6389 (N_6389,N_6138,N_6086);
nand U6390 (N_6390,N_6125,N_6148);
or U6391 (N_6391,N_6185,N_6182);
xnor U6392 (N_6392,N_6188,N_6140);
or U6393 (N_6393,N_6101,N_6131);
nor U6394 (N_6394,N_6228,N_6149);
nand U6395 (N_6395,N_6183,N_6195);
nor U6396 (N_6396,N_6101,N_6171);
xnor U6397 (N_6397,N_6190,N_6152);
or U6398 (N_6398,N_6178,N_6220);
or U6399 (N_6399,N_6134,N_6177);
nor U6400 (N_6400,N_6309,N_6324);
or U6401 (N_6401,N_6285,N_6364);
nand U6402 (N_6402,N_6359,N_6339);
nor U6403 (N_6403,N_6299,N_6263);
and U6404 (N_6404,N_6286,N_6280);
xor U6405 (N_6405,N_6396,N_6255);
nor U6406 (N_6406,N_6308,N_6321);
nand U6407 (N_6407,N_6391,N_6262);
xnor U6408 (N_6408,N_6294,N_6358);
nor U6409 (N_6409,N_6398,N_6272);
nor U6410 (N_6410,N_6245,N_6270);
and U6411 (N_6411,N_6352,N_6265);
and U6412 (N_6412,N_6283,N_6357);
nor U6413 (N_6413,N_6348,N_6292);
xor U6414 (N_6414,N_6327,N_6397);
nand U6415 (N_6415,N_6340,N_6378);
or U6416 (N_6416,N_6244,N_6363);
and U6417 (N_6417,N_6296,N_6287);
xnor U6418 (N_6418,N_6269,N_6304);
xor U6419 (N_6419,N_6344,N_6250);
nor U6420 (N_6420,N_6284,N_6356);
xor U6421 (N_6421,N_6350,N_6384);
nor U6422 (N_6422,N_6318,N_6257);
or U6423 (N_6423,N_6342,N_6277);
and U6424 (N_6424,N_6387,N_6249);
xor U6425 (N_6425,N_6345,N_6382);
and U6426 (N_6426,N_6389,N_6349);
and U6427 (N_6427,N_6298,N_6317);
nand U6428 (N_6428,N_6252,N_6275);
and U6429 (N_6429,N_6330,N_6376);
nor U6430 (N_6430,N_6328,N_6259);
or U6431 (N_6431,N_6331,N_6385);
xnor U6432 (N_6432,N_6315,N_6278);
or U6433 (N_6433,N_6251,N_6362);
or U6434 (N_6434,N_6370,N_6332);
nand U6435 (N_6435,N_6367,N_6288);
or U6436 (N_6436,N_6311,N_6386);
and U6437 (N_6437,N_6366,N_6291);
nand U6438 (N_6438,N_6347,N_6273);
or U6439 (N_6439,N_6394,N_6388);
nand U6440 (N_6440,N_6256,N_6258);
and U6441 (N_6441,N_6266,N_6374);
nand U6442 (N_6442,N_6240,N_6267);
and U6443 (N_6443,N_6390,N_6314);
nor U6444 (N_6444,N_6353,N_6329);
and U6445 (N_6445,N_6279,N_6320);
xnor U6446 (N_6446,N_6379,N_6253);
and U6447 (N_6447,N_6383,N_6241);
nor U6448 (N_6448,N_6268,N_6310);
and U6449 (N_6449,N_6305,N_6365);
or U6450 (N_6450,N_6351,N_6260);
nor U6451 (N_6451,N_6361,N_6246);
xor U6452 (N_6452,N_6316,N_6355);
nor U6453 (N_6453,N_6243,N_6335);
nand U6454 (N_6454,N_6334,N_6307);
and U6455 (N_6455,N_6302,N_6375);
nand U6456 (N_6456,N_6276,N_6271);
nor U6457 (N_6457,N_6282,N_6242);
or U6458 (N_6458,N_6261,N_6341);
nor U6459 (N_6459,N_6319,N_6338);
nor U6460 (N_6460,N_6336,N_6297);
and U6461 (N_6461,N_6368,N_6337);
xor U6462 (N_6462,N_6322,N_6295);
nor U6463 (N_6463,N_6306,N_6303);
nor U6464 (N_6464,N_6325,N_6333);
nor U6465 (N_6465,N_6343,N_6380);
or U6466 (N_6466,N_6393,N_6281);
and U6467 (N_6467,N_6290,N_6373);
nor U6468 (N_6468,N_6395,N_6293);
xnor U6469 (N_6469,N_6247,N_6399);
nand U6470 (N_6470,N_6274,N_6360);
xnor U6471 (N_6471,N_6264,N_6346);
and U6472 (N_6472,N_6371,N_6313);
nor U6473 (N_6473,N_6301,N_6392);
nor U6474 (N_6474,N_6326,N_6312);
nor U6475 (N_6475,N_6369,N_6381);
and U6476 (N_6476,N_6248,N_6254);
and U6477 (N_6477,N_6377,N_6323);
or U6478 (N_6478,N_6289,N_6354);
and U6479 (N_6479,N_6300,N_6372);
and U6480 (N_6480,N_6354,N_6392);
and U6481 (N_6481,N_6393,N_6389);
nand U6482 (N_6482,N_6308,N_6350);
nor U6483 (N_6483,N_6273,N_6267);
xor U6484 (N_6484,N_6389,N_6255);
xnor U6485 (N_6485,N_6383,N_6373);
and U6486 (N_6486,N_6287,N_6278);
and U6487 (N_6487,N_6324,N_6340);
nand U6488 (N_6488,N_6321,N_6270);
nand U6489 (N_6489,N_6382,N_6316);
or U6490 (N_6490,N_6384,N_6244);
or U6491 (N_6491,N_6393,N_6363);
or U6492 (N_6492,N_6343,N_6396);
and U6493 (N_6493,N_6266,N_6267);
or U6494 (N_6494,N_6385,N_6287);
and U6495 (N_6495,N_6330,N_6264);
nor U6496 (N_6496,N_6252,N_6314);
or U6497 (N_6497,N_6362,N_6329);
xor U6498 (N_6498,N_6319,N_6389);
or U6499 (N_6499,N_6329,N_6358);
and U6500 (N_6500,N_6246,N_6357);
or U6501 (N_6501,N_6307,N_6349);
or U6502 (N_6502,N_6269,N_6300);
or U6503 (N_6503,N_6376,N_6283);
nor U6504 (N_6504,N_6394,N_6361);
nand U6505 (N_6505,N_6373,N_6342);
nor U6506 (N_6506,N_6322,N_6336);
or U6507 (N_6507,N_6388,N_6372);
and U6508 (N_6508,N_6263,N_6393);
nor U6509 (N_6509,N_6359,N_6378);
or U6510 (N_6510,N_6320,N_6307);
nand U6511 (N_6511,N_6306,N_6247);
or U6512 (N_6512,N_6312,N_6395);
and U6513 (N_6513,N_6376,N_6265);
nand U6514 (N_6514,N_6345,N_6284);
nand U6515 (N_6515,N_6297,N_6344);
nor U6516 (N_6516,N_6256,N_6270);
nor U6517 (N_6517,N_6362,N_6289);
nor U6518 (N_6518,N_6258,N_6272);
and U6519 (N_6519,N_6359,N_6241);
nand U6520 (N_6520,N_6328,N_6387);
or U6521 (N_6521,N_6251,N_6286);
and U6522 (N_6522,N_6269,N_6343);
or U6523 (N_6523,N_6368,N_6256);
or U6524 (N_6524,N_6270,N_6349);
and U6525 (N_6525,N_6276,N_6382);
nand U6526 (N_6526,N_6387,N_6364);
nor U6527 (N_6527,N_6271,N_6368);
nor U6528 (N_6528,N_6335,N_6299);
nor U6529 (N_6529,N_6270,N_6288);
or U6530 (N_6530,N_6364,N_6287);
or U6531 (N_6531,N_6355,N_6349);
and U6532 (N_6532,N_6316,N_6265);
or U6533 (N_6533,N_6370,N_6286);
or U6534 (N_6534,N_6314,N_6330);
or U6535 (N_6535,N_6374,N_6397);
or U6536 (N_6536,N_6278,N_6336);
or U6537 (N_6537,N_6352,N_6324);
and U6538 (N_6538,N_6258,N_6248);
nor U6539 (N_6539,N_6349,N_6330);
nor U6540 (N_6540,N_6391,N_6342);
xnor U6541 (N_6541,N_6358,N_6312);
xor U6542 (N_6542,N_6283,N_6263);
and U6543 (N_6543,N_6351,N_6251);
or U6544 (N_6544,N_6394,N_6317);
and U6545 (N_6545,N_6325,N_6274);
or U6546 (N_6546,N_6330,N_6252);
nor U6547 (N_6547,N_6337,N_6303);
xnor U6548 (N_6548,N_6318,N_6363);
nand U6549 (N_6549,N_6356,N_6333);
nor U6550 (N_6550,N_6240,N_6330);
and U6551 (N_6551,N_6303,N_6396);
and U6552 (N_6552,N_6287,N_6244);
nand U6553 (N_6553,N_6304,N_6368);
nor U6554 (N_6554,N_6308,N_6369);
nor U6555 (N_6555,N_6343,N_6357);
nand U6556 (N_6556,N_6301,N_6370);
or U6557 (N_6557,N_6280,N_6305);
and U6558 (N_6558,N_6365,N_6261);
and U6559 (N_6559,N_6268,N_6284);
nor U6560 (N_6560,N_6434,N_6510);
xor U6561 (N_6561,N_6406,N_6403);
nor U6562 (N_6562,N_6550,N_6474);
nand U6563 (N_6563,N_6422,N_6426);
and U6564 (N_6564,N_6454,N_6452);
nand U6565 (N_6565,N_6525,N_6424);
xor U6566 (N_6566,N_6519,N_6472);
nand U6567 (N_6567,N_6529,N_6493);
nor U6568 (N_6568,N_6549,N_6523);
xor U6569 (N_6569,N_6536,N_6538);
nor U6570 (N_6570,N_6459,N_6524);
xor U6571 (N_6571,N_6543,N_6516);
and U6572 (N_6572,N_6436,N_6522);
or U6573 (N_6573,N_6464,N_6462);
nor U6574 (N_6574,N_6521,N_6421);
or U6575 (N_6575,N_6555,N_6554);
nor U6576 (N_6576,N_6502,N_6408);
nand U6577 (N_6577,N_6556,N_6495);
xor U6578 (N_6578,N_6540,N_6487);
xnor U6579 (N_6579,N_6476,N_6451);
nor U6580 (N_6580,N_6404,N_6435);
and U6581 (N_6581,N_6470,N_6409);
and U6582 (N_6582,N_6431,N_6558);
and U6583 (N_6583,N_6496,N_6445);
nor U6584 (N_6584,N_6506,N_6559);
or U6585 (N_6585,N_6507,N_6461);
nand U6586 (N_6586,N_6509,N_6534);
or U6587 (N_6587,N_6511,N_6450);
nand U6588 (N_6588,N_6444,N_6433);
nor U6589 (N_6589,N_6512,N_6475);
nor U6590 (N_6590,N_6465,N_6468);
nor U6591 (N_6591,N_6473,N_6477);
nor U6592 (N_6592,N_6427,N_6455);
and U6593 (N_6593,N_6539,N_6467);
nor U6594 (N_6594,N_6557,N_6417);
or U6595 (N_6595,N_6482,N_6407);
or U6596 (N_6596,N_6520,N_6537);
or U6597 (N_6597,N_6449,N_6479);
and U6598 (N_6598,N_6551,N_6527);
nand U6599 (N_6599,N_6514,N_6544);
and U6600 (N_6600,N_6548,N_6517);
or U6601 (N_6601,N_6504,N_6485);
nor U6602 (N_6602,N_6400,N_6508);
and U6603 (N_6603,N_6545,N_6518);
nand U6604 (N_6604,N_6469,N_6439);
nand U6605 (N_6605,N_6489,N_6552);
xor U6606 (N_6606,N_6492,N_6483);
nand U6607 (N_6607,N_6412,N_6505);
nand U6608 (N_6608,N_6478,N_6432);
nor U6609 (N_6609,N_6458,N_6447);
or U6610 (N_6610,N_6428,N_6443);
nor U6611 (N_6611,N_6532,N_6453);
nand U6612 (N_6612,N_6446,N_6430);
nand U6613 (N_6613,N_6415,N_6413);
and U6614 (N_6614,N_6530,N_6541);
nand U6615 (N_6615,N_6503,N_6440);
and U6616 (N_6616,N_6494,N_6429);
or U6617 (N_6617,N_6498,N_6526);
nor U6618 (N_6618,N_6515,N_6460);
or U6619 (N_6619,N_6471,N_6546);
and U6620 (N_6620,N_6491,N_6419);
xor U6621 (N_6621,N_6553,N_6410);
and U6622 (N_6622,N_6499,N_6463);
nand U6623 (N_6623,N_6488,N_6497);
nor U6624 (N_6624,N_6457,N_6438);
or U6625 (N_6625,N_6513,N_6425);
and U6626 (N_6626,N_6414,N_6420);
nand U6627 (N_6627,N_6528,N_6423);
and U6628 (N_6628,N_6535,N_6481);
or U6629 (N_6629,N_6411,N_6448);
or U6630 (N_6630,N_6547,N_6531);
nor U6631 (N_6631,N_6456,N_6486);
nand U6632 (N_6632,N_6441,N_6542);
or U6633 (N_6633,N_6437,N_6402);
nor U6634 (N_6634,N_6484,N_6501);
nor U6635 (N_6635,N_6500,N_6405);
nand U6636 (N_6636,N_6442,N_6466);
nor U6637 (N_6637,N_6480,N_6490);
or U6638 (N_6638,N_6416,N_6533);
nor U6639 (N_6639,N_6401,N_6418);
nand U6640 (N_6640,N_6462,N_6404);
nor U6641 (N_6641,N_6478,N_6410);
nand U6642 (N_6642,N_6530,N_6486);
nand U6643 (N_6643,N_6500,N_6496);
and U6644 (N_6644,N_6443,N_6476);
nand U6645 (N_6645,N_6535,N_6548);
or U6646 (N_6646,N_6460,N_6527);
and U6647 (N_6647,N_6540,N_6448);
nor U6648 (N_6648,N_6412,N_6495);
and U6649 (N_6649,N_6558,N_6457);
nand U6650 (N_6650,N_6511,N_6456);
or U6651 (N_6651,N_6540,N_6453);
or U6652 (N_6652,N_6465,N_6553);
nand U6653 (N_6653,N_6423,N_6483);
and U6654 (N_6654,N_6434,N_6465);
and U6655 (N_6655,N_6402,N_6457);
and U6656 (N_6656,N_6534,N_6443);
nor U6657 (N_6657,N_6518,N_6464);
nand U6658 (N_6658,N_6494,N_6473);
nand U6659 (N_6659,N_6412,N_6491);
or U6660 (N_6660,N_6457,N_6499);
nor U6661 (N_6661,N_6499,N_6525);
xnor U6662 (N_6662,N_6439,N_6473);
nand U6663 (N_6663,N_6547,N_6543);
and U6664 (N_6664,N_6553,N_6541);
nand U6665 (N_6665,N_6456,N_6514);
xor U6666 (N_6666,N_6538,N_6535);
nand U6667 (N_6667,N_6400,N_6493);
nand U6668 (N_6668,N_6525,N_6507);
and U6669 (N_6669,N_6498,N_6444);
or U6670 (N_6670,N_6497,N_6466);
or U6671 (N_6671,N_6529,N_6543);
or U6672 (N_6672,N_6527,N_6508);
nand U6673 (N_6673,N_6452,N_6520);
nand U6674 (N_6674,N_6449,N_6434);
nor U6675 (N_6675,N_6431,N_6531);
or U6676 (N_6676,N_6533,N_6448);
nand U6677 (N_6677,N_6496,N_6506);
or U6678 (N_6678,N_6521,N_6534);
nor U6679 (N_6679,N_6427,N_6471);
and U6680 (N_6680,N_6477,N_6459);
nand U6681 (N_6681,N_6457,N_6467);
xnor U6682 (N_6682,N_6530,N_6519);
and U6683 (N_6683,N_6464,N_6505);
nor U6684 (N_6684,N_6434,N_6496);
nor U6685 (N_6685,N_6424,N_6480);
and U6686 (N_6686,N_6421,N_6420);
or U6687 (N_6687,N_6514,N_6459);
or U6688 (N_6688,N_6407,N_6432);
xor U6689 (N_6689,N_6480,N_6446);
or U6690 (N_6690,N_6502,N_6418);
nand U6691 (N_6691,N_6503,N_6516);
nor U6692 (N_6692,N_6513,N_6472);
and U6693 (N_6693,N_6513,N_6532);
nand U6694 (N_6694,N_6431,N_6520);
nor U6695 (N_6695,N_6516,N_6525);
or U6696 (N_6696,N_6491,N_6473);
or U6697 (N_6697,N_6427,N_6529);
and U6698 (N_6698,N_6520,N_6501);
and U6699 (N_6699,N_6428,N_6411);
and U6700 (N_6700,N_6442,N_6418);
and U6701 (N_6701,N_6550,N_6515);
nor U6702 (N_6702,N_6559,N_6555);
or U6703 (N_6703,N_6549,N_6466);
or U6704 (N_6704,N_6440,N_6420);
nand U6705 (N_6705,N_6536,N_6559);
or U6706 (N_6706,N_6550,N_6452);
and U6707 (N_6707,N_6438,N_6500);
and U6708 (N_6708,N_6483,N_6464);
nor U6709 (N_6709,N_6493,N_6410);
nor U6710 (N_6710,N_6429,N_6412);
nor U6711 (N_6711,N_6470,N_6458);
and U6712 (N_6712,N_6424,N_6413);
and U6713 (N_6713,N_6490,N_6511);
or U6714 (N_6714,N_6554,N_6450);
and U6715 (N_6715,N_6500,N_6521);
and U6716 (N_6716,N_6511,N_6435);
and U6717 (N_6717,N_6556,N_6438);
and U6718 (N_6718,N_6444,N_6471);
and U6719 (N_6719,N_6505,N_6463);
and U6720 (N_6720,N_6711,N_6604);
or U6721 (N_6721,N_6713,N_6685);
nor U6722 (N_6722,N_6669,N_6617);
or U6723 (N_6723,N_6597,N_6632);
and U6724 (N_6724,N_6628,N_6702);
and U6725 (N_6725,N_6626,N_6661);
and U6726 (N_6726,N_6605,N_6687);
or U6727 (N_6727,N_6615,N_6660);
nor U6728 (N_6728,N_6718,N_6595);
and U6729 (N_6729,N_6643,N_6601);
nand U6730 (N_6730,N_6571,N_6693);
or U6731 (N_6731,N_6634,N_6649);
and U6732 (N_6732,N_6629,N_6588);
and U6733 (N_6733,N_6562,N_6635);
nor U6734 (N_6734,N_6619,N_6671);
nand U6735 (N_6735,N_6682,N_6621);
and U6736 (N_6736,N_6599,N_6662);
nand U6737 (N_6737,N_6624,N_6581);
or U6738 (N_6738,N_6659,N_6633);
or U6739 (N_6739,N_6677,N_6654);
xnor U6740 (N_6740,N_6701,N_6698);
or U6741 (N_6741,N_6564,N_6670);
nor U6742 (N_6742,N_6591,N_6692);
nor U6743 (N_6743,N_6576,N_6579);
nand U6744 (N_6744,N_6583,N_6610);
nor U6745 (N_6745,N_6612,N_6593);
and U6746 (N_6746,N_6714,N_6590);
nor U6747 (N_6747,N_6690,N_6676);
and U6748 (N_6748,N_6668,N_6574);
nand U6749 (N_6749,N_6691,N_6707);
nor U6750 (N_6750,N_6703,N_6607);
nand U6751 (N_6751,N_6697,N_6573);
and U6752 (N_6752,N_6704,N_6640);
or U6753 (N_6753,N_6715,N_6614);
and U6754 (N_6754,N_6567,N_6603);
and U6755 (N_6755,N_6561,N_6674);
xor U6756 (N_6756,N_6688,N_6686);
and U6757 (N_6757,N_6620,N_6608);
nor U6758 (N_6758,N_6577,N_6586);
or U6759 (N_6759,N_6710,N_6655);
nand U6760 (N_6760,N_6684,N_6596);
nor U6761 (N_6761,N_6664,N_6616);
nor U6762 (N_6762,N_6600,N_6652);
nor U6763 (N_6763,N_6566,N_6646);
nand U6764 (N_6764,N_6638,N_6694);
xnor U6765 (N_6765,N_6657,N_6584);
or U6766 (N_6766,N_6592,N_6630);
and U6767 (N_6767,N_6623,N_6611);
or U6768 (N_6768,N_6689,N_6631);
or U6769 (N_6769,N_6650,N_6705);
nand U6770 (N_6770,N_6667,N_6708);
and U6771 (N_6771,N_6666,N_6700);
nand U6772 (N_6772,N_6709,N_6602);
nand U6773 (N_6773,N_6589,N_6678);
or U6774 (N_6774,N_6706,N_6568);
or U6775 (N_6775,N_6647,N_6570);
nand U6776 (N_6776,N_6644,N_6642);
and U6777 (N_6777,N_6656,N_6675);
and U6778 (N_6778,N_6716,N_6613);
xnor U6779 (N_6779,N_6719,N_6578);
and U6780 (N_6780,N_6575,N_6637);
nand U6781 (N_6781,N_6622,N_6658);
or U6782 (N_6782,N_6585,N_6580);
and U6783 (N_6783,N_6653,N_6712);
nor U6784 (N_6784,N_6683,N_6618);
nor U6785 (N_6785,N_6673,N_6645);
nand U6786 (N_6786,N_6565,N_6641);
or U6787 (N_6787,N_6648,N_6681);
or U6788 (N_6788,N_6625,N_6587);
and U6789 (N_6789,N_6672,N_6665);
and U6790 (N_6790,N_6696,N_6598);
and U6791 (N_6791,N_6636,N_6651);
xor U6792 (N_6792,N_6569,N_6680);
and U6793 (N_6793,N_6606,N_6609);
nor U6794 (N_6794,N_6695,N_6572);
nand U6795 (N_6795,N_6582,N_6594);
nand U6796 (N_6796,N_6679,N_6639);
and U6797 (N_6797,N_6717,N_6563);
or U6798 (N_6798,N_6663,N_6627);
or U6799 (N_6799,N_6699,N_6560);
and U6800 (N_6800,N_6666,N_6685);
nor U6801 (N_6801,N_6626,N_6707);
and U6802 (N_6802,N_6707,N_6564);
and U6803 (N_6803,N_6689,N_6624);
nand U6804 (N_6804,N_6688,N_6588);
or U6805 (N_6805,N_6651,N_6673);
or U6806 (N_6806,N_6687,N_6571);
or U6807 (N_6807,N_6659,N_6578);
nor U6808 (N_6808,N_6635,N_6561);
or U6809 (N_6809,N_6711,N_6633);
nor U6810 (N_6810,N_6603,N_6661);
nand U6811 (N_6811,N_6656,N_6641);
nand U6812 (N_6812,N_6661,N_6657);
or U6813 (N_6813,N_6567,N_6657);
or U6814 (N_6814,N_6693,N_6573);
nor U6815 (N_6815,N_6560,N_6685);
or U6816 (N_6816,N_6573,N_6602);
nor U6817 (N_6817,N_6696,N_6564);
and U6818 (N_6818,N_6643,N_6662);
and U6819 (N_6819,N_6592,N_6571);
xor U6820 (N_6820,N_6564,N_6621);
or U6821 (N_6821,N_6600,N_6687);
or U6822 (N_6822,N_6718,N_6620);
nor U6823 (N_6823,N_6694,N_6601);
and U6824 (N_6824,N_6605,N_6626);
and U6825 (N_6825,N_6642,N_6670);
or U6826 (N_6826,N_6676,N_6651);
or U6827 (N_6827,N_6698,N_6622);
and U6828 (N_6828,N_6717,N_6632);
nor U6829 (N_6829,N_6705,N_6673);
and U6830 (N_6830,N_6565,N_6694);
and U6831 (N_6831,N_6698,N_6694);
or U6832 (N_6832,N_6621,N_6671);
or U6833 (N_6833,N_6673,N_6680);
nand U6834 (N_6834,N_6652,N_6689);
nand U6835 (N_6835,N_6590,N_6581);
nor U6836 (N_6836,N_6665,N_6651);
xor U6837 (N_6837,N_6669,N_6597);
and U6838 (N_6838,N_6586,N_6609);
nor U6839 (N_6839,N_6635,N_6717);
or U6840 (N_6840,N_6639,N_6702);
nand U6841 (N_6841,N_6694,N_6633);
nor U6842 (N_6842,N_6560,N_6713);
and U6843 (N_6843,N_6637,N_6652);
and U6844 (N_6844,N_6693,N_6668);
or U6845 (N_6845,N_6718,N_6664);
or U6846 (N_6846,N_6632,N_6571);
nand U6847 (N_6847,N_6561,N_6671);
xor U6848 (N_6848,N_6648,N_6673);
and U6849 (N_6849,N_6599,N_6694);
or U6850 (N_6850,N_6696,N_6615);
or U6851 (N_6851,N_6625,N_6693);
nand U6852 (N_6852,N_6661,N_6595);
and U6853 (N_6853,N_6595,N_6607);
nand U6854 (N_6854,N_6584,N_6586);
nor U6855 (N_6855,N_6581,N_6608);
nor U6856 (N_6856,N_6636,N_6632);
or U6857 (N_6857,N_6677,N_6697);
or U6858 (N_6858,N_6605,N_6563);
xor U6859 (N_6859,N_6704,N_6688);
or U6860 (N_6860,N_6653,N_6569);
nor U6861 (N_6861,N_6697,N_6648);
nand U6862 (N_6862,N_6673,N_6632);
nor U6863 (N_6863,N_6620,N_6715);
nand U6864 (N_6864,N_6658,N_6582);
nand U6865 (N_6865,N_6603,N_6578);
and U6866 (N_6866,N_6685,N_6706);
nor U6867 (N_6867,N_6573,N_6645);
nor U6868 (N_6868,N_6640,N_6586);
and U6869 (N_6869,N_6567,N_6707);
and U6870 (N_6870,N_6667,N_6586);
or U6871 (N_6871,N_6666,N_6578);
nor U6872 (N_6872,N_6616,N_6583);
nand U6873 (N_6873,N_6690,N_6637);
and U6874 (N_6874,N_6573,N_6596);
or U6875 (N_6875,N_6602,N_6584);
nand U6876 (N_6876,N_6576,N_6598);
and U6877 (N_6877,N_6621,N_6588);
nor U6878 (N_6878,N_6568,N_6667);
xnor U6879 (N_6879,N_6713,N_6698);
nand U6880 (N_6880,N_6803,N_6842);
xnor U6881 (N_6881,N_6869,N_6793);
nand U6882 (N_6882,N_6834,N_6815);
nand U6883 (N_6883,N_6742,N_6789);
or U6884 (N_6884,N_6765,N_6817);
xnor U6885 (N_6885,N_6788,N_6843);
or U6886 (N_6886,N_6854,N_6735);
nand U6887 (N_6887,N_6758,N_6727);
or U6888 (N_6888,N_6810,N_6874);
nand U6889 (N_6889,N_6802,N_6811);
or U6890 (N_6890,N_6736,N_6844);
nor U6891 (N_6891,N_6778,N_6739);
or U6892 (N_6892,N_6779,N_6744);
or U6893 (N_6893,N_6822,N_6777);
or U6894 (N_6894,N_6800,N_6865);
and U6895 (N_6895,N_6832,N_6805);
nor U6896 (N_6896,N_6850,N_6878);
and U6897 (N_6897,N_6857,N_6849);
and U6898 (N_6898,N_6785,N_6756);
or U6899 (N_6899,N_6771,N_6841);
nand U6900 (N_6900,N_6781,N_6753);
and U6901 (N_6901,N_6808,N_6858);
nor U6902 (N_6902,N_6792,N_6809);
xnor U6903 (N_6903,N_6795,N_6845);
and U6904 (N_6904,N_6864,N_6740);
nand U6905 (N_6905,N_6766,N_6859);
nor U6906 (N_6906,N_6784,N_6782);
nand U6907 (N_6907,N_6767,N_6720);
or U6908 (N_6908,N_6806,N_6732);
nand U6909 (N_6909,N_6791,N_6826);
or U6910 (N_6910,N_6745,N_6754);
or U6911 (N_6911,N_6746,N_6733);
or U6912 (N_6912,N_6728,N_6821);
and U6913 (N_6913,N_6751,N_6823);
and U6914 (N_6914,N_6867,N_6877);
and U6915 (N_6915,N_6731,N_6755);
or U6916 (N_6916,N_6723,N_6776);
and U6917 (N_6917,N_6737,N_6743);
nand U6918 (N_6918,N_6840,N_6798);
or U6919 (N_6919,N_6763,N_6856);
or U6920 (N_6920,N_6820,N_6761);
and U6921 (N_6921,N_6872,N_6773);
or U6922 (N_6922,N_6835,N_6870);
nand U6923 (N_6923,N_6830,N_6838);
nand U6924 (N_6924,N_6721,N_6871);
xnor U6925 (N_6925,N_6724,N_6768);
nor U6926 (N_6926,N_6819,N_6863);
nor U6927 (N_6927,N_6747,N_6879);
and U6928 (N_6928,N_6786,N_6734);
xor U6929 (N_6929,N_6799,N_6824);
nor U6930 (N_6930,N_6861,N_6770);
and U6931 (N_6931,N_6818,N_6796);
and U6932 (N_6932,N_6833,N_6760);
xor U6933 (N_6933,N_6836,N_6866);
and U6934 (N_6934,N_6847,N_6725);
or U6935 (N_6935,N_6730,N_6748);
or U6936 (N_6936,N_6868,N_6722);
nand U6937 (N_6937,N_6837,N_6813);
xor U6938 (N_6938,N_6875,N_6801);
nor U6939 (N_6939,N_6860,N_6853);
xnor U6940 (N_6940,N_6829,N_6816);
nand U6941 (N_6941,N_6828,N_6769);
nand U6942 (N_6942,N_6759,N_6873);
or U6943 (N_6943,N_6780,N_6839);
and U6944 (N_6944,N_6764,N_6750);
xor U6945 (N_6945,N_6807,N_6831);
and U6946 (N_6946,N_6797,N_6862);
nand U6947 (N_6947,N_6812,N_6804);
and U6948 (N_6948,N_6848,N_6852);
xnor U6949 (N_6949,N_6738,N_6774);
xor U6950 (N_6950,N_6855,N_6876);
nor U6951 (N_6951,N_6752,N_6794);
nor U6952 (N_6952,N_6729,N_6787);
xor U6953 (N_6953,N_6757,N_6772);
nor U6954 (N_6954,N_6851,N_6827);
nand U6955 (N_6955,N_6749,N_6726);
or U6956 (N_6956,N_6775,N_6762);
and U6957 (N_6957,N_6741,N_6846);
nand U6958 (N_6958,N_6783,N_6825);
or U6959 (N_6959,N_6790,N_6814);
and U6960 (N_6960,N_6733,N_6839);
and U6961 (N_6961,N_6847,N_6824);
nand U6962 (N_6962,N_6734,N_6796);
nand U6963 (N_6963,N_6873,N_6806);
nand U6964 (N_6964,N_6848,N_6850);
xnor U6965 (N_6965,N_6735,N_6816);
nor U6966 (N_6966,N_6801,N_6823);
and U6967 (N_6967,N_6801,N_6748);
nand U6968 (N_6968,N_6807,N_6797);
nand U6969 (N_6969,N_6825,N_6788);
nand U6970 (N_6970,N_6780,N_6740);
and U6971 (N_6971,N_6758,N_6830);
nand U6972 (N_6972,N_6771,N_6849);
xor U6973 (N_6973,N_6825,N_6733);
nor U6974 (N_6974,N_6874,N_6749);
or U6975 (N_6975,N_6766,N_6851);
nor U6976 (N_6976,N_6879,N_6805);
nand U6977 (N_6977,N_6785,N_6768);
or U6978 (N_6978,N_6829,N_6754);
nand U6979 (N_6979,N_6764,N_6844);
or U6980 (N_6980,N_6771,N_6791);
nand U6981 (N_6981,N_6840,N_6795);
nand U6982 (N_6982,N_6783,N_6810);
xor U6983 (N_6983,N_6829,N_6794);
nand U6984 (N_6984,N_6840,N_6742);
nor U6985 (N_6985,N_6874,N_6765);
nor U6986 (N_6986,N_6720,N_6799);
and U6987 (N_6987,N_6871,N_6874);
and U6988 (N_6988,N_6752,N_6807);
nor U6989 (N_6989,N_6833,N_6872);
xnor U6990 (N_6990,N_6878,N_6740);
nand U6991 (N_6991,N_6820,N_6818);
nand U6992 (N_6992,N_6827,N_6762);
nand U6993 (N_6993,N_6816,N_6828);
nor U6994 (N_6994,N_6807,N_6804);
or U6995 (N_6995,N_6765,N_6804);
nand U6996 (N_6996,N_6842,N_6743);
xor U6997 (N_6997,N_6811,N_6825);
nor U6998 (N_6998,N_6761,N_6876);
and U6999 (N_6999,N_6857,N_6742);
or U7000 (N_7000,N_6863,N_6833);
and U7001 (N_7001,N_6791,N_6738);
nor U7002 (N_7002,N_6751,N_6798);
nor U7003 (N_7003,N_6770,N_6846);
xnor U7004 (N_7004,N_6746,N_6857);
nand U7005 (N_7005,N_6729,N_6879);
or U7006 (N_7006,N_6814,N_6775);
or U7007 (N_7007,N_6732,N_6753);
nand U7008 (N_7008,N_6762,N_6745);
or U7009 (N_7009,N_6777,N_6814);
or U7010 (N_7010,N_6862,N_6867);
and U7011 (N_7011,N_6788,N_6727);
or U7012 (N_7012,N_6807,N_6811);
nor U7013 (N_7013,N_6830,N_6750);
nand U7014 (N_7014,N_6853,N_6722);
xor U7015 (N_7015,N_6745,N_6839);
and U7016 (N_7016,N_6725,N_6731);
and U7017 (N_7017,N_6847,N_6764);
nand U7018 (N_7018,N_6742,N_6725);
nor U7019 (N_7019,N_6745,N_6742);
or U7020 (N_7020,N_6813,N_6817);
xnor U7021 (N_7021,N_6802,N_6870);
or U7022 (N_7022,N_6796,N_6819);
and U7023 (N_7023,N_6808,N_6837);
xor U7024 (N_7024,N_6745,N_6856);
or U7025 (N_7025,N_6772,N_6730);
or U7026 (N_7026,N_6839,N_6746);
and U7027 (N_7027,N_6879,N_6808);
nor U7028 (N_7028,N_6873,N_6817);
or U7029 (N_7029,N_6813,N_6853);
nand U7030 (N_7030,N_6740,N_6851);
nand U7031 (N_7031,N_6872,N_6754);
and U7032 (N_7032,N_6752,N_6729);
nor U7033 (N_7033,N_6733,N_6801);
nand U7034 (N_7034,N_6804,N_6773);
nand U7035 (N_7035,N_6827,N_6786);
or U7036 (N_7036,N_6780,N_6747);
nor U7037 (N_7037,N_6740,N_6806);
nor U7038 (N_7038,N_6731,N_6749);
nand U7039 (N_7039,N_6856,N_6766);
and U7040 (N_7040,N_7010,N_7023);
or U7041 (N_7041,N_6990,N_7024);
or U7042 (N_7042,N_7012,N_6886);
nor U7043 (N_7043,N_6898,N_6890);
or U7044 (N_7044,N_6974,N_6925);
xnor U7045 (N_7045,N_7013,N_7032);
nand U7046 (N_7046,N_6911,N_6955);
nor U7047 (N_7047,N_6924,N_6888);
or U7048 (N_7048,N_6885,N_6940);
or U7049 (N_7049,N_6961,N_6973);
nand U7050 (N_7050,N_6893,N_6998);
nand U7051 (N_7051,N_6923,N_6906);
nor U7052 (N_7052,N_6986,N_6883);
or U7053 (N_7053,N_6944,N_6989);
or U7054 (N_7054,N_6930,N_6904);
nor U7055 (N_7055,N_6908,N_7033);
nand U7056 (N_7056,N_6945,N_7017);
and U7057 (N_7057,N_6987,N_6920);
or U7058 (N_7058,N_6912,N_6929);
and U7059 (N_7059,N_7036,N_7016);
nor U7060 (N_7060,N_6972,N_6982);
and U7061 (N_7061,N_7014,N_7038);
nor U7062 (N_7062,N_6960,N_7005);
nand U7063 (N_7063,N_7019,N_6969);
xor U7064 (N_7064,N_7003,N_6943);
nor U7065 (N_7065,N_7030,N_6900);
nand U7066 (N_7066,N_6976,N_6980);
or U7067 (N_7067,N_6951,N_7004);
nor U7068 (N_7068,N_7008,N_6915);
xor U7069 (N_7069,N_6958,N_6913);
or U7070 (N_7070,N_6947,N_7027);
nand U7071 (N_7071,N_6896,N_6884);
or U7072 (N_7072,N_6907,N_6899);
and U7073 (N_7073,N_6996,N_6950);
or U7074 (N_7074,N_7025,N_6952);
nand U7075 (N_7075,N_6891,N_6901);
xor U7076 (N_7076,N_6921,N_6934);
nor U7077 (N_7077,N_7000,N_6919);
or U7078 (N_7078,N_6916,N_7035);
nand U7079 (N_7079,N_6881,N_6948);
nand U7080 (N_7080,N_6882,N_7002);
or U7081 (N_7081,N_6931,N_6941);
and U7082 (N_7082,N_6939,N_6978);
nor U7083 (N_7083,N_6897,N_6932);
and U7084 (N_7084,N_6995,N_6964);
and U7085 (N_7085,N_6999,N_7031);
and U7086 (N_7086,N_6959,N_6968);
xnor U7087 (N_7087,N_6988,N_6917);
xnor U7088 (N_7088,N_6922,N_6966);
nor U7089 (N_7089,N_6981,N_7034);
xnor U7090 (N_7090,N_7039,N_6946);
nor U7091 (N_7091,N_6975,N_6895);
or U7092 (N_7092,N_6935,N_6927);
nand U7093 (N_7093,N_6994,N_6903);
nor U7094 (N_7094,N_7015,N_6909);
nand U7095 (N_7095,N_7011,N_6918);
nor U7096 (N_7096,N_6984,N_6954);
nand U7097 (N_7097,N_7026,N_6993);
nor U7098 (N_7098,N_7007,N_6991);
and U7099 (N_7099,N_6962,N_6992);
xnor U7100 (N_7100,N_6967,N_7020);
nor U7101 (N_7101,N_6985,N_6892);
xor U7102 (N_7102,N_6957,N_7001);
and U7103 (N_7103,N_6953,N_6938);
or U7104 (N_7104,N_6887,N_6889);
nand U7105 (N_7105,N_6933,N_6880);
or U7106 (N_7106,N_6905,N_6956);
xnor U7107 (N_7107,N_7029,N_6926);
nand U7108 (N_7108,N_6936,N_6937);
nand U7109 (N_7109,N_6910,N_6965);
nor U7110 (N_7110,N_7009,N_7028);
nand U7111 (N_7111,N_6970,N_7018);
and U7112 (N_7112,N_7006,N_6983);
nand U7113 (N_7113,N_7021,N_6914);
nand U7114 (N_7114,N_6997,N_7037);
nor U7115 (N_7115,N_6894,N_6963);
xor U7116 (N_7116,N_6902,N_6942);
and U7117 (N_7117,N_6971,N_6977);
nand U7118 (N_7118,N_6949,N_6979);
nor U7119 (N_7119,N_7022,N_6928);
nand U7120 (N_7120,N_6987,N_7036);
nand U7121 (N_7121,N_6961,N_6992);
or U7122 (N_7122,N_6963,N_7033);
and U7123 (N_7123,N_6978,N_6898);
or U7124 (N_7124,N_7034,N_6915);
nand U7125 (N_7125,N_6901,N_7028);
or U7126 (N_7126,N_7011,N_6931);
and U7127 (N_7127,N_7016,N_6910);
nand U7128 (N_7128,N_7027,N_6904);
nand U7129 (N_7129,N_6910,N_6983);
and U7130 (N_7130,N_6975,N_6922);
nand U7131 (N_7131,N_7031,N_6963);
and U7132 (N_7132,N_6995,N_6945);
nand U7133 (N_7133,N_6915,N_7019);
or U7134 (N_7134,N_6980,N_6946);
nor U7135 (N_7135,N_6969,N_6953);
nand U7136 (N_7136,N_6925,N_6984);
nand U7137 (N_7137,N_6920,N_6937);
nand U7138 (N_7138,N_6919,N_6936);
and U7139 (N_7139,N_7013,N_6899);
nor U7140 (N_7140,N_6956,N_6915);
nor U7141 (N_7141,N_6917,N_6921);
nor U7142 (N_7142,N_6897,N_7032);
nand U7143 (N_7143,N_6897,N_6902);
nand U7144 (N_7144,N_6890,N_6986);
or U7145 (N_7145,N_6926,N_7002);
nand U7146 (N_7146,N_6929,N_6996);
and U7147 (N_7147,N_6958,N_6939);
nand U7148 (N_7148,N_6954,N_6987);
nand U7149 (N_7149,N_6936,N_7014);
xnor U7150 (N_7150,N_7032,N_6880);
and U7151 (N_7151,N_6884,N_6996);
nand U7152 (N_7152,N_6906,N_6954);
or U7153 (N_7153,N_6907,N_7035);
and U7154 (N_7154,N_6970,N_6963);
xor U7155 (N_7155,N_6997,N_6931);
nand U7156 (N_7156,N_6888,N_6962);
nand U7157 (N_7157,N_6899,N_6971);
nor U7158 (N_7158,N_6967,N_6947);
nor U7159 (N_7159,N_6969,N_6991);
and U7160 (N_7160,N_7001,N_7034);
and U7161 (N_7161,N_7004,N_6892);
nand U7162 (N_7162,N_7001,N_7019);
or U7163 (N_7163,N_6899,N_6983);
nand U7164 (N_7164,N_6929,N_6880);
or U7165 (N_7165,N_6980,N_6943);
nor U7166 (N_7166,N_6993,N_6987);
or U7167 (N_7167,N_6958,N_7026);
nand U7168 (N_7168,N_6991,N_6952);
nor U7169 (N_7169,N_6982,N_7036);
nor U7170 (N_7170,N_6959,N_6912);
xnor U7171 (N_7171,N_6913,N_7033);
and U7172 (N_7172,N_7024,N_7010);
and U7173 (N_7173,N_7032,N_7031);
xor U7174 (N_7174,N_7031,N_7022);
nand U7175 (N_7175,N_6929,N_6909);
or U7176 (N_7176,N_6968,N_6945);
nand U7177 (N_7177,N_6947,N_7020);
or U7178 (N_7178,N_6934,N_7021);
and U7179 (N_7179,N_6887,N_6898);
xor U7180 (N_7180,N_7016,N_6959);
and U7181 (N_7181,N_6996,N_6958);
nand U7182 (N_7182,N_6946,N_6994);
nor U7183 (N_7183,N_6991,N_6880);
xor U7184 (N_7184,N_6944,N_6889);
and U7185 (N_7185,N_6908,N_6947);
xor U7186 (N_7186,N_6998,N_6914);
and U7187 (N_7187,N_6964,N_7029);
and U7188 (N_7188,N_6965,N_6998);
nand U7189 (N_7189,N_7023,N_7026);
nand U7190 (N_7190,N_6899,N_7023);
and U7191 (N_7191,N_6954,N_6971);
nand U7192 (N_7192,N_6979,N_6896);
and U7193 (N_7193,N_6885,N_7024);
xor U7194 (N_7194,N_6926,N_6991);
or U7195 (N_7195,N_7017,N_6907);
and U7196 (N_7196,N_7023,N_6881);
and U7197 (N_7197,N_6925,N_6976);
nand U7198 (N_7198,N_6899,N_6919);
or U7199 (N_7199,N_6950,N_7032);
xor U7200 (N_7200,N_7153,N_7048);
or U7201 (N_7201,N_7122,N_7086);
and U7202 (N_7202,N_7053,N_7192);
nand U7203 (N_7203,N_7098,N_7169);
or U7204 (N_7204,N_7066,N_7069);
nor U7205 (N_7205,N_7123,N_7171);
nor U7206 (N_7206,N_7149,N_7165);
and U7207 (N_7207,N_7185,N_7140);
nand U7208 (N_7208,N_7115,N_7116);
nor U7209 (N_7209,N_7143,N_7101);
and U7210 (N_7210,N_7159,N_7095);
and U7211 (N_7211,N_7162,N_7088);
and U7212 (N_7212,N_7135,N_7167);
or U7213 (N_7213,N_7194,N_7107);
nor U7214 (N_7214,N_7097,N_7172);
or U7215 (N_7215,N_7129,N_7184);
nor U7216 (N_7216,N_7133,N_7108);
nor U7217 (N_7217,N_7175,N_7073);
nor U7218 (N_7218,N_7064,N_7132);
or U7219 (N_7219,N_7154,N_7090);
xnor U7220 (N_7220,N_7081,N_7047);
nor U7221 (N_7221,N_7138,N_7104);
nor U7222 (N_7222,N_7144,N_7130);
nor U7223 (N_7223,N_7152,N_7114);
and U7224 (N_7224,N_7182,N_7043);
or U7225 (N_7225,N_7161,N_7062);
or U7226 (N_7226,N_7177,N_7075);
and U7227 (N_7227,N_7056,N_7134);
or U7228 (N_7228,N_7084,N_7045);
or U7229 (N_7229,N_7061,N_7102);
or U7230 (N_7230,N_7198,N_7199);
nor U7231 (N_7231,N_7174,N_7040);
or U7232 (N_7232,N_7176,N_7150);
and U7233 (N_7233,N_7189,N_7128);
and U7234 (N_7234,N_7119,N_7157);
or U7235 (N_7235,N_7118,N_7156);
nand U7236 (N_7236,N_7060,N_7050);
or U7237 (N_7237,N_7096,N_7059);
nor U7238 (N_7238,N_7186,N_7151);
or U7239 (N_7239,N_7079,N_7180);
nor U7240 (N_7240,N_7197,N_7137);
nand U7241 (N_7241,N_7058,N_7083);
and U7242 (N_7242,N_7044,N_7051);
or U7243 (N_7243,N_7136,N_7127);
nor U7244 (N_7244,N_7049,N_7042);
xor U7245 (N_7245,N_7109,N_7112);
or U7246 (N_7246,N_7077,N_7141);
nand U7247 (N_7247,N_7131,N_7093);
nor U7248 (N_7248,N_7147,N_7085);
nand U7249 (N_7249,N_7099,N_7160);
nor U7250 (N_7250,N_7052,N_7163);
and U7251 (N_7251,N_7046,N_7126);
or U7252 (N_7252,N_7074,N_7094);
nor U7253 (N_7253,N_7170,N_7193);
and U7254 (N_7254,N_7121,N_7195);
nor U7255 (N_7255,N_7181,N_7120);
and U7256 (N_7256,N_7071,N_7087);
nand U7257 (N_7257,N_7191,N_7117);
nor U7258 (N_7258,N_7113,N_7183);
nand U7259 (N_7259,N_7105,N_7124);
and U7260 (N_7260,N_7168,N_7110);
or U7261 (N_7261,N_7125,N_7196);
and U7262 (N_7262,N_7146,N_7103);
and U7263 (N_7263,N_7067,N_7055);
or U7264 (N_7264,N_7173,N_7080);
or U7265 (N_7265,N_7187,N_7188);
and U7266 (N_7266,N_7076,N_7068);
nor U7267 (N_7267,N_7091,N_7166);
or U7268 (N_7268,N_7082,N_7063);
nand U7269 (N_7269,N_7164,N_7089);
xor U7270 (N_7270,N_7078,N_7139);
and U7271 (N_7271,N_7106,N_7178);
and U7272 (N_7272,N_7065,N_7054);
nand U7273 (N_7273,N_7070,N_7100);
or U7274 (N_7274,N_7179,N_7190);
nor U7275 (N_7275,N_7041,N_7111);
or U7276 (N_7276,N_7145,N_7057);
or U7277 (N_7277,N_7142,N_7092);
nor U7278 (N_7278,N_7148,N_7072);
nand U7279 (N_7279,N_7158,N_7155);
xor U7280 (N_7280,N_7107,N_7095);
nor U7281 (N_7281,N_7123,N_7114);
nor U7282 (N_7282,N_7043,N_7175);
nand U7283 (N_7283,N_7173,N_7136);
and U7284 (N_7284,N_7187,N_7059);
nor U7285 (N_7285,N_7155,N_7100);
and U7286 (N_7286,N_7188,N_7054);
or U7287 (N_7287,N_7047,N_7052);
and U7288 (N_7288,N_7057,N_7168);
nor U7289 (N_7289,N_7188,N_7121);
nor U7290 (N_7290,N_7046,N_7153);
or U7291 (N_7291,N_7176,N_7093);
nor U7292 (N_7292,N_7079,N_7168);
and U7293 (N_7293,N_7066,N_7101);
and U7294 (N_7294,N_7085,N_7153);
nand U7295 (N_7295,N_7150,N_7058);
xor U7296 (N_7296,N_7090,N_7115);
or U7297 (N_7297,N_7146,N_7094);
or U7298 (N_7298,N_7071,N_7063);
and U7299 (N_7299,N_7164,N_7117);
or U7300 (N_7300,N_7089,N_7174);
or U7301 (N_7301,N_7144,N_7095);
nand U7302 (N_7302,N_7049,N_7061);
xnor U7303 (N_7303,N_7161,N_7054);
and U7304 (N_7304,N_7185,N_7156);
or U7305 (N_7305,N_7125,N_7169);
and U7306 (N_7306,N_7076,N_7118);
nand U7307 (N_7307,N_7040,N_7079);
nor U7308 (N_7308,N_7114,N_7185);
and U7309 (N_7309,N_7188,N_7194);
or U7310 (N_7310,N_7040,N_7047);
or U7311 (N_7311,N_7051,N_7088);
nand U7312 (N_7312,N_7101,N_7169);
nand U7313 (N_7313,N_7170,N_7197);
and U7314 (N_7314,N_7062,N_7118);
nand U7315 (N_7315,N_7195,N_7197);
nand U7316 (N_7316,N_7188,N_7110);
nand U7317 (N_7317,N_7158,N_7191);
nor U7318 (N_7318,N_7079,N_7132);
nor U7319 (N_7319,N_7120,N_7102);
and U7320 (N_7320,N_7048,N_7167);
and U7321 (N_7321,N_7163,N_7184);
nand U7322 (N_7322,N_7061,N_7056);
nor U7323 (N_7323,N_7198,N_7130);
or U7324 (N_7324,N_7199,N_7063);
nand U7325 (N_7325,N_7144,N_7153);
and U7326 (N_7326,N_7103,N_7101);
nor U7327 (N_7327,N_7189,N_7153);
or U7328 (N_7328,N_7052,N_7168);
and U7329 (N_7329,N_7170,N_7100);
or U7330 (N_7330,N_7169,N_7108);
and U7331 (N_7331,N_7119,N_7104);
xnor U7332 (N_7332,N_7073,N_7142);
or U7333 (N_7333,N_7150,N_7093);
or U7334 (N_7334,N_7080,N_7135);
nor U7335 (N_7335,N_7199,N_7187);
and U7336 (N_7336,N_7055,N_7096);
nand U7337 (N_7337,N_7113,N_7120);
xnor U7338 (N_7338,N_7125,N_7082);
nand U7339 (N_7339,N_7160,N_7196);
nor U7340 (N_7340,N_7184,N_7105);
nor U7341 (N_7341,N_7136,N_7177);
xor U7342 (N_7342,N_7189,N_7086);
nor U7343 (N_7343,N_7126,N_7156);
nor U7344 (N_7344,N_7061,N_7070);
and U7345 (N_7345,N_7102,N_7133);
nor U7346 (N_7346,N_7189,N_7120);
and U7347 (N_7347,N_7135,N_7095);
and U7348 (N_7348,N_7050,N_7092);
nand U7349 (N_7349,N_7199,N_7085);
and U7350 (N_7350,N_7137,N_7135);
nor U7351 (N_7351,N_7169,N_7184);
or U7352 (N_7352,N_7125,N_7100);
nor U7353 (N_7353,N_7106,N_7134);
nand U7354 (N_7354,N_7192,N_7075);
or U7355 (N_7355,N_7091,N_7110);
or U7356 (N_7356,N_7073,N_7113);
and U7357 (N_7357,N_7147,N_7060);
and U7358 (N_7358,N_7058,N_7194);
and U7359 (N_7359,N_7178,N_7058);
and U7360 (N_7360,N_7290,N_7275);
and U7361 (N_7361,N_7300,N_7356);
nand U7362 (N_7362,N_7246,N_7354);
nor U7363 (N_7363,N_7250,N_7210);
nor U7364 (N_7364,N_7332,N_7282);
or U7365 (N_7365,N_7264,N_7231);
nand U7366 (N_7366,N_7288,N_7317);
or U7367 (N_7367,N_7312,N_7348);
or U7368 (N_7368,N_7324,N_7223);
or U7369 (N_7369,N_7339,N_7285);
or U7370 (N_7370,N_7209,N_7306);
nand U7371 (N_7371,N_7315,N_7202);
nor U7372 (N_7372,N_7215,N_7353);
or U7373 (N_7373,N_7253,N_7232);
or U7374 (N_7374,N_7201,N_7345);
or U7375 (N_7375,N_7334,N_7293);
xor U7376 (N_7376,N_7239,N_7265);
nor U7377 (N_7377,N_7291,N_7270);
or U7378 (N_7378,N_7321,N_7298);
nand U7379 (N_7379,N_7355,N_7225);
xor U7380 (N_7380,N_7218,N_7257);
and U7381 (N_7381,N_7263,N_7295);
nand U7382 (N_7382,N_7279,N_7314);
nand U7383 (N_7383,N_7350,N_7220);
nor U7384 (N_7384,N_7203,N_7347);
and U7385 (N_7385,N_7338,N_7240);
nand U7386 (N_7386,N_7349,N_7242);
or U7387 (N_7387,N_7214,N_7292);
nor U7388 (N_7388,N_7262,N_7254);
nor U7389 (N_7389,N_7217,N_7258);
and U7390 (N_7390,N_7229,N_7247);
xnor U7391 (N_7391,N_7301,N_7322);
or U7392 (N_7392,N_7359,N_7278);
and U7393 (N_7393,N_7227,N_7319);
or U7394 (N_7394,N_7341,N_7261);
or U7395 (N_7395,N_7308,N_7234);
nand U7396 (N_7396,N_7336,N_7318);
nand U7397 (N_7397,N_7269,N_7200);
xnor U7398 (N_7398,N_7212,N_7329);
xnor U7399 (N_7399,N_7325,N_7309);
nand U7400 (N_7400,N_7273,N_7313);
nor U7401 (N_7401,N_7283,N_7274);
nor U7402 (N_7402,N_7284,N_7303);
or U7403 (N_7403,N_7287,N_7266);
or U7404 (N_7404,N_7304,N_7206);
and U7405 (N_7405,N_7259,N_7224);
or U7406 (N_7406,N_7245,N_7311);
or U7407 (N_7407,N_7249,N_7310);
nand U7408 (N_7408,N_7272,N_7236);
nor U7409 (N_7409,N_7277,N_7244);
or U7410 (N_7410,N_7328,N_7226);
nor U7411 (N_7411,N_7305,N_7228);
nor U7412 (N_7412,N_7219,N_7326);
nor U7413 (N_7413,N_7302,N_7343);
xor U7414 (N_7414,N_7280,N_7330);
nor U7415 (N_7415,N_7358,N_7297);
nor U7416 (N_7416,N_7316,N_7243);
and U7417 (N_7417,N_7237,N_7255);
nor U7418 (N_7418,N_7337,N_7331);
and U7419 (N_7419,N_7276,N_7251);
nand U7420 (N_7420,N_7267,N_7216);
nor U7421 (N_7421,N_7289,N_7213);
and U7422 (N_7422,N_7342,N_7238);
and U7423 (N_7423,N_7268,N_7204);
xnor U7424 (N_7424,N_7294,N_7222);
nand U7425 (N_7425,N_7296,N_7357);
nand U7426 (N_7426,N_7335,N_7351);
nand U7427 (N_7427,N_7281,N_7260);
nor U7428 (N_7428,N_7346,N_7299);
or U7429 (N_7429,N_7340,N_7333);
nand U7430 (N_7430,N_7271,N_7252);
or U7431 (N_7431,N_7256,N_7344);
or U7432 (N_7432,N_7286,N_7248);
or U7433 (N_7433,N_7207,N_7323);
and U7434 (N_7434,N_7241,N_7233);
xnor U7435 (N_7435,N_7221,N_7320);
and U7436 (N_7436,N_7352,N_7230);
nor U7437 (N_7437,N_7205,N_7327);
or U7438 (N_7438,N_7307,N_7235);
nand U7439 (N_7439,N_7211,N_7208);
xnor U7440 (N_7440,N_7201,N_7336);
xnor U7441 (N_7441,N_7296,N_7270);
nand U7442 (N_7442,N_7224,N_7262);
and U7443 (N_7443,N_7243,N_7308);
xor U7444 (N_7444,N_7345,N_7240);
nor U7445 (N_7445,N_7215,N_7242);
xor U7446 (N_7446,N_7205,N_7296);
and U7447 (N_7447,N_7350,N_7222);
or U7448 (N_7448,N_7307,N_7334);
or U7449 (N_7449,N_7343,N_7345);
and U7450 (N_7450,N_7349,N_7223);
nand U7451 (N_7451,N_7350,N_7205);
and U7452 (N_7452,N_7346,N_7203);
and U7453 (N_7453,N_7227,N_7275);
nand U7454 (N_7454,N_7204,N_7236);
nor U7455 (N_7455,N_7259,N_7253);
or U7456 (N_7456,N_7354,N_7228);
and U7457 (N_7457,N_7325,N_7227);
nand U7458 (N_7458,N_7330,N_7352);
and U7459 (N_7459,N_7283,N_7341);
or U7460 (N_7460,N_7295,N_7285);
nor U7461 (N_7461,N_7218,N_7304);
xnor U7462 (N_7462,N_7248,N_7344);
nor U7463 (N_7463,N_7205,N_7202);
and U7464 (N_7464,N_7249,N_7231);
or U7465 (N_7465,N_7263,N_7232);
nor U7466 (N_7466,N_7247,N_7235);
and U7467 (N_7467,N_7354,N_7355);
nand U7468 (N_7468,N_7206,N_7308);
or U7469 (N_7469,N_7357,N_7272);
and U7470 (N_7470,N_7324,N_7235);
and U7471 (N_7471,N_7327,N_7227);
nor U7472 (N_7472,N_7268,N_7310);
nor U7473 (N_7473,N_7344,N_7274);
nand U7474 (N_7474,N_7279,N_7229);
and U7475 (N_7475,N_7266,N_7305);
nand U7476 (N_7476,N_7258,N_7225);
nand U7477 (N_7477,N_7319,N_7206);
or U7478 (N_7478,N_7347,N_7335);
or U7479 (N_7479,N_7255,N_7298);
and U7480 (N_7480,N_7203,N_7276);
and U7481 (N_7481,N_7206,N_7218);
nor U7482 (N_7482,N_7241,N_7238);
xor U7483 (N_7483,N_7243,N_7333);
or U7484 (N_7484,N_7252,N_7312);
nor U7485 (N_7485,N_7219,N_7266);
nor U7486 (N_7486,N_7219,N_7272);
xnor U7487 (N_7487,N_7237,N_7210);
nor U7488 (N_7488,N_7307,N_7350);
and U7489 (N_7489,N_7212,N_7340);
nor U7490 (N_7490,N_7254,N_7305);
nor U7491 (N_7491,N_7305,N_7253);
and U7492 (N_7492,N_7297,N_7264);
or U7493 (N_7493,N_7240,N_7227);
and U7494 (N_7494,N_7264,N_7359);
nand U7495 (N_7495,N_7225,N_7288);
or U7496 (N_7496,N_7255,N_7273);
and U7497 (N_7497,N_7262,N_7340);
nor U7498 (N_7498,N_7277,N_7230);
or U7499 (N_7499,N_7352,N_7258);
nand U7500 (N_7500,N_7319,N_7291);
xnor U7501 (N_7501,N_7207,N_7200);
nand U7502 (N_7502,N_7215,N_7356);
nor U7503 (N_7503,N_7246,N_7211);
xor U7504 (N_7504,N_7266,N_7333);
nand U7505 (N_7505,N_7229,N_7287);
nor U7506 (N_7506,N_7241,N_7239);
or U7507 (N_7507,N_7327,N_7322);
and U7508 (N_7508,N_7357,N_7317);
xor U7509 (N_7509,N_7309,N_7216);
nand U7510 (N_7510,N_7299,N_7311);
or U7511 (N_7511,N_7333,N_7273);
nand U7512 (N_7512,N_7353,N_7232);
nand U7513 (N_7513,N_7246,N_7286);
nand U7514 (N_7514,N_7313,N_7268);
or U7515 (N_7515,N_7224,N_7231);
or U7516 (N_7516,N_7250,N_7327);
or U7517 (N_7517,N_7317,N_7200);
or U7518 (N_7518,N_7203,N_7206);
or U7519 (N_7519,N_7316,N_7204);
xor U7520 (N_7520,N_7404,N_7405);
xnor U7521 (N_7521,N_7444,N_7398);
or U7522 (N_7522,N_7454,N_7370);
nand U7523 (N_7523,N_7468,N_7461);
nor U7524 (N_7524,N_7396,N_7377);
and U7525 (N_7525,N_7425,N_7452);
or U7526 (N_7526,N_7515,N_7409);
nor U7527 (N_7527,N_7501,N_7448);
or U7528 (N_7528,N_7465,N_7428);
and U7529 (N_7529,N_7386,N_7446);
or U7530 (N_7530,N_7375,N_7419);
nand U7531 (N_7531,N_7391,N_7469);
nand U7532 (N_7532,N_7431,N_7488);
nor U7533 (N_7533,N_7441,N_7426);
xor U7534 (N_7534,N_7392,N_7407);
or U7535 (N_7535,N_7500,N_7487);
and U7536 (N_7536,N_7514,N_7373);
nor U7537 (N_7537,N_7421,N_7508);
and U7538 (N_7538,N_7434,N_7495);
nor U7539 (N_7539,N_7450,N_7474);
or U7540 (N_7540,N_7384,N_7477);
or U7541 (N_7541,N_7415,N_7463);
and U7542 (N_7542,N_7485,N_7466);
and U7543 (N_7543,N_7381,N_7363);
xnor U7544 (N_7544,N_7511,N_7453);
nand U7545 (N_7545,N_7516,N_7504);
nor U7546 (N_7546,N_7470,N_7494);
nor U7547 (N_7547,N_7395,N_7406);
nor U7548 (N_7548,N_7414,N_7483);
or U7549 (N_7549,N_7430,N_7365);
xnor U7550 (N_7550,N_7372,N_7418);
nor U7551 (N_7551,N_7481,N_7371);
nor U7552 (N_7552,N_7496,N_7394);
xnor U7553 (N_7553,N_7378,N_7459);
nor U7554 (N_7554,N_7423,N_7376);
nand U7555 (N_7555,N_7447,N_7507);
and U7556 (N_7556,N_7490,N_7369);
nand U7557 (N_7557,N_7416,N_7361);
nor U7558 (N_7558,N_7512,N_7429);
nor U7559 (N_7559,N_7438,N_7451);
xor U7560 (N_7560,N_7519,N_7517);
xor U7561 (N_7561,N_7368,N_7499);
nor U7562 (N_7562,N_7417,N_7367);
and U7563 (N_7563,N_7456,N_7445);
nor U7564 (N_7564,N_7401,N_7399);
nor U7565 (N_7565,N_7413,N_7506);
or U7566 (N_7566,N_7410,N_7390);
nor U7567 (N_7567,N_7482,N_7497);
xor U7568 (N_7568,N_7489,N_7433);
nor U7569 (N_7569,N_7412,N_7443);
and U7570 (N_7570,N_7440,N_7380);
or U7571 (N_7571,N_7389,N_7432);
nand U7572 (N_7572,N_7400,N_7436);
or U7573 (N_7573,N_7518,N_7364);
nand U7574 (N_7574,N_7422,N_7397);
or U7575 (N_7575,N_7472,N_7460);
nand U7576 (N_7576,N_7491,N_7437);
nor U7577 (N_7577,N_7493,N_7457);
nand U7578 (N_7578,N_7478,N_7484);
xnor U7579 (N_7579,N_7476,N_7479);
nor U7580 (N_7580,N_7435,N_7439);
nor U7581 (N_7581,N_7467,N_7374);
and U7582 (N_7582,N_7473,N_7360);
or U7583 (N_7583,N_7510,N_7403);
nor U7584 (N_7584,N_7480,N_7366);
nor U7585 (N_7585,N_7505,N_7402);
or U7586 (N_7586,N_7427,N_7408);
or U7587 (N_7587,N_7424,N_7502);
or U7588 (N_7588,N_7486,N_7509);
nor U7589 (N_7589,N_7420,N_7462);
or U7590 (N_7590,N_7379,N_7458);
and U7591 (N_7591,N_7475,N_7471);
nor U7592 (N_7592,N_7442,N_7464);
or U7593 (N_7593,N_7513,N_7383);
and U7594 (N_7594,N_7382,N_7498);
nand U7595 (N_7595,N_7385,N_7411);
nor U7596 (N_7596,N_7492,N_7387);
and U7597 (N_7597,N_7362,N_7503);
nor U7598 (N_7598,N_7449,N_7388);
nand U7599 (N_7599,N_7455,N_7393);
nor U7600 (N_7600,N_7396,N_7389);
nor U7601 (N_7601,N_7485,N_7491);
or U7602 (N_7602,N_7461,N_7492);
nand U7603 (N_7603,N_7427,N_7381);
or U7604 (N_7604,N_7469,N_7442);
nand U7605 (N_7605,N_7403,N_7459);
nor U7606 (N_7606,N_7510,N_7395);
and U7607 (N_7607,N_7503,N_7396);
nor U7608 (N_7608,N_7379,N_7382);
nand U7609 (N_7609,N_7503,N_7370);
nand U7610 (N_7610,N_7389,N_7368);
nor U7611 (N_7611,N_7481,N_7398);
nand U7612 (N_7612,N_7365,N_7479);
and U7613 (N_7613,N_7463,N_7416);
and U7614 (N_7614,N_7455,N_7373);
and U7615 (N_7615,N_7507,N_7512);
nor U7616 (N_7616,N_7457,N_7504);
nand U7617 (N_7617,N_7491,N_7488);
and U7618 (N_7618,N_7410,N_7363);
nand U7619 (N_7619,N_7507,N_7465);
nand U7620 (N_7620,N_7503,N_7424);
and U7621 (N_7621,N_7493,N_7477);
nor U7622 (N_7622,N_7405,N_7483);
nand U7623 (N_7623,N_7437,N_7477);
nand U7624 (N_7624,N_7395,N_7410);
or U7625 (N_7625,N_7452,N_7487);
or U7626 (N_7626,N_7451,N_7489);
nor U7627 (N_7627,N_7407,N_7372);
or U7628 (N_7628,N_7387,N_7457);
and U7629 (N_7629,N_7498,N_7499);
nor U7630 (N_7630,N_7507,N_7459);
or U7631 (N_7631,N_7497,N_7360);
or U7632 (N_7632,N_7423,N_7422);
nand U7633 (N_7633,N_7385,N_7395);
or U7634 (N_7634,N_7472,N_7517);
or U7635 (N_7635,N_7490,N_7502);
nor U7636 (N_7636,N_7403,N_7430);
and U7637 (N_7637,N_7444,N_7510);
nor U7638 (N_7638,N_7404,N_7459);
nor U7639 (N_7639,N_7461,N_7421);
xor U7640 (N_7640,N_7462,N_7487);
or U7641 (N_7641,N_7491,N_7374);
and U7642 (N_7642,N_7380,N_7450);
or U7643 (N_7643,N_7466,N_7481);
or U7644 (N_7644,N_7362,N_7420);
xnor U7645 (N_7645,N_7419,N_7371);
nor U7646 (N_7646,N_7440,N_7412);
xor U7647 (N_7647,N_7440,N_7360);
nor U7648 (N_7648,N_7448,N_7481);
xor U7649 (N_7649,N_7418,N_7377);
and U7650 (N_7650,N_7427,N_7461);
nand U7651 (N_7651,N_7454,N_7471);
nor U7652 (N_7652,N_7403,N_7437);
or U7653 (N_7653,N_7437,N_7449);
nand U7654 (N_7654,N_7437,N_7395);
and U7655 (N_7655,N_7471,N_7421);
nor U7656 (N_7656,N_7505,N_7416);
or U7657 (N_7657,N_7492,N_7372);
nand U7658 (N_7658,N_7469,N_7425);
nor U7659 (N_7659,N_7407,N_7425);
or U7660 (N_7660,N_7380,N_7397);
or U7661 (N_7661,N_7434,N_7468);
nand U7662 (N_7662,N_7504,N_7384);
nor U7663 (N_7663,N_7423,N_7435);
nand U7664 (N_7664,N_7421,N_7418);
or U7665 (N_7665,N_7399,N_7403);
or U7666 (N_7666,N_7508,N_7499);
or U7667 (N_7667,N_7496,N_7501);
nand U7668 (N_7668,N_7434,N_7441);
or U7669 (N_7669,N_7412,N_7505);
xor U7670 (N_7670,N_7488,N_7449);
and U7671 (N_7671,N_7377,N_7372);
or U7672 (N_7672,N_7376,N_7451);
or U7673 (N_7673,N_7369,N_7360);
nor U7674 (N_7674,N_7411,N_7434);
or U7675 (N_7675,N_7374,N_7453);
nor U7676 (N_7676,N_7386,N_7438);
or U7677 (N_7677,N_7473,N_7482);
nand U7678 (N_7678,N_7429,N_7441);
nor U7679 (N_7679,N_7481,N_7363);
nor U7680 (N_7680,N_7592,N_7596);
or U7681 (N_7681,N_7569,N_7588);
and U7682 (N_7682,N_7605,N_7616);
nand U7683 (N_7683,N_7527,N_7587);
nor U7684 (N_7684,N_7645,N_7671);
nand U7685 (N_7685,N_7624,N_7593);
nor U7686 (N_7686,N_7599,N_7563);
and U7687 (N_7687,N_7545,N_7608);
nor U7688 (N_7688,N_7555,N_7615);
and U7689 (N_7689,N_7613,N_7675);
xnor U7690 (N_7690,N_7576,N_7641);
or U7691 (N_7691,N_7667,N_7663);
nand U7692 (N_7692,N_7521,N_7558);
nand U7693 (N_7693,N_7551,N_7575);
nand U7694 (N_7694,N_7670,N_7535);
or U7695 (N_7695,N_7553,N_7620);
or U7696 (N_7696,N_7666,N_7570);
and U7697 (N_7697,N_7562,N_7656);
or U7698 (N_7698,N_7638,N_7533);
nor U7699 (N_7699,N_7600,N_7668);
nand U7700 (N_7700,N_7526,N_7590);
or U7701 (N_7701,N_7658,N_7578);
and U7702 (N_7702,N_7547,N_7665);
and U7703 (N_7703,N_7652,N_7660);
or U7704 (N_7704,N_7607,N_7540);
xor U7705 (N_7705,N_7612,N_7530);
nand U7706 (N_7706,N_7609,N_7617);
xor U7707 (N_7707,N_7522,N_7633);
nand U7708 (N_7708,N_7678,N_7618);
xor U7709 (N_7709,N_7661,N_7543);
and U7710 (N_7710,N_7669,N_7655);
or U7711 (N_7711,N_7647,N_7597);
or U7712 (N_7712,N_7623,N_7581);
and U7713 (N_7713,N_7525,N_7589);
and U7714 (N_7714,N_7546,N_7582);
nand U7715 (N_7715,N_7625,N_7603);
and U7716 (N_7716,N_7573,N_7559);
and U7717 (N_7717,N_7567,N_7637);
or U7718 (N_7718,N_7649,N_7614);
nand U7719 (N_7719,N_7564,N_7601);
nand U7720 (N_7720,N_7550,N_7536);
and U7721 (N_7721,N_7539,N_7561);
nand U7722 (N_7722,N_7523,N_7594);
nand U7723 (N_7723,N_7579,N_7586);
nand U7724 (N_7724,N_7664,N_7648);
xnor U7725 (N_7725,N_7548,N_7529);
and U7726 (N_7726,N_7630,N_7606);
nand U7727 (N_7727,N_7644,N_7532);
nand U7728 (N_7728,N_7534,N_7541);
or U7729 (N_7729,N_7676,N_7650);
and U7730 (N_7730,N_7574,N_7528);
or U7731 (N_7731,N_7677,N_7591);
nand U7732 (N_7732,N_7571,N_7626);
nor U7733 (N_7733,N_7556,N_7657);
or U7734 (N_7734,N_7572,N_7673);
nand U7735 (N_7735,N_7622,N_7674);
nand U7736 (N_7736,N_7628,N_7639);
nand U7737 (N_7737,N_7560,N_7544);
nand U7738 (N_7738,N_7679,N_7636);
and U7739 (N_7739,N_7610,N_7557);
nor U7740 (N_7740,N_7554,N_7542);
nor U7741 (N_7741,N_7565,N_7566);
and U7742 (N_7742,N_7659,N_7646);
nor U7743 (N_7743,N_7549,N_7584);
and U7744 (N_7744,N_7568,N_7619);
or U7745 (N_7745,N_7538,N_7524);
or U7746 (N_7746,N_7520,N_7662);
and U7747 (N_7747,N_7653,N_7577);
or U7748 (N_7748,N_7635,N_7643);
nand U7749 (N_7749,N_7611,N_7604);
and U7750 (N_7750,N_7627,N_7598);
or U7751 (N_7751,N_7629,N_7580);
nand U7752 (N_7752,N_7583,N_7632);
and U7753 (N_7753,N_7642,N_7531);
or U7754 (N_7754,N_7585,N_7672);
or U7755 (N_7755,N_7621,N_7640);
and U7756 (N_7756,N_7602,N_7634);
nor U7757 (N_7757,N_7631,N_7651);
xor U7758 (N_7758,N_7595,N_7552);
nor U7759 (N_7759,N_7654,N_7537);
nor U7760 (N_7760,N_7627,N_7658);
and U7761 (N_7761,N_7577,N_7630);
or U7762 (N_7762,N_7645,N_7585);
nor U7763 (N_7763,N_7631,N_7544);
nor U7764 (N_7764,N_7666,N_7542);
or U7765 (N_7765,N_7588,N_7619);
and U7766 (N_7766,N_7639,N_7575);
and U7767 (N_7767,N_7634,N_7542);
or U7768 (N_7768,N_7624,N_7598);
or U7769 (N_7769,N_7608,N_7562);
nor U7770 (N_7770,N_7604,N_7613);
xor U7771 (N_7771,N_7626,N_7648);
nand U7772 (N_7772,N_7574,N_7639);
and U7773 (N_7773,N_7655,N_7547);
nand U7774 (N_7774,N_7672,N_7646);
and U7775 (N_7775,N_7589,N_7665);
nor U7776 (N_7776,N_7543,N_7525);
and U7777 (N_7777,N_7615,N_7599);
nand U7778 (N_7778,N_7622,N_7660);
nand U7779 (N_7779,N_7612,N_7563);
and U7780 (N_7780,N_7660,N_7570);
nand U7781 (N_7781,N_7564,N_7617);
nor U7782 (N_7782,N_7569,N_7528);
nor U7783 (N_7783,N_7546,N_7529);
nand U7784 (N_7784,N_7584,N_7616);
nand U7785 (N_7785,N_7557,N_7568);
or U7786 (N_7786,N_7562,N_7537);
nor U7787 (N_7787,N_7524,N_7620);
and U7788 (N_7788,N_7661,N_7588);
nor U7789 (N_7789,N_7598,N_7569);
or U7790 (N_7790,N_7532,N_7641);
xor U7791 (N_7791,N_7634,N_7555);
or U7792 (N_7792,N_7648,N_7564);
xnor U7793 (N_7793,N_7640,N_7553);
or U7794 (N_7794,N_7650,N_7575);
nor U7795 (N_7795,N_7575,N_7583);
nor U7796 (N_7796,N_7634,N_7603);
or U7797 (N_7797,N_7573,N_7608);
nand U7798 (N_7798,N_7569,N_7589);
or U7799 (N_7799,N_7627,N_7629);
and U7800 (N_7800,N_7662,N_7660);
and U7801 (N_7801,N_7587,N_7649);
xor U7802 (N_7802,N_7540,N_7537);
or U7803 (N_7803,N_7562,N_7570);
and U7804 (N_7804,N_7654,N_7671);
or U7805 (N_7805,N_7621,N_7566);
nor U7806 (N_7806,N_7635,N_7608);
or U7807 (N_7807,N_7575,N_7632);
and U7808 (N_7808,N_7562,N_7544);
and U7809 (N_7809,N_7549,N_7658);
or U7810 (N_7810,N_7578,N_7650);
nand U7811 (N_7811,N_7536,N_7532);
or U7812 (N_7812,N_7613,N_7643);
and U7813 (N_7813,N_7545,N_7570);
nand U7814 (N_7814,N_7651,N_7625);
or U7815 (N_7815,N_7546,N_7579);
xor U7816 (N_7816,N_7656,N_7592);
or U7817 (N_7817,N_7652,N_7579);
xor U7818 (N_7818,N_7604,N_7585);
and U7819 (N_7819,N_7599,N_7606);
nand U7820 (N_7820,N_7625,N_7604);
and U7821 (N_7821,N_7589,N_7617);
nand U7822 (N_7822,N_7553,N_7582);
nor U7823 (N_7823,N_7625,N_7653);
and U7824 (N_7824,N_7656,N_7653);
nor U7825 (N_7825,N_7657,N_7520);
and U7826 (N_7826,N_7655,N_7584);
or U7827 (N_7827,N_7525,N_7569);
or U7828 (N_7828,N_7617,N_7652);
nand U7829 (N_7829,N_7591,N_7629);
nor U7830 (N_7830,N_7643,N_7671);
xor U7831 (N_7831,N_7674,N_7600);
nand U7832 (N_7832,N_7526,N_7675);
and U7833 (N_7833,N_7653,N_7655);
nor U7834 (N_7834,N_7525,N_7562);
nand U7835 (N_7835,N_7645,N_7637);
xnor U7836 (N_7836,N_7636,N_7524);
nor U7837 (N_7837,N_7658,N_7562);
or U7838 (N_7838,N_7597,N_7605);
and U7839 (N_7839,N_7571,N_7528);
nor U7840 (N_7840,N_7790,N_7837);
and U7841 (N_7841,N_7753,N_7823);
xor U7842 (N_7842,N_7736,N_7771);
or U7843 (N_7843,N_7698,N_7755);
and U7844 (N_7844,N_7706,N_7821);
and U7845 (N_7845,N_7718,N_7805);
xor U7846 (N_7846,N_7734,N_7731);
or U7847 (N_7847,N_7713,N_7686);
and U7848 (N_7848,N_7705,N_7722);
or U7849 (N_7849,N_7737,N_7817);
nand U7850 (N_7850,N_7785,N_7752);
nand U7851 (N_7851,N_7717,N_7779);
and U7852 (N_7852,N_7758,N_7830);
or U7853 (N_7853,N_7802,N_7723);
or U7854 (N_7854,N_7816,N_7749);
nand U7855 (N_7855,N_7747,N_7712);
and U7856 (N_7856,N_7738,N_7693);
or U7857 (N_7857,N_7794,N_7814);
nand U7858 (N_7858,N_7764,N_7746);
and U7859 (N_7859,N_7804,N_7715);
nand U7860 (N_7860,N_7766,N_7699);
and U7861 (N_7861,N_7768,N_7756);
xnor U7862 (N_7862,N_7739,N_7838);
or U7863 (N_7863,N_7819,N_7767);
nor U7864 (N_7864,N_7730,N_7743);
or U7865 (N_7865,N_7820,N_7694);
or U7866 (N_7866,N_7810,N_7789);
and U7867 (N_7867,N_7827,N_7726);
nor U7868 (N_7868,N_7772,N_7688);
nor U7869 (N_7869,N_7719,N_7782);
and U7870 (N_7870,N_7733,N_7702);
nor U7871 (N_7871,N_7806,N_7818);
or U7872 (N_7872,N_7711,N_7780);
nand U7873 (N_7873,N_7708,N_7799);
nand U7874 (N_7874,N_7788,N_7811);
nor U7875 (N_7875,N_7687,N_7696);
xor U7876 (N_7876,N_7689,N_7761);
nor U7877 (N_7877,N_7710,N_7792);
and U7878 (N_7878,N_7701,N_7833);
nand U7879 (N_7879,N_7783,N_7808);
nor U7880 (N_7880,N_7839,N_7815);
xnor U7881 (N_7881,N_7797,N_7685);
or U7882 (N_7882,N_7769,N_7728);
nor U7883 (N_7883,N_7742,N_7690);
nor U7884 (N_7884,N_7721,N_7732);
or U7885 (N_7885,N_7824,N_7709);
or U7886 (N_7886,N_7700,N_7703);
or U7887 (N_7887,N_7809,N_7750);
nand U7888 (N_7888,N_7781,N_7775);
nand U7889 (N_7889,N_7836,N_7727);
nor U7890 (N_7890,N_7751,N_7807);
nand U7891 (N_7891,N_7813,N_7759);
nand U7892 (N_7892,N_7812,N_7825);
and U7893 (N_7893,N_7692,N_7695);
nand U7894 (N_7894,N_7777,N_7828);
nor U7895 (N_7895,N_7822,N_7725);
nor U7896 (N_7896,N_7740,N_7757);
nand U7897 (N_7897,N_7795,N_7714);
and U7898 (N_7898,N_7691,N_7786);
nor U7899 (N_7899,N_7826,N_7791);
nand U7900 (N_7900,N_7720,N_7704);
or U7901 (N_7901,N_7716,N_7796);
and U7902 (N_7902,N_7697,N_7778);
or U7903 (N_7903,N_7798,N_7835);
nor U7904 (N_7904,N_7741,N_7776);
nand U7905 (N_7905,N_7801,N_7829);
nand U7906 (N_7906,N_7684,N_7682);
and U7907 (N_7907,N_7773,N_7770);
nand U7908 (N_7908,N_7831,N_7681);
or U7909 (N_7909,N_7793,N_7784);
nor U7910 (N_7910,N_7748,N_7832);
nand U7911 (N_7911,N_7765,N_7680);
nor U7912 (N_7912,N_7760,N_7724);
nor U7913 (N_7913,N_7735,N_7803);
nand U7914 (N_7914,N_7800,N_7744);
and U7915 (N_7915,N_7763,N_7774);
and U7916 (N_7916,N_7834,N_7707);
or U7917 (N_7917,N_7762,N_7729);
and U7918 (N_7918,N_7745,N_7754);
nor U7919 (N_7919,N_7683,N_7787);
nor U7920 (N_7920,N_7776,N_7687);
or U7921 (N_7921,N_7684,N_7764);
and U7922 (N_7922,N_7823,N_7772);
and U7923 (N_7923,N_7688,N_7817);
nor U7924 (N_7924,N_7794,N_7804);
and U7925 (N_7925,N_7801,N_7765);
nand U7926 (N_7926,N_7775,N_7696);
nand U7927 (N_7927,N_7685,N_7836);
nor U7928 (N_7928,N_7692,N_7839);
or U7929 (N_7929,N_7727,N_7724);
and U7930 (N_7930,N_7775,N_7731);
and U7931 (N_7931,N_7734,N_7783);
nor U7932 (N_7932,N_7720,N_7776);
nand U7933 (N_7933,N_7808,N_7810);
nand U7934 (N_7934,N_7709,N_7699);
nand U7935 (N_7935,N_7785,N_7684);
or U7936 (N_7936,N_7693,N_7683);
and U7937 (N_7937,N_7782,N_7833);
nand U7938 (N_7938,N_7762,N_7690);
nand U7939 (N_7939,N_7716,N_7686);
nor U7940 (N_7940,N_7819,N_7830);
or U7941 (N_7941,N_7708,N_7824);
nor U7942 (N_7942,N_7750,N_7711);
and U7943 (N_7943,N_7725,N_7763);
and U7944 (N_7944,N_7795,N_7832);
nand U7945 (N_7945,N_7723,N_7717);
nand U7946 (N_7946,N_7770,N_7826);
or U7947 (N_7947,N_7763,N_7785);
nor U7948 (N_7948,N_7716,N_7724);
nand U7949 (N_7949,N_7691,N_7827);
nor U7950 (N_7950,N_7726,N_7684);
nor U7951 (N_7951,N_7794,N_7698);
or U7952 (N_7952,N_7736,N_7699);
nor U7953 (N_7953,N_7755,N_7821);
nand U7954 (N_7954,N_7759,N_7824);
nand U7955 (N_7955,N_7800,N_7709);
xor U7956 (N_7956,N_7839,N_7827);
nor U7957 (N_7957,N_7736,N_7712);
nor U7958 (N_7958,N_7788,N_7707);
nor U7959 (N_7959,N_7758,N_7727);
nor U7960 (N_7960,N_7761,N_7781);
nor U7961 (N_7961,N_7687,N_7768);
xor U7962 (N_7962,N_7785,N_7764);
nor U7963 (N_7963,N_7730,N_7832);
nor U7964 (N_7964,N_7800,N_7742);
or U7965 (N_7965,N_7722,N_7696);
and U7966 (N_7966,N_7708,N_7800);
or U7967 (N_7967,N_7772,N_7807);
nand U7968 (N_7968,N_7788,N_7766);
nand U7969 (N_7969,N_7795,N_7680);
nor U7970 (N_7970,N_7729,N_7759);
nor U7971 (N_7971,N_7694,N_7794);
xnor U7972 (N_7972,N_7730,N_7751);
nor U7973 (N_7973,N_7759,N_7764);
or U7974 (N_7974,N_7707,N_7809);
nand U7975 (N_7975,N_7772,N_7744);
nand U7976 (N_7976,N_7729,N_7706);
nor U7977 (N_7977,N_7682,N_7685);
nand U7978 (N_7978,N_7686,N_7808);
nand U7979 (N_7979,N_7716,N_7698);
nor U7980 (N_7980,N_7684,N_7787);
nor U7981 (N_7981,N_7799,N_7814);
nor U7982 (N_7982,N_7801,N_7806);
and U7983 (N_7983,N_7774,N_7728);
and U7984 (N_7984,N_7827,N_7709);
nor U7985 (N_7985,N_7798,N_7765);
nor U7986 (N_7986,N_7705,N_7823);
nor U7987 (N_7987,N_7813,N_7832);
and U7988 (N_7988,N_7741,N_7705);
nor U7989 (N_7989,N_7813,N_7770);
xor U7990 (N_7990,N_7836,N_7805);
nand U7991 (N_7991,N_7717,N_7761);
xnor U7992 (N_7992,N_7702,N_7809);
nand U7993 (N_7993,N_7777,N_7681);
or U7994 (N_7994,N_7778,N_7785);
nor U7995 (N_7995,N_7729,N_7783);
nor U7996 (N_7996,N_7774,N_7720);
or U7997 (N_7997,N_7763,N_7748);
and U7998 (N_7998,N_7724,N_7711);
nor U7999 (N_7999,N_7790,N_7704);
nand U8000 (N_8000,N_7940,N_7867);
or U8001 (N_8001,N_7922,N_7987);
or U8002 (N_8002,N_7902,N_7928);
and U8003 (N_8003,N_7886,N_7926);
nand U8004 (N_8004,N_7997,N_7988);
and U8005 (N_8005,N_7854,N_7935);
and U8006 (N_8006,N_7893,N_7906);
and U8007 (N_8007,N_7876,N_7904);
xnor U8008 (N_8008,N_7979,N_7930);
and U8009 (N_8009,N_7934,N_7966);
nand U8010 (N_8010,N_7998,N_7957);
nand U8011 (N_8011,N_7980,N_7999);
or U8012 (N_8012,N_7950,N_7982);
or U8013 (N_8013,N_7941,N_7916);
nor U8014 (N_8014,N_7956,N_7905);
and U8015 (N_8015,N_7921,N_7967);
or U8016 (N_8016,N_7885,N_7920);
nand U8017 (N_8017,N_7910,N_7841);
and U8018 (N_8018,N_7970,N_7911);
and U8019 (N_8019,N_7960,N_7882);
and U8020 (N_8020,N_7949,N_7975);
and U8021 (N_8021,N_7874,N_7938);
or U8022 (N_8022,N_7881,N_7917);
nand U8023 (N_8023,N_7878,N_7986);
nor U8024 (N_8024,N_7851,N_7948);
nor U8025 (N_8025,N_7981,N_7984);
or U8026 (N_8026,N_7962,N_7945);
xor U8027 (N_8027,N_7925,N_7865);
nor U8028 (N_8028,N_7864,N_7844);
and U8029 (N_8029,N_7855,N_7872);
and U8030 (N_8030,N_7994,N_7860);
and U8031 (N_8031,N_7899,N_7900);
nor U8032 (N_8032,N_7908,N_7919);
or U8033 (N_8033,N_7840,N_7964);
or U8034 (N_8034,N_7901,N_7883);
or U8035 (N_8035,N_7850,N_7976);
nand U8036 (N_8036,N_7959,N_7863);
or U8037 (N_8037,N_7873,N_7869);
xor U8038 (N_8038,N_7858,N_7955);
nand U8039 (N_8039,N_7990,N_7870);
or U8040 (N_8040,N_7947,N_7965);
nor U8041 (N_8041,N_7845,N_7903);
xnor U8042 (N_8042,N_7862,N_7937);
or U8043 (N_8043,N_7857,N_7958);
nor U8044 (N_8044,N_7896,N_7961);
or U8045 (N_8045,N_7929,N_7952);
nor U8046 (N_8046,N_7932,N_7879);
nor U8047 (N_8047,N_7891,N_7871);
or U8048 (N_8048,N_7847,N_7996);
and U8049 (N_8049,N_7861,N_7924);
nor U8050 (N_8050,N_7907,N_7954);
nand U8051 (N_8051,N_7895,N_7927);
or U8052 (N_8052,N_7889,N_7985);
and U8053 (N_8053,N_7913,N_7969);
or U8054 (N_8054,N_7868,N_7993);
or U8055 (N_8055,N_7914,N_7953);
or U8056 (N_8056,N_7944,N_7973);
or U8057 (N_8057,N_7971,N_7888);
and U8058 (N_8058,N_7951,N_7892);
or U8059 (N_8059,N_7974,N_7897);
and U8060 (N_8060,N_7918,N_7848);
and U8061 (N_8061,N_7849,N_7912);
nand U8062 (N_8062,N_7936,N_7890);
or U8063 (N_8063,N_7853,N_7843);
and U8064 (N_8064,N_7931,N_7877);
and U8065 (N_8065,N_7842,N_7968);
and U8066 (N_8066,N_7946,N_7972);
xor U8067 (N_8067,N_7859,N_7866);
nand U8068 (N_8068,N_7939,N_7992);
nand U8069 (N_8069,N_7887,N_7923);
or U8070 (N_8070,N_7898,N_7909);
nor U8071 (N_8071,N_7991,N_7856);
or U8072 (N_8072,N_7942,N_7846);
or U8073 (N_8073,N_7943,N_7880);
nand U8074 (N_8074,N_7978,N_7915);
nand U8075 (N_8075,N_7989,N_7963);
or U8076 (N_8076,N_7977,N_7933);
and U8077 (N_8077,N_7852,N_7894);
nor U8078 (N_8078,N_7884,N_7995);
and U8079 (N_8079,N_7983,N_7875);
and U8080 (N_8080,N_7908,N_7996);
and U8081 (N_8081,N_7960,N_7876);
or U8082 (N_8082,N_7971,N_7952);
and U8083 (N_8083,N_7915,N_7896);
or U8084 (N_8084,N_7927,N_7955);
nor U8085 (N_8085,N_7848,N_7904);
and U8086 (N_8086,N_7905,N_7904);
nor U8087 (N_8087,N_7926,N_7929);
or U8088 (N_8088,N_7947,N_7909);
nand U8089 (N_8089,N_7970,N_7866);
and U8090 (N_8090,N_7961,N_7937);
xor U8091 (N_8091,N_7982,N_7893);
nand U8092 (N_8092,N_7982,N_7947);
nand U8093 (N_8093,N_7851,N_7895);
nor U8094 (N_8094,N_7860,N_7870);
nor U8095 (N_8095,N_7854,N_7872);
nor U8096 (N_8096,N_7970,N_7953);
and U8097 (N_8097,N_7926,N_7869);
xor U8098 (N_8098,N_7943,N_7913);
nor U8099 (N_8099,N_7923,N_7968);
nor U8100 (N_8100,N_7943,N_7879);
or U8101 (N_8101,N_7842,N_7939);
and U8102 (N_8102,N_7990,N_7989);
and U8103 (N_8103,N_7984,N_7977);
or U8104 (N_8104,N_7911,N_7961);
nand U8105 (N_8105,N_7869,N_7910);
nor U8106 (N_8106,N_7882,N_7845);
nand U8107 (N_8107,N_7968,N_7981);
or U8108 (N_8108,N_7908,N_7961);
or U8109 (N_8109,N_7973,N_7870);
nor U8110 (N_8110,N_7938,N_7840);
and U8111 (N_8111,N_7866,N_7844);
and U8112 (N_8112,N_7865,N_7910);
nand U8113 (N_8113,N_7934,N_7945);
nand U8114 (N_8114,N_7866,N_7849);
or U8115 (N_8115,N_7901,N_7906);
and U8116 (N_8116,N_7865,N_7974);
nor U8117 (N_8117,N_7878,N_7883);
xor U8118 (N_8118,N_7918,N_7995);
and U8119 (N_8119,N_7850,N_7844);
nor U8120 (N_8120,N_7859,N_7902);
and U8121 (N_8121,N_7880,N_7972);
nand U8122 (N_8122,N_7942,N_7930);
xor U8123 (N_8123,N_7973,N_7909);
nor U8124 (N_8124,N_7873,N_7902);
nor U8125 (N_8125,N_7955,N_7937);
or U8126 (N_8126,N_7947,N_7876);
or U8127 (N_8127,N_7910,N_7904);
nor U8128 (N_8128,N_7923,N_7877);
nand U8129 (N_8129,N_7914,N_7951);
or U8130 (N_8130,N_7877,N_7988);
nor U8131 (N_8131,N_7901,N_7848);
nor U8132 (N_8132,N_7910,N_7913);
nand U8133 (N_8133,N_7994,N_7996);
and U8134 (N_8134,N_7901,N_7853);
or U8135 (N_8135,N_7912,N_7851);
and U8136 (N_8136,N_7961,N_7900);
or U8137 (N_8137,N_7934,N_7841);
nor U8138 (N_8138,N_7944,N_7937);
and U8139 (N_8139,N_7856,N_7875);
nand U8140 (N_8140,N_7964,N_7928);
nand U8141 (N_8141,N_7964,N_7956);
nor U8142 (N_8142,N_7860,N_7962);
or U8143 (N_8143,N_7950,N_7957);
nand U8144 (N_8144,N_7871,N_7925);
nor U8145 (N_8145,N_7849,N_7956);
or U8146 (N_8146,N_7913,N_7898);
and U8147 (N_8147,N_7971,N_7899);
xor U8148 (N_8148,N_7967,N_7912);
or U8149 (N_8149,N_7855,N_7876);
and U8150 (N_8150,N_7901,N_7843);
or U8151 (N_8151,N_7941,N_7847);
and U8152 (N_8152,N_7914,N_7964);
nand U8153 (N_8153,N_7978,N_7961);
nor U8154 (N_8154,N_7973,N_7993);
and U8155 (N_8155,N_7940,N_7909);
nor U8156 (N_8156,N_7979,N_7952);
and U8157 (N_8157,N_7923,N_7866);
nand U8158 (N_8158,N_7938,N_7922);
nor U8159 (N_8159,N_7935,N_7941);
and U8160 (N_8160,N_8099,N_8101);
and U8161 (N_8161,N_8027,N_8014);
or U8162 (N_8162,N_8047,N_8147);
or U8163 (N_8163,N_8151,N_8034);
and U8164 (N_8164,N_8077,N_8007);
or U8165 (N_8165,N_8158,N_8030);
nand U8166 (N_8166,N_8136,N_8005);
xor U8167 (N_8167,N_8145,N_8066);
or U8168 (N_8168,N_8017,N_8002);
nand U8169 (N_8169,N_8056,N_8115);
nand U8170 (N_8170,N_8111,N_8092);
xnor U8171 (N_8171,N_8113,N_8057);
and U8172 (N_8172,N_8137,N_8024);
nor U8173 (N_8173,N_8094,N_8036);
and U8174 (N_8174,N_8029,N_8083);
and U8175 (N_8175,N_8001,N_8058);
or U8176 (N_8176,N_8096,N_8097);
or U8177 (N_8177,N_8100,N_8104);
nor U8178 (N_8178,N_8102,N_8045);
xor U8179 (N_8179,N_8086,N_8146);
xnor U8180 (N_8180,N_8084,N_8128);
and U8181 (N_8181,N_8125,N_8008);
nand U8182 (N_8182,N_8032,N_8148);
xnor U8183 (N_8183,N_8012,N_8078);
nand U8184 (N_8184,N_8043,N_8067);
or U8185 (N_8185,N_8103,N_8018);
xor U8186 (N_8186,N_8107,N_8031);
nand U8187 (N_8187,N_8140,N_8046);
or U8188 (N_8188,N_8009,N_8112);
nor U8189 (N_8189,N_8028,N_8091);
nand U8190 (N_8190,N_8124,N_8068);
or U8191 (N_8191,N_8055,N_8079);
nor U8192 (N_8192,N_8123,N_8120);
or U8193 (N_8193,N_8061,N_8116);
nor U8194 (N_8194,N_8042,N_8053);
nand U8195 (N_8195,N_8135,N_8082);
nor U8196 (N_8196,N_8114,N_8130);
nand U8197 (N_8197,N_8000,N_8073);
and U8198 (N_8198,N_8015,N_8011);
nand U8199 (N_8199,N_8003,N_8106);
or U8200 (N_8200,N_8022,N_8037);
and U8201 (N_8201,N_8155,N_8010);
and U8202 (N_8202,N_8087,N_8006);
nand U8203 (N_8203,N_8072,N_8150);
or U8204 (N_8204,N_8144,N_8133);
or U8205 (N_8205,N_8134,N_8059);
and U8206 (N_8206,N_8142,N_8090);
nor U8207 (N_8207,N_8019,N_8089);
nor U8208 (N_8208,N_8025,N_8095);
nand U8209 (N_8209,N_8063,N_8080);
nor U8210 (N_8210,N_8038,N_8035);
and U8211 (N_8211,N_8126,N_8052);
nor U8212 (N_8212,N_8121,N_8044);
nand U8213 (N_8213,N_8088,N_8143);
or U8214 (N_8214,N_8020,N_8051);
and U8215 (N_8215,N_8156,N_8153);
nor U8216 (N_8216,N_8039,N_8070);
nand U8217 (N_8217,N_8033,N_8081);
nand U8218 (N_8218,N_8131,N_8054);
nor U8219 (N_8219,N_8129,N_8064);
xnor U8220 (N_8220,N_8105,N_8050);
nand U8221 (N_8221,N_8074,N_8071);
nand U8222 (N_8222,N_8049,N_8085);
and U8223 (N_8223,N_8110,N_8118);
xnor U8224 (N_8224,N_8093,N_8023);
and U8225 (N_8225,N_8152,N_8139);
and U8226 (N_8226,N_8109,N_8119);
and U8227 (N_8227,N_8021,N_8108);
and U8228 (N_8228,N_8117,N_8157);
xnor U8229 (N_8229,N_8041,N_8076);
or U8230 (N_8230,N_8040,N_8138);
or U8231 (N_8231,N_8122,N_8069);
xnor U8232 (N_8232,N_8127,N_8149);
or U8233 (N_8233,N_8013,N_8065);
nor U8234 (N_8234,N_8154,N_8062);
or U8235 (N_8235,N_8048,N_8016);
nor U8236 (N_8236,N_8004,N_8141);
xor U8237 (N_8237,N_8075,N_8159);
or U8238 (N_8238,N_8098,N_8060);
nand U8239 (N_8239,N_8026,N_8132);
or U8240 (N_8240,N_8000,N_8047);
nor U8241 (N_8241,N_8039,N_8110);
nor U8242 (N_8242,N_8028,N_8023);
nor U8243 (N_8243,N_8149,N_8153);
nand U8244 (N_8244,N_8131,N_8107);
nor U8245 (N_8245,N_8047,N_8024);
and U8246 (N_8246,N_8104,N_8000);
xnor U8247 (N_8247,N_8068,N_8074);
xor U8248 (N_8248,N_8075,N_8066);
nor U8249 (N_8249,N_8023,N_8077);
and U8250 (N_8250,N_8072,N_8013);
nor U8251 (N_8251,N_8071,N_8136);
or U8252 (N_8252,N_8135,N_8079);
nor U8253 (N_8253,N_8026,N_8007);
nand U8254 (N_8254,N_8110,N_8073);
nand U8255 (N_8255,N_8054,N_8107);
or U8256 (N_8256,N_8015,N_8131);
xor U8257 (N_8257,N_8045,N_8018);
nor U8258 (N_8258,N_8035,N_8154);
nor U8259 (N_8259,N_8066,N_8131);
nand U8260 (N_8260,N_8134,N_8015);
nor U8261 (N_8261,N_8081,N_8013);
and U8262 (N_8262,N_8157,N_8014);
nand U8263 (N_8263,N_8025,N_8021);
and U8264 (N_8264,N_8021,N_8153);
nor U8265 (N_8265,N_8039,N_8078);
and U8266 (N_8266,N_8098,N_8037);
or U8267 (N_8267,N_8070,N_8096);
nor U8268 (N_8268,N_8075,N_8102);
or U8269 (N_8269,N_8132,N_8113);
and U8270 (N_8270,N_8095,N_8070);
xor U8271 (N_8271,N_8118,N_8074);
nand U8272 (N_8272,N_8064,N_8117);
xor U8273 (N_8273,N_8102,N_8132);
xnor U8274 (N_8274,N_8132,N_8057);
or U8275 (N_8275,N_8124,N_8110);
nand U8276 (N_8276,N_8150,N_8079);
or U8277 (N_8277,N_8107,N_8011);
or U8278 (N_8278,N_8042,N_8043);
or U8279 (N_8279,N_8001,N_8147);
nor U8280 (N_8280,N_8022,N_8024);
nor U8281 (N_8281,N_8010,N_8109);
and U8282 (N_8282,N_8159,N_8096);
xnor U8283 (N_8283,N_8080,N_8058);
and U8284 (N_8284,N_8032,N_8106);
nand U8285 (N_8285,N_8030,N_8012);
nand U8286 (N_8286,N_8111,N_8099);
nor U8287 (N_8287,N_8035,N_8119);
or U8288 (N_8288,N_8070,N_8136);
or U8289 (N_8289,N_8135,N_8061);
nand U8290 (N_8290,N_8036,N_8033);
or U8291 (N_8291,N_8159,N_8156);
nand U8292 (N_8292,N_8075,N_8030);
nand U8293 (N_8293,N_8099,N_8042);
nand U8294 (N_8294,N_8032,N_8019);
xor U8295 (N_8295,N_8000,N_8012);
or U8296 (N_8296,N_8018,N_8095);
or U8297 (N_8297,N_8038,N_8007);
nand U8298 (N_8298,N_8015,N_8056);
or U8299 (N_8299,N_8001,N_8146);
nand U8300 (N_8300,N_8123,N_8000);
nand U8301 (N_8301,N_8010,N_8065);
xnor U8302 (N_8302,N_8004,N_8135);
nand U8303 (N_8303,N_8027,N_8105);
nor U8304 (N_8304,N_8150,N_8157);
nand U8305 (N_8305,N_8149,N_8033);
nand U8306 (N_8306,N_8133,N_8086);
or U8307 (N_8307,N_8106,N_8063);
nor U8308 (N_8308,N_8139,N_8049);
and U8309 (N_8309,N_8090,N_8069);
or U8310 (N_8310,N_8068,N_8091);
nand U8311 (N_8311,N_8045,N_8021);
and U8312 (N_8312,N_8147,N_8025);
nor U8313 (N_8313,N_8150,N_8004);
nand U8314 (N_8314,N_8144,N_8090);
xor U8315 (N_8315,N_8116,N_8048);
and U8316 (N_8316,N_8002,N_8021);
nor U8317 (N_8317,N_8071,N_8086);
nand U8318 (N_8318,N_8144,N_8009);
or U8319 (N_8319,N_8125,N_8073);
nor U8320 (N_8320,N_8305,N_8215);
nor U8321 (N_8321,N_8198,N_8219);
and U8322 (N_8322,N_8265,N_8210);
and U8323 (N_8323,N_8310,N_8277);
and U8324 (N_8324,N_8254,N_8271);
nor U8325 (N_8325,N_8186,N_8161);
xor U8326 (N_8326,N_8239,N_8270);
nor U8327 (N_8327,N_8164,N_8311);
or U8328 (N_8328,N_8222,N_8168);
or U8329 (N_8329,N_8249,N_8292);
and U8330 (N_8330,N_8175,N_8267);
or U8331 (N_8331,N_8173,N_8163);
nand U8332 (N_8332,N_8225,N_8279);
and U8333 (N_8333,N_8274,N_8275);
nor U8334 (N_8334,N_8171,N_8309);
and U8335 (N_8335,N_8195,N_8188);
nor U8336 (N_8336,N_8204,N_8230);
xnor U8337 (N_8337,N_8276,N_8289);
nand U8338 (N_8338,N_8260,N_8201);
and U8339 (N_8339,N_8281,N_8308);
xnor U8340 (N_8340,N_8194,N_8211);
or U8341 (N_8341,N_8316,N_8257);
or U8342 (N_8342,N_8264,N_8262);
or U8343 (N_8343,N_8307,N_8256);
and U8344 (N_8344,N_8301,N_8174);
or U8345 (N_8345,N_8273,N_8224);
and U8346 (N_8346,N_8206,N_8191);
xnor U8347 (N_8347,N_8282,N_8231);
and U8348 (N_8348,N_8285,N_8169);
nor U8349 (N_8349,N_8218,N_8312);
and U8350 (N_8350,N_8314,N_8172);
nand U8351 (N_8351,N_8183,N_8248);
nor U8352 (N_8352,N_8226,N_8303);
and U8353 (N_8353,N_8207,N_8243);
and U8354 (N_8354,N_8295,N_8250);
or U8355 (N_8355,N_8227,N_8296);
nor U8356 (N_8356,N_8166,N_8306);
or U8357 (N_8357,N_8240,N_8208);
nand U8358 (N_8358,N_8290,N_8237);
and U8359 (N_8359,N_8181,N_8293);
or U8360 (N_8360,N_8203,N_8199);
nor U8361 (N_8361,N_8228,N_8286);
or U8362 (N_8362,N_8288,N_8300);
nor U8363 (N_8363,N_8266,N_8229);
nand U8364 (N_8364,N_8192,N_8200);
xnor U8365 (N_8365,N_8178,N_8269);
or U8366 (N_8366,N_8261,N_8244);
nor U8367 (N_8367,N_8189,N_8165);
or U8368 (N_8368,N_8193,N_8298);
nor U8369 (N_8369,N_8268,N_8187);
nor U8370 (N_8370,N_8223,N_8180);
nor U8371 (N_8371,N_8213,N_8182);
nor U8372 (N_8372,N_8160,N_8212);
and U8373 (N_8373,N_8235,N_8232);
nor U8374 (N_8374,N_8247,N_8253);
nand U8375 (N_8375,N_8297,N_8241);
nand U8376 (N_8376,N_8242,N_8278);
xor U8377 (N_8377,N_8233,N_8238);
nand U8378 (N_8378,N_8287,N_8283);
and U8379 (N_8379,N_8234,N_8318);
xor U8380 (N_8380,N_8177,N_8299);
nor U8381 (N_8381,N_8162,N_8255);
nand U8382 (N_8382,N_8304,N_8184);
and U8383 (N_8383,N_8220,N_8317);
nand U8384 (N_8384,N_8245,N_8170);
nor U8385 (N_8385,N_8252,N_8179);
and U8386 (N_8386,N_8280,N_8319);
and U8387 (N_8387,N_8315,N_8216);
nand U8388 (N_8388,N_8259,N_8291);
or U8389 (N_8389,N_8251,N_8167);
nor U8390 (N_8390,N_8258,N_8209);
or U8391 (N_8391,N_8313,N_8176);
or U8392 (N_8392,N_8217,N_8272);
nor U8393 (N_8393,N_8196,N_8221);
nor U8394 (N_8394,N_8246,N_8197);
or U8395 (N_8395,N_8284,N_8302);
nor U8396 (N_8396,N_8294,N_8236);
and U8397 (N_8397,N_8202,N_8190);
nand U8398 (N_8398,N_8263,N_8185);
and U8399 (N_8399,N_8214,N_8205);
nor U8400 (N_8400,N_8229,N_8163);
nor U8401 (N_8401,N_8232,N_8176);
nor U8402 (N_8402,N_8188,N_8184);
and U8403 (N_8403,N_8308,N_8239);
or U8404 (N_8404,N_8228,N_8188);
nor U8405 (N_8405,N_8282,N_8185);
and U8406 (N_8406,N_8160,N_8243);
or U8407 (N_8407,N_8242,N_8291);
xnor U8408 (N_8408,N_8229,N_8178);
xor U8409 (N_8409,N_8187,N_8225);
or U8410 (N_8410,N_8254,N_8264);
and U8411 (N_8411,N_8203,N_8317);
or U8412 (N_8412,N_8199,N_8212);
nand U8413 (N_8413,N_8218,N_8228);
nor U8414 (N_8414,N_8270,N_8212);
nand U8415 (N_8415,N_8289,N_8232);
nand U8416 (N_8416,N_8251,N_8182);
xor U8417 (N_8417,N_8247,N_8223);
or U8418 (N_8418,N_8224,N_8282);
and U8419 (N_8419,N_8266,N_8290);
or U8420 (N_8420,N_8166,N_8192);
nand U8421 (N_8421,N_8300,N_8209);
xnor U8422 (N_8422,N_8209,N_8297);
nor U8423 (N_8423,N_8280,N_8295);
or U8424 (N_8424,N_8176,N_8160);
nand U8425 (N_8425,N_8204,N_8165);
or U8426 (N_8426,N_8295,N_8316);
nand U8427 (N_8427,N_8193,N_8251);
xor U8428 (N_8428,N_8190,N_8285);
or U8429 (N_8429,N_8250,N_8271);
or U8430 (N_8430,N_8180,N_8214);
nand U8431 (N_8431,N_8253,N_8189);
and U8432 (N_8432,N_8204,N_8305);
nor U8433 (N_8433,N_8203,N_8169);
nand U8434 (N_8434,N_8302,N_8225);
and U8435 (N_8435,N_8234,N_8172);
nand U8436 (N_8436,N_8207,N_8222);
or U8437 (N_8437,N_8180,N_8313);
and U8438 (N_8438,N_8172,N_8219);
or U8439 (N_8439,N_8282,N_8275);
nor U8440 (N_8440,N_8171,N_8298);
or U8441 (N_8441,N_8257,N_8290);
nor U8442 (N_8442,N_8230,N_8177);
or U8443 (N_8443,N_8304,N_8172);
and U8444 (N_8444,N_8240,N_8173);
and U8445 (N_8445,N_8203,N_8239);
or U8446 (N_8446,N_8175,N_8305);
or U8447 (N_8447,N_8167,N_8163);
nand U8448 (N_8448,N_8217,N_8210);
nor U8449 (N_8449,N_8259,N_8175);
and U8450 (N_8450,N_8297,N_8220);
nor U8451 (N_8451,N_8271,N_8302);
or U8452 (N_8452,N_8317,N_8276);
and U8453 (N_8453,N_8246,N_8269);
xnor U8454 (N_8454,N_8225,N_8315);
nand U8455 (N_8455,N_8304,N_8299);
and U8456 (N_8456,N_8310,N_8299);
and U8457 (N_8457,N_8232,N_8274);
nor U8458 (N_8458,N_8266,N_8276);
nand U8459 (N_8459,N_8161,N_8182);
nand U8460 (N_8460,N_8191,N_8293);
nor U8461 (N_8461,N_8212,N_8304);
nor U8462 (N_8462,N_8277,N_8249);
or U8463 (N_8463,N_8317,N_8263);
and U8464 (N_8464,N_8175,N_8219);
nand U8465 (N_8465,N_8179,N_8203);
xor U8466 (N_8466,N_8230,N_8254);
nor U8467 (N_8467,N_8164,N_8172);
or U8468 (N_8468,N_8312,N_8170);
nor U8469 (N_8469,N_8185,N_8179);
nand U8470 (N_8470,N_8172,N_8257);
and U8471 (N_8471,N_8195,N_8254);
nand U8472 (N_8472,N_8163,N_8280);
xor U8473 (N_8473,N_8304,N_8235);
nand U8474 (N_8474,N_8250,N_8313);
nor U8475 (N_8475,N_8179,N_8312);
nand U8476 (N_8476,N_8272,N_8278);
nand U8477 (N_8477,N_8224,N_8207);
xor U8478 (N_8478,N_8312,N_8160);
and U8479 (N_8479,N_8173,N_8185);
xnor U8480 (N_8480,N_8427,N_8409);
and U8481 (N_8481,N_8449,N_8343);
and U8482 (N_8482,N_8397,N_8447);
and U8483 (N_8483,N_8378,N_8358);
nand U8484 (N_8484,N_8444,N_8347);
nand U8485 (N_8485,N_8329,N_8448);
and U8486 (N_8486,N_8426,N_8432);
and U8487 (N_8487,N_8415,N_8402);
nand U8488 (N_8488,N_8405,N_8390);
or U8489 (N_8489,N_8332,N_8424);
nand U8490 (N_8490,N_8451,N_8422);
and U8491 (N_8491,N_8418,N_8323);
or U8492 (N_8492,N_8472,N_8387);
and U8493 (N_8493,N_8429,N_8337);
nor U8494 (N_8494,N_8367,N_8435);
or U8495 (N_8495,N_8398,N_8438);
or U8496 (N_8496,N_8340,N_8396);
xor U8497 (N_8497,N_8363,N_8375);
and U8498 (N_8498,N_8454,N_8441);
and U8499 (N_8499,N_8453,N_8471);
and U8500 (N_8500,N_8380,N_8379);
nand U8501 (N_8501,N_8476,N_8404);
and U8502 (N_8502,N_8394,N_8348);
or U8503 (N_8503,N_8342,N_8320);
nor U8504 (N_8504,N_8467,N_8452);
xor U8505 (N_8505,N_8383,N_8351);
nor U8506 (N_8506,N_8456,N_8412);
or U8507 (N_8507,N_8339,N_8437);
or U8508 (N_8508,N_8391,N_8420);
or U8509 (N_8509,N_8346,N_8366);
and U8510 (N_8510,N_8419,N_8345);
and U8511 (N_8511,N_8468,N_8330);
and U8512 (N_8512,N_8369,N_8399);
and U8513 (N_8513,N_8459,N_8475);
nor U8514 (N_8514,N_8395,N_8474);
or U8515 (N_8515,N_8374,N_8362);
nor U8516 (N_8516,N_8368,N_8393);
nand U8517 (N_8517,N_8473,N_8478);
nor U8518 (N_8518,N_8357,N_8389);
and U8519 (N_8519,N_8333,N_8352);
and U8520 (N_8520,N_8463,N_8469);
and U8521 (N_8521,N_8353,N_8407);
nor U8522 (N_8522,N_8450,N_8410);
nor U8523 (N_8523,N_8336,N_8324);
nand U8524 (N_8524,N_8477,N_8406);
nand U8525 (N_8525,N_8359,N_8385);
nor U8526 (N_8526,N_8338,N_8372);
nor U8527 (N_8527,N_8423,N_8440);
nand U8528 (N_8528,N_8465,N_8377);
and U8529 (N_8529,N_8382,N_8443);
nand U8530 (N_8530,N_8411,N_8461);
nand U8531 (N_8531,N_8325,N_8327);
or U8532 (N_8532,N_8376,N_8392);
xor U8533 (N_8533,N_8350,N_8355);
nor U8534 (N_8534,N_8360,N_8328);
nand U8535 (N_8535,N_8408,N_8349);
nand U8536 (N_8536,N_8425,N_8416);
nor U8537 (N_8537,N_8458,N_8434);
nand U8538 (N_8538,N_8365,N_8470);
or U8539 (N_8539,N_8431,N_8462);
nor U8540 (N_8540,N_8401,N_8455);
or U8541 (N_8541,N_8403,N_8439);
xor U8542 (N_8542,N_8457,N_8433);
or U8543 (N_8543,N_8373,N_8335);
or U8544 (N_8544,N_8428,N_8445);
nand U8545 (N_8545,N_8341,N_8446);
and U8546 (N_8546,N_8386,N_8354);
and U8547 (N_8547,N_8442,N_8381);
and U8548 (N_8548,N_8326,N_8414);
or U8549 (N_8549,N_8400,N_8356);
nor U8550 (N_8550,N_8460,N_8364);
nand U8551 (N_8551,N_8464,N_8321);
xor U8552 (N_8552,N_8466,N_8371);
nand U8553 (N_8553,N_8413,N_8361);
or U8554 (N_8554,N_8479,N_8436);
nor U8555 (N_8555,N_8384,N_8388);
nor U8556 (N_8556,N_8331,N_8344);
and U8557 (N_8557,N_8322,N_8370);
nand U8558 (N_8558,N_8421,N_8417);
nor U8559 (N_8559,N_8334,N_8430);
or U8560 (N_8560,N_8325,N_8462);
or U8561 (N_8561,N_8426,N_8352);
nand U8562 (N_8562,N_8439,N_8371);
nor U8563 (N_8563,N_8393,N_8349);
nor U8564 (N_8564,N_8339,N_8424);
nor U8565 (N_8565,N_8358,N_8374);
and U8566 (N_8566,N_8379,N_8397);
xor U8567 (N_8567,N_8341,N_8402);
and U8568 (N_8568,N_8383,N_8370);
and U8569 (N_8569,N_8457,N_8423);
and U8570 (N_8570,N_8331,N_8475);
or U8571 (N_8571,N_8386,N_8448);
and U8572 (N_8572,N_8367,N_8426);
nor U8573 (N_8573,N_8396,N_8323);
or U8574 (N_8574,N_8448,N_8344);
nor U8575 (N_8575,N_8371,N_8425);
nand U8576 (N_8576,N_8466,N_8435);
nor U8577 (N_8577,N_8405,N_8327);
nand U8578 (N_8578,N_8366,N_8423);
xnor U8579 (N_8579,N_8471,N_8368);
nand U8580 (N_8580,N_8330,N_8475);
nand U8581 (N_8581,N_8360,N_8416);
nand U8582 (N_8582,N_8415,N_8372);
nor U8583 (N_8583,N_8413,N_8381);
or U8584 (N_8584,N_8345,N_8399);
or U8585 (N_8585,N_8342,N_8341);
nor U8586 (N_8586,N_8364,N_8367);
and U8587 (N_8587,N_8474,N_8330);
xnor U8588 (N_8588,N_8419,N_8462);
nor U8589 (N_8589,N_8374,N_8462);
or U8590 (N_8590,N_8337,N_8389);
nor U8591 (N_8591,N_8396,N_8381);
nor U8592 (N_8592,N_8448,N_8471);
and U8593 (N_8593,N_8427,N_8328);
and U8594 (N_8594,N_8446,N_8425);
and U8595 (N_8595,N_8475,N_8382);
nor U8596 (N_8596,N_8462,N_8465);
nand U8597 (N_8597,N_8357,N_8326);
nor U8598 (N_8598,N_8469,N_8404);
nand U8599 (N_8599,N_8375,N_8340);
and U8600 (N_8600,N_8466,N_8394);
or U8601 (N_8601,N_8423,N_8479);
nor U8602 (N_8602,N_8436,N_8449);
and U8603 (N_8603,N_8348,N_8382);
nand U8604 (N_8604,N_8365,N_8475);
or U8605 (N_8605,N_8472,N_8389);
nand U8606 (N_8606,N_8355,N_8321);
or U8607 (N_8607,N_8436,N_8420);
and U8608 (N_8608,N_8442,N_8399);
and U8609 (N_8609,N_8378,N_8464);
or U8610 (N_8610,N_8475,N_8462);
or U8611 (N_8611,N_8339,N_8426);
nor U8612 (N_8612,N_8360,N_8468);
and U8613 (N_8613,N_8348,N_8347);
nand U8614 (N_8614,N_8381,N_8406);
xnor U8615 (N_8615,N_8469,N_8432);
and U8616 (N_8616,N_8479,N_8352);
nor U8617 (N_8617,N_8439,N_8325);
nor U8618 (N_8618,N_8472,N_8344);
and U8619 (N_8619,N_8454,N_8388);
xor U8620 (N_8620,N_8418,N_8422);
nand U8621 (N_8621,N_8320,N_8394);
nand U8622 (N_8622,N_8472,N_8393);
nand U8623 (N_8623,N_8412,N_8345);
and U8624 (N_8624,N_8347,N_8479);
xnor U8625 (N_8625,N_8348,N_8357);
nor U8626 (N_8626,N_8431,N_8399);
and U8627 (N_8627,N_8418,N_8378);
xnor U8628 (N_8628,N_8400,N_8447);
or U8629 (N_8629,N_8405,N_8464);
xnor U8630 (N_8630,N_8354,N_8321);
and U8631 (N_8631,N_8479,N_8458);
nand U8632 (N_8632,N_8405,N_8344);
or U8633 (N_8633,N_8386,N_8375);
nor U8634 (N_8634,N_8413,N_8421);
and U8635 (N_8635,N_8417,N_8390);
nand U8636 (N_8636,N_8383,N_8452);
xor U8637 (N_8637,N_8360,N_8437);
nand U8638 (N_8638,N_8448,N_8412);
nand U8639 (N_8639,N_8334,N_8444);
and U8640 (N_8640,N_8552,N_8511);
nand U8641 (N_8641,N_8608,N_8484);
and U8642 (N_8642,N_8522,N_8521);
or U8643 (N_8643,N_8622,N_8575);
nor U8644 (N_8644,N_8585,N_8542);
or U8645 (N_8645,N_8482,N_8518);
nand U8646 (N_8646,N_8561,N_8512);
or U8647 (N_8647,N_8577,N_8540);
nor U8648 (N_8648,N_8544,N_8567);
nand U8649 (N_8649,N_8556,N_8593);
xnor U8650 (N_8650,N_8509,N_8582);
nor U8651 (N_8651,N_8553,N_8523);
or U8652 (N_8652,N_8500,N_8508);
or U8653 (N_8653,N_8617,N_8545);
nor U8654 (N_8654,N_8625,N_8524);
and U8655 (N_8655,N_8519,N_8637);
and U8656 (N_8656,N_8487,N_8539);
nand U8657 (N_8657,N_8565,N_8491);
nor U8658 (N_8658,N_8590,N_8525);
and U8659 (N_8659,N_8573,N_8498);
or U8660 (N_8660,N_8580,N_8572);
nand U8661 (N_8661,N_8592,N_8559);
nor U8662 (N_8662,N_8507,N_8581);
nor U8663 (N_8663,N_8570,N_8636);
nor U8664 (N_8664,N_8605,N_8492);
and U8665 (N_8665,N_8584,N_8633);
nor U8666 (N_8666,N_8602,N_8639);
nand U8667 (N_8667,N_8614,N_8558);
and U8668 (N_8668,N_8535,N_8624);
xor U8669 (N_8669,N_8549,N_8569);
nand U8670 (N_8670,N_8538,N_8486);
or U8671 (N_8671,N_8503,N_8514);
nor U8672 (N_8672,N_8609,N_8555);
nand U8673 (N_8673,N_8611,N_8557);
nor U8674 (N_8674,N_8586,N_8488);
and U8675 (N_8675,N_8620,N_8490);
and U8676 (N_8676,N_8613,N_8517);
and U8677 (N_8677,N_8571,N_8623);
nor U8678 (N_8678,N_8630,N_8594);
nand U8679 (N_8679,N_8497,N_8496);
nor U8680 (N_8680,N_8516,N_8604);
nand U8681 (N_8681,N_8493,N_8495);
or U8682 (N_8682,N_8531,N_8610);
xor U8683 (N_8683,N_8510,N_8520);
or U8684 (N_8684,N_8505,N_8591);
nand U8685 (N_8685,N_8528,N_8483);
and U8686 (N_8686,N_8627,N_8504);
or U8687 (N_8687,N_8621,N_8631);
and U8688 (N_8688,N_8626,N_8527);
and U8689 (N_8689,N_8615,N_8501);
and U8690 (N_8690,N_8506,N_8638);
nor U8691 (N_8691,N_8574,N_8601);
and U8692 (N_8692,N_8628,N_8485);
and U8693 (N_8693,N_8536,N_8600);
and U8694 (N_8694,N_8560,N_8513);
nor U8695 (N_8695,N_8499,N_8629);
or U8696 (N_8696,N_8599,N_8634);
or U8697 (N_8697,N_8480,N_8533);
nand U8698 (N_8698,N_8568,N_8619);
nand U8699 (N_8699,N_8537,N_8566);
nand U8700 (N_8700,N_8616,N_8534);
and U8701 (N_8701,N_8550,N_8578);
nand U8702 (N_8702,N_8564,N_8632);
and U8703 (N_8703,N_8583,N_8529);
nor U8704 (N_8704,N_8532,N_8579);
nand U8705 (N_8705,N_8588,N_8589);
or U8706 (N_8706,N_8494,N_8576);
xor U8707 (N_8707,N_8612,N_8595);
and U8708 (N_8708,N_8563,N_8526);
nor U8709 (N_8709,N_8515,N_8481);
and U8710 (N_8710,N_8598,N_8562);
nand U8711 (N_8711,N_8554,N_8603);
and U8712 (N_8712,N_8543,N_8606);
xor U8713 (N_8713,N_8489,N_8597);
nor U8714 (N_8714,N_8551,N_8618);
nor U8715 (N_8715,N_8547,N_8596);
and U8716 (N_8716,N_8607,N_8541);
nand U8717 (N_8717,N_8635,N_8546);
nand U8718 (N_8718,N_8587,N_8548);
or U8719 (N_8719,N_8502,N_8530);
nand U8720 (N_8720,N_8563,N_8585);
nor U8721 (N_8721,N_8553,N_8615);
or U8722 (N_8722,N_8513,N_8547);
nand U8723 (N_8723,N_8639,N_8517);
nor U8724 (N_8724,N_8545,N_8619);
nand U8725 (N_8725,N_8584,N_8636);
nor U8726 (N_8726,N_8629,N_8530);
or U8727 (N_8727,N_8575,N_8485);
xnor U8728 (N_8728,N_8608,N_8529);
nor U8729 (N_8729,N_8481,N_8615);
nor U8730 (N_8730,N_8546,N_8525);
xor U8731 (N_8731,N_8571,N_8609);
nor U8732 (N_8732,N_8590,N_8615);
nand U8733 (N_8733,N_8573,N_8541);
nand U8734 (N_8734,N_8539,N_8556);
nor U8735 (N_8735,N_8514,N_8500);
xor U8736 (N_8736,N_8552,N_8622);
or U8737 (N_8737,N_8599,N_8526);
nand U8738 (N_8738,N_8496,N_8543);
xor U8739 (N_8739,N_8494,N_8579);
nor U8740 (N_8740,N_8623,N_8607);
and U8741 (N_8741,N_8628,N_8538);
xnor U8742 (N_8742,N_8502,N_8595);
nor U8743 (N_8743,N_8612,N_8634);
or U8744 (N_8744,N_8517,N_8516);
and U8745 (N_8745,N_8629,N_8520);
and U8746 (N_8746,N_8518,N_8600);
nor U8747 (N_8747,N_8518,N_8596);
nand U8748 (N_8748,N_8593,N_8484);
nor U8749 (N_8749,N_8579,N_8600);
nand U8750 (N_8750,N_8574,N_8627);
nand U8751 (N_8751,N_8496,N_8585);
and U8752 (N_8752,N_8637,N_8552);
nand U8753 (N_8753,N_8565,N_8525);
nor U8754 (N_8754,N_8617,N_8530);
and U8755 (N_8755,N_8541,N_8564);
nand U8756 (N_8756,N_8509,N_8615);
xnor U8757 (N_8757,N_8614,N_8555);
nor U8758 (N_8758,N_8526,N_8535);
and U8759 (N_8759,N_8616,N_8598);
nor U8760 (N_8760,N_8533,N_8628);
nor U8761 (N_8761,N_8490,N_8524);
nand U8762 (N_8762,N_8513,N_8523);
and U8763 (N_8763,N_8571,N_8489);
and U8764 (N_8764,N_8596,N_8623);
or U8765 (N_8765,N_8584,N_8533);
nand U8766 (N_8766,N_8551,N_8578);
nor U8767 (N_8767,N_8598,N_8573);
and U8768 (N_8768,N_8597,N_8565);
nor U8769 (N_8769,N_8540,N_8529);
nor U8770 (N_8770,N_8576,N_8575);
or U8771 (N_8771,N_8571,N_8552);
xnor U8772 (N_8772,N_8571,N_8590);
and U8773 (N_8773,N_8596,N_8520);
nor U8774 (N_8774,N_8555,N_8528);
nand U8775 (N_8775,N_8480,N_8482);
or U8776 (N_8776,N_8615,N_8505);
nor U8777 (N_8777,N_8545,N_8561);
or U8778 (N_8778,N_8548,N_8530);
or U8779 (N_8779,N_8508,N_8629);
or U8780 (N_8780,N_8508,N_8546);
or U8781 (N_8781,N_8489,N_8613);
nor U8782 (N_8782,N_8586,N_8582);
nand U8783 (N_8783,N_8580,N_8615);
and U8784 (N_8784,N_8549,N_8614);
or U8785 (N_8785,N_8596,N_8606);
nand U8786 (N_8786,N_8612,N_8578);
or U8787 (N_8787,N_8584,N_8523);
and U8788 (N_8788,N_8591,N_8589);
nand U8789 (N_8789,N_8619,N_8531);
nor U8790 (N_8790,N_8555,N_8529);
nor U8791 (N_8791,N_8505,N_8552);
nand U8792 (N_8792,N_8571,N_8542);
nor U8793 (N_8793,N_8559,N_8576);
nor U8794 (N_8794,N_8487,N_8527);
or U8795 (N_8795,N_8606,N_8633);
xor U8796 (N_8796,N_8520,N_8514);
nand U8797 (N_8797,N_8619,N_8591);
nand U8798 (N_8798,N_8488,N_8611);
or U8799 (N_8799,N_8512,N_8534);
or U8800 (N_8800,N_8661,N_8749);
and U8801 (N_8801,N_8667,N_8717);
or U8802 (N_8802,N_8736,N_8723);
nand U8803 (N_8803,N_8788,N_8684);
or U8804 (N_8804,N_8644,N_8779);
xnor U8805 (N_8805,N_8765,N_8718);
xor U8806 (N_8806,N_8663,N_8735);
nor U8807 (N_8807,N_8796,N_8641);
nand U8808 (N_8808,N_8792,N_8654);
or U8809 (N_8809,N_8782,N_8769);
nand U8810 (N_8810,N_8737,N_8797);
nand U8811 (N_8811,N_8694,N_8703);
xor U8812 (N_8812,N_8730,N_8659);
nand U8813 (N_8813,N_8653,N_8768);
nand U8814 (N_8814,N_8655,N_8734);
or U8815 (N_8815,N_8773,N_8724);
or U8816 (N_8816,N_8760,N_8695);
or U8817 (N_8817,N_8698,N_8753);
or U8818 (N_8818,N_8795,N_8728);
nor U8819 (N_8819,N_8759,N_8692);
nand U8820 (N_8820,N_8721,N_8658);
or U8821 (N_8821,N_8770,N_8767);
nor U8822 (N_8822,N_8673,N_8651);
nor U8823 (N_8823,N_8758,N_8713);
or U8824 (N_8824,N_8714,N_8707);
nand U8825 (N_8825,N_8645,N_8742);
nand U8826 (N_8826,N_8669,N_8799);
xor U8827 (N_8827,N_8772,N_8647);
and U8828 (N_8828,N_8670,N_8783);
and U8829 (N_8829,N_8652,N_8640);
nor U8830 (N_8830,N_8764,N_8756);
nor U8831 (N_8831,N_8766,N_8757);
nand U8832 (N_8832,N_8738,N_8745);
nor U8833 (N_8833,N_8711,N_8729);
nand U8834 (N_8834,N_8789,N_8657);
nand U8835 (N_8835,N_8776,N_8660);
nand U8836 (N_8836,N_8708,N_8679);
or U8837 (N_8837,N_8682,N_8666);
or U8838 (N_8838,N_8676,N_8699);
and U8839 (N_8839,N_8650,N_8747);
or U8840 (N_8840,N_8681,N_8671);
nor U8841 (N_8841,N_8675,N_8793);
and U8842 (N_8842,N_8643,N_8668);
xnor U8843 (N_8843,N_8755,N_8775);
or U8844 (N_8844,N_8709,N_8794);
nor U8845 (N_8845,N_8710,N_8683);
nand U8846 (N_8846,N_8686,N_8697);
nor U8847 (N_8847,N_8751,N_8720);
or U8848 (N_8848,N_8726,N_8689);
nand U8849 (N_8849,N_8690,N_8781);
nor U8850 (N_8850,N_8740,N_8731);
and U8851 (N_8851,N_8688,N_8732);
or U8852 (N_8852,N_8787,N_8678);
nand U8853 (N_8853,N_8648,N_8763);
nor U8854 (N_8854,N_8680,N_8716);
and U8855 (N_8855,N_8696,N_8733);
nor U8856 (N_8856,N_8687,N_8741);
nor U8857 (N_8857,N_8691,N_8771);
nand U8858 (N_8858,N_8674,N_8791);
and U8859 (N_8859,N_8778,N_8784);
or U8860 (N_8860,N_8704,N_8748);
or U8861 (N_8861,N_8642,N_8656);
and U8862 (N_8862,N_8780,N_8762);
xor U8863 (N_8863,N_8701,N_8725);
nor U8864 (N_8864,N_8727,N_8744);
nor U8865 (N_8865,N_8646,N_8649);
nand U8866 (N_8866,N_8677,N_8662);
and U8867 (N_8867,N_8665,N_8706);
nor U8868 (N_8868,N_8743,N_8750);
or U8869 (N_8869,N_8722,N_8746);
xor U8870 (N_8870,N_8786,N_8785);
and U8871 (N_8871,N_8719,N_8739);
and U8872 (N_8872,N_8702,N_8777);
or U8873 (N_8873,N_8705,N_8774);
or U8874 (N_8874,N_8715,N_8754);
and U8875 (N_8875,N_8790,N_8693);
nand U8876 (N_8876,N_8752,N_8700);
nor U8877 (N_8877,N_8685,N_8664);
nor U8878 (N_8878,N_8761,N_8798);
or U8879 (N_8879,N_8712,N_8672);
nor U8880 (N_8880,N_8751,N_8773);
nor U8881 (N_8881,N_8787,N_8745);
nor U8882 (N_8882,N_8721,N_8759);
and U8883 (N_8883,N_8771,N_8645);
and U8884 (N_8884,N_8643,N_8663);
nand U8885 (N_8885,N_8643,N_8777);
nand U8886 (N_8886,N_8776,N_8761);
nand U8887 (N_8887,N_8687,N_8755);
and U8888 (N_8888,N_8740,N_8734);
xor U8889 (N_8889,N_8797,N_8651);
xnor U8890 (N_8890,N_8697,N_8753);
xor U8891 (N_8891,N_8676,N_8702);
nor U8892 (N_8892,N_8710,N_8665);
or U8893 (N_8893,N_8691,N_8670);
or U8894 (N_8894,N_8794,N_8740);
nor U8895 (N_8895,N_8649,N_8683);
nand U8896 (N_8896,N_8669,N_8743);
and U8897 (N_8897,N_8654,N_8714);
and U8898 (N_8898,N_8739,N_8706);
nor U8899 (N_8899,N_8753,N_8699);
nand U8900 (N_8900,N_8773,N_8681);
or U8901 (N_8901,N_8707,N_8678);
or U8902 (N_8902,N_8704,N_8657);
or U8903 (N_8903,N_8732,N_8687);
or U8904 (N_8904,N_8643,N_8722);
or U8905 (N_8905,N_8656,N_8663);
nor U8906 (N_8906,N_8724,N_8732);
nand U8907 (N_8907,N_8683,N_8753);
or U8908 (N_8908,N_8697,N_8701);
nand U8909 (N_8909,N_8796,N_8742);
or U8910 (N_8910,N_8786,N_8705);
nor U8911 (N_8911,N_8687,N_8652);
nand U8912 (N_8912,N_8710,N_8792);
or U8913 (N_8913,N_8646,N_8708);
and U8914 (N_8914,N_8763,N_8790);
nand U8915 (N_8915,N_8692,N_8765);
and U8916 (N_8916,N_8719,N_8762);
nor U8917 (N_8917,N_8797,N_8733);
nand U8918 (N_8918,N_8743,N_8667);
nor U8919 (N_8919,N_8761,N_8760);
or U8920 (N_8920,N_8772,N_8709);
nor U8921 (N_8921,N_8746,N_8665);
nand U8922 (N_8922,N_8700,N_8720);
nor U8923 (N_8923,N_8795,N_8771);
xor U8924 (N_8924,N_8651,N_8794);
nor U8925 (N_8925,N_8664,N_8778);
and U8926 (N_8926,N_8679,N_8760);
or U8927 (N_8927,N_8654,N_8790);
and U8928 (N_8928,N_8797,N_8700);
nor U8929 (N_8929,N_8756,N_8799);
and U8930 (N_8930,N_8759,N_8670);
nand U8931 (N_8931,N_8764,N_8681);
and U8932 (N_8932,N_8721,N_8747);
nand U8933 (N_8933,N_8699,N_8780);
nor U8934 (N_8934,N_8724,N_8717);
or U8935 (N_8935,N_8682,N_8704);
nor U8936 (N_8936,N_8791,N_8763);
and U8937 (N_8937,N_8705,N_8732);
or U8938 (N_8938,N_8726,N_8699);
and U8939 (N_8939,N_8698,N_8701);
and U8940 (N_8940,N_8694,N_8780);
and U8941 (N_8941,N_8683,N_8746);
nor U8942 (N_8942,N_8709,N_8665);
or U8943 (N_8943,N_8642,N_8787);
or U8944 (N_8944,N_8706,N_8640);
nand U8945 (N_8945,N_8763,N_8750);
or U8946 (N_8946,N_8727,N_8774);
xor U8947 (N_8947,N_8680,N_8738);
and U8948 (N_8948,N_8706,N_8719);
and U8949 (N_8949,N_8691,N_8721);
or U8950 (N_8950,N_8722,N_8726);
xor U8951 (N_8951,N_8686,N_8728);
nand U8952 (N_8952,N_8709,N_8731);
or U8953 (N_8953,N_8673,N_8703);
nand U8954 (N_8954,N_8743,N_8737);
nor U8955 (N_8955,N_8797,N_8665);
xor U8956 (N_8956,N_8733,N_8767);
or U8957 (N_8957,N_8721,N_8729);
or U8958 (N_8958,N_8758,N_8716);
xnor U8959 (N_8959,N_8641,N_8754);
and U8960 (N_8960,N_8847,N_8879);
nand U8961 (N_8961,N_8895,N_8841);
or U8962 (N_8962,N_8903,N_8829);
xor U8963 (N_8963,N_8830,N_8935);
nor U8964 (N_8964,N_8859,N_8881);
nor U8965 (N_8965,N_8912,N_8875);
nand U8966 (N_8966,N_8942,N_8833);
or U8967 (N_8967,N_8852,N_8925);
nand U8968 (N_8968,N_8948,N_8801);
nor U8969 (N_8969,N_8863,N_8826);
or U8970 (N_8970,N_8886,N_8933);
nor U8971 (N_8971,N_8921,N_8958);
and U8972 (N_8972,N_8943,N_8802);
xnor U8973 (N_8973,N_8810,N_8837);
and U8974 (N_8974,N_8865,N_8893);
nor U8975 (N_8975,N_8919,N_8855);
nor U8976 (N_8976,N_8930,N_8892);
xor U8977 (N_8977,N_8824,N_8896);
xnor U8978 (N_8978,N_8955,N_8805);
nand U8979 (N_8979,N_8809,N_8932);
xor U8980 (N_8980,N_8815,N_8936);
nor U8981 (N_8981,N_8928,N_8838);
xor U8982 (N_8982,N_8885,N_8938);
nand U8983 (N_8983,N_8915,N_8894);
and U8984 (N_8984,N_8853,N_8945);
nand U8985 (N_8985,N_8939,N_8911);
xor U8986 (N_8986,N_8880,N_8856);
or U8987 (N_8987,N_8828,N_8831);
nor U8988 (N_8988,N_8946,N_8926);
and U8989 (N_8989,N_8832,N_8884);
and U8990 (N_8990,N_8891,N_8887);
xnor U8991 (N_8991,N_8848,N_8819);
nor U8992 (N_8992,N_8934,N_8952);
xor U8993 (N_8993,N_8870,N_8806);
nor U8994 (N_8994,N_8873,N_8814);
and U8995 (N_8995,N_8866,N_8821);
nor U8996 (N_8996,N_8851,N_8920);
nor U8997 (N_8997,N_8864,N_8844);
nand U8998 (N_8998,N_8947,N_8840);
or U8999 (N_8999,N_8900,N_8825);
nor U9000 (N_9000,N_8929,N_8905);
nand U9001 (N_9001,N_8843,N_8868);
or U9002 (N_9002,N_8908,N_8872);
or U9003 (N_9003,N_8874,N_8924);
or U9004 (N_9004,N_8951,N_8835);
or U9005 (N_9005,N_8803,N_8842);
and U9006 (N_9006,N_8850,N_8807);
or U9007 (N_9007,N_8904,N_8822);
nand U9008 (N_9008,N_8922,N_8957);
and U9009 (N_9009,N_8914,N_8818);
and U9010 (N_9010,N_8916,N_8949);
nor U9011 (N_9011,N_8836,N_8858);
or U9012 (N_9012,N_8871,N_8906);
or U9013 (N_9013,N_8901,N_8827);
and U9014 (N_9014,N_8869,N_8804);
nand U9015 (N_9015,N_8909,N_8839);
and U9016 (N_9016,N_8917,N_8950);
xnor U9017 (N_9017,N_8846,N_8878);
or U9018 (N_9018,N_8862,N_8898);
and U9019 (N_9019,N_8854,N_8834);
nor U9020 (N_9020,N_8899,N_8913);
nand U9021 (N_9021,N_8857,N_8867);
nand U9022 (N_9022,N_8897,N_8845);
nor U9023 (N_9023,N_8937,N_8817);
or U9024 (N_9024,N_8800,N_8927);
and U9025 (N_9025,N_8883,N_8941);
nand U9026 (N_9026,N_8877,N_8944);
and U9027 (N_9027,N_8918,N_8931);
xnor U9028 (N_9028,N_8956,N_8820);
xor U9029 (N_9029,N_8816,N_8940);
nand U9030 (N_9030,N_8811,N_8888);
xnor U9031 (N_9031,N_8849,N_8902);
or U9032 (N_9032,N_8959,N_8808);
nor U9033 (N_9033,N_8910,N_8907);
nand U9034 (N_9034,N_8923,N_8882);
and U9035 (N_9035,N_8813,N_8823);
xor U9036 (N_9036,N_8954,N_8889);
nand U9037 (N_9037,N_8876,N_8953);
nor U9038 (N_9038,N_8860,N_8890);
nor U9039 (N_9039,N_8812,N_8861);
or U9040 (N_9040,N_8891,N_8829);
xor U9041 (N_9041,N_8903,N_8959);
and U9042 (N_9042,N_8866,N_8883);
nand U9043 (N_9043,N_8867,N_8898);
and U9044 (N_9044,N_8818,N_8820);
nor U9045 (N_9045,N_8959,N_8911);
xnor U9046 (N_9046,N_8826,N_8843);
nor U9047 (N_9047,N_8838,N_8890);
and U9048 (N_9048,N_8926,N_8899);
and U9049 (N_9049,N_8910,N_8809);
nor U9050 (N_9050,N_8908,N_8864);
nor U9051 (N_9051,N_8866,N_8805);
xnor U9052 (N_9052,N_8926,N_8882);
xor U9053 (N_9053,N_8953,N_8891);
and U9054 (N_9054,N_8845,N_8886);
and U9055 (N_9055,N_8892,N_8940);
or U9056 (N_9056,N_8953,N_8861);
nand U9057 (N_9057,N_8917,N_8875);
xnor U9058 (N_9058,N_8849,N_8907);
or U9059 (N_9059,N_8866,N_8913);
or U9060 (N_9060,N_8867,N_8833);
nor U9061 (N_9061,N_8843,N_8958);
or U9062 (N_9062,N_8805,N_8938);
and U9063 (N_9063,N_8882,N_8847);
nor U9064 (N_9064,N_8876,N_8884);
nand U9065 (N_9065,N_8914,N_8956);
xnor U9066 (N_9066,N_8853,N_8897);
and U9067 (N_9067,N_8950,N_8842);
or U9068 (N_9068,N_8812,N_8954);
xnor U9069 (N_9069,N_8933,N_8874);
and U9070 (N_9070,N_8907,N_8913);
or U9071 (N_9071,N_8931,N_8953);
nor U9072 (N_9072,N_8880,N_8838);
xor U9073 (N_9073,N_8854,N_8841);
or U9074 (N_9074,N_8817,N_8883);
nor U9075 (N_9075,N_8859,N_8889);
and U9076 (N_9076,N_8868,N_8833);
nand U9077 (N_9077,N_8943,N_8933);
or U9078 (N_9078,N_8870,N_8959);
and U9079 (N_9079,N_8868,N_8864);
nor U9080 (N_9080,N_8818,N_8885);
nor U9081 (N_9081,N_8872,N_8902);
nand U9082 (N_9082,N_8801,N_8917);
nand U9083 (N_9083,N_8810,N_8927);
or U9084 (N_9084,N_8954,N_8820);
and U9085 (N_9085,N_8866,N_8860);
nand U9086 (N_9086,N_8839,N_8827);
and U9087 (N_9087,N_8853,N_8935);
nand U9088 (N_9088,N_8929,N_8808);
or U9089 (N_9089,N_8930,N_8854);
and U9090 (N_9090,N_8864,N_8804);
nor U9091 (N_9091,N_8909,N_8936);
and U9092 (N_9092,N_8881,N_8899);
or U9093 (N_9093,N_8906,N_8920);
nor U9094 (N_9094,N_8896,N_8930);
and U9095 (N_9095,N_8946,N_8823);
nor U9096 (N_9096,N_8908,N_8951);
or U9097 (N_9097,N_8833,N_8821);
nand U9098 (N_9098,N_8854,N_8954);
or U9099 (N_9099,N_8883,N_8902);
nor U9100 (N_9100,N_8850,N_8924);
or U9101 (N_9101,N_8864,N_8914);
or U9102 (N_9102,N_8949,N_8860);
and U9103 (N_9103,N_8910,N_8814);
nand U9104 (N_9104,N_8902,N_8903);
or U9105 (N_9105,N_8811,N_8837);
and U9106 (N_9106,N_8946,N_8853);
or U9107 (N_9107,N_8959,N_8861);
and U9108 (N_9108,N_8926,N_8828);
nand U9109 (N_9109,N_8935,N_8820);
and U9110 (N_9110,N_8942,N_8838);
nor U9111 (N_9111,N_8835,N_8811);
or U9112 (N_9112,N_8911,N_8805);
nand U9113 (N_9113,N_8934,N_8916);
xor U9114 (N_9114,N_8891,N_8951);
and U9115 (N_9115,N_8959,N_8839);
or U9116 (N_9116,N_8822,N_8835);
and U9117 (N_9117,N_8917,N_8956);
nor U9118 (N_9118,N_8869,N_8830);
nor U9119 (N_9119,N_8863,N_8862);
nor U9120 (N_9120,N_8999,N_8963);
and U9121 (N_9121,N_9106,N_9068);
nor U9122 (N_9122,N_9094,N_8985);
nand U9123 (N_9123,N_9007,N_9118);
or U9124 (N_9124,N_8979,N_9032);
or U9125 (N_9125,N_9115,N_9024);
nand U9126 (N_9126,N_9053,N_9117);
and U9127 (N_9127,N_9021,N_9082);
nor U9128 (N_9128,N_9100,N_9033);
nor U9129 (N_9129,N_9116,N_9010);
nor U9130 (N_9130,N_9066,N_9113);
and U9131 (N_9131,N_9097,N_9070);
and U9132 (N_9132,N_9088,N_8996);
and U9133 (N_9133,N_9006,N_8973);
and U9134 (N_9134,N_8965,N_9040);
nor U9135 (N_9135,N_9076,N_9098);
nor U9136 (N_9136,N_9063,N_9083);
nor U9137 (N_9137,N_9016,N_9062);
nand U9138 (N_9138,N_9000,N_9004);
and U9139 (N_9139,N_8972,N_8988);
xnor U9140 (N_9140,N_9071,N_9031);
or U9141 (N_9141,N_9012,N_8993);
nand U9142 (N_9142,N_8960,N_9046);
and U9143 (N_9143,N_8971,N_9038);
nor U9144 (N_9144,N_9103,N_9056);
and U9145 (N_9145,N_9091,N_9022);
nor U9146 (N_9146,N_9084,N_8968);
and U9147 (N_9147,N_9002,N_9060);
nand U9148 (N_9148,N_9049,N_8970);
and U9149 (N_9149,N_9018,N_9042);
nor U9150 (N_9150,N_9073,N_8981);
xor U9151 (N_9151,N_9008,N_9023);
or U9152 (N_9152,N_9110,N_8978);
nand U9153 (N_9153,N_9048,N_8984);
or U9154 (N_9154,N_9111,N_8962);
and U9155 (N_9155,N_9041,N_9037);
nor U9156 (N_9156,N_9061,N_8964);
xnor U9157 (N_9157,N_8966,N_8980);
nor U9158 (N_9158,N_9054,N_9028);
nor U9159 (N_9159,N_8995,N_9064);
nand U9160 (N_9160,N_9090,N_9104);
and U9161 (N_9161,N_9001,N_9086);
nor U9162 (N_9162,N_9027,N_8998);
and U9163 (N_9163,N_9089,N_8987);
nand U9164 (N_9164,N_9107,N_9109);
nand U9165 (N_9165,N_9085,N_9087);
nor U9166 (N_9166,N_9003,N_9075);
or U9167 (N_9167,N_9036,N_9072);
nand U9168 (N_9168,N_9051,N_9029);
nor U9169 (N_9169,N_9030,N_9093);
nor U9170 (N_9170,N_9065,N_9047);
and U9171 (N_9171,N_8967,N_8961);
or U9172 (N_9172,N_8994,N_8977);
and U9173 (N_9173,N_9050,N_8990);
or U9174 (N_9174,N_9039,N_9005);
and U9175 (N_9175,N_9034,N_9044);
nor U9176 (N_9176,N_8969,N_9052);
nand U9177 (N_9177,N_9078,N_9017);
nand U9178 (N_9178,N_9092,N_9080);
and U9179 (N_9179,N_9020,N_9058);
nor U9180 (N_9180,N_8974,N_8975);
and U9181 (N_9181,N_8989,N_8991);
and U9182 (N_9182,N_9077,N_9067);
or U9183 (N_9183,N_8992,N_9043);
nand U9184 (N_9184,N_9081,N_9069);
and U9185 (N_9185,N_9079,N_8983);
or U9186 (N_9186,N_9045,N_9112);
xor U9187 (N_9187,N_9096,N_9095);
xnor U9188 (N_9188,N_9114,N_9102);
or U9189 (N_9189,N_8982,N_9119);
or U9190 (N_9190,N_9013,N_9059);
or U9191 (N_9191,N_9074,N_9014);
nor U9192 (N_9192,N_9057,N_9055);
nor U9193 (N_9193,N_9101,N_8997);
nand U9194 (N_9194,N_9011,N_8976);
nor U9195 (N_9195,N_9035,N_9015);
and U9196 (N_9196,N_9108,N_9099);
or U9197 (N_9197,N_9009,N_8986);
or U9198 (N_9198,N_9019,N_9025);
nor U9199 (N_9199,N_9105,N_9026);
xnor U9200 (N_9200,N_8990,N_9048);
and U9201 (N_9201,N_9029,N_9010);
or U9202 (N_9202,N_9032,N_9081);
or U9203 (N_9203,N_8986,N_9113);
and U9204 (N_9204,N_9047,N_9029);
xnor U9205 (N_9205,N_8989,N_9043);
nand U9206 (N_9206,N_8970,N_9050);
and U9207 (N_9207,N_9079,N_9114);
and U9208 (N_9208,N_9076,N_8989);
or U9209 (N_9209,N_9110,N_9048);
nor U9210 (N_9210,N_8985,N_9073);
or U9211 (N_9211,N_8964,N_9045);
or U9212 (N_9212,N_9008,N_8986);
nand U9213 (N_9213,N_8983,N_9070);
xor U9214 (N_9214,N_9013,N_9081);
or U9215 (N_9215,N_9070,N_9101);
nor U9216 (N_9216,N_8994,N_9016);
nor U9217 (N_9217,N_9059,N_8985);
nor U9218 (N_9218,N_9081,N_9108);
or U9219 (N_9219,N_9107,N_9030);
or U9220 (N_9220,N_8983,N_8968);
nand U9221 (N_9221,N_9017,N_9033);
nand U9222 (N_9222,N_8969,N_9076);
and U9223 (N_9223,N_8974,N_9007);
and U9224 (N_9224,N_9005,N_9085);
nor U9225 (N_9225,N_9022,N_9110);
and U9226 (N_9226,N_9080,N_9033);
nand U9227 (N_9227,N_9068,N_9075);
nand U9228 (N_9228,N_8982,N_9025);
and U9229 (N_9229,N_9082,N_9006);
xor U9230 (N_9230,N_8993,N_9018);
or U9231 (N_9231,N_9084,N_8997);
nand U9232 (N_9232,N_9061,N_8978);
nor U9233 (N_9233,N_9099,N_9113);
nand U9234 (N_9234,N_9099,N_9013);
xnor U9235 (N_9235,N_8994,N_8986);
xor U9236 (N_9236,N_9054,N_9118);
or U9237 (N_9237,N_9014,N_9025);
or U9238 (N_9238,N_8961,N_9068);
nand U9239 (N_9239,N_8979,N_9069);
nand U9240 (N_9240,N_8984,N_8967);
nor U9241 (N_9241,N_9013,N_9012);
nor U9242 (N_9242,N_9113,N_9053);
or U9243 (N_9243,N_8981,N_9084);
xor U9244 (N_9244,N_9116,N_8961);
or U9245 (N_9245,N_9101,N_9089);
nand U9246 (N_9246,N_8988,N_9013);
nand U9247 (N_9247,N_9115,N_9015);
nand U9248 (N_9248,N_8966,N_9102);
nor U9249 (N_9249,N_9080,N_9094);
nor U9250 (N_9250,N_9042,N_9075);
and U9251 (N_9251,N_9052,N_9026);
xor U9252 (N_9252,N_9024,N_9056);
nor U9253 (N_9253,N_9034,N_9042);
or U9254 (N_9254,N_9116,N_9013);
and U9255 (N_9255,N_8981,N_9032);
and U9256 (N_9256,N_8974,N_8965);
or U9257 (N_9257,N_8967,N_9029);
nor U9258 (N_9258,N_9091,N_8985);
nand U9259 (N_9259,N_9037,N_8991);
or U9260 (N_9260,N_8967,N_8962);
nand U9261 (N_9261,N_9050,N_8983);
nor U9262 (N_9262,N_8994,N_9000);
nand U9263 (N_9263,N_8978,N_8976);
nor U9264 (N_9264,N_9025,N_9093);
nand U9265 (N_9265,N_8977,N_9063);
or U9266 (N_9266,N_9058,N_8984);
and U9267 (N_9267,N_9078,N_9097);
and U9268 (N_9268,N_8967,N_9085);
nand U9269 (N_9269,N_9031,N_9088);
and U9270 (N_9270,N_9069,N_9034);
and U9271 (N_9271,N_8979,N_9100);
or U9272 (N_9272,N_9020,N_9112);
or U9273 (N_9273,N_9109,N_8970);
xor U9274 (N_9274,N_9048,N_8968);
nand U9275 (N_9275,N_9004,N_8998);
nand U9276 (N_9276,N_9048,N_9058);
or U9277 (N_9277,N_8986,N_9017);
nand U9278 (N_9278,N_9058,N_8979);
or U9279 (N_9279,N_9069,N_9038);
nand U9280 (N_9280,N_9131,N_9272);
or U9281 (N_9281,N_9278,N_9183);
xnor U9282 (N_9282,N_9144,N_9201);
nor U9283 (N_9283,N_9271,N_9134);
xor U9284 (N_9284,N_9178,N_9163);
and U9285 (N_9285,N_9152,N_9268);
nor U9286 (N_9286,N_9254,N_9232);
or U9287 (N_9287,N_9138,N_9259);
and U9288 (N_9288,N_9251,N_9182);
nand U9289 (N_9289,N_9124,N_9279);
or U9290 (N_9290,N_9154,N_9216);
or U9291 (N_9291,N_9175,N_9276);
or U9292 (N_9292,N_9247,N_9225);
nand U9293 (N_9293,N_9205,N_9160);
nor U9294 (N_9294,N_9132,N_9274);
nand U9295 (N_9295,N_9165,N_9212);
or U9296 (N_9296,N_9253,N_9136);
and U9297 (N_9297,N_9185,N_9224);
and U9298 (N_9298,N_9215,N_9244);
xnor U9299 (N_9299,N_9265,N_9248);
and U9300 (N_9300,N_9213,N_9208);
or U9301 (N_9301,N_9203,N_9191);
xor U9302 (N_9302,N_9167,N_9220);
xor U9303 (N_9303,N_9209,N_9153);
or U9304 (N_9304,N_9227,N_9200);
or U9305 (N_9305,N_9228,N_9266);
nor U9306 (N_9306,N_9229,N_9128);
nor U9307 (N_9307,N_9257,N_9158);
and U9308 (N_9308,N_9261,N_9173);
or U9309 (N_9309,N_9126,N_9240);
nand U9310 (N_9310,N_9189,N_9141);
or U9311 (N_9311,N_9249,N_9202);
and U9312 (N_9312,N_9255,N_9264);
nor U9313 (N_9313,N_9256,N_9149);
nand U9314 (N_9314,N_9198,N_9146);
nor U9315 (N_9315,N_9159,N_9135);
nand U9316 (N_9316,N_9219,N_9170);
and U9317 (N_9317,N_9190,N_9199);
nor U9318 (N_9318,N_9186,N_9211);
nor U9319 (N_9319,N_9207,N_9130);
nor U9320 (N_9320,N_9258,N_9193);
nor U9321 (N_9321,N_9127,N_9267);
and U9322 (N_9322,N_9218,N_9230);
and U9323 (N_9323,N_9226,N_9192);
nor U9324 (N_9324,N_9221,N_9273);
nor U9325 (N_9325,N_9243,N_9145);
nor U9326 (N_9326,N_9181,N_9140);
nor U9327 (N_9327,N_9239,N_9250);
xor U9328 (N_9328,N_9177,N_9179);
or U9329 (N_9329,N_9275,N_9142);
and U9330 (N_9330,N_9176,N_9242);
or U9331 (N_9331,N_9161,N_9166);
nand U9332 (N_9332,N_9204,N_9206);
xor U9333 (N_9333,N_9123,N_9125);
and U9334 (N_9334,N_9143,N_9133);
nor U9335 (N_9335,N_9139,N_9195);
nand U9336 (N_9336,N_9246,N_9252);
nor U9337 (N_9337,N_9120,N_9129);
or U9338 (N_9338,N_9162,N_9156);
nor U9339 (N_9339,N_9194,N_9151);
nor U9340 (N_9340,N_9222,N_9157);
or U9341 (N_9341,N_9270,N_9174);
and U9342 (N_9342,N_9188,N_9180);
nor U9343 (N_9343,N_9210,N_9234);
or U9344 (N_9344,N_9217,N_9262);
nand U9345 (N_9345,N_9223,N_9269);
nand U9346 (N_9346,N_9137,N_9184);
nor U9347 (N_9347,N_9263,N_9171);
or U9348 (N_9348,N_9238,N_9236);
nor U9349 (N_9349,N_9241,N_9121);
and U9350 (N_9350,N_9150,N_9277);
and U9351 (N_9351,N_9214,N_9172);
nand U9352 (N_9352,N_9148,N_9235);
and U9353 (N_9353,N_9168,N_9197);
nor U9354 (N_9354,N_9187,N_9122);
or U9355 (N_9355,N_9245,N_9169);
nor U9356 (N_9356,N_9155,N_9147);
nor U9357 (N_9357,N_9233,N_9164);
xor U9358 (N_9358,N_9260,N_9237);
xor U9359 (N_9359,N_9196,N_9231);
or U9360 (N_9360,N_9211,N_9227);
or U9361 (N_9361,N_9130,N_9216);
or U9362 (N_9362,N_9135,N_9126);
nand U9363 (N_9363,N_9269,N_9248);
or U9364 (N_9364,N_9145,N_9171);
xnor U9365 (N_9365,N_9144,N_9167);
and U9366 (N_9366,N_9129,N_9188);
nor U9367 (N_9367,N_9201,N_9186);
nor U9368 (N_9368,N_9166,N_9203);
and U9369 (N_9369,N_9149,N_9139);
nand U9370 (N_9370,N_9199,N_9243);
or U9371 (N_9371,N_9217,N_9226);
and U9372 (N_9372,N_9126,N_9143);
and U9373 (N_9373,N_9190,N_9276);
and U9374 (N_9374,N_9245,N_9225);
and U9375 (N_9375,N_9136,N_9185);
nor U9376 (N_9376,N_9244,N_9228);
or U9377 (N_9377,N_9220,N_9270);
or U9378 (N_9378,N_9130,N_9141);
xnor U9379 (N_9379,N_9260,N_9129);
and U9380 (N_9380,N_9172,N_9244);
xor U9381 (N_9381,N_9224,N_9269);
nor U9382 (N_9382,N_9120,N_9190);
and U9383 (N_9383,N_9239,N_9187);
nand U9384 (N_9384,N_9278,N_9162);
and U9385 (N_9385,N_9214,N_9198);
and U9386 (N_9386,N_9121,N_9233);
and U9387 (N_9387,N_9172,N_9211);
and U9388 (N_9388,N_9193,N_9215);
and U9389 (N_9389,N_9125,N_9252);
or U9390 (N_9390,N_9201,N_9217);
and U9391 (N_9391,N_9243,N_9247);
nor U9392 (N_9392,N_9262,N_9191);
or U9393 (N_9393,N_9186,N_9270);
nor U9394 (N_9394,N_9172,N_9202);
or U9395 (N_9395,N_9144,N_9184);
and U9396 (N_9396,N_9246,N_9262);
nor U9397 (N_9397,N_9128,N_9126);
or U9398 (N_9398,N_9237,N_9154);
xnor U9399 (N_9399,N_9142,N_9138);
nor U9400 (N_9400,N_9247,N_9251);
or U9401 (N_9401,N_9136,N_9218);
nor U9402 (N_9402,N_9220,N_9160);
or U9403 (N_9403,N_9120,N_9192);
nor U9404 (N_9404,N_9237,N_9120);
xor U9405 (N_9405,N_9224,N_9153);
nor U9406 (N_9406,N_9228,N_9158);
nand U9407 (N_9407,N_9197,N_9161);
nand U9408 (N_9408,N_9206,N_9238);
xor U9409 (N_9409,N_9248,N_9211);
and U9410 (N_9410,N_9264,N_9218);
nand U9411 (N_9411,N_9124,N_9249);
and U9412 (N_9412,N_9263,N_9164);
or U9413 (N_9413,N_9255,N_9166);
and U9414 (N_9414,N_9203,N_9184);
and U9415 (N_9415,N_9169,N_9197);
xnor U9416 (N_9416,N_9157,N_9166);
nor U9417 (N_9417,N_9130,N_9226);
nor U9418 (N_9418,N_9212,N_9201);
nor U9419 (N_9419,N_9248,N_9241);
nor U9420 (N_9420,N_9206,N_9256);
or U9421 (N_9421,N_9256,N_9120);
or U9422 (N_9422,N_9163,N_9162);
nor U9423 (N_9423,N_9183,N_9226);
and U9424 (N_9424,N_9194,N_9228);
nor U9425 (N_9425,N_9142,N_9209);
nand U9426 (N_9426,N_9259,N_9239);
nand U9427 (N_9427,N_9278,N_9217);
and U9428 (N_9428,N_9268,N_9158);
xnor U9429 (N_9429,N_9145,N_9211);
and U9430 (N_9430,N_9178,N_9239);
and U9431 (N_9431,N_9250,N_9164);
nand U9432 (N_9432,N_9208,N_9137);
nor U9433 (N_9433,N_9161,N_9160);
and U9434 (N_9434,N_9199,N_9257);
xor U9435 (N_9435,N_9130,N_9271);
nand U9436 (N_9436,N_9158,N_9146);
and U9437 (N_9437,N_9189,N_9146);
or U9438 (N_9438,N_9139,N_9279);
and U9439 (N_9439,N_9201,N_9276);
or U9440 (N_9440,N_9322,N_9287);
nor U9441 (N_9441,N_9370,N_9399);
or U9442 (N_9442,N_9437,N_9346);
nor U9443 (N_9443,N_9288,N_9353);
and U9444 (N_9444,N_9408,N_9335);
and U9445 (N_9445,N_9431,N_9415);
or U9446 (N_9446,N_9311,N_9356);
nand U9447 (N_9447,N_9386,N_9334);
or U9448 (N_9448,N_9319,N_9402);
and U9449 (N_9449,N_9298,N_9316);
and U9450 (N_9450,N_9403,N_9350);
and U9451 (N_9451,N_9348,N_9338);
or U9452 (N_9452,N_9329,N_9397);
nor U9453 (N_9453,N_9313,N_9331);
nor U9454 (N_9454,N_9336,N_9285);
and U9455 (N_9455,N_9365,N_9351);
and U9456 (N_9456,N_9339,N_9405);
nand U9457 (N_9457,N_9290,N_9379);
or U9458 (N_9458,N_9320,N_9326);
nor U9459 (N_9459,N_9284,N_9385);
and U9460 (N_9460,N_9304,N_9286);
and U9461 (N_9461,N_9376,N_9377);
nand U9462 (N_9462,N_9330,N_9315);
and U9463 (N_9463,N_9303,N_9400);
nand U9464 (N_9464,N_9325,N_9384);
or U9465 (N_9465,N_9395,N_9375);
or U9466 (N_9466,N_9404,N_9412);
nor U9467 (N_9467,N_9394,N_9372);
nor U9468 (N_9468,N_9436,N_9423);
and U9469 (N_9469,N_9439,N_9332);
or U9470 (N_9470,N_9411,N_9352);
xnor U9471 (N_9471,N_9307,N_9299);
nor U9472 (N_9472,N_9341,N_9396);
or U9473 (N_9473,N_9308,N_9294);
xnor U9474 (N_9474,N_9416,N_9433);
or U9475 (N_9475,N_9337,N_9327);
or U9476 (N_9476,N_9295,N_9310);
or U9477 (N_9477,N_9359,N_9419);
or U9478 (N_9478,N_9378,N_9301);
nand U9479 (N_9479,N_9318,N_9289);
nor U9480 (N_9480,N_9343,N_9417);
xor U9481 (N_9481,N_9393,N_9438);
or U9482 (N_9482,N_9398,N_9342);
and U9483 (N_9483,N_9354,N_9374);
and U9484 (N_9484,N_9418,N_9428);
and U9485 (N_9485,N_9383,N_9410);
and U9486 (N_9486,N_9409,N_9302);
nor U9487 (N_9487,N_9362,N_9373);
or U9488 (N_9488,N_9426,N_9382);
or U9489 (N_9489,N_9391,N_9407);
or U9490 (N_9490,N_9309,N_9363);
and U9491 (N_9491,N_9349,N_9435);
xor U9492 (N_9492,N_9371,N_9297);
nand U9493 (N_9493,N_9314,N_9280);
or U9494 (N_9494,N_9387,N_9317);
nand U9495 (N_9495,N_9357,N_9388);
nand U9496 (N_9496,N_9420,N_9392);
and U9497 (N_9497,N_9413,N_9324);
and U9498 (N_9498,N_9361,N_9340);
nand U9499 (N_9499,N_9425,N_9432);
nor U9500 (N_9500,N_9347,N_9283);
nand U9501 (N_9501,N_9305,N_9281);
and U9502 (N_9502,N_9366,N_9364);
xor U9503 (N_9503,N_9293,N_9380);
and U9504 (N_9504,N_9360,N_9424);
nand U9505 (N_9505,N_9355,N_9434);
xor U9506 (N_9506,N_9344,N_9381);
nor U9507 (N_9507,N_9389,N_9368);
or U9508 (N_9508,N_9367,N_9390);
and U9509 (N_9509,N_9328,N_9401);
nor U9510 (N_9510,N_9430,N_9421);
nand U9511 (N_9511,N_9427,N_9312);
and U9512 (N_9512,N_9323,N_9300);
nor U9513 (N_9513,N_9358,N_9333);
and U9514 (N_9514,N_9422,N_9292);
or U9515 (N_9515,N_9406,N_9306);
and U9516 (N_9516,N_9369,N_9282);
nor U9517 (N_9517,N_9291,N_9414);
xor U9518 (N_9518,N_9429,N_9345);
or U9519 (N_9519,N_9296,N_9321);
xor U9520 (N_9520,N_9348,N_9357);
nand U9521 (N_9521,N_9399,N_9347);
nor U9522 (N_9522,N_9406,N_9339);
or U9523 (N_9523,N_9282,N_9319);
nand U9524 (N_9524,N_9427,N_9382);
and U9525 (N_9525,N_9310,N_9326);
nand U9526 (N_9526,N_9353,N_9417);
nand U9527 (N_9527,N_9389,N_9316);
nand U9528 (N_9528,N_9343,N_9412);
and U9529 (N_9529,N_9358,N_9346);
nand U9530 (N_9530,N_9439,N_9379);
or U9531 (N_9531,N_9358,N_9406);
or U9532 (N_9532,N_9363,N_9351);
nand U9533 (N_9533,N_9305,N_9375);
nor U9534 (N_9534,N_9378,N_9401);
nor U9535 (N_9535,N_9424,N_9421);
and U9536 (N_9536,N_9401,N_9427);
or U9537 (N_9537,N_9362,N_9421);
or U9538 (N_9538,N_9281,N_9359);
and U9539 (N_9539,N_9366,N_9385);
xnor U9540 (N_9540,N_9316,N_9356);
and U9541 (N_9541,N_9299,N_9421);
and U9542 (N_9542,N_9414,N_9342);
nor U9543 (N_9543,N_9410,N_9419);
nand U9544 (N_9544,N_9317,N_9410);
xnor U9545 (N_9545,N_9381,N_9340);
xor U9546 (N_9546,N_9344,N_9437);
and U9547 (N_9547,N_9340,N_9327);
nand U9548 (N_9548,N_9380,N_9420);
or U9549 (N_9549,N_9365,N_9282);
and U9550 (N_9550,N_9312,N_9396);
nand U9551 (N_9551,N_9406,N_9321);
and U9552 (N_9552,N_9407,N_9412);
and U9553 (N_9553,N_9308,N_9394);
nor U9554 (N_9554,N_9411,N_9432);
and U9555 (N_9555,N_9410,N_9314);
or U9556 (N_9556,N_9384,N_9377);
nor U9557 (N_9557,N_9397,N_9405);
and U9558 (N_9558,N_9370,N_9326);
nor U9559 (N_9559,N_9338,N_9420);
nand U9560 (N_9560,N_9388,N_9394);
and U9561 (N_9561,N_9356,N_9310);
or U9562 (N_9562,N_9346,N_9420);
nand U9563 (N_9563,N_9312,N_9432);
nand U9564 (N_9564,N_9299,N_9384);
nor U9565 (N_9565,N_9310,N_9405);
or U9566 (N_9566,N_9406,N_9363);
nor U9567 (N_9567,N_9364,N_9290);
and U9568 (N_9568,N_9434,N_9415);
xor U9569 (N_9569,N_9349,N_9312);
xnor U9570 (N_9570,N_9307,N_9311);
nor U9571 (N_9571,N_9422,N_9406);
and U9572 (N_9572,N_9348,N_9437);
and U9573 (N_9573,N_9430,N_9358);
and U9574 (N_9574,N_9360,N_9418);
or U9575 (N_9575,N_9311,N_9342);
nor U9576 (N_9576,N_9293,N_9286);
or U9577 (N_9577,N_9427,N_9357);
nor U9578 (N_9578,N_9433,N_9355);
nor U9579 (N_9579,N_9404,N_9407);
nor U9580 (N_9580,N_9306,N_9325);
and U9581 (N_9581,N_9336,N_9416);
xor U9582 (N_9582,N_9383,N_9308);
or U9583 (N_9583,N_9381,N_9396);
or U9584 (N_9584,N_9405,N_9432);
and U9585 (N_9585,N_9357,N_9385);
and U9586 (N_9586,N_9345,N_9371);
and U9587 (N_9587,N_9299,N_9347);
and U9588 (N_9588,N_9304,N_9376);
and U9589 (N_9589,N_9395,N_9438);
or U9590 (N_9590,N_9393,N_9414);
and U9591 (N_9591,N_9406,N_9376);
and U9592 (N_9592,N_9324,N_9357);
nor U9593 (N_9593,N_9289,N_9383);
or U9594 (N_9594,N_9396,N_9284);
nor U9595 (N_9595,N_9357,N_9317);
nor U9596 (N_9596,N_9402,N_9344);
nor U9597 (N_9597,N_9426,N_9303);
nor U9598 (N_9598,N_9439,N_9362);
xor U9599 (N_9599,N_9417,N_9424);
xnor U9600 (N_9600,N_9441,N_9508);
nand U9601 (N_9601,N_9586,N_9447);
nor U9602 (N_9602,N_9524,N_9546);
nand U9603 (N_9603,N_9481,N_9555);
or U9604 (N_9604,N_9485,N_9495);
nor U9605 (N_9605,N_9476,N_9510);
and U9606 (N_9606,N_9507,N_9587);
nand U9607 (N_9607,N_9550,N_9489);
and U9608 (N_9608,N_9473,N_9558);
and U9609 (N_9609,N_9465,N_9482);
or U9610 (N_9610,N_9459,N_9458);
or U9611 (N_9611,N_9523,N_9514);
nor U9612 (N_9612,N_9486,N_9519);
nor U9613 (N_9613,N_9551,N_9528);
nand U9614 (N_9614,N_9454,N_9597);
nand U9615 (N_9615,N_9537,N_9569);
nand U9616 (N_9616,N_9502,N_9496);
xor U9617 (N_9617,N_9440,N_9517);
and U9618 (N_9618,N_9503,N_9491);
and U9619 (N_9619,N_9584,N_9563);
nand U9620 (N_9620,N_9548,N_9566);
nand U9621 (N_9621,N_9553,N_9543);
or U9622 (N_9622,N_9591,N_9544);
or U9623 (N_9623,N_9449,N_9515);
nor U9624 (N_9624,N_9444,N_9525);
xnor U9625 (N_9625,N_9590,N_9490);
and U9626 (N_9626,N_9534,N_9578);
nand U9627 (N_9627,N_9493,N_9469);
and U9628 (N_9628,N_9562,N_9451);
and U9629 (N_9629,N_9540,N_9512);
nand U9630 (N_9630,N_9560,N_9477);
nand U9631 (N_9631,N_9539,N_9588);
and U9632 (N_9632,N_9471,N_9554);
nand U9633 (N_9633,N_9463,N_9487);
nor U9634 (N_9634,N_9585,N_9498);
and U9635 (N_9635,N_9462,N_9509);
and U9636 (N_9636,N_9499,N_9567);
and U9637 (N_9637,N_9541,N_9466);
and U9638 (N_9638,N_9535,N_9580);
and U9639 (N_9639,N_9542,N_9522);
or U9640 (N_9640,N_9538,N_9595);
or U9641 (N_9641,N_9547,N_9470);
nand U9642 (N_9642,N_9531,N_9445);
or U9643 (N_9643,N_9474,N_9579);
and U9644 (N_9644,N_9518,N_9599);
and U9645 (N_9645,N_9483,N_9564);
nand U9646 (N_9646,N_9596,N_9526);
nand U9647 (N_9647,N_9573,N_9464);
nor U9648 (N_9648,N_9500,N_9501);
xor U9649 (N_9649,N_9468,N_9589);
nand U9650 (N_9650,N_9568,N_9576);
and U9651 (N_9651,N_9457,N_9571);
or U9652 (N_9652,N_9521,N_9479);
nor U9653 (N_9653,N_9565,N_9452);
or U9654 (N_9654,N_9533,N_9506);
nor U9655 (N_9655,N_9583,N_9442);
or U9656 (N_9656,N_9549,N_9581);
nor U9657 (N_9657,N_9575,N_9446);
nand U9658 (N_9658,N_9530,N_9572);
or U9659 (N_9659,N_9460,N_9594);
xor U9660 (N_9660,N_9545,N_9513);
and U9661 (N_9661,N_9574,N_9497);
nor U9662 (N_9662,N_9593,N_9520);
and U9663 (N_9663,N_9529,N_9480);
or U9664 (N_9664,N_9484,N_9582);
or U9665 (N_9665,N_9448,N_9552);
nor U9666 (N_9666,N_9488,N_9504);
nor U9667 (N_9667,N_9505,N_9577);
nor U9668 (N_9668,N_9461,N_9492);
or U9669 (N_9669,N_9557,N_9532);
and U9670 (N_9670,N_9556,N_9455);
and U9671 (N_9671,N_9598,N_9450);
and U9672 (N_9672,N_9475,N_9494);
nor U9673 (N_9673,N_9592,N_9527);
nand U9674 (N_9674,N_9511,N_9559);
nor U9675 (N_9675,N_9516,N_9472);
nor U9676 (N_9676,N_9536,N_9453);
or U9677 (N_9677,N_9561,N_9478);
or U9678 (N_9678,N_9570,N_9456);
or U9679 (N_9679,N_9443,N_9467);
nand U9680 (N_9680,N_9498,N_9573);
nor U9681 (N_9681,N_9470,N_9482);
or U9682 (N_9682,N_9485,N_9527);
and U9683 (N_9683,N_9463,N_9567);
nand U9684 (N_9684,N_9512,N_9516);
or U9685 (N_9685,N_9444,N_9595);
nor U9686 (N_9686,N_9549,N_9569);
nand U9687 (N_9687,N_9535,N_9494);
nand U9688 (N_9688,N_9591,N_9460);
and U9689 (N_9689,N_9463,N_9539);
nand U9690 (N_9690,N_9594,N_9549);
nand U9691 (N_9691,N_9578,N_9597);
or U9692 (N_9692,N_9471,N_9497);
xor U9693 (N_9693,N_9500,N_9523);
nor U9694 (N_9694,N_9518,N_9563);
nand U9695 (N_9695,N_9452,N_9521);
and U9696 (N_9696,N_9552,N_9536);
nand U9697 (N_9697,N_9492,N_9561);
and U9698 (N_9698,N_9482,N_9477);
nand U9699 (N_9699,N_9452,N_9560);
nor U9700 (N_9700,N_9514,N_9442);
or U9701 (N_9701,N_9577,N_9538);
xnor U9702 (N_9702,N_9500,N_9441);
or U9703 (N_9703,N_9515,N_9549);
or U9704 (N_9704,N_9450,N_9523);
or U9705 (N_9705,N_9579,N_9525);
and U9706 (N_9706,N_9450,N_9511);
nand U9707 (N_9707,N_9469,N_9574);
nand U9708 (N_9708,N_9486,N_9443);
nand U9709 (N_9709,N_9503,N_9504);
nand U9710 (N_9710,N_9469,N_9587);
or U9711 (N_9711,N_9483,N_9563);
or U9712 (N_9712,N_9594,N_9566);
nand U9713 (N_9713,N_9474,N_9534);
nand U9714 (N_9714,N_9502,N_9531);
nand U9715 (N_9715,N_9572,N_9557);
nor U9716 (N_9716,N_9474,N_9529);
nor U9717 (N_9717,N_9562,N_9575);
nor U9718 (N_9718,N_9502,N_9535);
nand U9719 (N_9719,N_9536,N_9502);
and U9720 (N_9720,N_9560,N_9555);
nor U9721 (N_9721,N_9461,N_9486);
or U9722 (N_9722,N_9527,N_9523);
or U9723 (N_9723,N_9503,N_9512);
and U9724 (N_9724,N_9599,N_9462);
or U9725 (N_9725,N_9466,N_9556);
nor U9726 (N_9726,N_9475,N_9456);
or U9727 (N_9727,N_9456,N_9503);
and U9728 (N_9728,N_9452,N_9524);
and U9729 (N_9729,N_9476,N_9503);
nor U9730 (N_9730,N_9529,N_9492);
or U9731 (N_9731,N_9534,N_9480);
nor U9732 (N_9732,N_9594,N_9547);
and U9733 (N_9733,N_9460,N_9476);
and U9734 (N_9734,N_9441,N_9506);
nand U9735 (N_9735,N_9540,N_9452);
nor U9736 (N_9736,N_9476,N_9523);
nor U9737 (N_9737,N_9477,N_9556);
nand U9738 (N_9738,N_9580,N_9563);
and U9739 (N_9739,N_9441,N_9483);
and U9740 (N_9740,N_9593,N_9453);
or U9741 (N_9741,N_9548,N_9462);
nand U9742 (N_9742,N_9471,N_9559);
and U9743 (N_9743,N_9542,N_9443);
nor U9744 (N_9744,N_9490,N_9582);
nor U9745 (N_9745,N_9594,N_9445);
xor U9746 (N_9746,N_9457,N_9446);
and U9747 (N_9747,N_9588,N_9535);
or U9748 (N_9748,N_9562,N_9504);
or U9749 (N_9749,N_9523,N_9516);
nor U9750 (N_9750,N_9510,N_9445);
xnor U9751 (N_9751,N_9564,N_9478);
nor U9752 (N_9752,N_9580,N_9492);
and U9753 (N_9753,N_9543,N_9583);
nor U9754 (N_9754,N_9548,N_9452);
and U9755 (N_9755,N_9459,N_9468);
nor U9756 (N_9756,N_9534,N_9475);
nand U9757 (N_9757,N_9490,N_9459);
nand U9758 (N_9758,N_9471,N_9465);
or U9759 (N_9759,N_9572,N_9480);
nor U9760 (N_9760,N_9649,N_9687);
and U9761 (N_9761,N_9636,N_9747);
and U9762 (N_9762,N_9658,N_9681);
nand U9763 (N_9763,N_9690,N_9624);
or U9764 (N_9764,N_9709,N_9744);
nor U9765 (N_9765,N_9610,N_9612);
or U9766 (N_9766,N_9736,N_9707);
nand U9767 (N_9767,N_9746,N_9609);
xnor U9768 (N_9768,N_9627,N_9685);
and U9769 (N_9769,N_9728,N_9640);
xnor U9770 (N_9770,N_9743,N_9712);
or U9771 (N_9771,N_9622,N_9625);
or U9772 (N_9772,N_9725,N_9650);
and U9773 (N_9773,N_9694,N_9734);
or U9774 (N_9774,N_9713,N_9715);
xor U9775 (N_9775,N_9710,N_9724);
nor U9776 (N_9776,N_9669,N_9684);
and U9777 (N_9777,N_9695,N_9623);
or U9778 (N_9778,N_9673,N_9702);
or U9779 (N_9779,N_9637,N_9708);
nand U9780 (N_9780,N_9641,N_9705);
or U9781 (N_9781,N_9675,N_9693);
or U9782 (N_9782,N_9654,N_9618);
and U9783 (N_9783,N_9602,N_9758);
xnor U9784 (N_9784,N_9737,N_9730);
and U9785 (N_9785,N_9601,N_9689);
xnor U9786 (N_9786,N_9635,N_9679);
or U9787 (N_9787,N_9677,N_9680);
nand U9788 (N_9788,N_9631,N_9671);
and U9789 (N_9789,N_9745,N_9750);
nor U9790 (N_9790,N_9757,N_9714);
and U9791 (N_9791,N_9605,N_9608);
and U9792 (N_9792,N_9692,N_9652);
nand U9793 (N_9793,N_9697,N_9616);
nand U9794 (N_9794,N_9666,N_9678);
nor U9795 (N_9795,N_9633,N_9756);
xor U9796 (N_9796,N_9629,N_9674);
or U9797 (N_9797,N_9600,N_9661);
and U9798 (N_9798,N_9759,N_9699);
xnor U9799 (N_9799,N_9613,N_9711);
or U9800 (N_9800,N_9651,N_9659);
nor U9801 (N_9801,N_9644,N_9646);
nand U9802 (N_9802,N_9755,N_9751);
or U9803 (N_9803,N_9620,N_9698);
nand U9804 (N_9804,N_9670,N_9749);
nand U9805 (N_9805,N_9683,N_9626);
nor U9806 (N_9806,N_9630,N_9628);
nor U9807 (N_9807,N_9723,N_9647);
or U9808 (N_9808,N_9682,N_9688);
nor U9809 (N_9809,N_9722,N_9603);
or U9810 (N_9810,N_9718,N_9726);
nor U9811 (N_9811,N_9721,N_9639);
nand U9812 (N_9812,N_9611,N_9754);
nand U9813 (N_9813,N_9732,N_9719);
or U9814 (N_9814,N_9606,N_9663);
xnor U9815 (N_9815,N_9735,N_9704);
nand U9816 (N_9816,N_9739,N_9655);
and U9817 (N_9817,N_9665,N_9664);
nand U9818 (N_9818,N_9700,N_9607);
nor U9819 (N_9819,N_9696,N_9741);
nand U9820 (N_9820,N_9738,N_9752);
and U9821 (N_9821,N_9615,N_9617);
and U9822 (N_9822,N_9642,N_9742);
and U9823 (N_9823,N_9619,N_9733);
and U9824 (N_9824,N_9740,N_9662);
and U9825 (N_9825,N_9668,N_9614);
nor U9826 (N_9826,N_9667,N_9653);
and U9827 (N_9827,N_9703,N_9645);
or U9828 (N_9828,N_9691,N_9720);
or U9829 (N_9829,N_9643,N_9604);
and U9830 (N_9830,N_9727,N_9676);
or U9831 (N_9831,N_9748,N_9632);
nor U9832 (N_9832,N_9701,N_9638);
and U9833 (N_9833,N_9706,N_9621);
or U9834 (N_9834,N_9656,N_9634);
nor U9835 (N_9835,N_9660,N_9731);
nor U9836 (N_9836,N_9729,N_9717);
and U9837 (N_9837,N_9686,N_9753);
nand U9838 (N_9838,N_9672,N_9657);
and U9839 (N_9839,N_9648,N_9716);
and U9840 (N_9840,N_9643,N_9733);
or U9841 (N_9841,N_9672,N_9661);
nor U9842 (N_9842,N_9747,N_9703);
nand U9843 (N_9843,N_9716,N_9671);
nor U9844 (N_9844,N_9642,N_9681);
nor U9845 (N_9845,N_9673,N_9753);
and U9846 (N_9846,N_9654,N_9745);
nor U9847 (N_9847,N_9628,N_9678);
nor U9848 (N_9848,N_9607,N_9627);
or U9849 (N_9849,N_9659,N_9638);
or U9850 (N_9850,N_9644,N_9637);
or U9851 (N_9851,N_9620,N_9639);
and U9852 (N_9852,N_9736,N_9726);
or U9853 (N_9853,N_9756,N_9747);
nor U9854 (N_9854,N_9724,N_9619);
nand U9855 (N_9855,N_9614,N_9617);
nand U9856 (N_9856,N_9696,N_9660);
nor U9857 (N_9857,N_9712,N_9676);
or U9858 (N_9858,N_9645,N_9675);
nor U9859 (N_9859,N_9708,N_9714);
nand U9860 (N_9860,N_9655,N_9692);
nor U9861 (N_9861,N_9711,N_9717);
nand U9862 (N_9862,N_9626,N_9687);
and U9863 (N_9863,N_9671,N_9715);
xnor U9864 (N_9864,N_9746,N_9692);
nor U9865 (N_9865,N_9698,N_9667);
nand U9866 (N_9866,N_9679,N_9744);
or U9867 (N_9867,N_9729,N_9666);
xor U9868 (N_9868,N_9602,N_9634);
nand U9869 (N_9869,N_9720,N_9689);
nor U9870 (N_9870,N_9625,N_9689);
and U9871 (N_9871,N_9651,N_9755);
and U9872 (N_9872,N_9699,N_9727);
and U9873 (N_9873,N_9747,N_9669);
and U9874 (N_9874,N_9686,N_9699);
nor U9875 (N_9875,N_9700,N_9705);
and U9876 (N_9876,N_9750,N_9601);
or U9877 (N_9877,N_9616,N_9727);
or U9878 (N_9878,N_9605,N_9689);
or U9879 (N_9879,N_9706,N_9613);
nor U9880 (N_9880,N_9683,N_9711);
nand U9881 (N_9881,N_9657,N_9744);
or U9882 (N_9882,N_9714,N_9681);
and U9883 (N_9883,N_9744,N_9644);
or U9884 (N_9884,N_9697,N_9700);
nand U9885 (N_9885,N_9759,N_9606);
nor U9886 (N_9886,N_9643,N_9691);
nor U9887 (N_9887,N_9700,N_9685);
and U9888 (N_9888,N_9704,N_9726);
nor U9889 (N_9889,N_9660,N_9750);
nor U9890 (N_9890,N_9672,N_9604);
nand U9891 (N_9891,N_9605,N_9666);
nand U9892 (N_9892,N_9756,N_9735);
and U9893 (N_9893,N_9721,N_9681);
xor U9894 (N_9894,N_9720,N_9609);
nand U9895 (N_9895,N_9657,N_9646);
or U9896 (N_9896,N_9632,N_9741);
nand U9897 (N_9897,N_9759,N_9612);
nor U9898 (N_9898,N_9726,N_9676);
or U9899 (N_9899,N_9684,N_9645);
nand U9900 (N_9900,N_9649,N_9704);
or U9901 (N_9901,N_9605,N_9724);
nor U9902 (N_9902,N_9702,N_9729);
nor U9903 (N_9903,N_9687,N_9706);
or U9904 (N_9904,N_9733,N_9701);
nor U9905 (N_9905,N_9690,N_9647);
and U9906 (N_9906,N_9610,N_9754);
and U9907 (N_9907,N_9749,N_9628);
and U9908 (N_9908,N_9723,N_9664);
nand U9909 (N_9909,N_9713,N_9725);
nor U9910 (N_9910,N_9687,N_9723);
xnor U9911 (N_9911,N_9676,N_9750);
and U9912 (N_9912,N_9650,N_9632);
or U9913 (N_9913,N_9659,N_9705);
and U9914 (N_9914,N_9733,N_9705);
nor U9915 (N_9915,N_9697,N_9620);
or U9916 (N_9916,N_9741,N_9620);
or U9917 (N_9917,N_9612,N_9601);
or U9918 (N_9918,N_9624,N_9725);
or U9919 (N_9919,N_9708,N_9651);
and U9920 (N_9920,N_9845,N_9892);
or U9921 (N_9921,N_9824,N_9847);
or U9922 (N_9922,N_9768,N_9861);
or U9923 (N_9923,N_9884,N_9797);
and U9924 (N_9924,N_9891,N_9841);
or U9925 (N_9925,N_9795,N_9881);
nor U9926 (N_9926,N_9802,N_9885);
xor U9927 (N_9927,N_9794,N_9904);
nor U9928 (N_9928,N_9886,N_9828);
nor U9929 (N_9929,N_9832,N_9830);
nor U9930 (N_9930,N_9809,N_9900);
and U9931 (N_9931,N_9798,N_9883);
nor U9932 (N_9932,N_9919,N_9868);
nor U9933 (N_9933,N_9829,N_9916);
or U9934 (N_9934,N_9858,N_9894);
xor U9935 (N_9935,N_9869,N_9889);
and U9936 (N_9936,N_9834,N_9862);
or U9937 (N_9937,N_9807,N_9875);
nand U9938 (N_9938,N_9872,N_9775);
nand U9939 (N_9939,N_9863,N_9910);
nor U9940 (N_9940,N_9903,N_9804);
and U9941 (N_9941,N_9827,N_9781);
or U9942 (N_9942,N_9866,N_9831);
nor U9943 (N_9943,N_9856,N_9851);
nand U9944 (N_9944,N_9770,N_9776);
nand U9945 (N_9945,N_9805,N_9819);
nand U9946 (N_9946,N_9810,N_9895);
nand U9947 (N_9947,N_9912,N_9906);
nor U9948 (N_9948,N_9865,N_9792);
or U9949 (N_9949,N_9901,N_9789);
nor U9950 (N_9950,N_9803,N_9821);
nor U9951 (N_9951,N_9762,N_9898);
and U9952 (N_9952,N_9835,N_9867);
xnor U9953 (N_9953,N_9913,N_9774);
nand U9954 (N_9954,N_9908,N_9849);
and U9955 (N_9955,N_9860,N_9769);
nand U9956 (N_9956,N_9837,N_9800);
nor U9957 (N_9957,N_9814,N_9779);
or U9958 (N_9958,N_9918,N_9820);
and U9959 (N_9959,N_9780,N_9811);
nand U9960 (N_9960,N_9764,N_9876);
nand U9961 (N_9961,N_9799,N_9907);
and U9962 (N_9962,N_9787,N_9772);
or U9963 (N_9963,N_9778,N_9888);
nand U9964 (N_9964,N_9890,N_9871);
nor U9965 (N_9965,N_9914,N_9822);
xor U9966 (N_9966,N_9878,N_9911);
xnor U9967 (N_9967,N_9760,N_9763);
nand U9968 (N_9968,N_9846,N_9844);
nor U9969 (N_9969,N_9817,N_9765);
nand U9970 (N_9970,N_9853,N_9816);
nand U9971 (N_9971,N_9761,N_9788);
and U9972 (N_9972,N_9796,N_9839);
nand U9973 (N_9973,N_9838,N_9897);
xor U9974 (N_9974,N_9859,N_9823);
xor U9975 (N_9975,N_9854,N_9899);
or U9976 (N_9976,N_9887,N_9777);
xor U9977 (N_9977,N_9842,N_9791);
or U9978 (N_9978,N_9812,N_9818);
or U9979 (N_9979,N_9893,N_9880);
nand U9980 (N_9980,N_9784,N_9833);
and U9981 (N_9981,N_9836,N_9909);
nand U9982 (N_9982,N_9857,N_9873);
nand U9983 (N_9983,N_9786,N_9840);
or U9984 (N_9984,N_9870,N_9783);
or U9985 (N_9985,N_9855,N_9917);
or U9986 (N_9986,N_9826,N_9848);
and U9987 (N_9987,N_9850,N_9773);
or U9988 (N_9988,N_9808,N_9843);
nand U9989 (N_9989,N_9801,N_9782);
or U9990 (N_9990,N_9813,N_9852);
and U9991 (N_9991,N_9806,N_9790);
nor U9992 (N_9992,N_9905,N_9793);
or U9993 (N_9993,N_9771,N_9879);
nor U9994 (N_9994,N_9896,N_9864);
xnor U9995 (N_9995,N_9874,N_9825);
nand U9996 (N_9996,N_9785,N_9767);
and U9997 (N_9997,N_9902,N_9877);
nand U9998 (N_9998,N_9766,N_9915);
and U9999 (N_9999,N_9815,N_9882);
and U10000 (N_10000,N_9818,N_9805);
xnor U10001 (N_10001,N_9895,N_9878);
and U10002 (N_10002,N_9840,N_9858);
nor U10003 (N_10003,N_9785,N_9823);
nand U10004 (N_10004,N_9798,N_9850);
and U10005 (N_10005,N_9816,N_9836);
nor U10006 (N_10006,N_9905,N_9774);
xor U10007 (N_10007,N_9874,N_9862);
or U10008 (N_10008,N_9784,N_9800);
nor U10009 (N_10009,N_9883,N_9864);
nand U10010 (N_10010,N_9770,N_9783);
and U10011 (N_10011,N_9764,N_9824);
nor U10012 (N_10012,N_9864,N_9829);
or U10013 (N_10013,N_9770,N_9854);
xnor U10014 (N_10014,N_9771,N_9893);
and U10015 (N_10015,N_9810,N_9842);
nor U10016 (N_10016,N_9815,N_9901);
nor U10017 (N_10017,N_9880,N_9776);
xnor U10018 (N_10018,N_9784,N_9875);
xnor U10019 (N_10019,N_9874,N_9892);
nand U10020 (N_10020,N_9847,N_9875);
or U10021 (N_10021,N_9899,N_9783);
or U10022 (N_10022,N_9905,N_9891);
nor U10023 (N_10023,N_9821,N_9771);
and U10024 (N_10024,N_9909,N_9797);
and U10025 (N_10025,N_9797,N_9786);
nor U10026 (N_10026,N_9768,N_9867);
nand U10027 (N_10027,N_9766,N_9872);
nand U10028 (N_10028,N_9900,N_9777);
nand U10029 (N_10029,N_9884,N_9898);
nand U10030 (N_10030,N_9826,N_9870);
nand U10031 (N_10031,N_9854,N_9780);
or U10032 (N_10032,N_9823,N_9841);
nor U10033 (N_10033,N_9876,N_9914);
or U10034 (N_10034,N_9799,N_9812);
or U10035 (N_10035,N_9860,N_9808);
nor U10036 (N_10036,N_9900,N_9868);
nand U10037 (N_10037,N_9856,N_9870);
or U10038 (N_10038,N_9785,N_9776);
or U10039 (N_10039,N_9782,N_9831);
xor U10040 (N_10040,N_9836,N_9820);
xnor U10041 (N_10041,N_9765,N_9782);
nor U10042 (N_10042,N_9828,N_9908);
nand U10043 (N_10043,N_9907,N_9798);
and U10044 (N_10044,N_9799,N_9882);
nand U10045 (N_10045,N_9771,N_9862);
or U10046 (N_10046,N_9768,N_9845);
nor U10047 (N_10047,N_9897,N_9910);
and U10048 (N_10048,N_9775,N_9856);
nor U10049 (N_10049,N_9822,N_9774);
and U10050 (N_10050,N_9777,N_9866);
and U10051 (N_10051,N_9850,N_9888);
and U10052 (N_10052,N_9789,N_9915);
xnor U10053 (N_10053,N_9862,N_9872);
and U10054 (N_10054,N_9785,N_9775);
nand U10055 (N_10055,N_9847,N_9761);
and U10056 (N_10056,N_9829,N_9781);
or U10057 (N_10057,N_9899,N_9853);
nor U10058 (N_10058,N_9847,N_9865);
nand U10059 (N_10059,N_9794,N_9841);
nor U10060 (N_10060,N_9843,N_9833);
or U10061 (N_10061,N_9888,N_9812);
or U10062 (N_10062,N_9843,N_9855);
or U10063 (N_10063,N_9840,N_9847);
nand U10064 (N_10064,N_9815,N_9818);
nand U10065 (N_10065,N_9820,N_9775);
and U10066 (N_10066,N_9767,N_9789);
xnor U10067 (N_10067,N_9847,N_9856);
and U10068 (N_10068,N_9817,N_9915);
nor U10069 (N_10069,N_9764,N_9761);
and U10070 (N_10070,N_9889,N_9844);
or U10071 (N_10071,N_9889,N_9769);
nor U10072 (N_10072,N_9822,N_9814);
xor U10073 (N_10073,N_9894,N_9884);
nand U10074 (N_10074,N_9843,N_9897);
or U10075 (N_10075,N_9876,N_9898);
and U10076 (N_10076,N_9768,N_9862);
nand U10077 (N_10077,N_9778,N_9791);
nor U10078 (N_10078,N_9875,N_9796);
nor U10079 (N_10079,N_9848,N_9835);
nor U10080 (N_10080,N_10040,N_10019);
nor U10081 (N_10081,N_10049,N_10069);
nand U10082 (N_10082,N_10060,N_9950);
nor U10083 (N_10083,N_10072,N_9952);
nand U10084 (N_10084,N_9995,N_10048);
nand U10085 (N_10085,N_9956,N_9961);
and U10086 (N_10086,N_10028,N_9979);
or U10087 (N_10087,N_10007,N_9970);
nor U10088 (N_10088,N_9944,N_10018);
xnor U10089 (N_10089,N_10043,N_10075);
and U10090 (N_10090,N_10071,N_9964);
xor U10091 (N_10091,N_10032,N_9984);
and U10092 (N_10092,N_9997,N_9982);
and U10093 (N_10093,N_9926,N_9991);
or U10094 (N_10094,N_9987,N_10027);
and U10095 (N_10095,N_10057,N_10065);
nand U10096 (N_10096,N_10066,N_9980);
and U10097 (N_10097,N_9953,N_9974);
xor U10098 (N_10098,N_10005,N_9972);
nand U10099 (N_10099,N_10003,N_9983);
or U10100 (N_10100,N_9999,N_9966);
or U10101 (N_10101,N_9958,N_9955);
nand U10102 (N_10102,N_9985,N_10045);
nor U10103 (N_10103,N_9921,N_10058);
and U10104 (N_10104,N_10041,N_9965);
nor U10105 (N_10105,N_10033,N_9925);
nand U10106 (N_10106,N_9920,N_9927);
and U10107 (N_10107,N_10036,N_10010);
or U10108 (N_10108,N_10001,N_9948);
and U10109 (N_10109,N_9969,N_10056);
and U10110 (N_10110,N_10012,N_9954);
nand U10111 (N_10111,N_10026,N_10011);
nand U10112 (N_10112,N_9986,N_10064);
or U10113 (N_10113,N_10031,N_10039);
and U10114 (N_10114,N_10046,N_10047);
or U10115 (N_10115,N_9988,N_10023);
xnor U10116 (N_10116,N_10067,N_10059);
nor U10117 (N_10117,N_10015,N_9942);
or U10118 (N_10118,N_9947,N_10037);
or U10119 (N_10119,N_9932,N_10034);
and U10120 (N_10120,N_9949,N_9992);
nor U10121 (N_10121,N_10020,N_10073);
xor U10122 (N_10122,N_9924,N_10044);
and U10123 (N_10123,N_10013,N_10070);
nand U10124 (N_10124,N_10055,N_10035);
xnor U10125 (N_10125,N_10008,N_9945);
xor U10126 (N_10126,N_10021,N_10022);
nor U10127 (N_10127,N_9989,N_9922);
nor U10128 (N_10128,N_10077,N_10006);
nand U10129 (N_10129,N_9994,N_9993);
xor U10130 (N_10130,N_10042,N_10025);
nor U10131 (N_10131,N_9998,N_10061);
xnor U10132 (N_10132,N_9946,N_9938);
nor U10133 (N_10133,N_10038,N_10052);
or U10134 (N_10134,N_9931,N_9976);
nand U10135 (N_10135,N_9973,N_10068);
or U10136 (N_10136,N_10074,N_10079);
or U10137 (N_10137,N_10014,N_9975);
xor U10138 (N_10138,N_10029,N_9951);
nor U10139 (N_10139,N_10024,N_9941);
nand U10140 (N_10140,N_9960,N_9967);
nand U10141 (N_10141,N_10062,N_9930);
nor U10142 (N_10142,N_10063,N_9957);
nor U10143 (N_10143,N_9939,N_10054);
nor U10144 (N_10144,N_10030,N_10002);
or U10145 (N_10145,N_9934,N_9959);
xnor U10146 (N_10146,N_9937,N_10051);
xnor U10147 (N_10147,N_9990,N_9940);
or U10148 (N_10148,N_9962,N_9936);
xnor U10149 (N_10149,N_10053,N_10004);
xnor U10150 (N_10150,N_9928,N_10016);
nor U10151 (N_10151,N_9963,N_9933);
xor U10152 (N_10152,N_9929,N_10017);
and U10153 (N_10153,N_10076,N_10009);
xor U10154 (N_10154,N_10000,N_9943);
nand U10155 (N_10155,N_9971,N_9977);
and U10156 (N_10156,N_9996,N_9923);
or U10157 (N_10157,N_9935,N_9968);
or U10158 (N_10158,N_10078,N_9978);
nor U10159 (N_10159,N_10050,N_9981);
or U10160 (N_10160,N_9933,N_10040);
and U10161 (N_10161,N_10043,N_9998);
and U10162 (N_10162,N_10061,N_9965);
nand U10163 (N_10163,N_10002,N_10016);
and U10164 (N_10164,N_10013,N_10020);
nor U10165 (N_10165,N_10048,N_10011);
nor U10166 (N_10166,N_10035,N_10016);
xnor U10167 (N_10167,N_9929,N_10044);
nor U10168 (N_10168,N_9926,N_10015);
xor U10169 (N_10169,N_10052,N_9992);
nor U10170 (N_10170,N_10038,N_10029);
and U10171 (N_10171,N_9942,N_9930);
nor U10172 (N_10172,N_9948,N_9922);
nor U10173 (N_10173,N_10070,N_9994);
nor U10174 (N_10174,N_9926,N_9933);
or U10175 (N_10175,N_10079,N_9962);
or U10176 (N_10176,N_10065,N_10031);
nand U10177 (N_10177,N_10036,N_10020);
or U10178 (N_10178,N_10020,N_9973);
nor U10179 (N_10179,N_9988,N_9931);
and U10180 (N_10180,N_10018,N_9952);
nor U10181 (N_10181,N_10020,N_10017);
or U10182 (N_10182,N_10030,N_9927);
nor U10183 (N_10183,N_9998,N_9981);
nand U10184 (N_10184,N_10029,N_9926);
nand U10185 (N_10185,N_9967,N_9932);
and U10186 (N_10186,N_9995,N_10036);
nor U10187 (N_10187,N_10016,N_9946);
nand U10188 (N_10188,N_9943,N_10019);
or U10189 (N_10189,N_9938,N_9988);
nor U10190 (N_10190,N_10056,N_9937);
xnor U10191 (N_10191,N_10079,N_9996);
nor U10192 (N_10192,N_10011,N_10052);
and U10193 (N_10193,N_9964,N_9965);
or U10194 (N_10194,N_10010,N_10018);
xnor U10195 (N_10195,N_9932,N_10069);
xor U10196 (N_10196,N_10008,N_9997);
or U10197 (N_10197,N_10000,N_10025);
nor U10198 (N_10198,N_10018,N_10011);
and U10199 (N_10199,N_9927,N_10034);
nand U10200 (N_10200,N_9982,N_10003);
or U10201 (N_10201,N_10059,N_10046);
or U10202 (N_10202,N_10057,N_9941);
nand U10203 (N_10203,N_9954,N_9936);
nor U10204 (N_10204,N_10029,N_9923);
nand U10205 (N_10205,N_9964,N_10013);
and U10206 (N_10206,N_10065,N_9925);
nand U10207 (N_10207,N_10065,N_9949);
nor U10208 (N_10208,N_10003,N_10079);
nor U10209 (N_10209,N_10057,N_10015);
nand U10210 (N_10210,N_10039,N_9975);
nand U10211 (N_10211,N_9941,N_10003);
or U10212 (N_10212,N_9966,N_9997);
nor U10213 (N_10213,N_10050,N_9975);
or U10214 (N_10214,N_10061,N_9959);
nand U10215 (N_10215,N_10016,N_9920);
or U10216 (N_10216,N_9985,N_9922);
and U10217 (N_10217,N_9986,N_9948);
or U10218 (N_10218,N_10008,N_10070);
xnor U10219 (N_10219,N_9925,N_10051);
nand U10220 (N_10220,N_9948,N_10028);
xor U10221 (N_10221,N_9961,N_10059);
and U10222 (N_10222,N_10031,N_9920);
nand U10223 (N_10223,N_9955,N_10018);
nand U10224 (N_10224,N_9973,N_9951);
and U10225 (N_10225,N_10033,N_10012);
nand U10226 (N_10226,N_9964,N_10022);
nand U10227 (N_10227,N_10014,N_9961);
or U10228 (N_10228,N_10063,N_10030);
nand U10229 (N_10229,N_10034,N_9964);
or U10230 (N_10230,N_9947,N_9941);
or U10231 (N_10231,N_10043,N_9942);
xor U10232 (N_10232,N_9934,N_10014);
nor U10233 (N_10233,N_9988,N_9973);
and U10234 (N_10234,N_9974,N_10022);
or U10235 (N_10235,N_10064,N_10059);
and U10236 (N_10236,N_10055,N_10006);
and U10237 (N_10237,N_9958,N_10025);
nor U10238 (N_10238,N_10017,N_9948);
nand U10239 (N_10239,N_9984,N_10038);
or U10240 (N_10240,N_10213,N_10154);
or U10241 (N_10241,N_10084,N_10157);
xnor U10242 (N_10242,N_10117,N_10080);
or U10243 (N_10243,N_10097,N_10189);
nor U10244 (N_10244,N_10208,N_10099);
nor U10245 (N_10245,N_10125,N_10120);
nand U10246 (N_10246,N_10138,N_10134);
and U10247 (N_10247,N_10082,N_10209);
nor U10248 (N_10248,N_10215,N_10128);
nand U10249 (N_10249,N_10229,N_10110);
nand U10250 (N_10250,N_10218,N_10196);
and U10251 (N_10251,N_10149,N_10224);
nor U10252 (N_10252,N_10091,N_10101);
and U10253 (N_10253,N_10234,N_10094);
xor U10254 (N_10254,N_10226,N_10121);
nand U10255 (N_10255,N_10201,N_10181);
or U10256 (N_10256,N_10102,N_10177);
xnor U10257 (N_10257,N_10190,N_10187);
nor U10258 (N_10258,N_10142,N_10170);
xor U10259 (N_10259,N_10087,N_10211);
and U10260 (N_10260,N_10219,N_10186);
nand U10261 (N_10261,N_10090,N_10147);
or U10262 (N_10262,N_10086,N_10115);
nor U10263 (N_10263,N_10162,N_10096);
nor U10264 (N_10264,N_10216,N_10169);
nor U10265 (N_10265,N_10118,N_10106);
or U10266 (N_10266,N_10098,N_10206);
nand U10267 (N_10267,N_10100,N_10220);
nor U10268 (N_10268,N_10127,N_10114);
nand U10269 (N_10269,N_10155,N_10119);
nor U10270 (N_10270,N_10109,N_10131);
or U10271 (N_10271,N_10159,N_10140);
or U10272 (N_10272,N_10158,N_10133);
and U10273 (N_10273,N_10184,N_10167);
nand U10274 (N_10274,N_10231,N_10092);
or U10275 (N_10275,N_10217,N_10108);
nand U10276 (N_10276,N_10198,N_10145);
xor U10277 (N_10277,N_10228,N_10152);
and U10278 (N_10278,N_10126,N_10183);
nor U10279 (N_10279,N_10174,N_10212);
and U10280 (N_10280,N_10095,N_10093);
and U10281 (N_10281,N_10081,N_10227);
or U10282 (N_10282,N_10089,N_10180);
nor U10283 (N_10283,N_10136,N_10179);
nand U10284 (N_10284,N_10104,N_10171);
or U10285 (N_10285,N_10124,N_10210);
xor U10286 (N_10286,N_10137,N_10141);
and U10287 (N_10287,N_10151,N_10193);
or U10288 (N_10288,N_10085,N_10178);
and U10289 (N_10289,N_10176,N_10144);
nor U10290 (N_10290,N_10192,N_10200);
and U10291 (N_10291,N_10112,N_10088);
nor U10292 (N_10292,N_10175,N_10204);
and U10293 (N_10293,N_10153,N_10236);
nor U10294 (N_10294,N_10199,N_10168);
nor U10295 (N_10295,N_10230,N_10164);
and U10296 (N_10296,N_10232,N_10116);
nand U10297 (N_10297,N_10107,N_10203);
and U10298 (N_10298,N_10103,N_10222);
or U10299 (N_10299,N_10113,N_10235);
nor U10300 (N_10300,N_10237,N_10233);
and U10301 (N_10301,N_10132,N_10225);
or U10302 (N_10302,N_10139,N_10165);
nand U10303 (N_10303,N_10188,N_10123);
and U10304 (N_10304,N_10135,N_10130);
or U10305 (N_10305,N_10173,N_10161);
xnor U10306 (N_10306,N_10166,N_10195);
and U10307 (N_10307,N_10122,N_10238);
or U10308 (N_10308,N_10143,N_10221);
nand U10309 (N_10309,N_10223,N_10160);
or U10310 (N_10310,N_10191,N_10129);
nor U10311 (N_10311,N_10148,N_10146);
xnor U10312 (N_10312,N_10172,N_10194);
nand U10313 (N_10313,N_10185,N_10105);
xnor U10314 (N_10314,N_10083,N_10202);
or U10315 (N_10315,N_10239,N_10150);
and U10316 (N_10316,N_10182,N_10111);
and U10317 (N_10317,N_10214,N_10207);
nand U10318 (N_10318,N_10197,N_10205);
xor U10319 (N_10319,N_10156,N_10163);
or U10320 (N_10320,N_10100,N_10173);
nor U10321 (N_10321,N_10187,N_10143);
nand U10322 (N_10322,N_10102,N_10150);
and U10323 (N_10323,N_10161,N_10167);
or U10324 (N_10324,N_10101,N_10186);
or U10325 (N_10325,N_10124,N_10201);
nand U10326 (N_10326,N_10098,N_10191);
nor U10327 (N_10327,N_10122,N_10161);
nor U10328 (N_10328,N_10201,N_10095);
and U10329 (N_10329,N_10131,N_10176);
and U10330 (N_10330,N_10127,N_10101);
or U10331 (N_10331,N_10123,N_10115);
and U10332 (N_10332,N_10133,N_10196);
or U10333 (N_10333,N_10146,N_10104);
nand U10334 (N_10334,N_10156,N_10151);
xor U10335 (N_10335,N_10193,N_10150);
and U10336 (N_10336,N_10194,N_10164);
and U10337 (N_10337,N_10083,N_10093);
nor U10338 (N_10338,N_10171,N_10089);
or U10339 (N_10339,N_10119,N_10148);
or U10340 (N_10340,N_10203,N_10104);
xnor U10341 (N_10341,N_10202,N_10091);
and U10342 (N_10342,N_10180,N_10216);
or U10343 (N_10343,N_10158,N_10101);
and U10344 (N_10344,N_10092,N_10109);
and U10345 (N_10345,N_10117,N_10086);
or U10346 (N_10346,N_10237,N_10232);
nand U10347 (N_10347,N_10107,N_10208);
nor U10348 (N_10348,N_10164,N_10219);
or U10349 (N_10349,N_10095,N_10181);
and U10350 (N_10350,N_10089,N_10135);
and U10351 (N_10351,N_10173,N_10128);
and U10352 (N_10352,N_10204,N_10104);
and U10353 (N_10353,N_10170,N_10165);
nand U10354 (N_10354,N_10163,N_10127);
or U10355 (N_10355,N_10200,N_10150);
and U10356 (N_10356,N_10111,N_10120);
and U10357 (N_10357,N_10096,N_10088);
nand U10358 (N_10358,N_10179,N_10183);
nor U10359 (N_10359,N_10087,N_10149);
nor U10360 (N_10360,N_10114,N_10113);
nor U10361 (N_10361,N_10125,N_10229);
nor U10362 (N_10362,N_10122,N_10085);
xnor U10363 (N_10363,N_10091,N_10115);
and U10364 (N_10364,N_10090,N_10130);
nand U10365 (N_10365,N_10222,N_10230);
nand U10366 (N_10366,N_10207,N_10209);
nor U10367 (N_10367,N_10132,N_10147);
or U10368 (N_10368,N_10234,N_10166);
or U10369 (N_10369,N_10132,N_10198);
nand U10370 (N_10370,N_10212,N_10107);
nor U10371 (N_10371,N_10141,N_10181);
and U10372 (N_10372,N_10187,N_10191);
or U10373 (N_10373,N_10159,N_10206);
nand U10374 (N_10374,N_10143,N_10149);
xor U10375 (N_10375,N_10175,N_10215);
nand U10376 (N_10376,N_10184,N_10204);
nor U10377 (N_10377,N_10225,N_10128);
and U10378 (N_10378,N_10190,N_10105);
and U10379 (N_10379,N_10109,N_10151);
nor U10380 (N_10380,N_10116,N_10100);
xnor U10381 (N_10381,N_10184,N_10152);
xor U10382 (N_10382,N_10234,N_10175);
nor U10383 (N_10383,N_10192,N_10219);
nand U10384 (N_10384,N_10115,N_10195);
nand U10385 (N_10385,N_10137,N_10112);
nand U10386 (N_10386,N_10110,N_10182);
and U10387 (N_10387,N_10121,N_10217);
and U10388 (N_10388,N_10220,N_10198);
nand U10389 (N_10389,N_10211,N_10199);
and U10390 (N_10390,N_10131,N_10118);
nor U10391 (N_10391,N_10236,N_10224);
nand U10392 (N_10392,N_10151,N_10167);
and U10393 (N_10393,N_10131,N_10230);
nor U10394 (N_10394,N_10143,N_10163);
nor U10395 (N_10395,N_10120,N_10220);
and U10396 (N_10396,N_10084,N_10134);
xor U10397 (N_10397,N_10184,N_10217);
nand U10398 (N_10398,N_10158,N_10229);
xor U10399 (N_10399,N_10175,N_10093);
and U10400 (N_10400,N_10357,N_10367);
and U10401 (N_10401,N_10392,N_10395);
nand U10402 (N_10402,N_10240,N_10343);
nand U10403 (N_10403,N_10364,N_10253);
and U10404 (N_10404,N_10321,N_10247);
or U10405 (N_10405,N_10269,N_10280);
nand U10406 (N_10406,N_10287,N_10241);
or U10407 (N_10407,N_10389,N_10373);
xor U10408 (N_10408,N_10265,N_10385);
nand U10409 (N_10409,N_10335,N_10306);
xor U10410 (N_10410,N_10371,N_10297);
xnor U10411 (N_10411,N_10366,N_10249);
or U10412 (N_10412,N_10279,N_10301);
and U10413 (N_10413,N_10259,N_10333);
and U10414 (N_10414,N_10302,N_10368);
nor U10415 (N_10415,N_10284,N_10362);
nand U10416 (N_10416,N_10319,N_10363);
or U10417 (N_10417,N_10376,N_10260);
nor U10418 (N_10418,N_10350,N_10310);
nand U10419 (N_10419,N_10289,N_10274);
nor U10420 (N_10420,N_10331,N_10291);
nand U10421 (N_10421,N_10345,N_10262);
nand U10422 (N_10422,N_10340,N_10353);
xnor U10423 (N_10423,N_10281,N_10318);
and U10424 (N_10424,N_10391,N_10347);
nor U10425 (N_10425,N_10258,N_10316);
xnor U10426 (N_10426,N_10369,N_10377);
nand U10427 (N_10427,N_10380,N_10268);
or U10428 (N_10428,N_10365,N_10255);
nor U10429 (N_10429,N_10242,N_10267);
xnor U10430 (N_10430,N_10352,N_10244);
nor U10431 (N_10431,N_10397,N_10320);
and U10432 (N_10432,N_10341,N_10271);
or U10433 (N_10433,N_10254,N_10325);
xnor U10434 (N_10434,N_10248,N_10379);
or U10435 (N_10435,N_10266,N_10322);
or U10436 (N_10436,N_10273,N_10337);
nand U10437 (N_10437,N_10275,N_10312);
nand U10438 (N_10438,N_10381,N_10382);
xnor U10439 (N_10439,N_10243,N_10272);
and U10440 (N_10440,N_10360,N_10278);
and U10441 (N_10441,N_10390,N_10326);
xor U10442 (N_10442,N_10388,N_10286);
or U10443 (N_10443,N_10256,N_10323);
nor U10444 (N_10444,N_10317,N_10394);
nor U10445 (N_10445,N_10358,N_10384);
nand U10446 (N_10446,N_10372,N_10299);
xor U10447 (N_10447,N_10300,N_10378);
nand U10448 (N_10448,N_10387,N_10339);
nand U10449 (N_10449,N_10294,N_10251);
or U10450 (N_10450,N_10313,N_10303);
or U10451 (N_10451,N_10257,N_10309);
and U10452 (N_10452,N_10295,N_10315);
and U10453 (N_10453,N_10370,N_10305);
nand U10454 (N_10454,N_10328,N_10330);
xnor U10455 (N_10455,N_10307,N_10288);
xnor U10456 (N_10456,N_10332,N_10329);
nand U10457 (N_10457,N_10349,N_10393);
nand U10458 (N_10458,N_10375,N_10324);
nand U10459 (N_10459,N_10277,N_10263);
or U10460 (N_10460,N_10264,N_10383);
xor U10461 (N_10461,N_10270,N_10276);
and U10462 (N_10462,N_10292,N_10308);
and U10463 (N_10463,N_10252,N_10304);
or U10464 (N_10464,N_10354,N_10336);
nand U10465 (N_10465,N_10355,N_10327);
nand U10466 (N_10466,N_10361,N_10396);
and U10467 (N_10467,N_10398,N_10344);
nor U10468 (N_10468,N_10296,N_10290);
or U10469 (N_10469,N_10399,N_10374);
or U10470 (N_10470,N_10334,N_10298);
nand U10471 (N_10471,N_10311,N_10386);
nor U10472 (N_10472,N_10293,N_10282);
and U10473 (N_10473,N_10348,N_10314);
and U10474 (N_10474,N_10261,N_10356);
nor U10475 (N_10475,N_10246,N_10342);
or U10476 (N_10476,N_10359,N_10285);
nand U10477 (N_10477,N_10338,N_10351);
and U10478 (N_10478,N_10346,N_10283);
nand U10479 (N_10479,N_10245,N_10250);
and U10480 (N_10480,N_10265,N_10311);
and U10481 (N_10481,N_10254,N_10286);
nor U10482 (N_10482,N_10247,N_10371);
nor U10483 (N_10483,N_10244,N_10295);
or U10484 (N_10484,N_10333,N_10340);
and U10485 (N_10485,N_10322,N_10279);
and U10486 (N_10486,N_10375,N_10267);
or U10487 (N_10487,N_10345,N_10265);
nand U10488 (N_10488,N_10391,N_10339);
nor U10489 (N_10489,N_10293,N_10360);
nand U10490 (N_10490,N_10381,N_10251);
xnor U10491 (N_10491,N_10319,N_10260);
nand U10492 (N_10492,N_10353,N_10330);
nand U10493 (N_10493,N_10248,N_10381);
nand U10494 (N_10494,N_10327,N_10370);
or U10495 (N_10495,N_10305,N_10336);
xnor U10496 (N_10496,N_10376,N_10243);
nand U10497 (N_10497,N_10282,N_10367);
xnor U10498 (N_10498,N_10389,N_10282);
xor U10499 (N_10499,N_10381,N_10336);
and U10500 (N_10500,N_10260,N_10254);
nand U10501 (N_10501,N_10387,N_10351);
or U10502 (N_10502,N_10317,N_10282);
nor U10503 (N_10503,N_10326,N_10289);
and U10504 (N_10504,N_10352,N_10398);
nand U10505 (N_10505,N_10293,N_10377);
nand U10506 (N_10506,N_10264,N_10268);
xnor U10507 (N_10507,N_10241,N_10376);
nor U10508 (N_10508,N_10377,N_10330);
or U10509 (N_10509,N_10323,N_10342);
nor U10510 (N_10510,N_10276,N_10321);
or U10511 (N_10511,N_10292,N_10386);
or U10512 (N_10512,N_10388,N_10279);
nand U10513 (N_10513,N_10399,N_10300);
nand U10514 (N_10514,N_10374,N_10351);
nor U10515 (N_10515,N_10246,N_10262);
nor U10516 (N_10516,N_10395,N_10250);
nand U10517 (N_10517,N_10277,N_10254);
and U10518 (N_10518,N_10360,N_10260);
and U10519 (N_10519,N_10278,N_10307);
nand U10520 (N_10520,N_10267,N_10393);
or U10521 (N_10521,N_10281,N_10333);
nor U10522 (N_10522,N_10340,N_10387);
and U10523 (N_10523,N_10275,N_10317);
nor U10524 (N_10524,N_10294,N_10244);
nand U10525 (N_10525,N_10281,N_10397);
or U10526 (N_10526,N_10242,N_10250);
or U10527 (N_10527,N_10261,N_10351);
and U10528 (N_10528,N_10394,N_10387);
or U10529 (N_10529,N_10287,N_10361);
and U10530 (N_10530,N_10244,N_10382);
or U10531 (N_10531,N_10263,N_10313);
nor U10532 (N_10532,N_10263,N_10366);
nor U10533 (N_10533,N_10392,N_10323);
and U10534 (N_10534,N_10395,N_10382);
or U10535 (N_10535,N_10251,N_10362);
or U10536 (N_10536,N_10363,N_10327);
and U10537 (N_10537,N_10303,N_10278);
and U10538 (N_10538,N_10350,N_10383);
or U10539 (N_10539,N_10244,N_10258);
or U10540 (N_10540,N_10276,N_10268);
xnor U10541 (N_10541,N_10289,N_10330);
xnor U10542 (N_10542,N_10329,N_10389);
nor U10543 (N_10543,N_10363,N_10368);
and U10544 (N_10544,N_10287,N_10373);
nand U10545 (N_10545,N_10286,N_10367);
or U10546 (N_10546,N_10244,N_10287);
and U10547 (N_10547,N_10379,N_10300);
nand U10548 (N_10548,N_10294,N_10344);
and U10549 (N_10549,N_10244,N_10325);
or U10550 (N_10550,N_10276,N_10304);
nor U10551 (N_10551,N_10299,N_10308);
nand U10552 (N_10552,N_10373,N_10350);
nor U10553 (N_10553,N_10297,N_10377);
and U10554 (N_10554,N_10322,N_10335);
nand U10555 (N_10555,N_10335,N_10385);
and U10556 (N_10556,N_10294,N_10307);
nand U10557 (N_10557,N_10329,N_10325);
or U10558 (N_10558,N_10240,N_10281);
and U10559 (N_10559,N_10376,N_10250);
or U10560 (N_10560,N_10556,N_10483);
and U10561 (N_10561,N_10451,N_10490);
nand U10562 (N_10562,N_10518,N_10533);
and U10563 (N_10563,N_10472,N_10406);
nand U10564 (N_10564,N_10548,N_10425);
or U10565 (N_10565,N_10487,N_10413);
nor U10566 (N_10566,N_10522,N_10508);
nand U10567 (N_10567,N_10496,N_10466);
nor U10568 (N_10568,N_10516,N_10478);
or U10569 (N_10569,N_10411,N_10550);
nor U10570 (N_10570,N_10510,N_10527);
or U10571 (N_10571,N_10464,N_10498);
and U10572 (N_10572,N_10538,N_10467);
nor U10573 (N_10573,N_10404,N_10446);
or U10574 (N_10574,N_10555,N_10485);
and U10575 (N_10575,N_10499,N_10403);
or U10576 (N_10576,N_10501,N_10428);
nand U10577 (N_10577,N_10427,N_10559);
xnor U10578 (N_10578,N_10459,N_10491);
and U10579 (N_10579,N_10494,N_10408);
xor U10580 (N_10580,N_10443,N_10462);
nand U10581 (N_10581,N_10468,N_10414);
or U10582 (N_10582,N_10455,N_10445);
and U10583 (N_10583,N_10471,N_10535);
nand U10584 (N_10584,N_10447,N_10405);
or U10585 (N_10585,N_10539,N_10452);
xnor U10586 (N_10586,N_10541,N_10409);
nand U10587 (N_10587,N_10453,N_10509);
xnor U10588 (N_10588,N_10407,N_10440);
or U10589 (N_10589,N_10422,N_10400);
and U10590 (N_10590,N_10461,N_10545);
nor U10591 (N_10591,N_10492,N_10517);
nand U10592 (N_10592,N_10526,N_10419);
and U10593 (N_10593,N_10540,N_10528);
nor U10594 (N_10594,N_10512,N_10434);
nand U10595 (N_10595,N_10534,N_10506);
nor U10596 (N_10596,N_10423,N_10463);
and U10597 (N_10597,N_10431,N_10514);
nor U10598 (N_10598,N_10531,N_10465);
or U10599 (N_10599,N_10544,N_10450);
nor U10600 (N_10600,N_10417,N_10457);
nor U10601 (N_10601,N_10504,N_10481);
and U10602 (N_10602,N_10458,N_10449);
xnor U10603 (N_10603,N_10418,N_10442);
and U10604 (N_10604,N_10489,N_10505);
nand U10605 (N_10605,N_10549,N_10437);
nor U10606 (N_10606,N_10537,N_10547);
nand U10607 (N_10607,N_10477,N_10523);
nand U10608 (N_10608,N_10495,N_10553);
nor U10609 (N_10609,N_10470,N_10476);
or U10610 (N_10610,N_10441,N_10554);
or U10611 (N_10611,N_10519,N_10435);
nor U10612 (N_10612,N_10436,N_10486);
nand U10613 (N_10613,N_10546,N_10480);
and U10614 (N_10614,N_10444,N_10421);
or U10615 (N_10615,N_10557,N_10497);
nand U10616 (N_10616,N_10503,N_10529);
or U10617 (N_10617,N_10484,N_10429);
nand U10618 (N_10618,N_10460,N_10524);
or U10619 (N_10619,N_10507,N_10488);
and U10620 (N_10620,N_10433,N_10530);
and U10621 (N_10621,N_10543,N_10402);
xor U10622 (N_10622,N_10479,N_10420);
and U10623 (N_10623,N_10511,N_10416);
or U10624 (N_10624,N_10410,N_10401);
xor U10625 (N_10625,N_10520,N_10454);
and U10626 (N_10626,N_10448,N_10439);
and U10627 (N_10627,N_10515,N_10551);
and U10628 (N_10628,N_10424,N_10475);
xor U10629 (N_10629,N_10513,N_10432);
nor U10630 (N_10630,N_10525,N_10521);
or U10631 (N_10631,N_10426,N_10415);
nor U10632 (N_10632,N_10456,N_10482);
nor U10633 (N_10633,N_10502,N_10469);
nand U10634 (N_10634,N_10493,N_10542);
or U10635 (N_10635,N_10532,N_10438);
xor U10636 (N_10636,N_10412,N_10558);
and U10637 (N_10637,N_10500,N_10473);
nand U10638 (N_10638,N_10552,N_10536);
nand U10639 (N_10639,N_10474,N_10430);
nand U10640 (N_10640,N_10440,N_10441);
or U10641 (N_10641,N_10412,N_10437);
and U10642 (N_10642,N_10461,N_10401);
xor U10643 (N_10643,N_10435,N_10490);
nor U10644 (N_10644,N_10446,N_10472);
nor U10645 (N_10645,N_10421,N_10540);
and U10646 (N_10646,N_10438,N_10496);
and U10647 (N_10647,N_10531,N_10510);
or U10648 (N_10648,N_10532,N_10482);
nor U10649 (N_10649,N_10488,N_10442);
nand U10650 (N_10650,N_10444,N_10448);
nand U10651 (N_10651,N_10498,N_10516);
nor U10652 (N_10652,N_10513,N_10524);
nor U10653 (N_10653,N_10529,N_10502);
and U10654 (N_10654,N_10454,N_10554);
or U10655 (N_10655,N_10482,N_10554);
nand U10656 (N_10656,N_10493,N_10528);
or U10657 (N_10657,N_10476,N_10467);
or U10658 (N_10658,N_10540,N_10544);
nor U10659 (N_10659,N_10504,N_10408);
nand U10660 (N_10660,N_10446,N_10468);
xor U10661 (N_10661,N_10535,N_10448);
nand U10662 (N_10662,N_10443,N_10497);
nand U10663 (N_10663,N_10465,N_10429);
and U10664 (N_10664,N_10406,N_10551);
and U10665 (N_10665,N_10418,N_10556);
and U10666 (N_10666,N_10420,N_10467);
nor U10667 (N_10667,N_10474,N_10492);
and U10668 (N_10668,N_10520,N_10548);
nand U10669 (N_10669,N_10527,N_10472);
or U10670 (N_10670,N_10497,N_10436);
and U10671 (N_10671,N_10425,N_10546);
and U10672 (N_10672,N_10480,N_10465);
or U10673 (N_10673,N_10504,N_10534);
nand U10674 (N_10674,N_10534,N_10520);
or U10675 (N_10675,N_10514,N_10536);
nor U10676 (N_10676,N_10559,N_10426);
xor U10677 (N_10677,N_10455,N_10558);
or U10678 (N_10678,N_10464,N_10460);
nor U10679 (N_10679,N_10450,N_10406);
and U10680 (N_10680,N_10464,N_10441);
nand U10681 (N_10681,N_10552,N_10521);
and U10682 (N_10682,N_10549,N_10530);
nand U10683 (N_10683,N_10553,N_10404);
nand U10684 (N_10684,N_10400,N_10427);
or U10685 (N_10685,N_10558,N_10550);
or U10686 (N_10686,N_10449,N_10483);
nor U10687 (N_10687,N_10480,N_10508);
and U10688 (N_10688,N_10456,N_10421);
or U10689 (N_10689,N_10471,N_10465);
or U10690 (N_10690,N_10515,N_10432);
or U10691 (N_10691,N_10434,N_10487);
and U10692 (N_10692,N_10541,N_10509);
and U10693 (N_10693,N_10504,N_10469);
xor U10694 (N_10694,N_10479,N_10542);
nand U10695 (N_10695,N_10498,N_10509);
nand U10696 (N_10696,N_10549,N_10472);
nand U10697 (N_10697,N_10490,N_10516);
nor U10698 (N_10698,N_10494,N_10435);
nand U10699 (N_10699,N_10475,N_10419);
or U10700 (N_10700,N_10467,N_10423);
and U10701 (N_10701,N_10457,N_10446);
and U10702 (N_10702,N_10550,N_10513);
and U10703 (N_10703,N_10507,N_10454);
and U10704 (N_10704,N_10508,N_10502);
and U10705 (N_10705,N_10460,N_10481);
nand U10706 (N_10706,N_10538,N_10507);
nor U10707 (N_10707,N_10514,N_10423);
and U10708 (N_10708,N_10488,N_10484);
xnor U10709 (N_10709,N_10507,N_10555);
and U10710 (N_10710,N_10449,N_10526);
and U10711 (N_10711,N_10427,N_10448);
nor U10712 (N_10712,N_10512,N_10410);
xor U10713 (N_10713,N_10546,N_10469);
or U10714 (N_10714,N_10410,N_10402);
or U10715 (N_10715,N_10423,N_10502);
nand U10716 (N_10716,N_10421,N_10525);
or U10717 (N_10717,N_10411,N_10450);
nand U10718 (N_10718,N_10515,N_10531);
xnor U10719 (N_10719,N_10484,N_10445);
or U10720 (N_10720,N_10676,N_10610);
and U10721 (N_10721,N_10650,N_10707);
nor U10722 (N_10722,N_10566,N_10624);
nor U10723 (N_10723,N_10597,N_10705);
nor U10724 (N_10724,N_10593,N_10651);
xor U10725 (N_10725,N_10679,N_10690);
nor U10726 (N_10726,N_10632,N_10659);
and U10727 (N_10727,N_10592,N_10681);
and U10728 (N_10728,N_10614,N_10661);
and U10729 (N_10729,N_10574,N_10668);
nand U10730 (N_10730,N_10584,N_10633);
nor U10731 (N_10731,N_10570,N_10649);
and U10732 (N_10732,N_10569,N_10629);
nor U10733 (N_10733,N_10682,N_10615);
and U10734 (N_10734,N_10577,N_10667);
xnor U10735 (N_10735,N_10670,N_10710);
and U10736 (N_10736,N_10709,N_10561);
or U10737 (N_10737,N_10598,N_10712);
and U10738 (N_10738,N_10616,N_10563);
nor U10739 (N_10739,N_10646,N_10700);
nor U10740 (N_10740,N_10639,N_10701);
nand U10741 (N_10741,N_10715,N_10609);
nor U10742 (N_10742,N_10613,N_10602);
nand U10743 (N_10743,N_10631,N_10608);
or U10744 (N_10744,N_10630,N_10678);
nor U10745 (N_10745,N_10666,N_10583);
or U10746 (N_10746,N_10687,N_10675);
nand U10747 (N_10747,N_10665,N_10594);
and U10748 (N_10748,N_10595,N_10647);
or U10749 (N_10749,N_10622,N_10662);
and U10750 (N_10750,N_10626,N_10587);
or U10751 (N_10751,N_10689,N_10601);
nand U10752 (N_10752,N_10605,N_10699);
xnor U10753 (N_10753,N_10644,N_10708);
nand U10754 (N_10754,N_10620,N_10655);
nor U10755 (N_10755,N_10713,N_10657);
and U10756 (N_10756,N_10565,N_10664);
xnor U10757 (N_10757,N_10562,N_10617);
and U10758 (N_10758,N_10599,N_10686);
or U10759 (N_10759,N_10645,N_10697);
and U10760 (N_10760,N_10704,N_10685);
or U10761 (N_10761,N_10693,N_10706);
and U10762 (N_10762,N_10684,N_10656);
or U10763 (N_10763,N_10611,N_10621);
or U10764 (N_10764,N_10692,N_10702);
and U10765 (N_10765,N_10683,N_10717);
nor U10766 (N_10766,N_10674,N_10603);
and U10767 (N_10767,N_10586,N_10677);
and U10768 (N_10768,N_10625,N_10694);
or U10769 (N_10769,N_10658,N_10591);
and U10770 (N_10770,N_10582,N_10568);
nor U10771 (N_10771,N_10572,N_10579);
nand U10772 (N_10772,N_10640,N_10634);
xor U10773 (N_10773,N_10688,N_10652);
xnor U10774 (N_10774,N_10627,N_10718);
xor U10775 (N_10775,N_10671,N_10576);
nand U10776 (N_10776,N_10567,N_10636);
or U10777 (N_10777,N_10635,N_10672);
nand U10778 (N_10778,N_10653,N_10691);
xor U10779 (N_10779,N_10711,N_10641);
or U10780 (N_10780,N_10606,N_10714);
and U10781 (N_10781,N_10607,N_10703);
nor U10782 (N_10782,N_10589,N_10560);
nor U10783 (N_10783,N_10719,N_10600);
nor U10784 (N_10784,N_10673,N_10680);
nor U10785 (N_10785,N_10573,N_10695);
nand U10786 (N_10786,N_10604,N_10648);
or U10787 (N_10787,N_10575,N_10642);
nand U10788 (N_10788,N_10623,N_10696);
and U10789 (N_10789,N_10564,N_10580);
nand U10790 (N_10790,N_10628,N_10663);
or U10791 (N_10791,N_10669,N_10618);
nor U10792 (N_10792,N_10578,N_10612);
nor U10793 (N_10793,N_10638,N_10596);
and U10794 (N_10794,N_10585,N_10637);
or U10795 (N_10795,N_10588,N_10571);
nand U10796 (N_10796,N_10716,N_10619);
nor U10797 (N_10797,N_10581,N_10654);
and U10798 (N_10798,N_10660,N_10698);
nand U10799 (N_10799,N_10643,N_10590);
nand U10800 (N_10800,N_10662,N_10714);
and U10801 (N_10801,N_10561,N_10670);
nand U10802 (N_10802,N_10619,N_10577);
nor U10803 (N_10803,N_10612,N_10670);
or U10804 (N_10804,N_10661,N_10564);
nor U10805 (N_10805,N_10564,N_10691);
xor U10806 (N_10806,N_10691,N_10574);
nor U10807 (N_10807,N_10622,N_10604);
nand U10808 (N_10808,N_10713,N_10593);
nor U10809 (N_10809,N_10637,N_10619);
and U10810 (N_10810,N_10682,N_10713);
and U10811 (N_10811,N_10614,N_10576);
and U10812 (N_10812,N_10705,N_10590);
and U10813 (N_10813,N_10576,N_10645);
and U10814 (N_10814,N_10566,N_10595);
or U10815 (N_10815,N_10644,N_10681);
xnor U10816 (N_10816,N_10662,N_10638);
or U10817 (N_10817,N_10622,N_10701);
nor U10818 (N_10818,N_10656,N_10577);
nand U10819 (N_10819,N_10631,N_10681);
nand U10820 (N_10820,N_10640,N_10689);
xnor U10821 (N_10821,N_10566,N_10590);
or U10822 (N_10822,N_10633,N_10714);
and U10823 (N_10823,N_10589,N_10635);
or U10824 (N_10824,N_10673,N_10716);
nor U10825 (N_10825,N_10693,N_10695);
or U10826 (N_10826,N_10710,N_10631);
and U10827 (N_10827,N_10645,N_10607);
nor U10828 (N_10828,N_10714,N_10646);
nand U10829 (N_10829,N_10615,N_10703);
or U10830 (N_10830,N_10612,N_10584);
nand U10831 (N_10831,N_10632,N_10627);
nor U10832 (N_10832,N_10711,N_10696);
nand U10833 (N_10833,N_10653,N_10679);
nor U10834 (N_10834,N_10690,N_10644);
or U10835 (N_10835,N_10689,N_10586);
and U10836 (N_10836,N_10593,N_10582);
nor U10837 (N_10837,N_10697,N_10626);
and U10838 (N_10838,N_10686,N_10716);
xnor U10839 (N_10839,N_10641,N_10597);
nor U10840 (N_10840,N_10562,N_10678);
nor U10841 (N_10841,N_10586,N_10657);
nor U10842 (N_10842,N_10704,N_10599);
nand U10843 (N_10843,N_10688,N_10689);
xnor U10844 (N_10844,N_10652,N_10638);
nor U10845 (N_10845,N_10634,N_10608);
or U10846 (N_10846,N_10595,N_10706);
nor U10847 (N_10847,N_10560,N_10706);
xor U10848 (N_10848,N_10562,N_10666);
or U10849 (N_10849,N_10563,N_10618);
nor U10850 (N_10850,N_10682,N_10573);
nor U10851 (N_10851,N_10664,N_10595);
nor U10852 (N_10852,N_10580,N_10691);
xnor U10853 (N_10853,N_10704,N_10640);
nor U10854 (N_10854,N_10668,N_10635);
and U10855 (N_10855,N_10710,N_10698);
and U10856 (N_10856,N_10637,N_10646);
xor U10857 (N_10857,N_10604,N_10621);
nor U10858 (N_10858,N_10564,N_10680);
nor U10859 (N_10859,N_10601,N_10565);
nor U10860 (N_10860,N_10570,N_10618);
and U10861 (N_10861,N_10603,N_10668);
and U10862 (N_10862,N_10615,N_10693);
nand U10863 (N_10863,N_10596,N_10617);
nand U10864 (N_10864,N_10646,N_10594);
nor U10865 (N_10865,N_10694,N_10640);
or U10866 (N_10866,N_10595,N_10650);
and U10867 (N_10867,N_10620,N_10695);
xnor U10868 (N_10868,N_10581,N_10615);
and U10869 (N_10869,N_10560,N_10623);
xor U10870 (N_10870,N_10662,N_10716);
or U10871 (N_10871,N_10708,N_10571);
nor U10872 (N_10872,N_10679,N_10590);
nand U10873 (N_10873,N_10640,N_10684);
or U10874 (N_10874,N_10692,N_10640);
and U10875 (N_10875,N_10707,N_10668);
xor U10876 (N_10876,N_10571,N_10578);
or U10877 (N_10877,N_10702,N_10627);
and U10878 (N_10878,N_10680,N_10611);
nand U10879 (N_10879,N_10701,N_10605);
or U10880 (N_10880,N_10834,N_10727);
nand U10881 (N_10881,N_10763,N_10873);
xor U10882 (N_10882,N_10786,N_10826);
nand U10883 (N_10883,N_10850,N_10722);
nand U10884 (N_10884,N_10764,N_10724);
nand U10885 (N_10885,N_10792,N_10747);
or U10886 (N_10886,N_10781,N_10846);
nand U10887 (N_10887,N_10867,N_10877);
and U10888 (N_10888,N_10729,N_10755);
nor U10889 (N_10889,N_10778,N_10738);
and U10890 (N_10890,N_10878,N_10825);
or U10891 (N_10891,N_10773,N_10766);
nand U10892 (N_10892,N_10734,N_10869);
and U10893 (N_10893,N_10720,N_10820);
or U10894 (N_10894,N_10762,N_10868);
or U10895 (N_10895,N_10783,N_10828);
xor U10896 (N_10896,N_10833,N_10874);
or U10897 (N_10897,N_10797,N_10802);
and U10898 (N_10898,N_10721,N_10823);
nor U10899 (N_10899,N_10803,N_10839);
and U10900 (N_10900,N_10723,N_10757);
and U10901 (N_10901,N_10875,N_10799);
nor U10902 (N_10902,N_10849,N_10739);
or U10903 (N_10903,N_10837,N_10855);
nor U10904 (N_10904,N_10819,N_10841);
and U10905 (N_10905,N_10812,N_10743);
or U10906 (N_10906,N_10827,N_10775);
or U10907 (N_10907,N_10821,N_10761);
nand U10908 (N_10908,N_10787,N_10838);
and U10909 (N_10909,N_10806,N_10798);
and U10910 (N_10910,N_10816,N_10831);
nor U10911 (N_10911,N_10733,N_10771);
nand U10912 (N_10912,N_10836,N_10796);
nand U10913 (N_10913,N_10843,N_10860);
nand U10914 (N_10914,N_10769,N_10845);
nor U10915 (N_10915,N_10815,N_10817);
nor U10916 (N_10916,N_10864,N_10751);
xnor U10917 (N_10917,N_10780,N_10732);
nand U10918 (N_10918,N_10726,N_10741);
nor U10919 (N_10919,N_10848,N_10744);
nand U10920 (N_10920,N_10731,N_10750);
or U10921 (N_10921,N_10840,N_10788);
nand U10922 (N_10922,N_10735,N_10805);
xnor U10923 (N_10923,N_10760,N_10772);
nor U10924 (N_10924,N_10856,N_10814);
nand U10925 (N_10925,N_10851,N_10862);
xnor U10926 (N_10926,N_10746,N_10765);
or U10927 (N_10927,N_10804,N_10793);
and U10928 (N_10928,N_10811,N_10777);
and U10929 (N_10929,N_10736,N_10871);
and U10930 (N_10930,N_10876,N_10865);
xnor U10931 (N_10931,N_10872,N_10794);
nor U10932 (N_10932,N_10842,N_10774);
xor U10933 (N_10933,N_10756,N_10776);
xor U10934 (N_10934,N_10742,N_10809);
xor U10935 (N_10935,N_10847,N_10844);
nor U10936 (N_10936,N_10835,N_10822);
and U10937 (N_10937,N_10866,N_10779);
and U10938 (N_10938,N_10784,N_10768);
or U10939 (N_10939,N_10863,N_10759);
or U10940 (N_10940,N_10859,N_10810);
or U10941 (N_10941,N_10824,N_10753);
and U10942 (N_10942,N_10879,N_10818);
nand U10943 (N_10943,N_10754,N_10807);
or U10944 (N_10944,N_10782,N_10758);
and U10945 (N_10945,N_10857,N_10740);
or U10946 (N_10946,N_10832,N_10748);
and U10947 (N_10947,N_10767,N_10745);
or U10948 (N_10948,N_10728,N_10791);
nand U10949 (N_10949,N_10854,N_10785);
nand U10950 (N_10950,N_10749,N_10853);
xnor U10951 (N_10951,N_10800,N_10737);
nand U10952 (N_10952,N_10813,N_10808);
nor U10953 (N_10953,N_10752,N_10830);
or U10954 (N_10954,N_10730,N_10790);
or U10955 (N_10955,N_10861,N_10725);
nor U10956 (N_10956,N_10829,N_10852);
and U10957 (N_10957,N_10795,N_10801);
and U10958 (N_10958,N_10789,N_10858);
nor U10959 (N_10959,N_10870,N_10770);
xor U10960 (N_10960,N_10800,N_10830);
xor U10961 (N_10961,N_10802,N_10760);
nand U10962 (N_10962,N_10803,N_10765);
and U10963 (N_10963,N_10868,N_10852);
nand U10964 (N_10964,N_10852,N_10846);
and U10965 (N_10965,N_10732,N_10749);
xor U10966 (N_10966,N_10753,N_10749);
and U10967 (N_10967,N_10733,N_10837);
or U10968 (N_10968,N_10745,N_10793);
and U10969 (N_10969,N_10840,N_10739);
nor U10970 (N_10970,N_10785,N_10736);
and U10971 (N_10971,N_10768,N_10832);
and U10972 (N_10972,N_10802,N_10824);
or U10973 (N_10973,N_10805,N_10743);
xor U10974 (N_10974,N_10844,N_10788);
and U10975 (N_10975,N_10825,N_10849);
nand U10976 (N_10976,N_10815,N_10721);
and U10977 (N_10977,N_10762,N_10851);
and U10978 (N_10978,N_10871,N_10758);
nand U10979 (N_10979,N_10807,N_10789);
and U10980 (N_10980,N_10821,N_10721);
nand U10981 (N_10981,N_10749,N_10862);
nand U10982 (N_10982,N_10741,N_10745);
nor U10983 (N_10983,N_10835,N_10764);
nand U10984 (N_10984,N_10861,N_10850);
xnor U10985 (N_10985,N_10818,N_10810);
nand U10986 (N_10986,N_10837,N_10866);
or U10987 (N_10987,N_10753,N_10780);
nor U10988 (N_10988,N_10742,N_10864);
and U10989 (N_10989,N_10875,N_10778);
nand U10990 (N_10990,N_10866,N_10764);
or U10991 (N_10991,N_10819,N_10774);
nor U10992 (N_10992,N_10873,N_10734);
and U10993 (N_10993,N_10724,N_10872);
nor U10994 (N_10994,N_10725,N_10781);
nor U10995 (N_10995,N_10777,N_10774);
nand U10996 (N_10996,N_10818,N_10752);
and U10997 (N_10997,N_10822,N_10840);
and U10998 (N_10998,N_10728,N_10800);
nand U10999 (N_10999,N_10835,N_10831);
nand U11000 (N_11000,N_10877,N_10757);
nand U11001 (N_11001,N_10799,N_10820);
nor U11002 (N_11002,N_10845,N_10801);
nor U11003 (N_11003,N_10875,N_10849);
and U11004 (N_11004,N_10872,N_10858);
or U11005 (N_11005,N_10742,N_10844);
nand U11006 (N_11006,N_10803,N_10727);
or U11007 (N_11007,N_10791,N_10720);
and U11008 (N_11008,N_10828,N_10737);
and U11009 (N_11009,N_10729,N_10773);
nor U11010 (N_11010,N_10851,N_10790);
and U11011 (N_11011,N_10821,N_10776);
or U11012 (N_11012,N_10815,N_10784);
or U11013 (N_11013,N_10740,N_10750);
nand U11014 (N_11014,N_10803,N_10771);
nand U11015 (N_11015,N_10839,N_10810);
and U11016 (N_11016,N_10747,N_10728);
and U11017 (N_11017,N_10736,N_10877);
nor U11018 (N_11018,N_10790,N_10761);
nor U11019 (N_11019,N_10875,N_10728);
nor U11020 (N_11020,N_10756,N_10767);
nor U11021 (N_11021,N_10807,N_10794);
and U11022 (N_11022,N_10824,N_10825);
nand U11023 (N_11023,N_10816,N_10734);
xor U11024 (N_11024,N_10769,N_10810);
nor U11025 (N_11025,N_10815,N_10874);
and U11026 (N_11026,N_10748,N_10742);
or U11027 (N_11027,N_10750,N_10732);
nand U11028 (N_11028,N_10725,N_10789);
or U11029 (N_11029,N_10807,N_10877);
nand U11030 (N_11030,N_10740,N_10741);
and U11031 (N_11031,N_10854,N_10759);
nor U11032 (N_11032,N_10760,N_10759);
xor U11033 (N_11033,N_10734,N_10868);
nor U11034 (N_11034,N_10720,N_10799);
and U11035 (N_11035,N_10736,N_10727);
xor U11036 (N_11036,N_10839,N_10813);
nand U11037 (N_11037,N_10809,N_10730);
nand U11038 (N_11038,N_10724,N_10744);
nor U11039 (N_11039,N_10791,N_10810);
or U11040 (N_11040,N_10889,N_10959);
xnor U11041 (N_11041,N_10973,N_10963);
nor U11042 (N_11042,N_11026,N_10992);
and U11043 (N_11043,N_10993,N_10900);
and U11044 (N_11044,N_10896,N_10933);
and U11045 (N_11045,N_10955,N_10936);
or U11046 (N_11046,N_10880,N_10966);
xnor U11047 (N_11047,N_10971,N_10989);
nand U11048 (N_11048,N_10906,N_11025);
or U11049 (N_11049,N_10912,N_11008);
or U11050 (N_11050,N_10930,N_11014);
nand U11051 (N_11051,N_10942,N_11019);
or U11052 (N_11052,N_10965,N_10911);
xor U11053 (N_11053,N_10988,N_10901);
nand U11054 (N_11054,N_10949,N_10970);
nor U11055 (N_11055,N_10897,N_11018);
nor U11056 (N_11056,N_10926,N_10997);
nor U11057 (N_11057,N_10932,N_10917);
xnor U11058 (N_11058,N_10996,N_10928);
nand U11059 (N_11059,N_10905,N_10931);
or U11060 (N_11060,N_10972,N_10894);
or U11061 (N_11061,N_11000,N_10999);
nor U11062 (N_11062,N_10893,N_10994);
xnor U11063 (N_11063,N_10916,N_10885);
nand U11064 (N_11064,N_10888,N_11037);
xor U11065 (N_11065,N_11020,N_10983);
and U11066 (N_11066,N_11028,N_10982);
or U11067 (N_11067,N_10943,N_10977);
and U11068 (N_11068,N_10991,N_10957);
or U11069 (N_11069,N_10946,N_10969);
nand U11070 (N_11070,N_10902,N_10924);
nor U11071 (N_11071,N_10937,N_10998);
nand U11072 (N_11072,N_11001,N_11033);
and U11073 (N_11073,N_10909,N_11027);
nand U11074 (N_11074,N_10881,N_11031);
and U11075 (N_11075,N_10979,N_10980);
or U11076 (N_11076,N_11012,N_10915);
nand U11077 (N_11077,N_11032,N_10985);
nor U11078 (N_11078,N_10923,N_10907);
nand U11079 (N_11079,N_10952,N_11017);
nand U11080 (N_11080,N_10995,N_10975);
or U11081 (N_11081,N_10913,N_10976);
xnor U11082 (N_11082,N_10986,N_10981);
nand U11083 (N_11083,N_10892,N_10882);
nor U11084 (N_11084,N_10904,N_11007);
or U11085 (N_11085,N_10960,N_11024);
or U11086 (N_11086,N_10978,N_11004);
and U11087 (N_11087,N_10964,N_10948);
and U11088 (N_11088,N_10984,N_11035);
nand U11089 (N_11089,N_10958,N_10927);
and U11090 (N_11090,N_10961,N_10962);
nor U11091 (N_11091,N_10954,N_10918);
nand U11092 (N_11092,N_11023,N_10953);
and U11093 (N_11093,N_11013,N_10919);
or U11094 (N_11094,N_10910,N_10908);
and U11095 (N_11095,N_10903,N_10884);
or U11096 (N_11096,N_10887,N_11006);
or U11097 (N_11097,N_11036,N_10940);
xnor U11098 (N_11098,N_10938,N_10968);
nand U11099 (N_11099,N_10914,N_10898);
and U11100 (N_11100,N_10895,N_10920);
or U11101 (N_11101,N_11038,N_10934);
or U11102 (N_11102,N_10987,N_10967);
xnor U11103 (N_11103,N_11015,N_11003);
or U11104 (N_11104,N_11002,N_11011);
xnor U11105 (N_11105,N_11022,N_10925);
nor U11106 (N_11106,N_11009,N_10941);
or U11107 (N_11107,N_10891,N_10890);
nor U11108 (N_11108,N_10944,N_10974);
xnor U11109 (N_11109,N_10922,N_10947);
nor U11110 (N_11110,N_10945,N_10939);
or U11111 (N_11111,N_11021,N_10883);
and U11112 (N_11112,N_10935,N_10899);
and U11113 (N_11113,N_10950,N_11016);
nand U11114 (N_11114,N_10929,N_11034);
nor U11115 (N_11115,N_10956,N_11010);
nand U11116 (N_11116,N_10951,N_11029);
or U11117 (N_11117,N_11030,N_10990);
nor U11118 (N_11118,N_11039,N_10886);
xor U11119 (N_11119,N_11005,N_10921);
nand U11120 (N_11120,N_10946,N_10980);
or U11121 (N_11121,N_10965,N_10881);
or U11122 (N_11122,N_10960,N_10907);
nor U11123 (N_11123,N_10929,N_10984);
or U11124 (N_11124,N_11016,N_10988);
nand U11125 (N_11125,N_11011,N_10895);
or U11126 (N_11126,N_11015,N_10920);
and U11127 (N_11127,N_10982,N_10933);
nand U11128 (N_11128,N_10975,N_10986);
nor U11129 (N_11129,N_10976,N_10958);
nor U11130 (N_11130,N_10934,N_11012);
or U11131 (N_11131,N_10924,N_10909);
nand U11132 (N_11132,N_10927,N_11000);
or U11133 (N_11133,N_11032,N_10903);
nor U11134 (N_11134,N_11018,N_10966);
and U11135 (N_11135,N_10969,N_10994);
and U11136 (N_11136,N_10904,N_11018);
or U11137 (N_11137,N_10970,N_10914);
or U11138 (N_11138,N_10997,N_10938);
nor U11139 (N_11139,N_10897,N_11003);
nor U11140 (N_11140,N_10978,N_11009);
nor U11141 (N_11141,N_10911,N_10995);
and U11142 (N_11142,N_10921,N_11036);
nor U11143 (N_11143,N_11026,N_10987);
and U11144 (N_11144,N_11011,N_10903);
xor U11145 (N_11145,N_10972,N_10974);
xnor U11146 (N_11146,N_10966,N_10950);
nor U11147 (N_11147,N_10998,N_10982);
nor U11148 (N_11148,N_10990,N_10899);
xor U11149 (N_11149,N_10937,N_10959);
nand U11150 (N_11150,N_11028,N_10900);
nor U11151 (N_11151,N_10993,N_10887);
and U11152 (N_11152,N_10982,N_10899);
xnor U11153 (N_11153,N_10920,N_10993);
nand U11154 (N_11154,N_10913,N_10926);
or U11155 (N_11155,N_10907,N_11016);
xnor U11156 (N_11156,N_10969,N_10899);
nor U11157 (N_11157,N_11017,N_10989);
nand U11158 (N_11158,N_10934,N_11023);
or U11159 (N_11159,N_10899,N_10907);
nor U11160 (N_11160,N_10928,N_10919);
nor U11161 (N_11161,N_11014,N_11022);
nor U11162 (N_11162,N_10979,N_10994);
or U11163 (N_11163,N_10909,N_10902);
and U11164 (N_11164,N_10898,N_10897);
or U11165 (N_11165,N_10957,N_10895);
nor U11166 (N_11166,N_10923,N_10904);
or U11167 (N_11167,N_10963,N_10906);
and U11168 (N_11168,N_10947,N_10892);
nor U11169 (N_11169,N_10901,N_10973);
or U11170 (N_11170,N_11016,N_10881);
and U11171 (N_11171,N_10997,N_11039);
nor U11172 (N_11172,N_11032,N_10999);
nor U11173 (N_11173,N_10994,N_10950);
and U11174 (N_11174,N_10882,N_11003);
or U11175 (N_11175,N_10975,N_10996);
or U11176 (N_11176,N_10974,N_11023);
and U11177 (N_11177,N_10951,N_10958);
or U11178 (N_11178,N_10906,N_10881);
or U11179 (N_11179,N_10940,N_11035);
and U11180 (N_11180,N_10977,N_10979);
and U11181 (N_11181,N_10935,N_11032);
nand U11182 (N_11182,N_11015,N_11030);
nor U11183 (N_11183,N_10979,N_11022);
nor U11184 (N_11184,N_11014,N_10993);
xnor U11185 (N_11185,N_11021,N_10905);
nand U11186 (N_11186,N_10979,N_10935);
nor U11187 (N_11187,N_10902,N_10957);
or U11188 (N_11188,N_10895,N_10970);
and U11189 (N_11189,N_10944,N_10967);
or U11190 (N_11190,N_11028,N_10966);
nand U11191 (N_11191,N_10943,N_10907);
and U11192 (N_11192,N_10961,N_11024);
or U11193 (N_11193,N_10909,N_10885);
or U11194 (N_11194,N_10977,N_11039);
nor U11195 (N_11195,N_10994,N_10947);
or U11196 (N_11196,N_11025,N_11014);
and U11197 (N_11197,N_11021,N_10950);
nor U11198 (N_11198,N_10919,N_11008);
or U11199 (N_11199,N_10888,N_10907);
and U11200 (N_11200,N_11187,N_11046);
and U11201 (N_11201,N_11040,N_11088);
and U11202 (N_11202,N_11041,N_11080);
xor U11203 (N_11203,N_11155,N_11182);
nand U11204 (N_11204,N_11196,N_11191);
or U11205 (N_11205,N_11141,N_11067);
nor U11206 (N_11206,N_11130,N_11045);
nand U11207 (N_11207,N_11127,N_11194);
nor U11208 (N_11208,N_11089,N_11079);
or U11209 (N_11209,N_11153,N_11148);
and U11210 (N_11210,N_11087,N_11048);
nor U11211 (N_11211,N_11096,N_11128);
nand U11212 (N_11212,N_11074,N_11103);
nor U11213 (N_11213,N_11177,N_11058);
nand U11214 (N_11214,N_11057,N_11171);
nand U11215 (N_11215,N_11181,N_11116);
or U11216 (N_11216,N_11053,N_11097);
and U11217 (N_11217,N_11161,N_11111);
nand U11218 (N_11218,N_11132,N_11082);
nor U11219 (N_11219,N_11185,N_11195);
nor U11220 (N_11220,N_11108,N_11061);
and U11221 (N_11221,N_11138,N_11174);
and U11222 (N_11222,N_11122,N_11193);
or U11223 (N_11223,N_11190,N_11152);
and U11224 (N_11224,N_11183,N_11077);
nor U11225 (N_11225,N_11140,N_11158);
nand U11226 (N_11226,N_11157,N_11094);
nand U11227 (N_11227,N_11118,N_11109);
and U11228 (N_11228,N_11102,N_11044);
nand U11229 (N_11229,N_11179,N_11124);
xor U11230 (N_11230,N_11099,N_11120);
or U11231 (N_11231,N_11106,N_11166);
nand U11232 (N_11232,N_11134,N_11121);
nand U11233 (N_11233,N_11112,N_11125);
nor U11234 (N_11234,N_11133,N_11107);
and U11235 (N_11235,N_11165,N_11160);
or U11236 (N_11236,N_11051,N_11150);
xor U11237 (N_11237,N_11123,N_11105);
nor U11238 (N_11238,N_11055,N_11085);
nor U11239 (N_11239,N_11081,N_11100);
or U11240 (N_11240,N_11135,N_11095);
nand U11241 (N_11241,N_11049,N_11101);
or U11242 (N_11242,N_11110,N_11064);
nand U11243 (N_11243,N_11042,N_11054);
or U11244 (N_11244,N_11199,N_11189);
nor U11245 (N_11245,N_11043,N_11151);
nand U11246 (N_11246,N_11163,N_11142);
or U11247 (N_11247,N_11068,N_11154);
nand U11248 (N_11248,N_11114,N_11076);
or U11249 (N_11249,N_11145,N_11070);
nand U11250 (N_11250,N_11178,N_11162);
or U11251 (N_11251,N_11078,N_11131);
or U11252 (N_11252,N_11091,N_11136);
nor U11253 (N_11253,N_11117,N_11168);
nand U11254 (N_11254,N_11146,N_11184);
or U11255 (N_11255,N_11113,N_11069);
or U11256 (N_11256,N_11188,N_11173);
and U11257 (N_11257,N_11056,N_11083);
nor U11258 (N_11258,N_11129,N_11197);
and U11259 (N_11259,N_11066,N_11119);
nor U11260 (N_11260,N_11050,N_11149);
or U11261 (N_11261,N_11167,N_11137);
nand U11262 (N_11262,N_11063,N_11198);
xnor U11263 (N_11263,N_11144,N_11084);
and U11264 (N_11264,N_11086,N_11075);
and U11265 (N_11265,N_11047,N_11175);
nand U11266 (N_11266,N_11172,N_11186);
or U11267 (N_11267,N_11071,N_11147);
nor U11268 (N_11268,N_11139,N_11126);
nand U11269 (N_11269,N_11170,N_11090);
nand U11270 (N_11270,N_11062,N_11159);
nand U11271 (N_11271,N_11192,N_11098);
nand U11272 (N_11272,N_11065,N_11164);
nand U11273 (N_11273,N_11104,N_11073);
nor U11274 (N_11274,N_11176,N_11143);
nor U11275 (N_11275,N_11156,N_11059);
or U11276 (N_11276,N_11169,N_11092);
and U11277 (N_11277,N_11060,N_11180);
nand U11278 (N_11278,N_11072,N_11115);
nand U11279 (N_11279,N_11093,N_11052);
nor U11280 (N_11280,N_11128,N_11082);
and U11281 (N_11281,N_11147,N_11162);
and U11282 (N_11282,N_11049,N_11156);
and U11283 (N_11283,N_11094,N_11162);
nor U11284 (N_11284,N_11099,N_11071);
and U11285 (N_11285,N_11103,N_11064);
nor U11286 (N_11286,N_11043,N_11075);
or U11287 (N_11287,N_11146,N_11156);
or U11288 (N_11288,N_11127,N_11153);
nand U11289 (N_11289,N_11082,N_11199);
or U11290 (N_11290,N_11173,N_11040);
nor U11291 (N_11291,N_11044,N_11137);
and U11292 (N_11292,N_11121,N_11056);
nand U11293 (N_11293,N_11136,N_11120);
nand U11294 (N_11294,N_11057,N_11100);
or U11295 (N_11295,N_11125,N_11042);
xor U11296 (N_11296,N_11136,N_11181);
nand U11297 (N_11297,N_11175,N_11165);
or U11298 (N_11298,N_11139,N_11190);
nand U11299 (N_11299,N_11137,N_11076);
nand U11300 (N_11300,N_11082,N_11186);
nand U11301 (N_11301,N_11123,N_11183);
and U11302 (N_11302,N_11089,N_11126);
xnor U11303 (N_11303,N_11083,N_11096);
or U11304 (N_11304,N_11181,N_11144);
nand U11305 (N_11305,N_11183,N_11141);
or U11306 (N_11306,N_11069,N_11068);
nand U11307 (N_11307,N_11140,N_11069);
nor U11308 (N_11308,N_11131,N_11194);
nand U11309 (N_11309,N_11043,N_11098);
or U11310 (N_11310,N_11186,N_11100);
or U11311 (N_11311,N_11086,N_11187);
nand U11312 (N_11312,N_11128,N_11097);
xor U11313 (N_11313,N_11150,N_11069);
nor U11314 (N_11314,N_11159,N_11138);
nor U11315 (N_11315,N_11142,N_11053);
and U11316 (N_11316,N_11179,N_11060);
nand U11317 (N_11317,N_11176,N_11118);
nand U11318 (N_11318,N_11087,N_11172);
and U11319 (N_11319,N_11101,N_11147);
or U11320 (N_11320,N_11046,N_11053);
nor U11321 (N_11321,N_11143,N_11088);
nor U11322 (N_11322,N_11174,N_11053);
xnor U11323 (N_11323,N_11112,N_11193);
nand U11324 (N_11324,N_11138,N_11124);
nand U11325 (N_11325,N_11087,N_11064);
nand U11326 (N_11326,N_11171,N_11113);
or U11327 (N_11327,N_11157,N_11091);
or U11328 (N_11328,N_11056,N_11125);
nor U11329 (N_11329,N_11053,N_11076);
and U11330 (N_11330,N_11104,N_11174);
nor U11331 (N_11331,N_11179,N_11056);
or U11332 (N_11332,N_11061,N_11157);
nand U11333 (N_11333,N_11069,N_11177);
nor U11334 (N_11334,N_11095,N_11177);
nor U11335 (N_11335,N_11122,N_11103);
and U11336 (N_11336,N_11186,N_11118);
or U11337 (N_11337,N_11160,N_11147);
nor U11338 (N_11338,N_11164,N_11117);
nand U11339 (N_11339,N_11187,N_11042);
and U11340 (N_11340,N_11165,N_11128);
or U11341 (N_11341,N_11128,N_11130);
nand U11342 (N_11342,N_11052,N_11154);
or U11343 (N_11343,N_11143,N_11140);
nor U11344 (N_11344,N_11056,N_11168);
or U11345 (N_11345,N_11046,N_11064);
and U11346 (N_11346,N_11050,N_11104);
and U11347 (N_11347,N_11196,N_11099);
nand U11348 (N_11348,N_11109,N_11133);
or U11349 (N_11349,N_11121,N_11172);
nand U11350 (N_11350,N_11158,N_11069);
nand U11351 (N_11351,N_11095,N_11174);
nor U11352 (N_11352,N_11168,N_11064);
or U11353 (N_11353,N_11062,N_11124);
nor U11354 (N_11354,N_11149,N_11065);
nand U11355 (N_11355,N_11178,N_11166);
nor U11356 (N_11356,N_11082,N_11137);
or U11357 (N_11357,N_11089,N_11180);
and U11358 (N_11358,N_11117,N_11097);
and U11359 (N_11359,N_11040,N_11104);
nor U11360 (N_11360,N_11291,N_11275);
nand U11361 (N_11361,N_11348,N_11238);
and U11362 (N_11362,N_11264,N_11265);
nor U11363 (N_11363,N_11303,N_11230);
nor U11364 (N_11364,N_11294,N_11331);
and U11365 (N_11365,N_11352,N_11269);
and U11366 (N_11366,N_11274,N_11340);
nand U11367 (N_11367,N_11245,N_11217);
nor U11368 (N_11368,N_11214,N_11358);
or U11369 (N_11369,N_11308,N_11244);
nand U11370 (N_11370,N_11304,N_11225);
nand U11371 (N_11371,N_11322,N_11270);
nor U11372 (N_11372,N_11278,N_11239);
xnor U11373 (N_11373,N_11281,N_11353);
and U11374 (N_11374,N_11356,N_11237);
or U11375 (N_11375,N_11295,N_11272);
or U11376 (N_11376,N_11288,N_11207);
or U11377 (N_11377,N_11203,N_11341);
xor U11378 (N_11378,N_11250,N_11211);
nand U11379 (N_11379,N_11226,N_11209);
or U11380 (N_11380,N_11307,N_11325);
and U11381 (N_11381,N_11316,N_11280);
nand U11382 (N_11382,N_11247,N_11345);
nor U11383 (N_11383,N_11219,N_11333);
nand U11384 (N_11384,N_11285,N_11227);
or U11385 (N_11385,N_11204,N_11259);
nor U11386 (N_11386,N_11201,N_11231);
nor U11387 (N_11387,N_11208,N_11327);
and U11388 (N_11388,N_11344,N_11235);
nor U11389 (N_11389,N_11215,N_11292);
nand U11390 (N_11390,N_11228,N_11324);
xor U11391 (N_11391,N_11357,N_11262);
or U11392 (N_11392,N_11266,N_11284);
nor U11393 (N_11393,N_11260,N_11351);
nand U11394 (N_11394,N_11205,N_11317);
or U11395 (N_11395,N_11218,N_11242);
nand U11396 (N_11396,N_11290,N_11305);
and U11397 (N_11397,N_11301,N_11349);
nor U11398 (N_11398,N_11233,N_11306);
and U11399 (N_11399,N_11343,N_11334);
nor U11400 (N_11400,N_11330,N_11271);
nand U11401 (N_11401,N_11312,N_11256);
nor U11402 (N_11402,N_11213,N_11246);
or U11403 (N_11403,N_11296,N_11293);
or U11404 (N_11404,N_11252,N_11309);
xnor U11405 (N_11405,N_11321,N_11243);
nor U11406 (N_11406,N_11354,N_11241);
and U11407 (N_11407,N_11254,N_11313);
and U11408 (N_11408,N_11240,N_11223);
nand U11409 (N_11409,N_11332,N_11279);
xnor U11410 (N_11410,N_11314,N_11319);
and U11411 (N_11411,N_11210,N_11336);
nor U11412 (N_11412,N_11287,N_11328);
or U11413 (N_11413,N_11224,N_11297);
nand U11414 (N_11414,N_11346,N_11326);
nor U11415 (N_11415,N_11335,N_11206);
xor U11416 (N_11416,N_11236,N_11249);
nand U11417 (N_11417,N_11299,N_11255);
or U11418 (N_11418,N_11323,N_11282);
and U11419 (N_11419,N_11277,N_11248);
nor U11420 (N_11420,N_11251,N_11359);
or U11421 (N_11421,N_11222,N_11355);
nor U11422 (N_11422,N_11283,N_11232);
and U11423 (N_11423,N_11258,N_11273);
and U11424 (N_11424,N_11257,N_11276);
nor U11425 (N_11425,N_11310,N_11315);
nand U11426 (N_11426,N_11261,N_11342);
xnor U11427 (N_11427,N_11347,N_11339);
and U11428 (N_11428,N_11318,N_11229);
nor U11429 (N_11429,N_11300,N_11220);
and U11430 (N_11430,N_11329,N_11200);
or U11431 (N_11431,N_11298,N_11212);
nor U11432 (N_11432,N_11286,N_11289);
and U11433 (N_11433,N_11253,N_11267);
and U11434 (N_11434,N_11337,N_11234);
xor U11435 (N_11435,N_11216,N_11268);
or U11436 (N_11436,N_11263,N_11302);
and U11437 (N_11437,N_11320,N_11202);
nor U11438 (N_11438,N_11350,N_11338);
nor U11439 (N_11439,N_11221,N_11311);
nor U11440 (N_11440,N_11329,N_11315);
nor U11441 (N_11441,N_11247,N_11226);
or U11442 (N_11442,N_11262,N_11249);
nand U11443 (N_11443,N_11287,N_11314);
or U11444 (N_11444,N_11333,N_11265);
nand U11445 (N_11445,N_11244,N_11351);
nand U11446 (N_11446,N_11258,N_11299);
or U11447 (N_11447,N_11293,N_11207);
nand U11448 (N_11448,N_11267,N_11212);
and U11449 (N_11449,N_11300,N_11297);
nor U11450 (N_11450,N_11264,N_11206);
or U11451 (N_11451,N_11216,N_11227);
and U11452 (N_11452,N_11340,N_11349);
nor U11453 (N_11453,N_11215,N_11330);
nor U11454 (N_11454,N_11263,N_11207);
nand U11455 (N_11455,N_11220,N_11321);
nor U11456 (N_11456,N_11322,N_11284);
or U11457 (N_11457,N_11350,N_11262);
nor U11458 (N_11458,N_11349,N_11265);
nand U11459 (N_11459,N_11331,N_11327);
nand U11460 (N_11460,N_11333,N_11278);
and U11461 (N_11461,N_11314,N_11313);
and U11462 (N_11462,N_11284,N_11282);
and U11463 (N_11463,N_11203,N_11326);
nand U11464 (N_11464,N_11213,N_11289);
xnor U11465 (N_11465,N_11336,N_11237);
xor U11466 (N_11466,N_11208,N_11299);
or U11467 (N_11467,N_11310,N_11313);
xnor U11468 (N_11468,N_11346,N_11269);
and U11469 (N_11469,N_11258,N_11356);
nand U11470 (N_11470,N_11217,N_11279);
nand U11471 (N_11471,N_11358,N_11308);
and U11472 (N_11472,N_11341,N_11301);
or U11473 (N_11473,N_11256,N_11296);
or U11474 (N_11474,N_11200,N_11325);
nor U11475 (N_11475,N_11293,N_11359);
or U11476 (N_11476,N_11218,N_11261);
nor U11477 (N_11477,N_11227,N_11206);
and U11478 (N_11478,N_11285,N_11256);
nand U11479 (N_11479,N_11258,N_11349);
and U11480 (N_11480,N_11338,N_11255);
nor U11481 (N_11481,N_11344,N_11269);
and U11482 (N_11482,N_11226,N_11314);
nand U11483 (N_11483,N_11284,N_11341);
nand U11484 (N_11484,N_11342,N_11266);
nand U11485 (N_11485,N_11337,N_11307);
nor U11486 (N_11486,N_11312,N_11221);
nand U11487 (N_11487,N_11220,N_11348);
and U11488 (N_11488,N_11283,N_11335);
nor U11489 (N_11489,N_11326,N_11259);
nor U11490 (N_11490,N_11257,N_11295);
and U11491 (N_11491,N_11204,N_11330);
nand U11492 (N_11492,N_11232,N_11326);
nor U11493 (N_11493,N_11287,N_11234);
and U11494 (N_11494,N_11256,N_11238);
or U11495 (N_11495,N_11334,N_11210);
xor U11496 (N_11496,N_11354,N_11226);
nor U11497 (N_11497,N_11351,N_11279);
or U11498 (N_11498,N_11217,N_11259);
nand U11499 (N_11499,N_11313,N_11343);
and U11500 (N_11500,N_11348,N_11329);
and U11501 (N_11501,N_11301,N_11256);
and U11502 (N_11502,N_11209,N_11221);
nor U11503 (N_11503,N_11303,N_11316);
and U11504 (N_11504,N_11297,N_11320);
or U11505 (N_11505,N_11262,N_11247);
or U11506 (N_11506,N_11289,N_11264);
and U11507 (N_11507,N_11301,N_11241);
or U11508 (N_11508,N_11242,N_11244);
and U11509 (N_11509,N_11310,N_11258);
nand U11510 (N_11510,N_11225,N_11319);
nor U11511 (N_11511,N_11309,N_11354);
and U11512 (N_11512,N_11298,N_11202);
nor U11513 (N_11513,N_11308,N_11233);
nor U11514 (N_11514,N_11308,N_11354);
nor U11515 (N_11515,N_11296,N_11297);
nor U11516 (N_11516,N_11299,N_11201);
and U11517 (N_11517,N_11316,N_11319);
nand U11518 (N_11518,N_11214,N_11224);
or U11519 (N_11519,N_11273,N_11231);
nand U11520 (N_11520,N_11390,N_11428);
or U11521 (N_11521,N_11397,N_11442);
or U11522 (N_11522,N_11519,N_11394);
or U11523 (N_11523,N_11376,N_11367);
nor U11524 (N_11524,N_11371,N_11464);
xor U11525 (N_11525,N_11506,N_11384);
or U11526 (N_11526,N_11459,N_11372);
nand U11527 (N_11527,N_11495,N_11424);
and U11528 (N_11528,N_11493,N_11409);
nand U11529 (N_11529,N_11518,N_11425);
or U11530 (N_11530,N_11448,N_11415);
nor U11531 (N_11531,N_11422,N_11412);
and U11532 (N_11532,N_11414,N_11482);
xor U11533 (N_11533,N_11435,N_11444);
and U11534 (N_11534,N_11366,N_11417);
nor U11535 (N_11535,N_11392,N_11423);
and U11536 (N_11536,N_11381,N_11514);
nand U11537 (N_11537,N_11496,N_11515);
and U11538 (N_11538,N_11445,N_11395);
nand U11539 (N_11539,N_11396,N_11512);
or U11540 (N_11540,N_11454,N_11465);
and U11541 (N_11541,N_11455,N_11360);
xor U11542 (N_11542,N_11449,N_11481);
nor U11543 (N_11543,N_11447,N_11473);
and U11544 (N_11544,N_11386,N_11452);
or U11545 (N_11545,N_11374,N_11499);
xnor U11546 (N_11546,N_11420,N_11504);
or U11547 (N_11547,N_11438,N_11403);
nor U11548 (N_11548,N_11461,N_11468);
xnor U11549 (N_11549,N_11382,N_11483);
nand U11550 (N_11550,N_11370,N_11404);
nand U11551 (N_11551,N_11439,N_11432);
nand U11552 (N_11552,N_11470,N_11511);
nor U11553 (N_11553,N_11475,N_11410);
and U11554 (N_11554,N_11491,N_11385);
nor U11555 (N_11555,N_11413,N_11467);
nand U11556 (N_11556,N_11457,N_11436);
or U11557 (N_11557,N_11469,N_11365);
or U11558 (N_11558,N_11517,N_11479);
nand U11559 (N_11559,N_11474,N_11485);
nor U11560 (N_11560,N_11437,N_11492);
nor U11561 (N_11561,N_11490,N_11362);
and U11562 (N_11562,N_11378,N_11472);
and U11563 (N_11563,N_11383,N_11426);
nand U11564 (N_11564,N_11480,N_11487);
nand U11565 (N_11565,N_11489,N_11380);
nand U11566 (N_11566,N_11393,N_11476);
or U11567 (N_11567,N_11443,N_11401);
and U11568 (N_11568,N_11434,N_11373);
nor U11569 (N_11569,N_11471,N_11456);
or U11570 (N_11570,N_11451,N_11418);
or U11571 (N_11571,N_11405,N_11377);
or U11572 (N_11572,N_11458,N_11497);
and U11573 (N_11573,N_11513,N_11363);
or U11574 (N_11574,N_11398,N_11509);
nand U11575 (N_11575,N_11391,N_11399);
or U11576 (N_11576,N_11441,N_11488);
nand U11577 (N_11577,N_11368,N_11501);
and U11578 (N_11578,N_11505,N_11498);
nand U11579 (N_11579,N_11388,N_11389);
and U11580 (N_11580,N_11494,N_11419);
and U11581 (N_11581,N_11433,N_11407);
or U11582 (N_11582,N_11361,N_11431);
nor U11583 (N_11583,N_11446,N_11379);
nor U11584 (N_11584,N_11400,N_11430);
and U11585 (N_11585,N_11421,N_11402);
nand U11586 (N_11586,N_11450,N_11460);
nor U11587 (N_11587,N_11500,N_11406);
and U11588 (N_11588,N_11516,N_11440);
nand U11589 (N_11589,N_11369,N_11387);
nor U11590 (N_11590,N_11427,N_11486);
nor U11591 (N_11591,N_11411,N_11466);
or U11592 (N_11592,N_11484,N_11502);
nand U11593 (N_11593,N_11478,N_11507);
xnor U11594 (N_11594,N_11408,N_11453);
or U11595 (N_11595,N_11462,N_11463);
or U11596 (N_11596,N_11503,N_11375);
nor U11597 (N_11597,N_11510,N_11364);
nor U11598 (N_11598,N_11477,N_11429);
nand U11599 (N_11599,N_11508,N_11416);
or U11600 (N_11600,N_11410,N_11456);
nand U11601 (N_11601,N_11404,N_11506);
nor U11602 (N_11602,N_11401,N_11474);
and U11603 (N_11603,N_11474,N_11377);
or U11604 (N_11604,N_11482,N_11507);
xor U11605 (N_11605,N_11418,N_11392);
or U11606 (N_11606,N_11425,N_11477);
or U11607 (N_11607,N_11500,N_11391);
or U11608 (N_11608,N_11495,N_11398);
and U11609 (N_11609,N_11463,N_11458);
nand U11610 (N_11610,N_11495,N_11406);
or U11611 (N_11611,N_11516,N_11419);
nor U11612 (N_11612,N_11383,N_11473);
nor U11613 (N_11613,N_11421,N_11446);
and U11614 (N_11614,N_11462,N_11446);
or U11615 (N_11615,N_11401,N_11430);
nor U11616 (N_11616,N_11447,N_11439);
or U11617 (N_11617,N_11446,N_11455);
nand U11618 (N_11618,N_11369,N_11478);
or U11619 (N_11619,N_11382,N_11450);
xor U11620 (N_11620,N_11399,N_11433);
and U11621 (N_11621,N_11454,N_11473);
nand U11622 (N_11622,N_11385,N_11427);
or U11623 (N_11623,N_11505,N_11422);
xnor U11624 (N_11624,N_11511,N_11390);
nand U11625 (N_11625,N_11518,N_11481);
xor U11626 (N_11626,N_11422,N_11444);
nand U11627 (N_11627,N_11364,N_11471);
and U11628 (N_11628,N_11401,N_11470);
nor U11629 (N_11629,N_11446,N_11514);
and U11630 (N_11630,N_11374,N_11447);
or U11631 (N_11631,N_11510,N_11372);
and U11632 (N_11632,N_11439,N_11436);
or U11633 (N_11633,N_11473,N_11364);
and U11634 (N_11634,N_11383,N_11367);
or U11635 (N_11635,N_11437,N_11424);
and U11636 (N_11636,N_11362,N_11376);
nand U11637 (N_11637,N_11453,N_11393);
nand U11638 (N_11638,N_11364,N_11402);
nand U11639 (N_11639,N_11420,N_11430);
nor U11640 (N_11640,N_11372,N_11451);
and U11641 (N_11641,N_11387,N_11438);
nand U11642 (N_11642,N_11448,N_11374);
or U11643 (N_11643,N_11462,N_11374);
and U11644 (N_11644,N_11498,N_11485);
and U11645 (N_11645,N_11454,N_11494);
and U11646 (N_11646,N_11471,N_11386);
or U11647 (N_11647,N_11432,N_11422);
nor U11648 (N_11648,N_11465,N_11435);
nand U11649 (N_11649,N_11441,N_11442);
nor U11650 (N_11650,N_11464,N_11488);
and U11651 (N_11651,N_11403,N_11497);
or U11652 (N_11652,N_11441,N_11492);
nand U11653 (N_11653,N_11461,N_11462);
nor U11654 (N_11654,N_11427,N_11463);
nand U11655 (N_11655,N_11483,N_11461);
xnor U11656 (N_11656,N_11363,N_11380);
nor U11657 (N_11657,N_11455,N_11511);
nand U11658 (N_11658,N_11374,N_11439);
nor U11659 (N_11659,N_11461,N_11374);
nor U11660 (N_11660,N_11482,N_11448);
and U11661 (N_11661,N_11478,N_11514);
and U11662 (N_11662,N_11509,N_11474);
and U11663 (N_11663,N_11445,N_11367);
xor U11664 (N_11664,N_11444,N_11456);
nand U11665 (N_11665,N_11491,N_11394);
nor U11666 (N_11666,N_11395,N_11382);
or U11667 (N_11667,N_11438,N_11463);
and U11668 (N_11668,N_11503,N_11400);
nand U11669 (N_11669,N_11502,N_11489);
nand U11670 (N_11670,N_11483,N_11389);
and U11671 (N_11671,N_11444,N_11377);
nor U11672 (N_11672,N_11459,N_11431);
or U11673 (N_11673,N_11439,N_11396);
nor U11674 (N_11674,N_11458,N_11515);
nor U11675 (N_11675,N_11424,N_11444);
nor U11676 (N_11676,N_11374,N_11455);
and U11677 (N_11677,N_11470,N_11379);
nor U11678 (N_11678,N_11394,N_11402);
nand U11679 (N_11679,N_11418,N_11383);
or U11680 (N_11680,N_11564,N_11580);
or U11681 (N_11681,N_11577,N_11582);
and U11682 (N_11682,N_11553,N_11669);
nor U11683 (N_11683,N_11609,N_11575);
or U11684 (N_11684,N_11572,N_11654);
and U11685 (N_11685,N_11657,N_11560);
nor U11686 (N_11686,N_11624,N_11653);
nand U11687 (N_11687,N_11635,N_11673);
and U11688 (N_11688,N_11588,N_11570);
nor U11689 (N_11689,N_11583,N_11576);
nor U11690 (N_11690,N_11594,N_11550);
and U11691 (N_11691,N_11662,N_11574);
or U11692 (N_11692,N_11539,N_11631);
and U11693 (N_11693,N_11530,N_11658);
xor U11694 (N_11694,N_11619,N_11677);
nor U11695 (N_11695,N_11533,N_11532);
and U11696 (N_11696,N_11573,N_11674);
nand U11697 (N_11697,N_11663,N_11610);
and U11698 (N_11698,N_11651,N_11650);
nor U11699 (N_11699,N_11640,N_11642);
or U11700 (N_11700,N_11527,N_11634);
or U11701 (N_11701,N_11656,N_11523);
and U11702 (N_11702,N_11679,N_11558);
nor U11703 (N_11703,N_11628,N_11639);
nand U11704 (N_11704,N_11648,N_11551);
nor U11705 (N_11705,N_11602,N_11557);
xnor U11706 (N_11706,N_11544,N_11615);
or U11707 (N_11707,N_11562,N_11621);
and U11708 (N_11708,N_11637,N_11659);
or U11709 (N_11709,N_11596,N_11591);
nor U11710 (N_11710,N_11548,N_11566);
nand U11711 (N_11711,N_11606,N_11625);
or U11712 (N_11712,N_11525,N_11571);
or U11713 (N_11713,N_11668,N_11647);
nand U11714 (N_11714,N_11529,N_11526);
xnor U11715 (N_11715,N_11528,N_11641);
xnor U11716 (N_11716,N_11652,N_11604);
or U11717 (N_11717,N_11569,N_11620);
or U11718 (N_11718,N_11541,N_11617);
nor U11719 (N_11719,N_11630,N_11599);
and U11720 (N_11720,N_11535,N_11540);
nor U11721 (N_11721,N_11590,N_11531);
nand U11722 (N_11722,N_11586,N_11678);
nand U11723 (N_11723,N_11549,N_11556);
xor U11724 (N_11724,N_11600,N_11534);
or U11725 (N_11725,N_11660,N_11675);
nand U11726 (N_11726,N_11633,N_11643);
and U11727 (N_11727,N_11536,N_11649);
and U11728 (N_11728,N_11595,N_11584);
nand U11729 (N_11729,N_11589,N_11665);
nor U11730 (N_11730,N_11598,N_11612);
nor U11731 (N_11731,N_11538,N_11622);
and U11732 (N_11732,N_11608,N_11626);
nor U11733 (N_11733,N_11547,N_11567);
or U11734 (N_11734,N_11607,N_11616);
nor U11735 (N_11735,N_11592,N_11542);
and U11736 (N_11736,N_11644,N_11618);
or U11737 (N_11737,N_11629,N_11655);
or U11738 (N_11738,N_11554,N_11537);
xor U11739 (N_11739,N_11614,N_11520);
or U11740 (N_11740,N_11524,N_11676);
or U11741 (N_11741,N_11543,N_11632);
nor U11742 (N_11742,N_11667,N_11568);
nand U11743 (N_11743,N_11552,N_11579);
nor U11744 (N_11744,N_11578,N_11585);
nand U11745 (N_11745,N_11581,N_11672);
and U11746 (N_11746,N_11593,N_11623);
nand U11747 (N_11747,N_11664,N_11646);
and U11748 (N_11748,N_11613,N_11587);
nor U11749 (N_11749,N_11670,N_11522);
or U11750 (N_11750,N_11605,N_11671);
nor U11751 (N_11751,N_11638,N_11661);
nor U11752 (N_11752,N_11555,N_11521);
xnor U11753 (N_11753,N_11645,N_11546);
nand U11754 (N_11754,N_11565,N_11627);
and U11755 (N_11755,N_11559,N_11563);
or U11756 (N_11756,N_11603,N_11545);
nor U11757 (N_11757,N_11601,N_11611);
and U11758 (N_11758,N_11636,N_11561);
nand U11759 (N_11759,N_11666,N_11597);
and U11760 (N_11760,N_11534,N_11552);
and U11761 (N_11761,N_11581,N_11643);
xor U11762 (N_11762,N_11655,N_11575);
nor U11763 (N_11763,N_11530,N_11537);
or U11764 (N_11764,N_11546,N_11584);
nand U11765 (N_11765,N_11571,N_11626);
and U11766 (N_11766,N_11638,N_11586);
nand U11767 (N_11767,N_11652,N_11619);
and U11768 (N_11768,N_11657,N_11569);
or U11769 (N_11769,N_11657,N_11606);
nand U11770 (N_11770,N_11573,N_11565);
and U11771 (N_11771,N_11661,N_11595);
nor U11772 (N_11772,N_11615,N_11584);
nor U11773 (N_11773,N_11611,N_11633);
nor U11774 (N_11774,N_11615,N_11643);
nand U11775 (N_11775,N_11649,N_11658);
xor U11776 (N_11776,N_11556,N_11637);
nor U11777 (N_11777,N_11647,N_11591);
nor U11778 (N_11778,N_11641,N_11614);
xor U11779 (N_11779,N_11564,N_11586);
or U11780 (N_11780,N_11658,N_11667);
xnor U11781 (N_11781,N_11591,N_11637);
or U11782 (N_11782,N_11550,N_11657);
and U11783 (N_11783,N_11576,N_11546);
nor U11784 (N_11784,N_11546,N_11550);
nor U11785 (N_11785,N_11545,N_11541);
or U11786 (N_11786,N_11553,N_11663);
nand U11787 (N_11787,N_11572,N_11536);
or U11788 (N_11788,N_11614,N_11531);
nand U11789 (N_11789,N_11675,N_11583);
nand U11790 (N_11790,N_11600,N_11572);
nand U11791 (N_11791,N_11607,N_11528);
or U11792 (N_11792,N_11663,N_11533);
or U11793 (N_11793,N_11668,N_11521);
and U11794 (N_11794,N_11618,N_11664);
xnor U11795 (N_11795,N_11639,N_11528);
or U11796 (N_11796,N_11609,N_11539);
nor U11797 (N_11797,N_11534,N_11643);
nand U11798 (N_11798,N_11616,N_11540);
nand U11799 (N_11799,N_11643,N_11533);
nor U11800 (N_11800,N_11614,N_11643);
nor U11801 (N_11801,N_11603,N_11576);
xnor U11802 (N_11802,N_11606,N_11635);
nand U11803 (N_11803,N_11535,N_11568);
nand U11804 (N_11804,N_11609,N_11577);
nor U11805 (N_11805,N_11624,N_11571);
and U11806 (N_11806,N_11622,N_11576);
and U11807 (N_11807,N_11596,N_11675);
or U11808 (N_11808,N_11587,N_11580);
nand U11809 (N_11809,N_11665,N_11549);
nor U11810 (N_11810,N_11648,N_11539);
or U11811 (N_11811,N_11576,N_11637);
and U11812 (N_11812,N_11550,N_11553);
xor U11813 (N_11813,N_11532,N_11543);
nor U11814 (N_11814,N_11590,N_11627);
and U11815 (N_11815,N_11607,N_11633);
and U11816 (N_11816,N_11603,N_11601);
nand U11817 (N_11817,N_11665,N_11655);
and U11818 (N_11818,N_11644,N_11568);
or U11819 (N_11819,N_11623,N_11611);
xnor U11820 (N_11820,N_11549,N_11608);
and U11821 (N_11821,N_11592,N_11611);
or U11822 (N_11822,N_11535,N_11571);
xor U11823 (N_11823,N_11602,N_11547);
or U11824 (N_11824,N_11550,N_11636);
and U11825 (N_11825,N_11641,N_11654);
and U11826 (N_11826,N_11627,N_11671);
xnor U11827 (N_11827,N_11552,N_11520);
nand U11828 (N_11828,N_11664,N_11677);
and U11829 (N_11829,N_11626,N_11587);
xor U11830 (N_11830,N_11536,N_11545);
and U11831 (N_11831,N_11604,N_11654);
xor U11832 (N_11832,N_11614,N_11602);
or U11833 (N_11833,N_11539,N_11577);
nand U11834 (N_11834,N_11545,N_11657);
xnor U11835 (N_11835,N_11678,N_11624);
nor U11836 (N_11836,N_11627,N_11664);
and U11837 (N_11837,N_11565,N_11539);
and U11838 (N_11838,N_11565,N_11649);
nand U11839 (N_11839,N_11590,N_11565);
nor U11840 (N_11840,N_11836,N_11718);
nand U11841 (N_11841,N_11719,N_11767);
nor U11842 (N_11842,N_11765,N_11820);
nand U11843 (N_11843,N_11737,N_11753);
and U11844 (N_11844,N_11796,N_11808);
nor U11845 (N_11845,N_11746,N_11742);
nand U11846 (N_11846,N_11698,N_11739);
and U11847 (N_11847,N_11838,N_11747);
xnor U11848 (N_11848,N_11735,N_11793);
and U11849 (N_11849,N_11734,N_11809);
or U11850 (N_11850,N_11811,N_11807);
and U11851 (N_11851,N_11689,N_11815);
nor U11852 (N_11852,N_11721,N_11789);
or U11853 (N_11853,N_11818,N_11712);
nor U11854 (N_11854,N_11794,N_11696);
nor U11855 (N_11855,N_11821,N_11764);
nand U11856 (N_11856,N_11711,N_11837);
nand U11857 (N_11857,N_11705,N_11830);
xor U11858 (N_11858,N_11740,N_11706);
nor U11859 (N_11859,N_11833,N_11701);
nand U11860 (N_11860,N_11800,N_11795);
and U11861 (N_11861,N_11730,N_11806);
or U11862 (N_11862,N_11693,N_11741);
and U11863 (N_11863,N_11814,N_11702);
nor U11864 (N_11864,N_11697,N_11781);
nand U11865 (N_11865,N_11690,N_11716);
xor U11866 (N_11866,N_11812,N_11726);
nor U11867 (N_11867,N_11825,N_11715);
nor U11868 (N_11868,N_11788,N_11770);
and U11869 (N_11869,N_11688,N_11752);
and U11870 (N_11870,N_11723,N_11816);
or U11871 (N_11871,N_11801,N_11805);
nor U11872 (N_11872,N_11729,N_11839);
nor U11873 (N_11873,N_11835,N_11762);
nand U11874 (N_11874,N_11738,N_11754);
nor U11875 (N_11875,N_11819,N_11687);
xor U11876 (N_11876,N_11680,N_11758);
nand U11877 (N_11877,N_11803,N_11763);
or U11878 (N_11878,N_11755,N_11695);
nand U11879 (N_11879,N_11778,N_11757);
nor U11880 (N_11880,N_11694,N_11744);
nor U11881 (N_11881,N_11745,N_11787);
nand U11882 (N_11882,N_11792,N_11728);
nor U11883 (N_11883,N_11713,N_11736);
or U11884 (N_11884,N_11699,N_11710);
xor U11885 (N_11885,N_11724,N_11759);
and U11886 (N_11886,N_11722,N_11828);
nand U11887 (N_11887,N_11683,N_11727);
nor U11888 (N_11888,N_11760,N_11691);
nor U11889 (N_11889,N_11834,N_11799);
nor U11890 (N_11890,N_11817,N_11810);
nor U11891 (N_11891,N_11772,N_11766);
nand U11892 (N_11892,N_11751,N_11829);
and U11893 (N_11893,N_11733,N_11720);
and U11894 (N_11894,N_11783,N_11804);
and U11895 (N_11895,N_11826,N_11824);
or U11896 (N_11896,N_11703,N_11813);
or U11897 (N_11897,N_11775,N_11748);
nand U11898 (N_11898,N_11776,N_11774);
nor U11899 (N_11899,N_11769,N_11802);
or U11900 (N_11900,N_11692,N_11750);
xor U11901 (N_11901,N_11827,N_11798);
and U11902 (N_11902,N_11771,N_11832);
xnor U11903 (N_11903,N_11682,N_11700);
or U11904 (N_11904,N_11749,N_11707);
and U11905 (N_11905,N_11784,N_11717);
or U11906 (N_11906,N_11786,N_11681);
or U11907 (N_11907,N_11785,N_11823);
nand U11908 (N_11908,N_11708,N_11684);
and U11909 (N_11909,N_11777,N_11686);
nor U11910 (N_11910,N_11761,N_11768);
and U11911 (N_11911,N_11780,N_11782);
nand U11912 (N_11912,N_11822,N_11831);
and U11913 (N_11913,N_11704,N_11685);
and U11914 (N_11914,N_11756,N_11725);
and U11915 (N_11915,N_11714,N_11743);
nor U11916 (N_11916,N_11732,N_11779);
nor U11917 (N_11917,N_11797,N_11731);
nor U11918 (N_11918,N_11773,N_11791);
nand U11919 (N_11919,N_11709,N_11790);
or U11920 (N_11920,N_11716,N_11689);
and U11921 (N_11921,N_11738,N_11820);
and U11922 (N_11922,N_11765,N_11736);
nand U11923 (N_11923,N_11828,N_11692);
xor U11924 (N_11924,N_11770,N_11820);
nand U11925 (N_11925,N_11752,N_11749);
xnor U11926 (N_11926,N_11689,N_11821);
xnor U11927 (N_11927,N_11788,N_11789);
nand U11928 (N_11928,N_11693,N_11714);
and U11929 (N_11929,N_11689,N_11756);
and U11930 (N_11930,N_11757,N_11809);
or U11931 (N_11931,N_11745,N_11773);
nor U11932 (N_11932,N_11685,N_11813);
nor U11933 (N_11933,N_11828,N_11734);
or U11934 (N_11934,N_11775,N_11684);
or U11935 (N_11935,N_11829,N_11697);
or U11936 (N_11936,N_11777,N_11804);
nand U11937 (N_11937,N_11791,N_11763);
and U11938 (N_11938,N_11800,N_11753);
nand U11939 (N_11939,N_11729,N_11773);
nor U11940 (N_11940,N_11716,N_11733);
nand U11941 (N_11941,N_11815,N_11690);
nor U11942 (N_11942,N_11833,N_11739);
or U11943 (N_11943,N_11820,N_11714);
nor U11944 (N_11944,N_11719,N_11831);
or U11945 (N_11945,N_11811,N_11745);
xnor U11946 (N_11946,N_11806,N_11822);
nor U11947 (N_11947,N_11820,N_11710);
nand U11948 (N_11948,N_11828,N_11794);
or U11949 (N_11949,N_11723,N_11690);
and U11950 (N_11950,N_11770,N_11760);
nor U11951 (N_11951,N_11731,N_11832);
nor U11952 (N_11952,N_11784,N_11760);
or U11953 (N_11953,N_11780,N_11746);
and U11954 (N_11954,N_11829,N_11766);
nor U11955 (N_11955,N_11752,N_11786);
or U11956 (N_11956,N_11712,N_11837);
and U11957 (N_11957,N_11748,N_11744);
and U11958 (N_11958,N_11785,N_11782);
and U11959 (N_11959,N_11751,N_11755);
nor U11960 (N_11960,N_11737,N_11822);
or U11961 (N_11961,N_11715,N_11805);
or U11962 (N_11962,N_11708,N_11832);
or U11963 (N_11963,N_11766,N_11822);
or U11964 (N_11964,N_11681,N_11749);
or U11965 (N_11965,N_11815,N_11682);
and U11966 (N_11966,N_11813,N_11694);
or U11967 (N_11967,N_11687,N_11700);
or U11968 (N_11968,N_11717,N_11698);
or U11969 (N_11969,N_11790,N_11737);
nand U11970 (N_11970,N_11719,N_11811);
xor U11971 (N_11971,N_11718,N_11838);
xor U11972 (N_11972,N_11720,N_11775);
or U11973 (N_11973,N_11694,N_11765);
and U11974 (N_11974,N_11744,N_11720);
or U11975 (N_11975,N_11792,N_11707);
and U11976 (N_11976,N_11697,N_11826);
and U11977 (N_11977,N_11748,N_11817);
nand U11978 (N_11978,N_11748,N_11792);
and U11979 (N_11979,N_11802,N_11809);
nand U11980 (N_11980,N_11758,N_11697);
and U11981 (N_11981,N_11698,N_11690);
nand U11982 (N_11982,N_11780,N_11839);
and U11983 (N_11983,N_11753,N_11838);
nor U11984 (N_11984,N_11827,N_11794);
and U11985 (N_11985,N_11742,N_11789);
nand U11986 (N_11986,N_11801,N_11744);
xnor U11987 (N_11987,N_11688,N_11815);
or U11988 (N_11988,N_11721,N_11689);
and U11989 (N_11989,N_11684,N_11750);
or U11990 (N_11990,N_11696,N_11786);
nand U11991 (N_11991,N_11684,N_11769);
nand U11992 (N_11992,N_11731,N_11720);
nand U11993 (N_11993,N_11825,N_11833);
or U11994 (N_11994,N_11713,N_11705);
nand U11995 (N_11995,N_11757,N_11831);
and U11996 (N_11996,N_11779,N_11752);
nand U11997 (N_11997,N_11715,N_11747);
nand U11998 (N_11998,N_11706,N_11702);
nand U11999 (N_11999,N_11700,N_11784);
nor U12000 (N_12000,N_11993,N_11957);
or U12001 (N_12001,N_11934,N_11919);
nor U12002 (N_12002,N_11987,N_11867);
nand U12003 (N_12003,N_11865,N_11971);
and U12004 (N_12004,N_11899,N_11861);
xor U12005 (N_12005,N_11958,N_11984);
nor U12006 (N_12006,N_11901,N_11983);
or U12007 (N_12007,N_11959,N_11851);
and U12008 (N_12008,N_11963,N_11908);
or U12009 (N_12009,N_11939,N_11858);
nor U12010 (N_12010,N_11859,N_11956);
nand U12011 (N_12011,N_11954,N_11863);
and U12012 (N_12012,N_11970,N_11889);
nand U12013 (N_12013,N_11853,N_11887);
or U12014 (N_12014,N_11982,N_11903);
nor U12015 (N_12015,N_11906,N_11857);
and U12016 (N_12016,N_11980,N_11904);
and U12017 (N_12017,N_11967,N_11925);
xor U12018 (N_12018,N_11926,N_11900);
nand U12019 (N_12019,N_11913,N_11989);
nor U12020 (N_12020,N_11948,N_11860);
or U12021 (N_12021,N_11888,N_11879);
nand U12022 (N_12022,N_11930,N_11933);
nand U12023 (N_12023,N_11931,N_11975);
nor U12024 (N_12024,N_11940,N_11920);
nor U12025 (N_12025,N_11877,N_11962);
nor U12026 (N_12026,N_11976,N_11952);
and U12027 (N_12027,N_11870,N_11951);
and U12028 (N_12028,N_11949,N_11884);
and U12029 (N_12029,N_11872,N_11946);
nor U12030 (N_12030,N_11849,N_11895);
and U12031 (N_12031,N_11922,N_11856);
or U12032 (N_12032,N_11994,N_11846);
or U12033 (N_12033,N_11936,N_11923);
nand U12034 (N_12034,N_11862,N_11950);
nand U12035 (N_12035,N_11842,N_11937);
nor U12036 (N_12036,N_11897,N_11912);
nor U12037 (N_12037,N_11938,N_11964);
xor U12038 (N_12038,N_11840,N_11921);
or U12039 (N_12039,N_11845,N_11990);
and U12040 (N_12040,N_11969,N_11942);
nand U12041 (N_12041,N_11972,N_11960);
nor U12042 (N_12042,N_11896,N_11978);
and U12043 (N_12043,N_11916,N_11991);
nor U12044 (N_12044,N_11873,N_11911);
or U12045 (N_12045,N_11875,N_11947);
and U12046 (N_12046,N_11915,N_11876);
nor U12047 (N_12047,N_11979,N_11905);
or U12048 (N_12048,N_11881,N_11910);
nor U12049 (N_12049,N_11974,N_11883);
nand U12050 (N_12050,N_11882,N_11848);
or U12051 (N_12051,N_11965,N_11924);
or U12052 (N_12052,N_11986,N_11866);
nor U12053 (N_12053,N_11927,N_11995);
or U12054 (N_12054,N_11850,N_11894);
xnor U12055 (N_12055,N_11932,N_11885);
and U12056 (N_12056,N_11941,N_11855);
nand U12057 (N_12057,N_11907,N_11854);
and U12058 (N_12058,N_11868,N_11878);
and U12059 (N_12059,N_11988,N_11928);
xor U12060 (N_12060,N_11852,N_11944);
and U12061 (N_12061,N_11869,N_11871);
or U12062 (N_12062,N_11893,N_11918);
and U12063 (N_12063,N_11945,N_11841);
nand U12064 (N_12064,N_11968,N_11917);
nor U12065 (N_12065,N_11864,N_11890);
nand U12066 (N_12066,N_11953,N_11955);
xnor U12067 (N_12067,N_11847,N_11935);
xnor U12068 (N_12068,N_11909,N_11898);
nor U12069 (N_12069,N_11996,N_11843);
xor U12070 (N_12070,N_11985,N_11943);
nand U12071 (N_12071,N_11844,N_11929);
xor U12072 (N_12072,N_11966,N_11914);
nor U12073 (N_12073,N_11902,N_11973);
nand U12074 (N_12074,N_11981,N_11977);
or U12075 (N_12075,N_11997,N_11892);
and U12076 (N_12076,N_11961,N_11886);
or U12077 (N_12077,N_11891,N_11999);
nand U12078 (N_12078,N_11992,N_11998);
nor U12079 (N_12079,N_11880,N_11874);
nor U12080 (N_12080,N_11943,N_11879);
or U12081 (N_12081,N_11952,N_11897);
and U12082 (N_12082,N_11892,N_11999);
and U12083 (N_12083,N_11845,N_11956);
nor U12084 (N_12084,N_11922,N_11984);
nor U12085 (N_12085,N_11932,N_11902);
and U12086 (N_12086,N_11994,N_11954);
nor U12087 (N_12087,N_11845,N_11890);
xor U12088 (N_12088,N_11990,N_11853);
xor U12089 (N_12089,N_11890,N_11936);
and U12090 (N_12090,N_11910,N_11913);
nor U12091 (N_12091,N_11878,N_11894);
nor U12092 (N_12092,N_11998,N_11934);
xnor U12093 (N_12093,N_11965,N_11876);
nor U12094 (N_12094,N_11919,N_11859);
nor U12095 (N_12095,N_11912,N_11899);
nand U12096 (N_12096,N_11864,N_11971);
nor U12097 (N_12097,N_11942,N_11977);
nand U12098 (N_12098,N_11873,N_11868);
or U12099 (N_12099,N_11904,N_11915);
xor U12100 (N_12100,N_11884,N_11875);
nor U12101 (N_12101,N_11865,N_11937);
nand U12102 (N_12102,N_11942,N_11862);
and U12103 (N_12103,N_11993,N_11863);
nand U12104 (N_12104,N_11913,N_11856);
and U12105 (N_12105,N_11917,N_11846);
nor U12106 (N_12106,N_11950,N_11969);
and U12107 (N_12107,N_11957,N_11848);
and U12108 (N_12108,N_11850,N_11911);
xor U12109 (N_12109,N_11885,N_11874);
nand U12110 (N_12110,N_11877,N_11840);
nor U12111 (N_12111,N_11933,N_11881);
nor U12112 (N_12112,N_11907,N_11903);
nand U12113 (N_12113,N_11878,N_11984);
nor U12114 (N_12114,N_11878,N_11870);
or U12115 (N_12115,N_11907,N_11884);
and U12116 (N_12116,N_11849,N_11969);
or U12117 (N_12117,N_11878,N_11917);
nand U12118 (N_12118,N_11996,N_11980);
or U12119 (N_12119,N_11934,N_11945);
nand U12120 (N_12120,N_11850,N_11865);
xor U12121 (N_12121,N_11888,N_11992);
or U12122 (N_12122,N_11887,N_11979);
nand U12123 (N_12123,N_11938,N_11999);
or U12124 (N_12124,N_11852,N_11967);
nand U12125 (N_12125,N_11953,N_11945);
nand U12126 (N_12126,N_11961,N_11993);
nor U12127 (N_12127,N_11940,N_11858);
nand U12128 (N_12128,N_11945,N_11954);
nand U12129 (N_12129,N_11847,N_11939);
and U12130 (N_12130,N_11990,N_11968);
nor U12131 (N_12131,N_11939,N_11927);
or U12132 (N_12132,N_11855,N_11930);
nand U12133 (N_12133,N_11907,N_11883);
nor U12134 (N_12134,N_11958,N_11898);
nand U12135 (N_12135,N_11938,N_11849);
nor U12136 (N_12136,N_11903,N_11988);
nor U12137 (N_12137,N_11946,N_11843);
nand U12138 (N_12138,N_11927,N_11969);
nor U12139 (N_12139,N_11995,N_11982);
or U12140 (N_12140,N_11858,N_11930);
nor U12141 (N_12141,N_11942,N_11974);
or U12142 (N_12142,N_11938,N_11887);
and U12143 (N_12143,N_11988,N_11865);
nand U12144 (N_12144,N_11964,N_11986);
nor U12145 (N_12145,N_11914,N_11872);
nor U12146 (N_12146,N_11951,N_11904);
nand U12147 (N_12147,N_11891,N_11853);
nor U12148 (N_12148,N_11960,N_11874);
or U12149 (N_12149,N_11928,N_11884);
or U12150 (N_12150,N_11867,N_11953);
and U12151 (N_12151,N_11923,N_11998);
nor U12152 (N_12152,N_11947,N_11962);
nor U12153 (N_12153,N_11996,N_11904);
and U12154 (N_12154,N_11868,N_11965);
nor U12155 (N_12155,N_11922,N_11885);
xnor U12156 (N_12156,N_11962,N_11860);
xnor U12157 (N_12157,N_11840,N_11941);
nand U12158 (N_12158,N_11905,N_11906);
nand U12159 (N_12159,N_11881,N_11861);
or U12160 (N_12160,N_12004,N_12149);
nor U12161 (N_12161,N_12124,N_12054);
and U12162 (N_12162,N_12001,N_12013);
and U12163 (N_12163,N_12040,N_12112);
nand U12164 (N_12164,N_12121,N_12016);
nor U12165 (N_12165,N_12103,N_12147);
nor U12166 (N_12166,N_12085,N_12025);
or U12167 (N_12167,N_12041,N_12074);
or U12168 (N_12168,N_12106,N_12063);
xnor U12169 (N_12169,N_12023,N_12066);
and U12170 (N_12170,N_12120,N_12032);
and U12171 (N_12171,N_12005,N_12044);
or U12172 (N_12172,N_12037,N_12102);
xnor U12173 (N_12173,N_12104,N_12077);
and U12174 (N_12174,N_12086,N_12030);
and U12175 (N_12175,N_12158,N_12123);
xnor U12176 (N_12176,N_12056,N_12081);
and U12177 (N_12177,N_12118,N_12130);
or U12178 (N_12178,N_12003,N_12115);
and U12179 (N_12179,N_12065,N_12072);
nand U12180 (N_12180,N_12026,N_12052);
and U12181 (N_12181,N_12034,N_12138);
xor U12182 (N_12182,N_12092,N_12133);
or U12183 (N_12183,N_12129,N_12036);
nand U12184 (N_12184,N_12064,N_12159);
or U12185 (N_12185,N_12020,N_12101);
and U12186 (N_12186,N_12019,N_12084);
and U12187 (N_12187,N_12117,N_12058);
or U12188 (N_12188,N_12132,N_12039);
nor U12189 (N_12189,N_12009,N_12049);
nor U12190 (N_12190,N_12154,N_12038);
or U12191 (N_12191,N_12057,N_12151);
xor U12192 (N_12192,N_12033,N_12119);
nand U12193 (N_12193,N_12015,N_12135);
nand U12194 (N_12194,N_12029,N_12073);
nand U12195 (N_12195,N_12091,N_12035);
xnor U12196 (N_12196,N_12126,N_12143);
and U12197 (N_12197,N_12137,N_12122);
and U12198 (N_12198,N_12002,N_12146);
nor U12199 (N_12199,N_12097,N_12078);
or U12200 (N_12200,N_12110,N_12024);
nor U12201 (N_12201,N_12080,N_12082);
or U12202 (N_12202,N_12067,N_12021);
nand U12203 (N_12203,N_12145,N_12141);
or U12204 (N_12204,N_12107,N_12155);
and U12205 (N_12205,N_12087,N_12150);
nor U12206 (N_12206,N_12089,N_12042);
nand U12207 (N_12207,N_12010,N_12014);
and U12208 (N_12208,N_12060,N_12047);
xor U12209 (N_12209,N_12051,N_12006);
and U12210 (N_12210,N_12157,N_12027);
xnor U12211 (N_12211,N_12144,N_12011);
nor U12212 (N_12212,N_12093,N_12070);
or U12213 (N_12213,N_12007,N_12045);
or U12214 (N_12214,N_12125,N_12152);
or U12215 (N_12215,N_12094,N_12055);
nor U12216 (N_12216,N_12140,N_12053);
or U12217 (N_12217,N_12090,N_12127);
or U12218 (N_12218,N_12068,N_12088);
nor U12219 (N_12219,N_12156,N_12018);
nor U12220 (N_12220,N_12069,N_12031);
and U12221 (N_12221,N_12075,N_12100);
xor U12222 (N_12222,N_12028,N_12142);
nand U12223 (N_12223,N_12062,N_12043);
and U12224 (N_12224,N_12046,N_12134);
and U12225 (N_12225,N_12048,N_12083);
and U12226 (N_12226,N_12061,N_12079);
nor U12227 (N_12227,N_12012,N_12113);
xor U12228 (N_12228,N_12099,N_12116);
nand U12229 (N_12229,N_12153,N_12059);
and U12230 (N_12230,N_12095,N_12131);
or U12231 (N_12231,N_12096,N_12111);
nor U12232 (N_12232,N_12109,N_12105);
nand U12233 (N_12233,N_12050,N_12128);
nor U12234 (N_12234,N_12071,N_12136);
xor U12235 (N_12235,N_12108,N_12139);
and U12236 (N_12236,N_12076,N_12000);
nand U12237 (N_12237,N_12148,N_12008);
and U12238 (N_12238,N_12022,N_12098);
nand U12239 (N_12239,N_12114,N_12017);
or U12240 (N_12240,N_12058,N_12033);
and U12241 (N_12241,N_12153,N_12117);
or U12242 (N_12242,N_12020,N_12118);
and U12243 (N_12243,N_12137,N_12073);
nor U12244 (N_12244,N_12121,N_12109);
nor U12245 (N_12245,N_12138,N_12123);
nand U12246 (N_12246,N_12031,N_12014);
xnor U12247 (N_12247,N_12133,N_12130);
nand U12248 (N_12248,N_12059,N_12156);
and U12249 (N_12249,N_12068,N_12143);
xor U12250 (N_12250,N_12009,N_12034);
nand U12251 (N_12251,N_12014,N_12016);
xor U12252 (N_12252,N_12147,N_12102);
or U12253 (N_12253,N_12028,N_12076);
nor U12254 (N_12254,N_12051,N_12078);
xnor U12255 (N_12255,N_12088,N_12041);
nand U12256 (N_12256,N_12019,N_12063);
and U12257 (N_12257,N_12098,N_12044);
xnor U12258 (N_12258,N_12041,N_12022);
nor U12259 (N_12259,N_12115,N_12035);
xor U12260 (N_12260,N_12149,N_12071);
nand U12261 (N_12261,N_12106,N_12089);
and U12262 (N_12262,N_12057,N_12102);
nand U12263 (N_12263,N_12072,N_12015);
nor U12264 (N_12264,N_12107,N_12149);
nand U12265 (N_12265,N_12120,N_12117);
nor U12266 (N_12266,N_12143,N_12019);
and U12267 (N_12267,N_12149,N_12104);
nor U12268 (N_12268,N_12126,N_12055);
nand U12269 (N_12269,N_12013,N_12123);
nor U12270 (N_12270,N_12143,N_12061);
xor U12271 (N_12271,N_12040,N_12093);
and U12272 (N_12272,N_12073,N_12080);
nand U12273 (N_12273,N_12122,N_12002);
and U12274 (N_12274,N_12123,N_12050);
nand U12275 (N_12275,N_12069,N_12030);
nand U12276 (N_12276,N_12004,N_12120);
or U12277 (N_12277,N_12129,N_12052);
or U12278 (N_12278,N_12128,N_12001);
or U12279 (N_12279,N_12126,N_12022);
nand U12280 (N_12280,N_12107,N_12147);
or U12281 (N_12281,N_12075,N_12055);
and U12282 (N_12282,N_12114,N_12005);
nor U12283 (N_12283,N_12004,N_12023);
or U12284 (N_12284,N_12053,N_12146);
or U12285 (N_12285,N_12132,N_12023);
or U12286 (N_12286,N_12068,N_12013);
nand U12287 (N_12287,N_12057,N_12007);
and U12288 (N_12288,N_12092,N_12121);
and U12289 (N_12289,N_12107,N_12078);
nand U12290 (N_12290,N_12077,N_12066);
nor U12291 (N_12291,N_12058,N_12018);
nor U12292 (N_12292,N_12132,N_12122);
and U12293 (N_12293,N_12106,N_12147);
or U12294 (N_12294,N_12123,N_12093);
nor U12295 (N_12295,N_12129,N_12011);
or U12296 (N_12296,N_12137,N_12023);
xnor U12297 (N_12297,N_12005,N_12020);
and U12298 (N_12298,N_12113,N_12060);
nor U12299 (N_12299,N_12018,N_12013);
or U12300 (N_12300,N_12010,N_12002);
nand U12301 (N_12301,N_12107,N_12023);
or U12302 (N_12302,N_12009,N_12014);
and U12303 (N_12303,N_12084,N_12151);
nor U12304 (N_12304,N_12110,N_12084);
nor U12305 (N_12305,N_12039,N_12032);
or U12306 (N_12306,N_12023,N_12094);
nand U12307 (N_12307,N_12118,N_12045);
and U12308 (N_12308,N_12001,N_12125);
nand U12309 (N_12309,N_12063,N_12069);
and U12310 (N_12310,N_12145,N_12060);
or U12311 (N_12311,N_12104,N_12006);
or U12312 (N_12312,N_12120,N_12072);
and U12313 (N_12313,N_12158,N_12009);
or U12314 (N_12314,N_12154,N_12153);
nor U12315 (N_12315,N_12106,N_12141);
xnor U12316 (N_12316,N_12119,N_12131);
and U12317 (N_12317,N_12152,N_12046);
xor U12318 (N_12318,N_12020,N_12030);
and U12319 (N_12319,N_12121,N_12028);
or U12320 (N_12320,N_12307,N_12186);
nor U12321 (N_12321,N_12274,N_12257);
and U12322 (N_12322,N_12208,N_12210);
and U12323 (N_12323,N_12271,N_12230);
and U12324 (N_12324,N_12308,N_12213);
nor U12325 (N_12325,N_12317,N_12223);
nand U12326 (N_12326,N_12225,N_12215);
nor U12327 (N_12327,N_12286,N_12184);
and U12328 (N_12328,N_12233,N_12236);
nor U12329 (N_12329,N_12250,N_12194);
or U12330 (N_12330,N_12174,N_12240);
nor U12331 (N_12331,N_12277,N_12221);
xor U12332 (N_12332,N_12243,N_12259);
or U12333 (N_12333,N_12183,N_12193);
nor U12334 (N_12334,N_12198,N_12226);
or U12335 (N_12335,N_12246,N_12217);
nor U12336 (N_12336,N_12278,N_12241);
nand U12337 (N_12337,N_12216,N_12310);
and U12338 (N_12338,N_12173,N_12172);
nor U12339 (N_12339,N_12202,N_12228);
or U12340 (N_12340,N_12290,N_12287);
nand U12341 (N_12341,N_12247,N_12268);
xor U12342 (N_12342,N_12197,N_12251);
nand U12343 (N_12343,N_12249,N_12199);
xor U12344 (N_12344,N_12205,N_12179);
nor U12345 (N_12345,N_12220,N_12315);
xor U12346 (N_12346,N_12188,N_12176);
or U12347 (N_12347,N_12298,N_12244);
xnor U12348 (N_12348,N_12314,N_12185);
nand U12349 (N_12349,N_12239,N_12235);
xnor U12350 (N_12350,N_12304,N_12171);
or U12351 (N_12351,N_12201,N_12309);
nor U12352 (N_12352,N_12252,N_12165);
and U12353 (N_12353,N_12318,N_12262);
and U12354 (N_12354,N_12245,N_12264);
nand U12355 (N_12355,N_12203,N_12311);
nor U12356 (N_12356,N_12234,N_12196);
and U12357 (N_12357,N_12238,N_12276);
and U12358 (N_12358,N_12182,N_12285);
or U12359 (N_12359,N_12232,N_12167);
nor U12360 (N_12360,N_12207,N_12316);
or U12361 (N_12361,N_12218,N_12248);
or U12362 (N_12362,N_12283,N_12296);
and U12363 (N_12363,N_12293,N_12253);
and U12364 (N_12364,N_12229,N_12260);
or U12365 (N_12365,N_12291,N_12195);
or U12366 (N_12366,N_12168,N_12255);
or U12367 (N_12367,N_12180,N_12292);
xnor U12368 (N_12368,N_12279,N_12200);
and U12369 (N_12369,N_12313,N_12222);
xnor U12370 (N_12370,N_12164,N_12319);
nor U12371 (N_12371,N_12299,N_12281);
xnor U12372 (N_12372,N_12302,N_12206);
nor U12373 (N_12373,N_12219,N_12161);
nor U12374 (N_12374,N_12270,N_12288);
and U12375 (N_12375,N_12231,N_12294);
nand U12376 (N_12376,N_12312,N_12263);
xor U12377 (N_12377,N_12160,N_12211);
nor U12378 (N_12378,N_12190,N_12178);
nand U12379 (N_12379,N_12169,N_12297);
and U12380 (N_12380,N_12191,N_12181);
and U12381 (N_12381,N_12162,N_12212);
nand U12382 (N_12382,N_12300,N_12187);
nor U12383 (N_12383,N_12204,N_12289);
and U12384 (N_12384,N_12306,N_12258);
nor U12385 (N_12385,N_12166,N_12273);
nor U12386 (N_12386,N_12192,N_12254);
nor U12387 (N_12387,N_12267,N_12177);
or U12388 (N_12388,N_12280,N_12242);
or U12389 (N_12389,N_12284,N_12275);
nor U12390 (N_12390,N_12256,N_12269);
nand U12391 (N_12391,N_12301,N_12261);
and U12392 (N_12392,N_12272,N_12305);
or U12393 (N_12393,N_12170,N_12209);
and U12394 (N_12394,N_12189,N_12237);
and U12395 (N_12395,N_12266,N_12214);
nand U12396 (N_12396,N_12295,N_12265);
xnor U12397 (N_12397,N_12163,N_12175);
nor U12398 (N_12398,N_12282,N_12303);
nand U12399 (N_12399,N_12224,N_12227);
nor U12400 (N_12400,N_12206,N_12229);
nand U12401 (N_12401,N_12184,N_12160);
nand U12402 (N_12402,N_12306,N_12196);
nor U12403 (N_12403,N_12298,N_12166);
xnor U12404 (N_12404,N_12280,N_12217);
or U12405 (N_12405,N_12278,N_12236);
and U12406 (N_12406,N_12229,N_12304);
and U12407 (N_12407,N_12289,N_12279);
or U12408 (N_12408,N_12300,N_12279);
or U12409 (N_12409,N_12248,N_12295);
and U12410 (N_12410,N_12258,N_12277);
and U12411 (N_12411,N_12162,N_12280);
nor U12412 (N_12412,N_12223,N_12256);
or U12413 (N_12413,N_12238,N_12211);
xor U12414 (N_12414,N_12187,N_12227);
nor U12415 (N_12415,N_12247,N_12210);
and U12416 (N_12416,N_12193,N_12218);
xor U12417 (N_12417,N_12239,N_12224);
nand U12418 (N_12418,N_12219,N_12223);
nand U12419 (N_12419,N_12242,N_12199);
or U12420 (N_12420,N_12309,N_12193);
nand U12421 (N_12421,N_12240,N_12239);
nor U12422 (N_12422,N_12185,N_12287);
nand U12423 (N_12423,N_12255,N_12160);
nand U12424 (N_12424,N_12249,N_12248);
nand U12425 (N_12425,N_12218,N_12264);
nor U12426 (N_12426,N_12217,N_12238);
or U12427 (N_12427,N_12304,N_12240);
nand U12428 (N_12428,N_12193,N_12317);
or U12429 (N_12429,N_12302,N_12192);
nand U12430 (N_12430,N_12309,N_12165);
and U12431 (N_12431,N_12214,N_12228);
nand U12432 (N_12432,N_12275,N_12240);
xnor U12433 (N_12433,N_12299,N_12170);
nor U12434 (N_12434,N_12297,N_12192);
and U12435 (N_12435,N_12267,N_12309);
and U12436 (N_12436,N_12244,N_12176);
or U12437 (N_12437,N_12197,N_12261);
nand U12438 (N_12438,N_12262,N_12309);
or U12439 (N_12439,N_12200,N_12171);
or U12440 (N_12440,N_12254,N_12315);
nor U12441 (N_12441,N_12220,N_12219);
xnor U12442 (N_12442,N_12231,N_12187);
or U12443 (N_12443,N_12204,N_12288);
and U12444 (N_12444,N_12318,N_12298);
and U12445 (N_12445,N_12282,N_12182);
nand U12446 (N_12446,N_12278,N_12287);
nor U12447 (N_12447,N_12198,N_12189);
xnor U12448 (N_12448,N_12292,N_12290);
nor U12449 (N_12449,N_12270,N_12316);
and U12450 (N_12450,N_12241,N_12283);
nor U12451 (N_12451,N_12160,N_12218);
nand U12452 (N_12452,N_12262,N_12161);
or U12453 (N_12453,N_12249,N_12177);
or U12454 (N_12454,N_12212,N_12176);
nor U12455 (N_12455,N_12258,N_12299);
nand U12456 (N_12456,N_12173,N_12311);
and U12457 (N_12457,N_12256,N_12317);
nand U12458 (N_12458,N_12259,N_12278);
and U12459 (N_12459,N_12280,N_12265);
or U12460 (N_12460,N_12254,N_12308);
nor U12461 (N_12461,N_12280,N_12240);
nand U12462 (N_12462,N_12195,N_12286);
and U12463 (N_12463,N_12187,N_12258);
nand U12464 (N_12464,N_12272,N_12299);
and U12465 (N_12465,N_12271,N_12169);
nand U12466 (N_12466,N_12195,N_12308);
nor U12467 (N_12467,N_12212,N_12181);
and U12468 (N_12468,N_12226,N_12247);
nand U12469 (N_12469,N_12312,N_12229);
nand U12470 (N_12470,N_12207,N_12308);
xor U12471 (N_12471,N_12232,N_12198);
or U12472 (N_12472,N_12204,N_12196);
nor U12473 (N_12473,N_12246,N_12185);
or U12474 (N_12474,N_12302,N_12300);
or U12475 (N_12475,N_12290,N_12275);
nor U12476 (N_12476,N_12184,N_12266);
and U12477 (N_12477,N_12262,N_12185);
or U12478 (N_12478,N_12163,N_12236);
or U12479 (N_12479,N_12248,N_12250);
or U12480 (N_12480,N_12331,N_12328);
and U12481 (N_12481,N_12424,N_12341);
xnor U12482 (N_12482,N_12324,N_12459);
nor U12483 (N_12483,N_12445,N_12414);
and U12484 (N_12484,N_12373,N_12405);
and U12485 (N_12485,N_12332,N_12382);
or U12486 (N_12486,N_12327,N_12384);
and U12487 (N_12487,N_12419,N_12329);
nand U12488 (N_12488,N_12475,N_12379);
xor U12489 (N_12489,N_12348,N_12362);
nand U12490 (N_12490,N_12385,N_12444);
nor U12491 (N_12491,N_12374,N_12402);
nor U12492 (N_12492,N_12342,N_12352);
nor U12493 (N_12493,N_12432,N_12418);
xnor U12494 (N_12494,N_12359,N_12433);
or U12495 (N_12495,N_12410,N_12389);
or U12496 (N_12496,N_12467,N_12436);
or U12497 (N_12497,N_12361,N_12322);
xor U12498 (N_12498,N_12453,N_12439);
nand U12499 (N_12499,N_12372,N_12425);
nand U12500 (N_12500,N_12451,N_12360);
nor U12501 (N_12501,N_12441,N_12465);
and U12502 (N_12502,N_12367,N_12429);
xor U12503 (N_12503,N_12466,N_12357);
and U12504 (N_12504,N_12407,N_12428);
nand U12505 (N_12505,N_12448,N_12371);
nor U12506 (N_12506,N_12469,N_12454);
or U12507 (N_12507,N_12394,N_12447);
nand U12508 (N_12508,N_12399,N_12345);
nand U12509 (N_12509,N_12411,N_12435);
nor U12510 (N_12510,N_12395,N_12350);
or U12511 (N_12511,N_12463,N_12403);
or U12512 (N_12512,N_12438,N_12416);
nor U12513 (N_12513,N_12449,N_12380);
nand U12514 (N_12514,N_12366,N_12386);
or U12515 (N_12515,N_12381,N_12456);
nand U12516 (N_12516,N_12458,N_12423);
xor U12517 (N_12517,N_12408,N_12370);
or U12518 (N_12518,N_12337,N_12471);
or U12519 (N_12519,N_12462,N_12404);
nand U12520 (N_12520,N_12461,N_12434);
nor U12521 (N_12521,N_12457,N_12479);
and U12522 (N_12522,N_12363,N_12365);
xnor U12523 (N_12523,N_12338,N_12476);
nor U12524 (N_12524,N_12412,N_12356);
and U12525 (N_12525,N_12427,N_12358);
nand U12526 (N_12526,N_12344,N_12392);
and U12527 (N_12527,N_12450,N_12452);
nor U12528 (N_12528,N_12478,N_12325);
nand U12529 (N_12529,N_12470,N_12472);
and U12530 (N_12530,N_12406,N_12323);
and U12531 (N_12531,N_12383,N_12354);
nor U12532 (N_12532,N_12388,N_12368);
nor U12533 (N_12533,N_12340,N_12473);
or U12534 (N_12534,N_12339,N_12378);
and U12535 (N_12535,N_12398,N_12376);
xnor U12536 (N_12536,N_12443,N_12336);
and U12537 (N_12537,N_12349,N_12417);
nor U12538 (N_12538,N_12431,N_12377);
nor U12539 (N_12539,N_12421,N_12397);
nand U12540 (N_12540,N_12330,N_12364);
and U12541 (N_12541,N_12415,N_12477);
nor U12542 (N_12542,N_12334,N_12353);
and U12543 (N_12543,N_12321,N_12369);
or U12544 (N_12544,N_12326,N_12440);
nand U12545 (N_12545,N_12375,N_12346);
and U12546 (N_12546,N_12409,N_12468);
and U12547 (N_12547,N_12347,N_12400);
nor U12548 (N_12548,N_12355,N_12442);
nor U12549 (N_12549,N_12396,N_12420);
nor U12550 (N_12550,N_12430,N_12446);
or U12551 (N_12551,N_12401,N_12391);
nor U12552 (N_12552,N_12455,N_12474);
or U12553 (N_12553,N_12437,N_12343);
nand U12554 (N_12554,N_12460,N_12351);
or U12555 (N_12555,N_12387,N_12390);
nand U12556 (N_12556,N_12422,N_12335);
xnor U12557 (N_12557,N_12320,N_12393);
nor U12558 (N_12558,N_12413,N_12333);
nor U12559 (N_12559,N_12426,N_12464);
or U12560 (N_12560,N_12461,N_12421);
nor U12561 (N_12561,N_12448,N_12387);
nand U12562 (N_12562,N_12395,N_12399);
nor U12563 (N_12563,N_12475,N_12463);
nor U12564 (N_12564,N_12342,N_12351);
and U12565 (N_12565,N_12472,N_12330);
nor U12566 (N_12566,N_12427,N_12340);
xnor U12567 (N_12567,N_12354,N_12438);
xor U12568 (N_12568,N_12477,N_12381);
and U12569 (N_12569,N_12431,N_12475);
or U12570 (N_12570,N_12326,N_12365);
nand U12571 (N_12571,N_12408,N_12448);
nand U12572 (N_12572,N_12338,N_12441);
nor U12573 (N_12573,N_12428,N_12430);
nor U12574 (N_12574,N_12437,N_12422);
nor U12575 (N_12575,N_12456,N_12394);
and U12576 (N_12576,N_12346,N_12411);
nor U12577 (N_12577,N_12369,N_12408);
xnor U12578 (N_12578,N_12475,N_12453);
nor U12579 (N_12579,N_12370,N_12336);
or U12580 (N_12580,N_12359,N_12426);
or U12581 (N_12581,N_12445,N_12444);
and U12582 (N_12582,N_12399,N_12420);
and U12583 (N_12583,N_12413,N_12345);
and U12584 (N_12584,N_12445,N_12434);
or U12585 (N_12585,N_12450,N_12374);
nand U12586 (N_12586,N_12402,N_12430);
or U12587 (N_12587,N_12381,N_12414);
and U12588 (N_12588,N_12370,N_12414);
xnor U12589 (N_12589,N_12346,N_12407);
nor U12590 (N_12590,N_12366,N_12404);
and U12591 (N_12591,N_12440,N_12467);
and U12592 (N_12592,N_12413,N_12455);
nor U12593 (N_12593,N_12464,N_12453);
or U12594 (N_12594,N_12359,N_12377);
and U12595 (N_12595,N_12364,N_12353);
and U12596 (N_12596,N_12329,N_12415);
or U12597 (N_12597,N_12433,N_12437);
nor U12598 (N_12598,N_12337,N_12462);
or U12599 (N_12599,N_12432,N_12421);
or U12600 (N_12600,N_12382,N_12467);
nand U12601 (N_12601,N_12445,N_12385);
nor U12602 (N_12602,N_12446,N_12394);
nand U12603 (N_12603,N_12338,N_12333);
nand U12604 (N_12604,N_12347,N_12391);
nor U12605 (N_12605,N_12447,N_12401);
or U12606 (N_12606,N_12409,N_12440);
or U12607 (N_12607,N_12431,N_12386);
and U12608 (N_12608,N_12460,N_12391);
and U12609 (N_12609,N_12425,N_12460);
nor U12610 (N_12610,N_12391,N_12350);
nor U12611 (N_12611,N_12479,N_12341);
or U12612 (N_12612,N_12345,N_12429);
or U12613 (N_12613,N_12344,N_12454);
and U12614 (N_12614,N_12356,N_12436);
and U12615 (N_12615,N_12435,N_12384);
nor U12616 (N_12616,N_12412,N_12346);
nor U12617 (N_12617,N_12440,N_12367);
nor U12618 (N_12618,N_12330,N_12347);
nor U12619 (N_12619,N_12370,N_12335);
or U12620 (N_12620,N_12456,N_12345);
nand U12621 (N_12621,N_12464,N_12391);
and U12622 (N_12622,N_12328,N_12400);
nand U12623 (N_12623,N_12355,N_12429);
nor U12624 (N_12624,N_12409,N_12343);
or U12625 (N_12625,N_12331,N_12321);
or U12626 (N_12626,N_12361,N_12473);
nand U12627 (N_12627,N_12385,N_12379);
and U12628 (N_12628,N_12355,N_12330);
nand U12629 (N_12629,N_12424,N_12440);
and U12630 (N_12630,N_12419,N_12388);
xor U12631 (N_12631,N_12353,N_12345);
nor U12632 (N_12632,N_12425,N_12391);
or U12633 (N_12633,N_12357,N_12380);
or U12634 (N_12634,N_12349,N_12334);
or U12635 (N_12635,N_12409,N_12320);
nor U12636 (N_12636,N_12406,N_12351);
nand U12637 (N_12637,N_12438,N_12358);
nor U12638 (N_12638,N_12458,N_12330);
or U12639 (N_12639,N_12442,N_12430);
nor U12640 (N_12640,N_12495,N_12589);
xnor U12641 (N_12641,N_12578,N_12590);
nand U12642 (N_12642,N_12569,N_12546);
nor U12643 (N_12643,N_12605,N_12595);
or U12644 (N_12644,N_12586,N_12513);
nor U12645 (N_12645,N_12549,N_12585);
nor U12646 (N_12646,N_12543,N_12524);
and U12647 (N_12647,N_12512,N_12594);
or U12648 (N_12648,N_12529,N_12542);
nor U12649 (N_12649,N_12591,N_12628);
nand U12650 (N_12650,N_12631,N_12550);
nand U12651 (N_12651,N_12532,N_12600);
or U12652 (N_12652,N_12526,N_12564);
and U12653 (N_12653,N_12519,N_12567);
nand U12654 (N_12654,N_12575,N_12560);
xor U12655 (N_12655,N_12622,N_12563);
or U12656 (N_12656,N_12619,N_12566);
nor U12657 (N_12657,N_12593,N_12584);
nor U12658 (N_12658,N_12485,N_12573);
nand U12659 (N_12659,N_12535,N_12638);
nor U12660 (N_12660,N_12603,N_12636);
and U12661 (N_12661,N_12576,N_12557);
or U12662 (N_12662,N_12499,N_12506);
and U12663 (N_12663,N_12612,N_12624);
and U12664 (N_12664,N_12606,N_12553);
nor U12665 (N_12665,N_12486,N_12497);
or U12666 (N_12666,N_12551,N_12601);
nor U12667 (N_12667,N_12492,N_12599);
nand U12668 (N_12668,N_12500,N_12637);
nor U12669 (N_12669,N_12533,N_12587);
nor U12670 (N_12670,N_12487,N_12579);
and U12671 (N_12671,N_12490,N_12496);
xnor U12672 (N_12672,N_12536,N_12608);
and U12673 (N_12673,N_12482,N_12534);
nor U12674 (N_12674,N_12583,N_12558);
nor U12675 (N_12675,N_12607,N_12616);
nand U12676 (N_12676,N_12507,N_12597);
nand U12677 (N_12677,N_12627,N_12484);
nor U12678 (N_12678,N_12625,N_12538);
and U12679 (N_12679,N_12555,N_12531);
xnor U12680 (N_12680,N_12503,N_12525);
and U12681 (N_12681,N_12633,N_12509);
and U12682 (N_12682,N_12618,N_12632);
and U12683 (N_12683,N_12494,N_12518);
nand U12684 (N_12684,N_12491,N_12520);
and U12685 (N_12685,N_12515,N_12611);
or U12686 (N_12686,N_12489,N_12565);
nor U12687 (N_12687,N_12604,N_12562);
nand U12688 (N_12688,N_12544,N_12545);
or U12689 (N_12689,N_12623,N_12501);
nand U12690 (N_12690,N_12556,N_12571);
or U12691 (N_12691,N_12615,N_12630);
and U12692 (N_12692,N_12480,N_12559);
or U12693 (N_12693,N_12554,N_12626);
or U12694 (N_12694,N_12514,N_12521);
and U12695 (N_12695,N_12592,N_12580);
nand U12696 (N_12696,N_12613,N_12481);
and U12697 (N_12697,N_12523,N_12629);
nor U12698 (N_12698,N_12537,N_12602);
or U12699 (N_12699,N_12541,N_12504);
nand U12700 (N_12700,N_12539,N_12547);
nor U12701 (N_12701,N_12570,N_12548);
xor U12702 (N_12702,N_12530,N_12483);
nand U12703 (N_12703,N_12510,N_12634);
nor U12704 (N_12704,N_12540,N_12517);
nor U12705 (N_12705,N_12528,N_12614);
or U12706 (N_12706,N_12582,N_12561);
nand U12707 (N_12707,N_12516,N_12498);
and U12708 (N_12708,N_12493,N_12572);
or U12709 (N_12709,N_12598,N_12635);
or U12710 (N_12710,N_12488,N_12621);
or U12711 (N_12711,N_12505,N_12596);
or U12712 (N_12712,N_12609,N_12522);
nand U12713 (N_12713,N_12508,N_12502);
nand U12714 (N_12714,N_12617,N_12511);
and U12715 (N_12715,N_12574,N_12610);
or U12716 (N_12716,N_12577,N_12568);
nor U12717 (N_12717,N_12620,N_12552);
nor U12718 (N_12718,N_12527,N_12581);
nor U12719 (N_12719,N_12639,N_12588);
or U12720 (N_12720,N_12560,N_12493);
nor U12721 (N_12721,N_12622,N_12609);
nand U12722 (N_12722,N_12621,N_12597);
xor U12723 (N_12723,N_12550,N_12500);
or U12724 (N_12724,N_12613,N_12558);
nor U12725 (N_12725,N_12633,N_12494);
and U12726 (N_12726,N_12505,N_12549);
or U12727 (N_12727,N_12580,N_12562);
and U12728 (N_12728,N_12621,N_12535);
and U12729 (N_12729,N_12576,N_12510);
or U12730 (N_12730,N_12633,N_12620);
nand U12731 (N_12731,N_12612,N_12638);
and U12732 (N_12732,N_12549,N_12566);
or U12733 (N_12733,N_12495,N_12631);
nor U12734 (N_12734,N_12494,N_12504);
or U12735 (N_12735,N_12576,N_12599);
nor U12736 (N_12736,N_12590,N_12522);
or U12737 (N_12737,N_12575,N_12534);
or U12738 (N_12738,N_12595,N_12616);
nor U12739 (N_12739,N_12566,N_12499);
nand U12740 (N_12740,N_12509,N_12571);
xor U12741 (N_12741,N_12615,N_12574);
nor U12742 (N_12742,N_12607,N_12633);
nand U12743 (N_12743,N_12486,N_12569);
and U12744 (N_12744,N_12600,N_12530);
nand U12745 (N_12745,N_12635,N_12607);
nand U12746 (N_12746,N_12510,N_12589);
nor U12747 (N_12747,N_12622,N_12565);
and U12748 (N_12748,N_12628,N_12506);
nor U12749 (N_12749,N_12568,N_12538);
or U12750 (N_12750,N_12612,N_12632);
or U12751 (N_12751,N_12530,N_12569);
nor U12752 (N_12752,N_12625,N_12628);
or U12753 (N_12753,N_12517,N_12570);
xnor U12754 (N_12754,N_12549,N_12514);
or U12755 (N_12755,N_12611,N_12604);
nor U12756 (N_12756,N_12589,N_12609);
and U12757 (N_12757,N_12618,N_12627);
and U12758 (N_12758,N_12618,N_12547);
and U12759 (N_12759,N_12575,N_12594);
and U12760 (N_12760,N_12550,N_12504);
or U12761 (N_12761,N_12638,N_12617);
or U12762 (N_12762,N_12608,N_12488);
nand U12763 (N_12763,N_12558,N_12592);
and U12764 (N_12764,N_12529,N_12634);
nor U12765 (N_12765,N_12606,N_12498);
and U12766 (N_12766,N_12540,N_12608);
or U12767 (N_12767,N_12486,N_12512);
and U12768 (N_12768,N_12625,N_12634);
and U12769 (N_12769,N_12508,N_12498);
nand U12770 (N_12770,N_12571,N_12589);
nor U12771 (N_12771,N_12489,N_12560);
nor U12772 (N_12772,N_12540,N_12593);
xor U12773 (N_12773,N_12534,N_12524);
or U12774 (N_12774,N_12549,N_12551);
nand U12775 (N_12775,N_12583,N_12528);
nor U12776 (N_12776,N_12571,N_12630);
and U12777 (N_12777,N_12514,N_12486);
or U12778 (N_12778,N_12565,N_12628);
nor U12779 (N_12779,N_12494,N_12521);
nand U12780 (N_12780,N_12547,N_12573);
nand U12781 (N_12781,N_12549,N_12632);
or U12782 (N_12782,N_12637,N_12499);
nand U12783 (N_12783,N_12564,N_12532);
nor U12784 (N_12784,N_12556,N_12617);
xnor U12785 (N_12785,N_12598,N_12601);
or U12786 (N_12786,N_12488,N_12494);
nand U12787 (N_12787,N_12484,N_12521);
and U12788 (N_12788,N_12626,N_12589);
nand U12789 (N_12789,N_12540,N_12636);
and U12790 (N_12790,N_12627,N_12557);
nor U12791 (N_12791,N_12637,N_12531);
and U12792 (N_12792,N_12570,N_12567);
and U12793 (N_12793,N_12599,N_12504);
nand U12794 (N_12794,N_12482,N_12491);
nor U12795 (N_12795,N_12597,N_12516);
xnor U12796 (N_12796,N_12544,N_12540);
or U12797 (N_12797,N_12514,N_12594);
xor U12798 (N_12798,N_12626,N_12507);
or U12799 (N_12799,N_12636,N_12495);
and U12800 (N_12800,N_12789,N_12787);
nand U12801 (N_12801,N_12710,N_12716);
and U12802 (N_12802,N_12644,N_12717);
or U12803 (N_12803,N_12677,N_12664);
nor U12804 (N_12804,N_12676,N_12701);
nor U12805 (N_12805,N_12674,N_12654);
xnor U12806 (N_12806,N_12776,N_12779);
xor U12807 (N_12807,N_12780,N_12679);
or U12808 (N_12808,N_12788,N_12772);
nand U12809 (N_12809,N_12689,N_12724);
nand U12810 (N_12810,N_12775,N_12680);
nand U12811 (N_12811,N_12687,N_12798);
xnor U12812 (N_12812,N_12762,N_12714);
or U12813 (N_12813,N_12665,N_12698);
nand U12814 (N_12814,N_12731,N_12748);
or U12815 (N_12815,N_12795,N_12756);
nand U12816 (N_12816,N_12704,N_12686);
or U12817 (N_12817,N_12666,N_12688);
and U12818 (N_12818,N_12723,N_12784);
or U12819 (N_12819,N_12722,N_12759);
and U12820 (N_12820,N_12671,N_12659);
nand U12821 (N_12821,N_12738,N_12643);
and U12822 (N_12822,N_12729,N_12754);
and U12823 (N_12823,N_12708,N_12725);
nand U12824 (N_12824,N_12733,N_12650);
and U12825 (N_12825,N_12757,N_12763);
or U12826 (N_12826,N_12736,N_12790);
nand U12827 (N_12827,N_12669,N_12764);
xnor U12828 (N_12828,N_12656,N_12690);
or U12829 (N_12829,N_12750,N_12770);
nor U12830 (N_12830,N_12660,N_12767);
nor U12831 (N_12831,N_12672,N_12663);
xor U12832 (N_12832,N_12778,N_12658);
nand U12833 (N_12833,N_12715,N_12673);
or U12834 (N_12834,N_12781,N_12683);
nand U12835 (N_12835,N_12703,N_12728);
and U12836 (N_12836,N_12766,N_12734);
and U12837 (N_12837,N_12651,N_12700);
nand U12838 (N_12838,N_12765,N_12670);
and U12839 (N_12839,N_12694,N_12743);
nand U12840 (N_12840,N_12758,N_12741);
or U12841 (N_12841,N_12642,N_12735);
nand U12842 (N_12842,N_12768,N_12684);
nand U12843 (N_12843,N_12773,N_12792);
or U12844 (N_12844,N_12713,N_12727);
and U12845 (N_12845,N_12719,N_12760);
nor U12846 (N_12846,N_12691,N_12712);
nor U12847 (N_12847,N_12747,N_12783);
nor U12848 (N_12848,N_12799,N_12678);
nor U12849 (N_12849,N_12706,N_12797);
and U12850 (N_12850,N_12681,N_12675);
or U12851 (N_12851,N_12696,N_12753);
or U12852 (N_12852,N_12705,N_12782);
and U12853 (N_12853,N_12702,N_12761);
xor U12854 (N_12854,N_12697,N_12661);
or U12855 (N_12855,N_12793,N_12737);
or U12856 (N_12856,N_12742,N_12657);
nor U12857 (N_12857,N_12796,N_12721);
and U12858 (N_12858,N_12777,N_12641);
nor U12859 (N_12859,N_12751,N_12769);
nor U12860 (N_12860,N_12682,N_12699);
and U12861 (N_12861,N_12655,N_12695);
nor U12862 (N_12862,N_12667,N_12692);
nand U12863 (N_12863,N_12653,N_12744);
and U12864 (N_12864,N_12648,N_12649);
nand U12865 (N_12865,N_12739,N_12693);
or U12866 (N_12866,N_12745,N_12640);
nand U12867 (N_12867,N_12645,N_12771);
nor U12868 (N_12868,N_12732,N_12709);
nand U12869 (N_12869,N_12749,N_12662);
and U12870 (N_12870,N_12652,N_12685);
or U12871 (N_12871,N_12752,N_12730);
nand U12872 (N_12872,N_12646,N_12740);
nand U12873 (N_12873,N_12791,N_12794);
or U12874 (N_12874,N_12755,N_12668);
and U12875 (N_12875,N_12746,N_12718);
or U12876 (N_12876,N_12726,N_12711);
and U12877 (N_12877,N_12720,N_12786);
nor U12878 (N_12878,N_12707,N_12647);
and U12879 (N_12879,N_12774,N_12785);
nand U12880 (N_12880,N_12741,N_12744);
and U12881 (N_12881,N_12690,N_12686);
nor U12882 (N_12882,N_12735,N_12750);
nand U12883 (N_12883,N_12792,N_12668);
nand U12884 (N_12884,N_12655,N_12672);
and U12885 (N_12885,N_12694,N_12652);
nand U12886 (N_12886,N_12731,N_12648);
or U12887 (N_12887,N_12642,N_12695);
nor U12888 (N_12888,N_12720,N_12774);
nand U12889 (N_12889,N_12684,N_12696);
and U12890 (N_12890,N_12727,N_12735);
or U12891 (N_12891,N_12678,N_12641);
and U12892 (N_12892,N_12686,N_12792);
nand U12893 (N_12893,N_12740,N_12662);
nor U12894 (N_12894,N_12657,N_12705);
nand U12895 (N_12895,N_12656,N_12789);
and U12896 (N_12896,N_12775,N_12793);
or U12897 (N_12897,N_12731,N_12728);
xnor U12898 (N_12898,N_12677,N_12759);
nor U12899 (N_12899,N_12664,N_12668);
nor U12900 (N_12900,N_12687,N_12796);
xnor U12901 (N_12901,N_12713,N_12663);
and U12902 (N_12902,N_12713,N_12706);
and U12903 (N_12903,N_12758,N_12648);
and U12904 (N_12904,N_12780,N_12666);
or U12905 (N_12905,N_12665,N_12786);
nand U12906 (N_12906,N_12682,N_12693);
nand U12907 (N_12907,N_12793,N_12798);
nand U12908 (N_12908,N_12694,N_12701);
nand U12909 (N_12909,N_12742,N_12680);
or U12910 (N_12910,N_12710,N_12769);
and U12911 (N_12911,N_12665,N_12719);
and U12912 (N_12912,N_12748,N_12674);
and U12913 (N_12913,N_12767,N_12745);
or U12914 (N_12914,N_12720,N_12665);
nor U12915 (N_12915,N_12707,N_12675);
nand U12916 (N_12916,N_12722,N_12690);
nor U12917 (N_12917,N_12640,N_12785);
and U12918 (N_12918,N_12784,N_12687);
or U12919 (N_12919,N_12736,N_12711);
nand U12920 (N_12920,N_12737,N_12710);
xnor U12921 (N_12921,N_12795,N_12743);
or U12922 (N_12922,N_12726,N_12752);
nor U12923 (N_12923,N_12682,N_12684);
and U12924 (N_12924,N_12758,N_12743);
nand U12925 (N_12925,N_12652,N_12660);
or U12926 (N_12926,N_12646,N_12788);
xor U12927 (N_12927,N_12666,N_12733);
or U12928 (N_12928,N_12749,N_12719);
or U12929 (N_12929,N_12666,N_12658);
and U12930 (N_12930,N_12778,N_12665);
and U12931 (N_12931,N_12763,N_12751);
or U12932 (N_12932,N_12658,N_12651);
nand U12933 (N_12933,N_12659,N_12647);
xor U12934 (N_12934,N_12645,N_12769);
nor U12935 (N_12935,N_12756,N_12725);
nor U12936 (N_12936,N_12640,N_12765);
and U12937 (N_12937,N_12748,N_12694);
nor U12938 (N_12938,N_12690,N_12685);
xnor U12939 (N_12939,N_12777,N_12704);
nor U12940 (N_12940,N_12642,N_12665);
or U12941 (N_12941,N_12767,N_12659);
xnor U12942 (N_12942,N_12683,N_12764);
and U12943 (N_12943,N_12744,N_12758);
nand U12944 (N_12944,N_12713,N_12704);
and U12945 (N_12945,N_12660,N_12698);
and U12946 (N_12946,N_12743,N_12740);
and U12947 (N_12947,N_12751,N_12766);
nand U12948 (N_12948,N_12654,N_12787);
or U12949 (N_12949,N_12751,N_12745);
nand U12950 (N_12950,N_12692,N_12702);
and U12951 (N_12951,N_12701,N_12647);
nor U12952 (N_12952,N_12656,N_12724);
or U12953 (N_12953,N_12642,N_12691);
nand U12954 (N_12954,N_12775,N_12686);
nor U12955 (N_12955,N_12727,N_12700);
or U12956 (N_12956,N_12799,N_12772);
nand U12957 (N_12957,N_12762,N_12684);
nand U12958 (N_12958,N_12698,N_12646);
nor U12959 (N_12959,N_12657,N_12754);
and U12960 (N_12960,N_12850,N_12878);
nor U12961 (N_12961,N_12806,N_12862);
nor U12962 (N_12962,N_12934,N_12804);
xor U12963 (N_12963,N_12838,N_12815);
nand U12964 (N_12964,N_12914,N_12887);
and U12965 (N_12965,N_12879,N_12866);
nor U12966 (N_12966,N_12821,N_12864);
or U12967 (N_12967,N_12946,N_12933);
nor U12968 (N_12968,N_12876,N_12855);
nand U12969 (N_12969,N_12834,N_12955);
and U12970 (N_12970,N_12936,N_12863);
nand U12971 (N_12971,N_12822,N_12883);
or U12972 (N_12972,N_12803,N_12836);
nor U12973 (N_12973,N_12837,N_12924);
nand U12974 (N_12974,N_12894,N_12811);
nor U12975 (N_12975,N_12886,N_12865);
and U12976 (N_12976,N_12890,N_12920);
and U12977 (N_12977,N_12927,N_12945);
and U12978 (N_12978,N_12938,N_12948);
and U12979 (N_12979,N_12958,N_12841);
or U12980 (N_12980,N_12859,N_12868);
or U12981 (N_12981,N_12832,N_12826);
nor U12982 (N_12982,N_12930,N_12800);
nand U12983 (N_12983,N_12901,N_12949);
or U12984 (N_12984,N_12898,N_12856);
nand U12985 (N_12985,N_12954,N_12919);
xnor U12986 (N_12986,N_12869,N_12851);
nor U12987 (N_12987,N_12881,N_12874);
or U12988 (N_12988,N_12932,N_12854);
and U12989 (N_12989,N_12833,N_12842);
or U12990 (N_12990,N_12951,N_12912);
nor U12991 (N_12991,N_12873,N_12861);
xor U12992 (N_12992,N_12817,N_12923);
nand U12993 (N_12993,N_12899,N_12950);
nand U12994 (N_12994,N_12902,N_12942);
nor U12995 (N_12995,N_12947,N_12889);
xor U12996 (N_12996,N_12952,N_12840);
and U12997 (N_12997,N_12896,N_12807);
nor U12998 (N_12998,N_12922,N_12845);
nand U12999 (N_12999,N_12941,N_12925);
and U13000 (N_13000,N_12805,N_12953);
or U13001 (N_13001,N_12904,N_12911);
nor U13002 (N_13002,N_12935,N_12944);
nor U13003 (N_13003,N_12929,N_12910);
nand U13004 (N_13004,N_12915,N_12839);
nand U13005 (N_13005,N_12956,N_12917);
and U13006 (N_13006,N_12875,N_12888);
and U13007 (N_13007,N_12957,N_12918);
and U13008 (N_13008,N_12885,N_12871);
xor U13009 (N_13009,N_12931,N_12870);
and U13010 (N_13010,N_12897,N_12816);
and U13011 (N_13011,N_12926,N_12843);
and U13012 (N_13012,N_12895,N_12823);
and U13013 (N_13013,N_12849,N_12846);
nand U13014 (N_13014,N_12882,N_12907);
nor U13015 (N_13015,N_12905,N_12893);
and U13016 (N_13016,N_12857,N_12891);
nor U13017 (N_13017,N_12858,N_12853);
or U13018 (N_13018,N_12808,N_12937);
and U13019 (N_13019,N_12872,N_12900);
and U13020 (N_13020,N_12818,N_12909);
nand U13021 (N_13021,N_12852,N_12814);
and U13022 (N_13022,N_12829,N_12892);
and U13023 (N_13023,N_12844,N_12880);
nand U13024 (N_13024,N_12802,N_12813);
nor U13025 (N_13025,N_12916,N_12903);
nor U13026 (N_13026,N_12809,N_12913);
nand U13027 (N_13027,N_12831,N_12820);
nor U13028 (N_13028,N_12908,N_12812);
xnor U13029 (N_13029,N_12928,N_12860);
or U13030 (N_13030,N_12847,N_12848);
nor U13031 (N_13031,N_12906,N_12825);
and U13032 (N_13032,N_12877,N_12835);
or U13033 (N_13033,N_12828,N_12819);
or U13034 (N_13034,N_12943,N_12867);
xnor U13035 (N_13035,N_12827,N_12921);
or U13036 (N_13036,N_12939,N_12824);
xor U13037 (N_13037,N_12810,N_12830);
nor U13038 (N_13038,N_12959,N_12940);
nand U13039 (N_13039,N_12884,N_12801);
nand U13040 (N_13040,N_12908,N_12909);
or U13041 (N_13041,N_12820,N_12911);
nor U13042 (N_13042,N_12860,N_12939);
and U13043 (N_13043,N_12839,N_12862);
xnor U13044 (N_13044,N_12946,N_12945);
nand U13045 (N_13045,N_12864,N_12860);
nand U13046 (N_13046,N_12888,N_12825);
nand U13047 (N_13047,N_12860,N_12917);
or U13048 (N_13048,N_12925,N_12910);
or U13049 (N_13049,N_12851,N_12842);
and U13050 (N_13050,N_12809,N_12802);
xor U13051 (N_13051,N_12813,N_12848);
and U13052 (N_13052,N_12832,N_12912);
nor U13053 (N_13053,N_12940,N_12924);
nor U13054 (N_13054,N_12855,N_12937);
nand U13055 (N_13055,N_12890,N_12906);
or U13056 (N_13056,N_12822,N_12918);
and U13057 (N_13057,N_12889,N_12812);
nand U13058 (N_13058,N_12869,N_12953);
nor U13059 (N_13059,N_12830,N_12951);
nand U13060 (N_13060,N_12915,N_12908);
or U13061 (N_13061,N_12920,N_12939);
nand U13062 (N_13062,N_12825,N_12882);
and U13063 (N_13063,N_12911,N_12818);
or U13064 (N_13064,N_12941,N_12949);
xor U13065 (N_13065,N_12808,N_12930);
or U13066 (N_13066,N_12879,N_12841);
and U13067 (N_13067,N_12809,N_12903);
xnor U13068 (N_13068,N_12827,N_12911);
xor U13069 (N_13069,N_12860,N_12831);
and U13070 (N_13070,N_12830,N_12923);
nand U13071 (N_13071,N_12934,N_12933);
or U13072 (N_13072,N_12956,N_12947);
xnor U13073 (N_13073,N_12861,N_12823);
or U13074 (N_13074,N_12939,N_12952);
nand U13075 (N_13075,N_12939,N_12874);
xor U13076 (N_13076,N_12835,N_12867);
nand U13077 (N_13077,N_12913,N_12836);
nor U13078 (N_13078,N_12950,N_12941);
nor U13079 (N_13079,N_12919,N_12849);
and U13080 (N_13080,N_12938,N_12829);
or U13081 (N_13081,N_12903,N_12847);
and U13082 (N_13082,N_12936,N_12939);
nor U13083 (N_13083,N_12851,N_12841);
nor U13084 (N_13084,N_12824,N_12883);
or U13085 (N_13085,N_12850,N_12839);
nand U13086 (N_13086,N_12848,N_12873);
or U13087 (N_13087,N_12827,N_12925);
and U13088 (N_13088,N_12867,N_12908);
nor U13089 (N_13089,N_12886,N_12835);
nor U13090 (N_13090,N_12911,N_12941);
xnor U13091 (N_13091,N_12870,N_12845);
and U13092 (N_13092,N_12951,N_12904);
nor U13093 (N_13093,N_12803,N_12864);
or U13094 (N_13094,N_12939,N_12921);
nor U13095 (N_13095,N_12950,N_12822);
nor U13096 (N_13096,N_12888,N_12871);
nand U13097 (N_13097,N_12919,N_12915);
and U13098 (N_13098,N_12825,N_12876);
nor U13099 (N_13099,N_12950,N_12815);
or U13100 (N_13100,N_12839,N_12874);
and U13101 (N_13101,N_12868,N_12882);
nor U13102 (N_13102,N_12873,N_12937);
xnor U13103 (N_13103,N_12813,N_12943);
and U13104 (N_13104,N_12917,N_12821);
nor U13105 (N_13105,N_12940,N_12902);
and U13106 (N_13106,N_12833,N_12930);
nor U13107 (N_13107,N_12805,N_12819);
nand U13108 (N_13108,N_12815,N_12914);
nand U13109 (N_13109,N_12862,N_12869);
nor U13110 (N_13110,N_12864,N_12826);
nand U13111 (N_13111,N_12926,N_12943);
or U13112 (N_13112,N_12900,N_12843);
nor U13113 (N_13113,N_12909,N_12925);
nand U13114 (N_13114,N_12837,N_12951);
nor U13115 (N_13115,N_12909,N_12911);
or U13116 (N_13116,N_12930,N_12907);
or U13117 (N_13117,N_12933,N_12853);
and U13118 (N_13118,N_12861,N_12855);
nand U13119 (N_13119,N_12930,N_12820);
nand U13120 (N_13120,N_12998,N_13113);
nor U13121 (N_13121,N_13070,N_13063);
nand U13122 (N_13122,N_13056,N_13037);
nand U13123 (N_13123,N_12963,N_13031);
xnor U13124 (N_13124,N_13071,N_13006);
or U13125 (N_13125,N_13099,N_13042);
or U13126 (N_13126,N_13021,N_12971);
nand U13127 (N_13127,N_12975,N_12972);
nand U13128 (N_13128,N_13030,N_13036);
nand U13129 (N_13129,N_13053,N_13047);
or U13130 (N_13130,N_13003,N_13092);
nand U13131 (N_13131,N_13107,N_13111);
nand U13132 (N_13132,N_13109,N_13067);
and U13133 (N_13133,N_13068,N_13011);
xnor U13134 (N_13134,N_13075,N_13094);
and U13135 (N_13135,N_12996,N_13052);
nor U13136 (N_13136,N_13086,N_12987);
or U13137 (N_13137,N_13103,N_13096);
or U13138 (N_13138,N_13046,N_13110);
or U13139 (N_13139,N_13015,N_13022);
nor U13140 (N_13140,N_13088,N_13090);
xnor U13141 (N_13141,N_13023,N_13080);
nor U13142 (N_13142,N_12974,N_13095);
nand U13143 (N_13143,N_13084,N_12993);
nor U13144 (N_13144,N_13079,N_13027);
xnor U13145 (N_13145,N_13033,N_13007);
nand U13146 (N_13146,N_13106,N_13116);
or U13147 (N_13147,N_13093,N_13065);
and U13148 (N_13148,N_12967,N_13062);
and U13149 (N_13149,N_13041,N_13057);
nand U13150 (N_13150,N_13034,N_13004);
or U13151 (N_13151,N_13073,N_13016);
nand U13152 (N_13152,N_13100,N_13098);
nand U13153 (N_13153,N_13012,N_13118);
and U13154 (N_13154,N_13025,N_13104);
and U13155 (N_13155,N_13044,N_12976);
or U13156 (N_13156,N_12979,N_12997);
or U13157 (N_13157,N_13020,N_12983);
nand U13158 (N_13158,N_12981,N_13010);
xnor U13159 (N_13159,N_13069,N_13097);
nand U13160 (N_13160,N_12966,N_13089);
nand U13161 (N_13161,N_13051,N_13038);
or U13162 (N_13162,N_12962,N_12980);
or U13163 (N_13163,N_13039,N_12977);
nand U13164 (N_13164,N_13018,N_12984);
and U13165 (N_13165,N_13064,N_13074);
and U13166 (N_13166,N_12989,N_13055);
nand U13167 (N_13167,N_13017,N_12999);
nand U13168 (N_13168,N_13009,N_13028);
nor U13169 (N_13169,N_12968,N_12994);
nor U13170 (N_13170,N_13005,N_13066);
and U13171 (N_13171,N_12991,N_13061);
nand U13172 (N_13172,N_13117,N_12970);
nor U13173 (N_13173,N_12990,N_13058);
and U13174 (N_13174,N_13108,N_13008);
and U13175 (N_13175,N_13076,N_13019);
or U13176 (N_13176,N_13043,N_12964);
nor U13177 (N_13177,N_13082,N_12978);
nor U13178 (N_13178,N_13059,N_13002);
or U13179 (N_13179,N_13085,N_12973);
and U13180 (N_13180,N_13045,N_13081);
and U13181 (N_13181,N_13050,N_13013);
or U13182 (N_13182,N_13102,N_13014);
nor U13183 (N_13183,N_13035,N_13091);
or U13184 (N_13184,N_12992,N_13101);
nand U13185 (N_13185,N_12961,N_13114);
and U13186 (N_13186,N_13072,N_13077);
nor U13187 (N_13187,N_13078,N_13083);
or U13188 (N_13188,N_12969,N_13029);
nand U13189 (N_13189,N_13087,N_12982);
or U13190 (N_13190,N_13119,N_13049);
xor U13191 (N_13191,N_13032,N_13040);
nor U13192 (N_13192,N_12995,N_12985);
and U13193 (N_13193,N_13112,N_12986);
nor U13194 (N_13194,N_13105,N_12960);
nand U13195 (N_13195,N_13054,N_13060);
xnor U13196 (N_13196,N_13001,N_12988);
or U13197 (N_13197,N_13000,N_13115);
or U13198 (N_13198,N_13048,N_13026);
and U13199 (N_13199,N_13024,N_12965);
xor U13200 (N_13200,N_13036,N_13024);
or U13201 (N_13201,N_13116,N_13033);
nand U13202 (N_13202,N_13083,N_13022);
and U13203 (N_13203,N_13061,N_13073);
xnor U13204 (N_13204,N_13102,N_13105);
nor U13205 (N_13205,N_12995,N_13089);
and U13206 (N_13206,N_13030,N_12974);
or U13207 (N_13207,N_13061,N_13052);
xor U13208 (N_13208,N_13038,N_13058);
nor U13209 (N_13209,N_13089,N_12972);
or U13210 (N_13210,N_13097,N_12962);
nor U13211 (N_13211,N_13105,N_12982);
xor U13212 (N_13212,N_12981,N_13073);
xnor U13213 (N_13213,N_12993,N_13103);
nor U13214 (N_13214,N_12970,N_12999);
or U13215 (N_13215,N_13063,N_13069);
nor U13216 (N_13216,N_12993,N_13018);
xnor U13217 (N_13217,N_13110,N_13042);
xnor U13218 (N_13218,N_13076,N_13035);
or U13219 (N_13219,N_13051,N_13113);
nor U13220 (N_13220,N_13082,N_13050);
xnor U13221 (N_13221,N_13007,N_13004);
and U13222 (N_13222,N_13092,N_13078);
and U13223 (N_13223,N_13092,N_13008);
xnor U13224 (N_13224,N_13045,N_13009);
or U13225 (N_13225,N_13072,N_13003);
nand U13226 (N_13226,N_13081,N_12961);
and U13227 (N_13227,N_13017,N_13095);
and U13228 (N_13228,N_13086,N_13051);
nor U13229 (N_13229,N_12975,N_13066);
nand U13230 (N_13230,N_12997,N_12996);
or U13231 (N_13231,N_12968,N_13037);
nand U13232 (N_13232,N_13111,N_13070);
and U13233 (N_13233,N_13090,N_13092);
and U13234 (N_13234,N_13045,N_12995);
nand U13235 (N_13235,N_13048,N_12974);
nand U13236 (N_13236,N_13069,N_13108);
xnor U13237 (N_13237,N_13000,N_13080);
nand U13238 (N_13238,N_13071,N_13068);
nor U13239 (N_13239,N_13010,N_12967);
or U13240 (N_13240,N_13066,N_12994);
or U13241 (N_13241,N_13024,N_13083);
and U13242 (N_13242,N_12982,N_13042);
nor U13243 (N_13243,N_12986,N_13091);
nand U13244 (N_13244,N_12976,N_13114);
nor U13245 (N_13245,N_12980,N_12964);
nor U13246 (N_13246,N_12975,N_13007);
or U13247 (N_13247,N_12996,N_13072);
xor U13248 (N_13248,N_13003,N_13098);
and U13249 (N_13249,N_13118,N_13024);
nand U13250 (N_13250,N_12963,N_13010);
nand U13251 (N_13251,N_13101,N_13102);
nand U13252 (N_13252,N_13074,N_12996);
nand U13253 (N_13253,N_13105,N_13001);
and U13254 (N_13254,N_13002,N_13006);
or U13255 (N_13255,N_13035,N_12999);
and U13256 (N_13256,N_13105,N_13096);
or U13257 (N_13257,N_13044,N_12960);
or U13258 (N_13258,N_12960,N_13018);
and U13259 (N_13259,N_13044,N_12996);
xor U13260 (N_13260,N_13012,N_13113);
and U13261 (N_13261,N_12994,N_13009);
nand U13262 (N_13262,N_13071,N_12997);
nand U13263 (N_13263,N_13110,N_12977);
and U13264 (N_13264,N_13070,N_13112);
nand U13265 (N_13265,N_13096,N_13090);
nor U13266 (N_13266,N_13026,N_12980);
nor U13267 (N_13267,N_12980,N_12991);
xor U13268 (N_13268,N_12989,N_13078);
or U13269 (N_13269,N_13004,N_13038);
xor U13270 (N_13270,N_12992,N_13003);
nor U13271 (N_13271,N_13113,N_13052);
nor U13272 (N_13272,N_13090,N_13087);
nor U13273 (N_13273,N_13116,N_13107);
or U13274 (N_13274,N_13020,N_13111);
nor U13275 (N_13275,N_13036,N_13003);
nand U13276 (N_13276,N_13091,N_13010);
and U13277 (N_13277,N_12971,N_13030);
xor U13278 (N_13278,N_13059,N_13000);
and U13279 (N_13279,N_12962,N_13037);
and U13280 (N_13280,N_13215,N_13228);
nor U13281 (N_13281,N_13192,N_13128);
or U13282 (N_13282,N_13256,N_13237);
or U13283 (N_13283,N_13172,N_13243);
and U13284 (N_13284,N_13229,N_13168);
and U13285 (N_13285,N_13261,N_13241);
nand U13286 (N_13286,N_13236,N_13197);
nor U13287 (N_13287,N_13154,N_13270);
xnor U13288 (N_13288,N_13213,N_13247);
nor U13289 (N_13289,N_13159,N_13239);
nand U13290 (N_13290,N_13124,N_13169);
or U13291 (N_13291,N_13202,N_13186);
nand U13292 (N_13292,N_13240,N_13195);
or U13293 (N_13293,N_13269,N_13177);
nand U13294 (N_13294,N_13238,N_13178);
nor U13295 (N_13295,N_13259,N_13255);
nor U13296 (N_13296,N_13176,N_13250);
nor U13297 (N_13297,N_13164,N_13245);
nor U13298 (N_13298,N_13158,N_13127);
nor U13299 (N_13299,N_13218,N_13142);
and U13300 (N_13300,N_13140,N_13180);
xor U13301 (N_13301,N_13193,N_13149);
or U13302 (N_13302,N_13212,N_13184);
nand U13303 (N_13303,N_13258,N_13174);
and U13304 (N_13304,N_13225,N_13143);
nand U13305 (N_13305,N_13166,N_13147);
nor U13306 (N_13306,N_13226,N_13254);
nor U13307 (N_13307,N_13252,N_13221);
nand U13308 (N_13308,N_13201,N_13189);
nand U13309 (N_13309,N_13133,N_13220);
nand U13310 (N_13310,N_13151,N_13191);
and U13311 (N_13311,N_13146,N_13279);
or U13312 (N_13312,N_13262,N_13224);
nand U13313 (N_13313,N_13249,N_13181);
nand U13314 (N_13314,N_13182,N_13162);
and U13315 (N_13315,N_13260,N_13275);
xor U13316 (N_13316,N_13138,N_13185);
and U13317 (N_13317,N_13205,N_13131);
or U13318 (N_13318,N_13246,N_13200);
or U13319 (N_13319,N_13217,N_13208);
nand U13320 (N_13320,N_13242,N_13155);
nor U13321 (N_13321,N_13223,N_13126);
and U13322 (N_13322,N_13219,N_13165);
xnor U13323 (N_13323,N_13139,N_13244);
nand U13324 (N_13324,N_13125,N_13263);
nor U13325 (N_13325,N_13179,N_13264);
nor U13326 (N_13326,N_13257,N_13231);
nor U13327 (N_13327,N_13134,N_13227);
and U13328 (N_13328,N_13167,N_13235);
nand U13329 (N_13329,N_13253,N_13265);
and U13330 (N_13330,N_13230,N_13276);
and U13331 (N_13331,N_13190,N_13204);
nand U13332 (N_13332,N_13267,N_13123);
or U13333 (N_13333,N_13203,N_13187);
nor U13334 (N_13334,N_13175,N_13161);
nor U13335 (N_13335,N_13170,N_13183);
xnor U13336 (N_13336,N_13157,N_13129);
xor U13337 (N_13337,N_13122,N_13141);
xnor U13338 (N_13338,N_13199,N_13173);
nor U13339 (N_13339,N_13278,N_13188);
and U13340 (N_13340,N_13194,N_13266);
and U13341 (N_13341,N_13274,N_13136);
nand U13342 (N_13342,N_13132,N_13135);
nor U13343 (N_13343,N_13198,N_13216);
or U13344 (N_13344,N_13234,N_13120);
nand U13345 (N_13345,N_13233,N_13271);
and U13346 (N_13346,N_13145,N_13153);
or U13347 (N_13347,N_13121,N_13211);
nor U13348 (N_13348,N_13163,N_13251);
and U13349 (N_13349,N_13248,N_13207);
or U13350 (N_13350,N_13210,N_13277);
nor U13351 (N_13351,N_13273,N_13206);
or U13352 (N_13352,N_13130,N_13222);
nor U13353 (N_13353,N_13209,N_13156);
xnor U13354 (N_13354,N_13152,N_13214);
nor U13355 (N_13355,N_13268,N_13144);
and U13356 (N_13356,N_13196,N_13160);
xor U13357 (N_13357,N_13272,N_13232);
nand U13358 (N_13358,N_13171,N_13148);
or U13359 (N_13359,N_13137,N_13150);
nor U13360 (N_13360,N_13122,N_13209);
and U13361 (N_13361,N_13222,N_13124);
nor U13362 (N_13362,N_13239,N_13237);
nor U13363 (N_13363,N_13193,N_13150);
and U13364 (N_13364,N_13261,N_13191);
or U13365 (N_13365,N_13267,N_13149);
and U13366 (N_13366,N_13240,N_13276);
xor U13367 (N_13367,N_13126,N_13241);
and U13368 (N_13368,N_13190,N_13182);
nand U13369 (N_13369,N_13214,N_13167);
nor U13370 (N_13370,N_13148,N_13157);
or U13371 (N_13371,N_13278,N_13187);
nor U13372 (N_13372,N_13221,N_13135);
or U13373 (N_13373,N_13244,N_13196);
or U13374 (N_13374,N_13213,N_13195);
nor U13375 (N_13375,N_13176,N_13174);
nor U13376 (N_13376,N_13138,N_13158);
and U13377 (N_13377,N_13169,N_13123);
or U13378 (N_13378,N_13241,N_13164);
or U13379 (N_13379,N_13182,N_13205);
nor U13380 (N_13380,N_13253,N_13205);
xor U13381 (N_13381,N_13164,N_13236);
and U13382 (N_13382,N_13137,N_13218);
or U13383 (N_13383,N_13241,N_13173);
nor U13384 (N_13384,N_13263,N_13210);
nor U13385 (N_13385,N_13267,N_13206);
nor U13386 (N_13386,N_13165,N_13272);
nand U13387 (N_13387,N_13171,N_13248);
or U13388 (N_13388,N_13169,N_13178);
xor U13389 (N_13389,N_13278,N_13176);
or U13390 (N_13390,N_13275,N_13136);
nand U13391 (N_13391,N_13279,N_13245);
nand U13392 (N_13392,N_13278,N_13259);
and U13393 (N_13393,N_13158,N_13163);
nor U13394 (N_13394,N_13225,N_13279);
and U13395 (N_13395,N_13162,N_13191);
nor U13396 (N_13396,N_13213,N_13143);
nand U13397 (N_13397,N_13228,N_13218);
nand U13398 (N_13398,N_13180,N_13216);
nor U13399 (N_13399,N_13153,N_13277);
or U13400 (N_13400,N_13172,N_13191);
or U13401 (N_13401,N_13220,N_13249);
nor U13402 (N_13402,N_13234,N_13173);
or U13403 (N_13403,N_13278,N_13169);
and U13404 (N_13404,N_13243,N_13213);
xnor U13405 (N_13405,N_13257,N_13220);
nand U13406 (N_13406,N_13187,N_13211);
nor U13407 (N_13407,N_13245,N_13150);
and U13408 (N_13408,N_13239,N_13227);
and U13409 (N_13409,N_13232,N_13239);
and U13410 (N_13410,N_13267,N_13204);
and U13411 (N_13411,N_13271,N_13236);
xor U13412 (N_13412,N_13171,N_13258);
nor U13413 (N_13413,N_13126,N_13203);
nand U13414 (N_13414,N_13236,N_13152);
and U13415 (N_13415,N_13246,N_13172);
nand U13416 (N_13416,N_13196,N_13267);
nand U13417 (N_13417,N_13200,N_13127);
and U13418 (N_13418,N_13162,N_13158);
or U13419 (N_13419,N_13270,N_13175);
or U13420 (N_13420,N_13149,N_13206);
nor U13421 (N_13421,N_13137,N_13207);
nand U13422 (N_13422,N_13221,N_13169);
or U13423 (N_13423,N_13162,N_13173);
nand U13424 (N_13424,N_13159,N_13190);
and U13425 (N_13425,N_13139,N_13171);
and U13426 (N_13426,N_13136,N_13160);
or U13427 (N_13427,N_13179,N_13276);
nor U13428 (N_13428,N_13130,N_13247);
and U13429 (N_13429,N_13265,N_13150);
or U13430 (N_13430,N_13253,N_13273);
nand U13431 (N_13431,N_13141,N_13165);
nor U13432 (N_13432,N_13207,N_13177);
xor U13433 (N_13433,N_13200,N_13239);
nand U13434 (N_13434,N_13264,N_13210);
and U13435 (N_13435,N_13230,N_13234);
nor U13436 (N_13436,N_13234,N_13213);
and U13437 (N_13437,N_13182,N_13279);
or U13438 (N_13438,N_13207,N_13216);
nor U13439 (N_13439,N_13167,N_13259);
nor U13440 (N_13440,N_13416,N_13317);
nand U13441 (N_13441,N_13350,N_13364);
and U13442 (N_13442,N_13379,N_13315);
and U13443 (N_13443,N_13335,N_13285);
or U13444 (N_13444,N_13357,N_13420);
and U13445 (N_13445,N_13381,N_13319);
nor U13446 (N_13446,N_13328,N_13289);
and U13447 (N_13447,N_13287,N_13311);
or U13448 (N_13448,N_13434,N_13331);
and U13449 (N_13449,N_13325,N_13297);
xnor U13450 (N_13450,N_13329,N_13399);
and U13451 (N_13451,N_13436,N_13382);
or U13452 (N_13452,N_13341,N_13378);
xnor U13453 (N_13453,N_13375,N_13418);
and U13454 (N_13454,N_13344,N_13322);
or U13455 (N_13455,N_13389,N_13403);
or U13456 (N_13456,N_13430,N_13283);
or U13457 (N_13457,N_13307,N_13345);
and U13458 (N_13458,N_13310,N_13295);
nand U13459 (N_13459,N_13334,N_13305);
nor U13460 (N_13460,N_13414,N_13313);
or U13461 (N_13461,N_13431,N_13327);
nor U13462 (N_13462,N_13300,N_13404);
or U13463 (N_13463,N_13318,N_13304);
or U13464 (N_13464,N_13419,N_13354);
and U13465 (N_13465,N_13290,N_13383);
or U13466 (N_13466,N_13369,N_13401);
and U13467 (N_13467,N_13308,N_13337);
xnor U13468 (N_13468,N_13323,N_13347);
or U13469 (N_13469,N_13306,N_13284);
or U13470 (N_13470,N_13362,N_13405);
and U13471 (N_13471,N_13426,N_13400);
or U13472 (N_13472,N_13407,N_13370);
nand U13473 (N_13473,N_13393,N_13312);
nor U13474 (N_13474,N_13371,N_13439);
and U13475 (N_13475,N_13372,N_13348);
and U13476 (N_13476,N_13366,N_13338);
nand U13477 (N_13477,N_13423,N_13406);
or U13478 (N_13478,N_13298,N_13361);
nand U13479 (N_13479,N_13320,N_13346);
nand U13480 (N_13480,N_13373,N_13351);
and U13481 (N_13481,N_13294,N_13422);
nor U13482 (N_13482,N_13392,N_13415);
nor U13483 (N_13483,N_13425,N_13359);
and U13484 (N_13484,N_13360,N_13394);
nand U13485 (N_13485,N_13293,N_13377);
xnor U13486 (N_13486,N_13291,N_13428);
or U13487 (N_13487,N_13286,N_13367);
nand U13488 (N_13488,N_13299,N_13376);
and U13489 (N_13489,N_13356,N_13332);
or U13490 (N_13490,N_13316,N_13303);
nand U13491 (N_13491,N_13437,N_13363);
and U13492 (N_13492,N_13336,N_13358);
and U13493 (N_13493,N_13349,N_13339);
and U13494 (N_13494,N_13280,N_13408);
nor U13495 (N_13495,N_13413,N_13386);
nor U13496 (N_13496,N_13435,N_13296);
or U13497 (N_13497,N_13340,N_13421);
and U13498 (N_13498,N_13330,N_13391);
xor U13499 (N_13499,N_13302,N_13396);
xor U13500 (N_13500,N_13292,N_13380);
or U13501 (N_13501,N_13402,N_13433);
and U13502 (N_13502,N_13333,N_13282);
nor U13503 (N_13503,N_13390,N_13324);
and U13504 (N_13504,N_13321,N_13301);
and U13505 (N_13505,N_13412,N_13353);
xnor U13506 (N_13506,N_13398,N_13281);
and U13507 (N_13507,N_13429,N_13374);
nand U13508 (N_13508,N_13409,N_13410);
and U13509 (N_13509,N_13342,N_13309);
and U13510 (N_13510,N_13384,N_13352);
and U13511 (N_13511,N_13424,N_13438);
and U13512 (N_13512,N_13365,N_13355);
xnor U13513 (N_13513,N_13385,N_13288);
and U13514 (N_13514,N_13314,N_13368);
nand U13515 (N_13515,N_13427,N_13411);
nor U13516 (N_13516,N_13388,N_13395);
or U13517 (N_13517,N_13326,N_13387);
or U13518 (N_13518,N_13432,N_13397);
or U13519 (N_13519,N_13417,N_13343);
xnor U13520 (N_13520,N_13401,N_13388);
or U13521 (N_13521,N_13356,N_13369);
nor U13522 (N_13522,N_13393,N_13287);
xnor U13523 (N_13523,N_13387,N_13414);
and U13524 (N_13524,N_13331,N_13332);
xor U13525 (N_13525,N_13317,N_13398);
nand U13526 (N_13526,N_13353,N_13400);
nor U13527 (N_13527,N_13327,N_13282);
or U13528 (N_13528,N_13304,N_13395);
or U13529 (N_13529,N_13416,N_13373);
or U13530 (N_13530,N_13393,N_13345);
nand U13531 (N_13531,N_13413,N_13402);
or U13532 (N_13532,N_13426,N_13340);
and U13533 (N_13533,N_13354,N_13370);
and U13534 (N_13534,N_13411,N_13378);
or U13535 (N_13535,N_13401,N_13419);
or U13536 (N_13536,N_13348,N_13346);
nand U13537 (N_13537,N_13379,N_13292);
and U13538 (N_13538,N_13292,N_13400);
or U13539 (N_13539,N_13312,N_13339);
nor U13540 (N_13540,N_13385,N_13370);
nand U13541 (N_13541,N_13305,N_13369);
and U13542 (N_13542,N_13329,N_13376);
and U13543 (N_13543,N_13343,N_13436);
nor U13544 (N_13544,N_13282,N_13344);
or U13545 (N_13545,N_13313,N_13318);
nor U13546 (N_13546,N_13377,N_13362);
nand U13547 (N_13547,N_13385,N_13304);
xor U13548 (N_13548,N_13415,N_13327);
nor U13549 (N_13549,N_13329,N_13367);
nor U13550 (N_13550,N_13348,N_13362);
nand U13551 (N_13551,N_13316,N_13352);
or U13552 (N_13552,N_13425,N_13321);
nor U13553 (N_13553,N_13415,N_13293);
and U13554 (N_13554,N_13340,N_13373);
nand U13555 (N_13555,N_13329,N_13307);
or U13556 (N_13556,N_13391,N_13329);
nor U13557 (N_13557,N_13280,N_13331);
nand U13558 (N_13558,N_13307,N_13378);
and U13559 (N_13559,N_13402,N_13373);
and U13560 (N_13560,N_13386,N_13415);
or U13561 (N_13561,N_13290,N_13293);
xnor U13562 (N_13562,N_13374,N_13399);
or U13563 (N_13563,N_13378,N_13308);
nand U13564 (N_13564,N_13329,N_13434);
nor U13565 (N_13565,N_13360,N_13432);
and U13566 (N_13566,N_13417,N_13380);
nand U13567 (N_13567,N_13356,N_13297);
nand U13568 (N_13568,N_13426,N_13399);
or U13569 (N_13569,N_13417,N_13318);
and U13570 (N_13570,N_13287,N_13425);
or U13571 (N_13571,N_13384,N_13302);
or U13572 (N_13572,N_13377,N_13411);
xnor U13573 (N_13573,N_13404,N_13385);
or U13574 (N_13574,N_13348,N_13306);
xnor U13575 (N_13575,N_13309,N_13327);
nor U13576 (N_13576,N_13385,N_13335);
or U13577 (N_13577,N_13317,N_13337);
and U13578 (N_13578,N_13403,N_13343);
nand U13579 (N_13579,N_13299,N_13389);
nor U13580 (N_13580,N_13290,N_13346);
nand U13581 (N_13581,N_13381,N_13424);
xor U13582 (N_13582,N_13432,N_13344);
nor U13583 (N_13583,N_13410,N_13360);
and U13584 (N_13584,N_13323,N_13390);
and U13585 (N_13585,N_13307,N_13311);
xor U13586 (N_13586,N_13388,N_13429);
and U13587 (N_13587,N_13371,N_13343);
and U13588 (N_13588,N_13335,N_13419);
nor U13589 (N_13589,N_13410,N_13298);
or U13590 (N_13590,N_13307,N_13313);
and U13591 (N_13591,N_13337,N_13287);
and U13592 (N_13592,N_13407,N_13381);
nand U13593 (N_13593,N_13397,N_13433);
nand U13594 (N_13594,N_13292,N_13373);
or U13595 (N_13595,N_13397,N_13413);
nor U13596 (N_13596,N_13365,N_13423);
nand U13597 (N_13597,N_13289,N_13294);
and U13598 (N_13598,N_13377,N_13360);
nand U13599 (N_13599,N_13287,N_13363);
nand U13600 (N_13600,N_13445,N_13560);
nand U13601 (N_13601,N_13551,N_13498);
nand U13602 (N_13602,N_13567,N_13499);
and U13603 (N_13603,N_13591,N_13563);
or U13604 (N_13604,N_13585,N_13529);
nor U13605 (N_13605,N_13516,N_13497);
nor U13606 (N_13606,N_13474,N_13441);
nand U13607 (N_13607,N_13475,N_13577);
xor U13608 (N_13608,N_13599,N_13448);
nand U13609 (N_13609,N_13472,N_13575);
or U13610 (N_13610,N_13571,N_13576);
nor U13611 (N_13611,N_13520,N_13579);
and U13612 (N_13612,N_13538,N_13452);
nand U13613 (N_13613,N_13527,N_13542);
or U13614 (N_13614,N_13528,N_13589);
nor U13615 (N_13615,N_13590,N_13550);
nor U13616 (N_13616,N_13453,N_13487);
and U13617 (N_13617,N_13457,N_13491);
nor U13618 (N_13618,N_13496,N_13565);
nand U13619 (N_13619,N_13443,N_13588);
nor U13620 (N_13620,N_13476,N_13488);
xnor U13621 (N_13621,N_13500,N_13471);
nand U13622 (N_13622,N_13592,N_13581);
nand U13623 (N_13623,N_13568,N_13489);
and U13624 (N_13624,N_13522,N_13572);
nand U13625 (N_13625,N_13503,N_13477);
xor U13626 (N_13626,N_13587,N_13544);
nand U13627 (N_13627,N_13524,N_13597);
nor U13628 (N_13628,N_13548,N_13552);
or U13629 (N_13629,N_13549,N_13501);
nor U13630 (N_13630,N_13458,N_13468);
nand U13631 (N_13631,N_13546,N_13456);
nand U13632 (N_13632,N_13534,N_13557);
nor U13633 (N_13633,N_13515,N_13482);
nand U13634 (N_13634,N_13554,N_13469);
and U13635 (N_13635,N_13532,N_13533);
nand U13636 (N_13636,N_13519,N_13493);
nand U13637 (N_13637,N_13479,N_13555);
and U13638 (N_13638,N_13566,N_13574);
nor U13639 (N_13639,N_13570,N_13478);
or U13640 (N_13640,N_13483,N_13460);
nor U13641 (N_13641,N_13523,N_13543);
or U13642 (N_13642,N_13530,N_13440);
and U13643 (N_13643,N_13485,N_13473);
and U13644 (N_13644,N_13513,N_13514);
nand U13645 (N_13645,N_13598,N_13505);
xor U13646 (N_13646,N_13451,N_13517);
nand U13647 (N_13647,N_13518,N_13525);
nand U13648 (N_13648,N_13512,N_13596);
nor U13649 (N_13649,N_13464,N_13578);
and U13650 (N_13650,N_13508,N_13461);
or U13651 (N_13651,N_13442,N_13494);
nand U13652 (N_13652,N_13526,N_13446);
nand U13653 (N_13653,N_13536,N_13454);
nand U13654 (N_13654,N_13511,N_13480);
nand U13655 (N_13655,N_13559,N_13495);
nor U13656 (N_13656,N_13558,N_13492);
nor U13657 (N_13657,N_13466,N_13450);
nor U13658 (N_13658,N_13481,N_13547);
nor U13659 (N_13659,N_13502,N_13449);
or U13660 (N_13660,N_13583,N_13467);
nor U13661 (N_13661,N_13541,N_13510);
or U13662 (N_13662,N_13507,N_13564);
nand U13663 (N_13663,N_13539,N_13594);
nand U13664 (N_13664,N_13531,N_13582);
and U13665 (N_13665,N_13540,N_13486);
and U13666 (N_13666,N_13573,N_13506);
nor U13667 (N_13667,N_13521,N_13484);
nand U13668 (N_13668,N_13553,N_13586);
xor U13669 (N_13669,N_13462,N_13580);
nor U13670 (N_13670,N_13562,N_13490);
and U13671 (N_13671,N_13509,N_13535);
or U13672 (N_13672,N_13545,N_13463);
nor U13673 (N_13673,N_13459,N_13537);
or U13674 (N_13674,N_13561,N_13593);
and U13675 (N_13675,N_13584,N_13556);
nand U13676 (N_13676,N_13444,N_13504);
or U13677 (N_13677,N_13465,N_13447);
nand U13678 (N_13678,N_13595,N_13569);
or U13679 (N_13679,N_13455,N_13470);
and U13680 (N_13680,N_13545,N_13530);
and U13681 (N_13681,N_13539,N_13484);
nand U13682 (N_13682,N_13441,N_13468);
nand U13683 (N_13683,N_13581,N_13465);
nor U13684 (N_13684,N_13477,N_13521);
and U13685 (N_13685,N_13486,N_13592);
or U13686 (N_13686,N_13547,N_13575);
or U13687 (N_13687,N_13516,N_13444);
nor U13688 (N_13688,N_13590,N_13490);
nor U13689 (N_13689,N_13581,N_13554);
and U13690 (N_13690,N_13444,N_13483);
nor U13691 (N_13691,N_13583,N_13496);
nand U13692 (N_13692,N_13586,N_13455);
xor U13693 (N_13693,N_13535,N_13443);
nand U13694 (N_13694,N_13509,N_13521);
or U13695 (N_13695,N_13580,N_13553);
nand U13696 (N_13696,N_13571,N_13506);
and U13697 (N_13697,N_13552,N_13556);
nor U13698 (N_13698,N_13492,N_13442);
nor U13699 (N_13699,N_13502,N_13453);
and U13700 (N_13700,N_13496,N_13468);
nor U13701 (N_13701,N_13533,N_13494);
nand U13702 (N_13702,N_13471,N_13463);
nand U13703 (N_13703,N_13549,N_13589);
or U13704 (N_13704,N_13498,N_13442);
nor U13705 (N_13705,N_13468,N_13585);
nor U13706 (N_13706,N_13513,N_13536);
nand U13707 (N_13707,N_13465,N_13569);
nor U13708 (N_13708,N_13512,N_13457);
and U13709 (N_13709,N_13503,N_13578);
xor U13710 (N_13710,N_13463,N_13519);
nor U13711 (N_13711,N_13459,N_13567);
and U13712 (N_13712,N_13513,N_13477);
nor U13713 (N_13713,N_13514,N_13445);
nor U13714 (N_13714,N_13484,N_13532);
xnor U13715 (N_13715,N_13566,N_13482);
and U13716 (N_13716,N_13491,N_13470);
nand U13717 (N_13717,N_13502,N_13537);
nor U13718 (N_13718,N_13451,N_13560);
xor U13719 (N_13719,N_13495,N_13466);
nand U13720 (N_13720,N_13573,N_13557);
or U13721 (N_13721,N_13522,N_13529);
and U13722 (N_13722,N_13471,N_13576);
nor U13723 (N_13723,N_13470,N_13440);
or U13724 (N_13724,N_13588,N_13449);
and U13725 (N_13725,N_13529,N_13483);
and U13726 (N_13726,N_13505,N_13514);
nand U13727 (N_13727,N_13463,N_13561);
nor U13728 (N_13728,N_13509,N_13446);
nor U13729 (N_13729,N_13563,N_13443);
or U13730 (N_13730,N_13533,N_13553);
nor U13731 (N_13731,N_13502,N_13446);
or U13732 (N_13732,N_13584,N_13496);
and U13733 (N_13733,N_13476,N_13550);
and U13734 (N_13734,N_13585,N_13554);
and U13735 (N_13735,N_13456,N_13462);
nor U13736 (N_13736,N_13489,N_13554);
nand U13737 (N_13737,N_13556,N_13485);
nand U13738 (N_13738,N_13542,N_13548);
or U13739 (N_13739,N_13591,N_13530);
nand U13740 (N_13740,N_13534,N_13547);
nor U13741 (N_13741,N_13494,N_13479);
or U13742 (N_13742,N_13498,N_13495);
nor U13743 (N_13743,N_13451,N_13550);
nand U13744 (N_13744,N_13486,N_13454);
nand U13745 (N_13745,N_13536,N_13558);
and U13746 (N_13746,N_13553,N_13502);
and U13747 (N_13747,N_13595,N_13590);
or U13748 (N_13748,N_13551,N_13464);
or U13749 (N_13749,N_13526,N_13589);
nor U13750 (N_13750,N_13584,N_13512);
xnor U13751 (N_13751,N_13533,N_13564);
nand U13752 (N_13752,N_13445,N_13540);
or U13753 (N_13753,N_13588,N_13477);
nor U13754 (N_13754,N_13591,N_13449);
and U13755 (N_13755,N_13577,N_13517);
and U13756 (N_13756,N_13471,N_13457);
nor U13757 (N_13757,N_13584,N_13508);
nor U13758 (N_13758,N_13499,N_13446);
nor U13759 (N_13759,N_13588,N_13551);
or U13760 (N_13760,N_13663,N_13755);
nand U13761 (N_13761,N_13741,N_13724);
or U13762 (N_13762,N_13701,N_13679);
xor U13763 (N_13763,N_13604,N_13707);
nor U13764 (N_13764,N_13716,N_13734);
nor U13765 (N_13765,N_13635,N_13631);
or U13766 (N_13766,N_13620,N_13752);
or U13767 (N_13767,N_13633,N_13643);
xor U13768 (N_13768,N_13736,N_13756);
or U13769 (N_13769,N_13743,N_13615);
or U13770 (N_13770,N_13652,N_13758);
or U13771 (N_13771,N_13727,N_13626);
and U13772 (N_13772,N_13644,N_13618);
nand U13773 (N_13773,N_13738,N_13739);
nor U13774 (N_13774,N_13668,N_13737);
xnor U13775 (N_13775,N_13649,N_13702);
nor U13776 (N_13776,N_13711,N_13753);
and U13777 (N_13777,N_13748,N_13669);
and U13778 (N_13778,N_13732,N_13715);
nand U13779 (N_13779,N_13640,N_13697);
and U13780 (N_13780,N_13689,N_13609);
nand U13781 (N_13781,N_13693,N_13726);
and U13782 (N_13782,N_13645,N_13720);
and U13783 (N_13783,N_13657,N_13634);
nand U13784 (N_13784,N_13642,N_13641);
or U13785 (N_13785,N_13664,N_13613);
nor U13786 (N_13786,N_13606,N_13612);
xor U13787 (N_13787,N_13696,N_13754);
and U13788 (N_13788,N_13654,N_13623);
nor U13789 (N_13789,N_13718,N_13690);
or U13790 (N_13790,N_13617,N_13710);
and U13791 (N_13791,N_13608,N_13719);
or U13792 (N_13792,N_13600,N_13750);
or U13793 (N_13793,N_13673,N_13630);
or U13794 (N_13794,N_13667,N_13682);
nand U13795 (N_13795,N_13694,N_13735);
or U13796 (N_13796,N_13636,N_13611);
xor U13797 (N_13797,N_13699,N_13603);
nand U13798 (N_13798,N_13751,N_13629);
and U13799 (N_13799,N_13733,N_13681);
and U13800 (N_13800,N_13757,N_13647);
and U13801 (N_13801,N_13601,N_13685);
nor U13802 (N_13802,N_13674,N_13723);
nor U13803 (N_13803,N_13714,N_13703);
nor U13804 (N_13804,N_13605,N_13709);
or U13805 (N_13805,N_13680,N_13659);
and U13806 (N_13806,N_13725,N_13622);
nor U13807 (N_13807,N_13687,N_13672);
and U13808 (N_13808,N_13713,N_13650);
nor U13809 (N_13809,N_13717,N_13721);
nand U13810 (N_13810,N_13730,N_13651);
and U13811 (N_13811,N_13678,N_13648);
or U13812 (N_13812,N_13602,N_13653);
and U13813 (N_13813,N_13661,N_13621);
or U13814 (N_13814,N_13662,N_13671);
nand U13815 (N_13815,N_13684,N_13692);
or U13816 (N_13816,N_13700,N_13656);
nor U13817 (N_13817,N_13676,N_13759);
nor U13818 (N_13818,N_13638,N_13686);
or U13819 (N_13819,N_13675,N_13744);
nand U13820 (N_13820,N_13731,N_13670);
and U13821 (N_13821,N_13614,N_13708);
nand U13822 (N_13822,N_13722,N_13746);
nand U13823 (N_13823,N_13666,N_13660);
xnor U13824 (N_13824,N_13742,N_13616);
and U13825 (N_13825,N_13695,N_13698);
xnor U13826 (N_13826,N_13655,N_13691);
or U13827 (N_13827,N_13607,N_13658);
nand U13828 (N_13828,N_13665,N_13749);
xnor U13829 (N_13829,N_13627,N_13745);
nand U13830 (N_13830,N_13619,N_13632);
nand U13831 (N_13831,N_13712,N_13683);
nand U13832 (N_13832,N_13706,N_13704);
nand U13833 (N_13833,N_13610,N_13639);
nand U13834 (N_13834,N_13705,N_13646);
and U13835 (N_13835,N_13637,N_13729);
nand U13836 (N_13836,N_13677,N_13747);
or U13837 (N_13837,N_13740,N_13628);
or U13838 (N_13838,N_13688,N_13624);
nand U13839 (N_13839,N_13625,N_13728);
and U13840 (N_13840,N_13676,N_13670);
and U13841 (N_13841,N_13655,N_13726);
and U13842 (N_13842,N_13689,N_13757);
or U13843 (N_13843,N_13709,N_13711);
and U13844 (N_13844,N_13600,N_13718);
and U13845 (N_13845,N_13742,N_13657);
or U13846 (N_13846,N_13619,N_13626);
xor U13847 (N_13847,N_13677,N_13684);
nor U13848 (N_13848,N_13671,N_13742);
xor U13849 (N_13849,N_13670,N_13675);
nor U13850 (N_13850,N_13726,N_13674);
and U13851 (N_13851,N_13619,N_13731);
or U13852 (N_13852,N_13607,N_13677);
or U13853 (N_13853,N_13691,N_13621);
nor U13854 (N_13854,N_13745,N_13632);
and U13855 (N_13855,N_13609,N_13721);
nor U13856 (N_13856,N_13688,N_13745);
nor U13857 (N_13857,N_13691,N_13623);
or U13858 (N_13858,N_13604,N_13634);
nor U13859 (N_13859,N_13733,N_13690);
xnor U13860 (N_13860,N_13714,N_13731);
and U13861 (N_13861,N_13655,N_13732);
or U13862 (N_13862,N_13609,N_13620);
or U13863 (N_13863,N_13610,N_13635);
nand U13864 (N_13864,N_13629,N_13759);
nand U13865 (N_13865,N_13695,N_13758);
nor U13866 (N_13866,N_13603,N_13756);
and U13867 (N_13867,N_13648,N_13623);
and U13868 (N_13868,N_13734,N_13654);
or U13869 (N_13869,N_13725,N_13687);
and U13870 (N_13870,N_13640,N_13674);
or U13871 (N_13871,N_13631,N_13734);
and U13872 (N_13872,N_13710,N_13603);
nand U13873 (N_13873,N_13618,N_13759);
nor U13874 (N_13874,N_13748,N_13709);
or U13875 (N_13875,N_13732,N_13716);
nor U13876 (N_13876,N_13623,N_13645);
or U13877 (N_13877,N_13626,N_13644);
and U13878 (N_13878,N_13693,N_13736);
and U13879 (N_13879,N_13617,N_13752);
and U13880 (N_13880,N_13627,N_13755);
nand U13881 (N_13881,N_13690,N_13723);
nor U13882 (N_13882,N_13602,N_13711);
nor U13883 (N_13883,N_13702,N_13712);
and U13884 (N_13884,N_13669,N_13758);
xor U13885 (N_13885,N_13646,N_13718);
nand U13886 (N_13886,N_13701,N_13704);
and U13887 (N_13887,N_13707,N_13709);
nor U13888 (N_13888,N_13750,N_13646);
nand U13889 (N_13889,N_13752,N_13608);
nor U13890 (N_13890,N_13730,N_13628);
nor U13891 (N_13891,N_13644,N_13603);
nor U13892 (N_13892,N_13730,N_13746);
nor U13893 (N_13893,N_13628,N_13661);
nor U13894 (N_13894,N_13602,N_13656);
and U13895 (N_13895,N_13621,N_13711);
and U13896 (N_13896,N_13677,N_13638);
nand U13897 (N_13897,N_13735,N_13713);
nor U13898 (N_13898,N_13605,N_13680);
nor U13899 (N_13899,N_13616,N_13612);
or U13900 (N_13900,N_13609,N_13752);
and U13901 (N_13901,N_13733,N_13703);
nor U13902 (N_13902,N_13668,N_13616);
or U13903 (N_13903,N_13676,N_13623);
nand U13904 (N_13904,N_13737,N_13603);
nand U13905 (N_13905,N_13601,N_13675);
or U13906 (N_13906,N_13673,N_13750);
and U13907 (N_13907,N_13746,N_13628);
nor U13908 (N_13908,N_13702,N_13601);
nor U13909 (N_13909,N_13624,N_13751);
nand U13910 (N_13910,N_13748,N_13696);
and U13911 (N_13911,N_13746,N_13656);
and U13912 (N_13912,N_13690,N_13652);
nand U13913 (N_13913,N_13733,N_13686);
and U13914 (N_13914,N_13713,N_13678);
and U13915 (N_13915,N_13709,N_13621);
or U13916 (N_13916,N_13694,N_13610);
nor U13917 (N_13917,N_13656,N_13607);
nand U13918 (N_13918,N_13664,N_13723);
nor U13919 (N_13919,N_13699,N_13731);
or U13920 (N_13920,N_13810,N_13782);
nand U13921 (N_13921,N_13898,N_13902);
and U13922 (N_13922,N_13788,N_13907);
nand U13923 (N_13923,N_13796,N_13904);
nor U13924 (N_13924,N_13883,N_13849);
and U13925 (N_13925,N_13803,N_13834);
and U13926 (N_13926,N_13801,N_13760);
and U13927 (N_13927,N_13843,N_13808);
xnor U13928 (N_13928,N_13888,N_13900);
nor U13929 (N_13929,N_13766,N_13890);
and U13930 (N_13930,N_13761,N_13807);
and U13931 (N_13931,N_13762,N_13845);
nor U13932 (N_13932,N_13910,N_13781);
nand U13933 (N_13933,N_13826,N_13859);
and U13934 (N_13934,N_13866,N_13800);
and U13935 (N_13935,N_13897,N_13881);
nand U13936 (N_13936,N_13794,N_13893);
nand U13937 (N_13937,N_13817,N_13916);
nand U13938 (N_13938,N_13822,N_13863);
nor U13939 (N_13939,N_13769,N_13790);
or U13940 (N_13940,N_13870,N_13797);
nor U13941 (N_13941,N_13798,N_13799);
and U13942 (N_13942,N_13789,N_13909);
nand U13943 (N_13943,N_13835,N_13889);
nand U13944 (N_13944,N_13885,N_13786);
and U13945 (N_13945,N_13855,N_13873);
nand U13946 (N_13946,N_13857,N_13765);
and U13947 (N_13947,N_13830,N_13896);
or U13948 (N_13948,N_13846,N_13811);
and U13949 (N_13949,N_13886,N_13805);
nor U13950 (N_13950,N_13787,N_13812);
or U13951 (N_13951,N_13836,N_13824);
nor U13952 (N_13952,N_13869,N_13793);
or U13953 (N_13953,N_13819,N_13813);
and U13954 (N_13954,N_13784,N_13841);
nor U13955 (N_13955,N_13816,N_13785);
or U13956 (N_13956,N_13844,N_13908);
or U13957 (N_13957,N_13776,N_13878);
xnor U13958 (N_13958,N_13771,N_13795);
nand U13959 (N_13959,N_13792,N_13850);
and U13960 (N_13960,N_13828,N_13767);
nor U13961 (N_13961,N_13778,N_13818);
nand U13962 (N_13962,N_13854,N_13763);
or U13963 (N_13963,N_13880,N_13864);
or U13964 (N_13964,N_13825,N_13851);
nor U13965 (N_13965,N_13842,N_13783);
or U13966 (N_13966,N_13839,N_13877);
nand U13967 (N_13967,N_13852,N_13874);
and U13968 (N_13968,N_13901,N_13871);
or U13969 (N_13969,N_13780,N_13906);
nand U13970 (N_13970,N_13882,N_13768);
or U13971 (N_13971,N_13861,N_13838);
nor U13972 (N_13972,N_13875,N_13829);
or U13973 (N_13973,N_13831,N_13837);
and U13974 (N_13974,N_13876,N_13821);
or U13975 (N_13975,N_13804,N_13892);
nand U13976 (N_13976,N_13802,N_13853);
and U13977 (N_13977,N_13894,N_13775);
and U13978 (N_13978,N_13779,N_13791);
or U13979 (N_13979,N_13858,N_13777);
or U13980 (N_13980,N_13879,N_13905);
nor U13981 (N_13981,N_13823,N_13764);
nand U13982 (N_13982,N_13914,N_13911);
nor U13983 (N_13983,N_13860,N_13809);
xor U13984 (N_13984,N_13915,N_13865);
nand U13985 (N_13985,N_13919,N_13827);
and U13986 (N_13986,N_13806,N_13847);
or U13987 (N_13987,N_13867,N_13918);
xnor U13988 (N_13988,N_13772,N_13884);
or U13989 (N_13989,N_13895,N_13773);
and U13990 (N_13990,N_13872,N_13833);
nand U13991 (N_13991,N_13868,N_13903);
nand U13992 (N_13992,N_13887,N_13848);
nand U13993 (N_13993,N_13856,N_13862);
nand U13994 (N_13994,N_13774,N_13912);
nor U13995 (N_13995,N_13840,N_13820);
nand U13996 (N_13996,N_13814,N_13832);
nor U13997 (N_13997,N_13913,N_13815);
and U13998 (N_13998,N_13891,N_13917);
or U13999 (N_13999,N_13899,N_13770);
nand U14000 (N_14000,N_13914,N_13867);
nor U14001 (N_14001,N_13771,N_13830);
or U14002 (N_14002,N_13818,N_13835);
or U14003 (N_14003,N_13768,N_13870);
or U14004 (N_14004,N_13917,N_13821);
or U14005 (N_14005,N_13786,N_13803);
xor U14006 (N_14006,N_13813,N_13918);
nor U14007 (N_14007,N_13762,N_13833);
nand U14008 (N_14008,N_13847,N_13834);
and U14009 (N_14009,N_13784,N_13782);
nand U14010 (N_14010,N_13886,N_13817);
or U14011 (N_14011,N_13819,N_13816);
and U14012 (N_14012,N_13912,N_13895);
nand U14013 (N_14013,N_13857,N_13864);
nor U14014 (N_14014,N_13887,N_13850);
nor U14015 (N_14015,N_13910,N_13908);
xor U14016 (N_14016,N_13878,N_13840);
nor U14017 (N_14017,N_13882,N_13790);
or U14018 (N_14018,N_13780,N_13831);
xnor U14019 (N_14019,N_13915,N_13918);
or U14020 (N_14020,N_13862,N_13822);
and U14021 (N_14021,N_13816,N_13830);
or U14022 (N_14022,N_13845,N_13829);
or U14023 (N_14023,N_13912,N_13785);
xnor U14024 (N_14024,N_13867,N_13848);
and U14025 (N_14025,N_13905,N_13861);
nor U14026 (N_14026,N_13778,N_13904);
xor U14027 (N_14027,N_13905,N_13779);
or U14028 (N_14028,N_13857,N_13858);
xnor U14029 (N_14029,N_13864,N_13888);
nand U14030 (N_14030,N_13886,N_13769);
or U14031 (N_14031,N_13862,N_13888);
and U14032 (N_14032,N_13890,N_13843);
xor U14033 (N_14033,N_13844,N_13879);
nand U14034 (N_14034,N_13801,N_13904);
xor U14035 (N_14035,N_13771,N_13760);
and U14036 (N_14036,N_13837,N_13760);
and U14037 (N_14037,N_13824,N_13852);
or U14038 (N_14038,N_13775,N_13872);
nand U14039 (N_14039,N_13914,N_13912);
nand U14040 (N_14040,N_13808,N_13773);
and U14041 (N_14041,N_13761,N_13901);
and U14042 (N_14042,N_13895,N_13785);
nor U14043 (N_14043,N_13891,N_13805);
and U14044 (N_14044,N_13784,N_13761);
or U14045 (N_14045,N_13892,N_13816);
or U14046 (N_14046,N_13895,N_13822);
nor U14047 (N_14047,N_13790,N_13868);
nand U14048 (N_14048,N_13775,N_13844);
nor U14049 (N_14049,N_13917,N_13852);
nand U14050 (N_14050,N_13795,N_13885);
xor U14051 (N_14051,N_13781,N_13821);
nand U14052 (N_14052,N_13827,N_13810);
or U14053 (N_14053,N_13818,N_13794);
and U14054 (N_14054,N_13829,N_13814);
nor U14055 (N_14055,N_13909,N_13881);
nor U14056 (N_14056,N_13817,N_13783);
and U14057 (N_14057,N_13858,N_13852);
and U14058 (N_14058,N_13872,N_13802);
and U14059 (N_14059,N_13806,N_13892);
nand U14060 (N_14060,N_13864,N_13829);
and U14061 (N_14061,N_13824,N_13909);
nor U14062 (N_14062,N_13791,N_13864);
nand U14063 (N_14063,N_13869,N_13832);
or U14064 (N_14064,N_13834,N_13767);
nand U14065 (N_14065,N_13775,N_13831);
nand U14066 (N_14066,N_13805,N_13839);
xor U14067 (N_14067,N_13782,N_13809);
and U14068 (N_14068,N_13909,N_13790);
nor U14069 (N_14069,N_13882,N_13831);
nor U14070 (N_14070,N_13883,N_13890);
and U14071 (N_14071,N_13864,N_13870);
or U14072 (N_14072,N_13803,N_13767);
xnor U14073 (N_14073,N_13854,N_13881);
nand U14074 (N_14074,N_13867,N_13849);
xor U14075 (N_14075,N_13824,N_13913);
xor U14076 (N_14076,N_13786,N_13782);
nor U14077 (N_14077,N_13889,N_13912);
nor U14078 (N_14078,N_13794,N_13790);
nor U14079 (N_14079,N_13788,N_13882);
nor U14080 (N_14080,N_14015,N_13987);
nand U14081 (N_14081,N_14065,N_13945);
nor U14082 (N_14082,N_14055,N_14064);
and U14083 (N_14083,N_14025,N_13946);
nand U14084 (N_14084,N_13973,N_14007);
nor U14085 (N_14085,N_14073,N_13934);
or U14086 (N_14086,N_14059,N_14012);
and U14087 (N_14087,N_13927,N_14057);
or U14088 (N_14088,N_14056,N_14001);
and U14089 (N_14089,N_14027,N_14078);
or U14090 (N_14090,N_13920,N_13979);
nand U14091 (N_14091,N_14032,N_13921);
or U14092 (N_14092,N_14010,N_14069);
and U14093 (N_14093,N_14058,N_14009);
nand U14094 (N_14094,N_13931,N_13955);
or U14095 (N_14095,N_14017,N_13977);
nor U14096 (N_14096,N_13962,N_13952);
xnor U14097 (N_14097,N_14049,N_13970);
xnor U14098 (N_14098,N_13999,N_14014);
nand U14099 (N_14099,N_13997,N_14076);
xor U14100 (N_14100,N_13942,N_13922);
xnor U14101 (N_14101,N_14040,N_14011);
nor U14102 (N_14102,N_14039,N_14074);
and U14103 (N_14103,N_13939,N_14060);
or U14104 (N_14104,N_13943,N_14061);
and U14105 (N_14105,N_13930,N_14041);
nor U14106 (N_14106,N_14072,N_14063);
or U14107 (N_14107,N_13954,N_13948);
xnor U14108 (N_14108,N_13972,N_14045);
nor U14109 (N_14109,N_13996,N_14034);
nand U14110 (N_14110,N_13981,N_14043);
nand U14111 (N_14111,N_14024,N_14044);
nor U14112 (N_14112,N_13992,N_14022);
and U14113 (N_14113,N_13960,N_13933);
xnor U14114 (N_14114,N_13951,N_13963);
nand U14115 (N_14115,N_14030,N_13988);
or U14116 (N_14116,N_14038,N_13941);
nand U14117 (N_14117,N_14062,N_13984);
nor U14118 (N_14118,N_13953,N_14036);
nor U14119 (N_14119,N_14079,N_14071);
xnor U14120 (N_14120,N_13998,N_13976);
xor U14121 (N_14121,N_14006,N_14028);
xor U14122 (N_14122,N_14037,N_13949);
nand U14123 (N_14123,N_14000,N_14046);
or U14124 (N_14124,N_14067,N_14051);
or U14125 (N_14125,N_13932,N_14016);
or U14126 (N_14126,N_13989,N_13985);
or U14127 (N_14127,N_13971,N_14068);
or U14128 (N_14128,N_13947,N_13964);
or U14129 (N_14129,N_14066,N_14029);
xnor U14130 (N_14130,N_13958,N_14023);
nand U14131 (N_14131,N_14070,N_13966);
nand U14132 (N_14132,N_13990,N_13978);
nor U14133 (N_14133,N_13991,N_13994);
and U14134 (N_14134,N_13928,N_13968);
nor U14135 (N_14135,N_13969,N_13929);
nand U14136 (N_14136,N_14033,N_13944);
or U14137 (N_14137,N_14053,N_14021);
nor U14138 (N_14138,N_13923,N_13957);
nor U14139 (N_14139,N_14002,N_14047);
nor U14140 (N_14140,N_14008,N_14075);
or U14141 (N_14141,N_13956,N_14005);
and U14142 (N_14142,N_13924,N_13995);
nor U14143 (N_14143,N_13961,N_13936);
or U14144 (N_14144,N_13975,N_13993);
nand U14145 (N_14145,N_13983,N_14018);
nor U14146 (N_14146,N_14020,N_13980);
nor U14147 (N_14147,N_14048,N_14077);
nand U14148 (N_14148,N_13938,N_13935);
nor U14149 (N_14149,N_14050,N_13982);
and U14150 (N_14150,N_14035,N_13965);
and U14151 (N_14151,N_13940,N_14013);
xnor U14152 (N_14152,N_13959,N_14052);
and U14153 (N_14153,N_13974,N_13937);
and U14154 (N_14154,N_13926,N_14004);
and U14155 (N_14155,N_14019,N_13986);
nor U14156 (N_14156,N_13950,N_14003);
nor U14157 (N_14157,N_13967,N_13925);
nand U14158 (N_14158,N_14026,N_14031);
or U14159 (N_14159,N_14054,N_14042);
nand U14160 (N_14160,N_13942,N_13997);
and U14161 (N_14161,N_13929,N_13981);
nor U14162 (N_14162,N_14000,N_13972);
nand U14163 (N_14163,N_13937,N_13934);
xor U14164 (N_14164,N_13998,N_14032);
nor U14165 (N_14165,N_14054,N_13970);
or U14166 (N_14166,N_13970,N_14020);
nor U14167 (N_14167,N_13953,N_14071);
nand U14168 (N_14168,N_14042,N_14055);
and U14169 (N_14169,N_13948,N_13991);
or U14170 (N_14170,N_14020,N_14027);
nand U14171 (N_14171,N_14055,N_14019);
or U14172 (N_14172,N_14071,N_13933);
nand U14173 (N_14173,N_13954,N_13955);
nor U14174 (N_14174,N_14065,N_14079);
nand U14175 (N_14175,N_13941,N_14058);
and U14176 (N_14176,N_13934,N_14014);
xnor U14177 (N_14177,N_14058,N_14044);
nor U14178 (N_14178,N_14037,N_14043);
nand U14179 (N_14179,N_14015,N_13951);
nor U14180 (N_14180,N_13950,N_14067);
nand U14181 (N_14181,N_13926,N_14003);
nand U14182 (N_14182,N_13938,N_13991);
xnor U14183 (N_14183,N_14054,N_14018);
xor U14184 (N_14184,N_14004,N_13978);
or U14185 (N_14185,N_13920,N_14019);
nor U14186 (N_14186,N_13944,N_13983);
and U14187 (N_14187,N_13970,N_13960);
or U14188 (N_14188,N_14027,N_13983);
nor U14189 (N_14189,N_14043,N_14040);
nor U14190 (N_14190,N_14011,N_13947);
nand U14191 (N_14191,N_13937,N_13975);
nor U14192 (N_14192,N_14073,N_13931);
nor U14193 (N_14193,N_13942,N_14052);
or U14194 (N_14194,N_14070,N_13993);
or U14195 (N_14195,N_14065,N_14050);
nand U14196 (N_14196,N_14073,N_14006);
nor U14197 (N_14197,N_14057,N_14055);
nand U14198 (N_14198,N_13942,N_14068);
nand U14199 (N_14199,N_13925,N_13956);
or U14200 (N_14200,N_14025,N_13936);
and U14201 (N_14201,N_14022,N_13960);
nor U14202 (N_14202,N_14045,N_13944);
and U14203 (N_14203,N_14066,N_14045);
xor U14204 (N_14204,N_14014,N_13970);
or U14205 (N_14205,N_14029,N_14006);
and U14206 (N_14206,N_13923,N_13971);
nand U14207 (N_14207,N_14070,N_14074);
nand U14208 (N_14208,N_13942,N_14069);
and U14209 (N_14209,N_14056,N_13948);
and U14210 (N_14210,N_13983,N_13938);
nand U14211 (N_14211,N_14068,N_14025);
nor U14212 (N_14212,N_14030,N_14058);
nand U14213 (N_14213,N_13946,N_13942);
nor U14214 (N_14214,N_13996,N_14008);
or U14215 (N_14215,N_14042,N_13982);
nand U14216 (N_14216,N_14006,N_14017);
or U14217 (N_14217,N_14009,N_13975);
and U14218 (N_14218,N_14018,N_13973);
nand U14219 (N_14219,N_13973,N_13958);
or U14220 (N_14220,N_13948,N_14079);
or U14221 (N_14221,N_14061,N_13981);
or U14222 (N_14222,N_13960,N_14015);
or U14223 (N_14223,N_13956,N_13950);
nor U14224 (N_14224,N_14033,N_14067);
xor U14225 (N_14225,N_13950,N_14062);
nand U14226 (N_14226,N_13976,N_13935);
nor U14227 (N_14227,N_14013,N_14051);
and U14228 (N_14228,N_14020,N_13990);
or U14229 (N_14229,N_13981,N_14025);
and U14230 (N_14230,N_13927,N_13987);
xor U14231 (N_14231,N_14037,N_13989);
nor U14232 (N_14232,N_13959,N_14025);
or U14233 (N_14233,N_14028,N_14019);
nand U14234 (N_14234,N_13940,N_14000);
and U14235 (N_14235,N_13969,N_13927);
or U14236 (N_14236,N_13929,N_14006);
and U14237 (N_14237,N_13995,N_14064);
nor U14238 (N_14238,N_14063,N_13946);
xor U14239 (N_14239,N_14043,N_14058);
or U14240 (N_14240,N_14141,N_14221);
and U14241 (N_14241,N_14101,N_14229);
or U14242 (N_14242,N_14124,N_14119);
nand U14243 (N_14243,N_14239,N_14127);
xnor U14244 (N_14244,N_14179,N_14205);
nor U14245 (N_14245,N_14184,N_14129);
or U14246 (N_14246,N_14202,N_14181);
xor U14247 (N_14247,N_14210,N_14152);
or U14248 (N_14248,N_14168,N_14180);
nor U14249 (N_14249,N_14234,N_14106);
nand U14250 (N_14250,N_14102,N_14148);
and U14251 (N_14251,N_14143,N_14169);
or U14252 (N_14252,N_14084,N_14140);
and U14253 (N_14253,N_14235,N_14081);
and U14254 (N_14254,N_14236,N_14134);
nand U14255 (N_14255,N_14216,N_14147);
or U14256 (N_14256,N_14135,N_14155);
or U14257 (N_14257,N_14122,N_14186);
nand U14258 (N_14258,N_14201,N_14218);
nor U14259 (N_14259,N_14104,N_14196);
or U14260 (N_14260,N_14220,N_14142);
nand U14261 (N_14261,N_14080,N_14174);
or U14262 (N_14262,N_14172,N_14118);
nand U14263 (N_14263,N_14232,N_14161);
and U14264 (N_14264,N_14099,N_14092);
and U14265 (N_14265,N_14123,N_14146);
or U14266 (N_14266,N_14108,N_14165);
xor U14267 (N_14267,N_14219,N_14194);
nor U14268 (N_14268,N_14206,N_14215);
and U14269 (N_14269,N_14237,N_14111);
nand U14270 (N_14270,N_14187,N_14208);
or U14271 (N_14271,N_14126,N_14082);
xnor U14272 (N_14272,N_14109,N_14233);
or U14273 (N_14273,N_14191,N_14149);
and U14274 (N_14274,N_14125,N_14110);
nor U14275 (N_14275,N_14224,N_14089);
nor U14276 (N_14276,N_14093,N_14188);
nand U14277 (N_14277,N_14153,N_14200);
and U14278 (N_14278,N_14217,N_14226);
nor U14279 (N_14279,N_14199,N_14204);
xor U14280 (N_14280,N_14213,N_14107);
nor U14281 (N_14281,N_14171,N_14158);
and U14282 (N_14282,N_14098,N_14103);
or U14283 (N_14283,N_14223,N_14182);
nand U14284 (N_14284,N_14214,N_14130);
and U14285 (N_14285,N_14160,N_14162);
or U14286 (N_14286,N_14231,N_14116);
nand U14287 (N_14287,N_14090,N_14085);
nor U14288 (N_14288,N_14238,N_14139);
and U14289 (N_14289,N_14121,N_14193);
nand U14290 (N_14290,N_14156,N_14225);
nand U14291 (N_14291,N_14207,N_14173);
or U14292 (N_14292,N_14227,N_14151);
and U14293 (N_14293,N_14209,N_14211);
nand U14294 (N_14294,N_14203,N_14176);
or U14295 (N_14295,N_14100,N_14131);
and U14296 (N_14296,N_14138,N_14097);
xnor U14297 (N_14297,N_14178,N_14167);
nor U14298 (N_14298,N_14185,N_14163);
xnor U14299 (N_14299,N_14195,N_14112);
or U14300 (N_14300,N_14136,N_14132);
nand U14301 (N_14301,N_14159,N_14094);
nor U14302 (N_14302,N_14230,N_14177);
xnor U14303 (N_14303,N_14095,N_14166);
or U14304 (N_14304,N_14087,N_14189);
or U14305 (N_14305,N_14192,N_14133);
nand U14306 (N_14306,N_14114,N_14088);
and U14307 (N_14307,N_14120,N_14170);
nor U14308 (N_14308,N_14175,N_14150);
or U14309 (N_14309,N_14117,N_14190);
and U14310 (N_14310,N_14105,N_14086);
nor U14311 (N_14311,N_14083,N_14183);
xor U14312 (N_14312,N_14113,N_14137);
nand U14313 (N_14313,N_14145,N_14197);
and U14314 (N_14314,N_14154,N_14096);
nand U14315 (N_14315,N_14228,N_14164);
nand U14316 (N_14316,N_14222,N_14115);
nand U14317 (N_14317,N_14128,N_14212);
nand U14318 (N_14318,N_14091,N_14198);
or U14319 (N_14319,N_14144,N_14157);
nor U14320 (N_14320,N_14118,N_14134);
xor U14321 (N_14321,N_14148,N_14092);
xnor U14322 (N_14322,N_14130,N_14236);
or U14323 (N_14323,N_14185,N_14090);
and U14324 (N_14324,N_14162,N_14106);
or U14325 (N_14325,N_14082,N_14238);
or U14326 (N_14326,N_14096,N_14176);
nor U14327 (N_14327,N_14094,N_14183);
or U14328 (N_14328,N_14235,N_14139);
nor U14329 (N_14329,N_14131,N_14188);
and U14330 (N_14330,N_14180,N_14205);
or U14331 (N_14331,N_14207,N_14216);
nand U14332 (N_14332,N_14081,N_14119);
xnor U14333 (N_14333,N_14083,N_14150);
nand U14334 (N_14334,N_14164,N_14110);
nand U14335 (N_14335,N_14111,N_14104);
and U14336 (N_14336,N_14084,N_14081);
nor U14337 (N_14337,N_14186,N_14108);
nand U14338 (N_14338,N_14092,N_14086);
or U14339 (N_14339,N_14229,N_14087);
nor U14340 (N_14340,N_14230,N_14091);
or U14341 (N_14341,N_14096,N_14237);
and U14342 (N_14342,N_14143,N_14171);
nand U14343 (N_14343,N_14105,N_14236);
and U14344 (N_14344,N_14148,N_14097);
nor U14345 (N_14345,N_14114,N_14221);
nor U14346 (N_14346,N_14174,N_14082);
and U14347 (N_14347,N_14106,N_14123);
nor U14348 (N_14348,N_14145,N_14128);
nand U14349 (N_14349,N_14215,N_14130);
nand U14350 (N_14350,N_14159,N_14228);
nor U14351 (N_14351,N_14130,N_14126);
xor U14352 (N_14352,N_14115,N_14201);
nor U14353 (N_14353,N_14226,N_14150);
xnor U14354 (N_14354,N_14227,N_14206);
and U14355 (N_14355,N_14233,N_14144);
xnor U14356 (N_14356,N_14125,N_14119);
nor U14357 (N_14357,N_14172,N_14083);
nand U14358 (N_14358,N_14227,N_14237);
or U14359 (N_14359,N_14232,N_14117);
nor U14360 (N_14360,N_14210,N_14101);
xnor U14361 (N_14361,N_14151,N_14139);
xor U14362 (N_14362,N_14166,N_14235);
nand U14363 (N_14363,N_14105,N_14121);
nor U14364 (N_14364,N_14165,N_14115);
and U14365 (N_14365,N_14224,N_14132);
or U14366 (N_14366,N_14102,N_14181);
nor U14367 (N_14367,N_14146,N_14230);
nand U14368 (N_14368,N_14173,N_14171);
xor U14369 (N_14369,N_14186,N_14091);
nor U14370 (N_14370,N_14126,N_14169);
and U14371 (N_14371,N_14207,N_14215);
or U14372 (N_14372,N_14233,N_14234);
nor U14373 (N_14373,N_14208,N_14205);
and U14374 (N_14374,N_14115,N_14168);
or U14375 (N_14375,N_14217,N_14237);
nand U14376 (N_14376,N_14218,N_14207);
xor U14377 (N_14377,N_14196,N_14218);
nand U14378 (N_14378,N_14151,N_14145);
and U14379 (N_14379,N_14209,N_14080);
and U14380 (N_14380,N_14120,N_14111);
xor U14381 (N_14381,N_14225,N_14145);
xnor U14382 (N_14382,N_14166,N_14218);
and U14383 (N_14383,N_14223,N_14129);
xnor U14384 (N_14384,N_14131,N_14138);
nor U14385 (N_14385,N_14239,N_14165);
and U14386 (N_14386,N_14124,N_14212);
or U14387 (N_14387,N_14148,N_14108);
nand U14388 (N_14388,N_14200,N_14157);
nor U14389 (N_14389,N_14179,N_14144);
nor U14390 (N_14390,N_14146,N_14191);
nor U14391 (N_14391,N_14210,N_14206);
nor U14392 (N_14392,N_14088,N_14174);
and U14393 (N_14393,N_14205,N_14100);
nand U14394 (N_14394,N_14127,N_14169);
or U14395 (N_14395,N_14093,N_14109);
and U14396 (N_14396,N_14145,N_14120);
nor U14397 (N_14397,N_14191,N_14090);
and U14398 (N_14398,N_14183,N_14200);
nand U14399 (N_14399,N_14177,N_14142);
and U14400 (N_14400,N_14340,N_14302);
or U14401 (N_14401,N_14353,N_14263);
nand U14402 (N_14402,N_14283,N_14316);
or U14403 (N_14403,N_14355,N_14265);
and U14404 (N_14404,N_14275,N_14284);
nor U14405 (N_14405,N_14245,N_14240);
and U14406 (N_14406,N_14242,N_14325);
or U14407 (N_14407,N_14329,N_14369);
nand U14408 (N_14408,N_14333,N_14346);
nor U14409 (N_14409,N_14248,N_14247);
nand U14410 (N_14410,N_14380,N_14388);
or U14411 (N_14411,N_14313,N_14330);
or U14412 (N_14412,N_14326,N_14290);
xor U14413 (N_14413,N_14393,N_14269);
xor U14414 (N_14414,N_14251,N_14331);
xor U14415 (N_14415,N_14304,N_14366);
xor U14416 (N_14416,N_14334,N_14339);
nor U14417 (N_14417,N_14305,N_14252);
and U14418 (N_14418,N_14282,N_14322);
and U14419 (N_14419,N_14266,N_14387);
and U14420 (N_14420,N_14382,N_14389);
nor U14421 (N_14421,N_14364,N_14376);
or U14422 (N_14422,N_14273,N_14286);
nor U14423 (N_14423,N_14289,N_14394);
xnor U14424 (N_14424,N_14362,N_14395);
xnor U14425 (N_14425,N_14292,N_14390);
and U14426 (N_14426,N_14320,N_14259);
or U14427 (N_14427,N_14391,N_14371);
nand U14428 (N_14428,N_14349,N_14250);
nor U14429 (N_14429,N_14351,N_14295);
and U14430 (N_14430,N_14354,N_14293);
nand U14431 (N_14431,N_14379,N_14314);
nor U14432 (N_14432,N_14297,N_14370);
and U14433 (N_14433,N_14398,N_14299);
nand U14434 (N_14434,N_14285,N_14246);
or U14435 (N_14435,N_14257,N_14274);
and U14436 (N_14436,N_14298,N_14287);
and U14437 (N_14437,N_14310,N_14308);
or U14438 (N_14438,N_14291,N_14323);
or U14439 (N_14439,N_14350,N_14241);
and U14440 (N_14440,N_14397,N_14359);
nand U14441 (N_14441,N_14312,N_14279);
nor U14442 (N_14442,N_14328,N_14317);
nor U14443 (N_14443,N_14352,N_14319);
or U14444 (N_14444,N_14262,N_14309);
and U14445 (N_14445,N_14300,N_14321);
and U14446 (N_14446,N_14344,N_14336);
xor U14447 (N_14447,N_14356,N_14303);
and U14448 (N_14448,N_14341,N_14253);
nand U14449 (N_14449,N_14375,N_14374);
nand U14450 (N_14450,N_14377,N_14244);
nor U14451 (N_14451,N_14381,N_14347);
nand U14452 (N_14452,N_14307,N_14365);
or U14453 (N_14453,N_14243,N_14343);
or U14454 (N_14454,N_14392,N_14361);
and U14455 (N_14455,N_14260,N_14383);
and U14456 (N_14456,N_14386,N_14288);
nor U14457 (N_14457,N_14271,N_14335);
nand U14458 (N_14458,N_14296,N_14278);
xnor U14459 (N_14459,N_14268,N_14384);
or U14460 (N_14460,N_14327,N_14280);
nor U14461 (N_14461,N_14255,N_14272);
and U14462 (N_14462,N_14311,N_14264);
or U14463 (N_14463,N_14276,N_14254);
or U14464 (N_14464,N_14363,N_14368);
xor U14465 (N_14465,N_14358,N_14270);
nand U14466 (N_14466,N_14396,N_14261);
nor U14467 (N_14467,N_14385,N_14306);
or U14468 (N_14468,N_14357,N_14348);
nand U14469 (N_14469,N_14378,N_14342);
nand U14470 (N_14470,N_14256,N_14372);
nand U14471 (N_14471,N_14318,N_14258);
or U14472 (N_14472,N_14324,N_14332);
or U14473 (N_14473,N_14367,N_14277);
xnor U14474 (N_14474,N_14281,N_14360);
or U14475 (N_14475,N_14301,N_14345);
and U14476 (N_14476,N_14294,N_14399);
nor U14477 (N_14477,N_14338,N_14373);
nor U14478 (N_14478,N_14337,N_14267);
nor U14479 (N_14479,N_14315,N_14249);
nand U14480 (N_14480,N_14245,N_14387);
or U14481 (N_14481,N_14396,N_14269);
nand U14482 (N_14482,N_14386,N_14268);
nor U14483 (N_14483,N_14351,N_14358);
nand U14484 (N_14484,N_14327,N_14290);
nand U14485 (N_14485,N_14310,N_14299);
and U14486 (N_14486,N_14314,N_14375);
and U14487 (N_14487,N_14312,N_14355);
and U14488 (N_14488,N_14351,N_14292);
and U14489 (N_14489,N_14322,N_14305);
nor U14490 (N_14490,N_14332,N_14330);
nand U14491 (N_14491,N_14279,N_14314);
or U14492 (N_14492,N_14310,N_14279);
and U14493 (N_14493,N_14305,N_14254);
or U14494 (N_14494,N_14261,N_14259);
nand U14495 (N_14495,N_14252,N_14287);
nand U14496 (N_14496,N_14386,N_14279);
nand U14497 (N_14497,N_14363,N_14322);
or U14498 (N_14498,N_14249,N_14285);
and U14499 (N_14499,N_14304,N_14375);
nand U14500 (N_14500,N_14253,N_14287);
nor U14501 (N_14501,N_14347,N_14387);
or U14502 (N_14502,N_14332,N_14365);
nand U14503 (N_14503,N_14264,N_14297);
nor U14504 (N_14504,N_14282,N_14350);
and U14505 (N_14505,N_14332,N_14373);
nor U14506 (N_14506,N_14306,N_14305);
nand U14507 (N_14507,N_14289,N_14264);
nor U14508 (N_14508,N_14334,N_14319);
nor U14509 (N_14509,N_14328,N_14292);
nor U14510 (N_14510,N_14281,N_14358);
xor U14511 (N_14511,N_14389,N_14250);
nand U14512 (N_14512,N_14396,N_14322);
nor U14513 (N_14513,N_14271,N_14388);
nor U14514 (N_14514,N_14383,N_14386);
and U14515 (N_14515,N_14248,N_14299);
and U14516 (N_14516,N_14246,N_14304);
or U14517 (N_14517,N_14395,N_14262);
xor U14518 (N_14518,N_14385,N_14338);
nand U14519 (N_14519,N_14275,N_14334);
or U14520 (N_14520,N_14341,N_14398);
and U14521 (N_14521,N_14326,N_14349);
or U14522 (N_14522,N_14324,N_14277);
nor U14523 (N_14523,N_14252,N_14318);
xor U14524 (N_14524,N_14319,N_14372);
or U14525 (N_14525,N_14344,N_14368);
nand U14526 (N_14526,N_14241,N_14322);
nor U14527 (N_14527,N_14277,N_14378);
nor U14528 (N_14528,N_14353,N_14288);
nand U14529 (N_14529,N_14301,N_14294);
nor U14530 (N_14530,N_14280,N_14291);
nor U14531 (N_14531,N_14365,N_14302);
or U14532 (N_14532,N_14331,N_14396);
and U14533 (N_14533,N_14246,N_14320);
or U14534 (N_14534,N_14379,N_14293);
and U14535 (N_14535,N_14361,N_14272);
or U14536 (N_14536,N_14260,N_14300);
nand U14537 (N_14537,N_14318,N_14267);
and U14538 (N_14538,N_14247,N_14386);
or U14539 (N_14539,N_14259,N_14389);
nor U14540 (N_14540,N_14270,N_14394);
nor U14541 (N_14541,N_14306,N_14245);
nand U14542 (N_14542,N_14357,N_14302);
nand U14543 (N_14543,N_14255,N_14317);
nand U14544 (N_14544,N_14285,N_14340);
nand U14545 (N_14545,N_14254,N_14290);
or U14546 (N_14546,N_14375,N_14387);
or U14547 (N_14547,N_14292,N_14362);
or U14548 (N_14548,N_14304,N_14333);
nor U14549 (N_14549,N_14362,N_14342);
nor U14550 (N_14550,N_14387,N_14390);
nor U14551 (N_14551,N_14327,N_14325);
and U14552 (N_14552,N_14380,N_14305);
or U14553 (N_14553,N_14348,N_14326);
or U14554 (N_14554,N_14369,N_14379);
nand U14555 (N_14555,N_14249,N_14331);
nand U14556 (N_14556,N_14291,N_14264);
or U14557 (N_14557,N_14269,N_14288);
nor U14558 (N_14558,N_14334,N_14361);
or U14559 (N_14559,N_14366,N_14384);
nand U14560 (N_14560,N_14554,N_14499);
or U14561 (N_14561,N_14416,N_14501);
nand U14562 (N_14562,N_14502,N_14506);
nand U14563 (N_14563,N_14507,N_14513);
nor U14564 (N_14564,N_14504,N_14412);
nand U14565 (N_14565,N_14445,N_14505);
nor U14566 (N_14566,N_14411,N_14444);
nor U14567 (N_14567,N_14531,N_14438);
and U14568 (N_14568,N_14521,N_14529);
and U14569 (N_14569,N_14403,N_14417);
or U14570 (N_14570,N_14485,N_14460);
nor U14571 (N_14571,N_14545,N_14463);
or U14572 (N_14572,N_14518,N_14449);
nand U14573 (N_14573,N_14436,N_14489);
nor U14574 (N_14574,N_14400,N_14469);
nand U14575 (N_14575,N_14483,N_14523);
or U14576 (N_14576,N_14555,N_14420);
nor U14577 (N_14577,N_14527,N_14495);
nor U14578 (N_14578,N_14433,N_14440);
nor U14579 (N_14579,N_14404,N_14522);
xor U14580 (N_14580,N_14421,N_14496);
and U14581 (N_14581,N_14426,N_14544);
and U14582 (N_14582,N_14480,N_14556);
xor U14583 (N_14583,N_14516,N_14481);
nor U14584 (N_14584,N_14487,N_14455);
or U14585 (N_14585,N_14541,N_14540);
or U14586 (N_14586,N_14430,N_14539);
or U14587 (N_14587,N_14464,N_14549);
and U14588 (N_14588,N_14410,N_14405);
nor U14589 (N_14589,N_14450,N_14446);
and U14590 (N_14590,N_14431,N_14402);
or U14591 (N_14591,N_14401,N_14466);
or U14592 (N_14592,N_14482,N_14478);
or U14593 (N_14593,N_14439,N_14550);
and U14594 (N_14594,N_14418,N_14476);
nor U14595 (N_14595,N_14508,N_14465);
nand U14596 (N_14596,N_14517,N_14414);
nand U14597 (N_14597,N_14461,N_14519);
xnor U14598 (N_14598,N_14468,N_14427);
nand U14599 (N_14599,N_14472,N_14543);
nor U14600 (N_14600,N_14479,N_14553);
nor U14601 (N_14601,N_14434,N_14406);
nand U14602 (N_14602,N_14520,N_14490);
nor U14603 (N_14603,N_14526,N_14515);
or U14604 (N_14604,N_14477,N_14530);
and U14605 (N_14605,N_14524,N_14511);
or U14606 (N_14606,N_14413,N_14408);
or U14607 (N_14607,N_14494,N_14533);
or U14608 (N_14608,N_14457,N_14443);
and U14609 (N_14609,N_14467,N_14558);
xnor U14610 (N_14610,N_14422,N_14497);
nor U14611 (N_14611,N_14459,N_14452);
nand U14612 (N_14612,N_14491,N_14498);
and U14613 (N_14613,N_14528,N_14538);
and U14614 (N_14614,N_14419,N_14536);
and U14615 (N_14615,N_14429,N_14500);
and U14616 (N_14616,N_14470,N_14547);
nor U14617 (N_14617,N_14514,N_14510);
and U14618 (N_14618,N_14447,N_14407);
and U14619 (N_14619,N_14432,N_14509);
xor U14620 (N_14620,N_14473,N_14548);
nand U14621 (N_14621,N_14441,N_14409);
nand U14622 (N_14622,N_14546,N_14486);
nor U14623 (N_14623,N_14458,N_14503);
and U14624 (N_14624,N_14471,N_14424);
nand U14625 (N_14625,N_14425,N_14512);
and U14626 (N_14626,N_14552,N_14428);
nand U14627 (N_14627,N_14456,N_14535);
xor U14628 (N_14628,N_14448,N_14453);
or U14629 (N_14629,N_14475,N_14525);
nand U14630 (N_14630,N_14423,N_14451);
and U14631 (N_14631,N_14454,N_14474);
nor U14632 (N_14632,N_14484,N_14493);
nor U14633 (N_14633,N_14551,N_14415);
nor U14634 (N_14634,N_14442,N_14492);
xor U14635 (N_14635,N_14559,N_14488);
or U14636 (N_14636,N_14534,N_14537);
nor U14637 (N_14637,N_14542,N_14532);
or U14638 (N_14638,N_14437,N_14557);
or U14639 (N_14639,N_14462,N_14435);
nor U14640 (N_14640,N_14455,N_14518);
nand U14641 (N_14641,N_14555,N_14531);
or U14642 (N_14642,N_14405,N_14558);
or U14643 (N_14643,N_14559,N_14404);
xnor U14644 (N_14644,N_14526,N_14450);
xnor U14645 (N_14645,N_14406,N_14512);
and U14646 (N_14646,N_14434,N_14450);
xor U14647 (N_14647,N_14415,N_14475);
and U14648 (N_14648,N_14473,N_14402);
nand U14649 (N_14649,N_14495,N_14506);
nor U14650 (N_14650,N_14504,N_14502);
nor U14651 (N_14651,N_14400,N_14405);
and U14652 (N_14652,N_14460,N_14414);
nand U14653 (N_14653,N_14490,N_14402);
and U14654 (N_14654,N_14541,N_14401);
nand U14655 (N_14655,N_14421,N_14409);
nand U14656 (N_14656,N_14536,N_14469);
or U14657 (N_14657,N_14462,N_14415);
nand U14658 (N_14658,N_14550,N_14415);
or U14659 (N_14659,N_14557,N_14524);
nor U14660 (N_14660,N_14466,N_14554);
nor U14661 (N_14661,N_14433,N_14551);
nor U14662 (N_14662,N_14532,N_14509);
xnor U14663 (N_14663,N_14412,N_14523);
nand U14664 (N_14664,N_14491,N_14553);
or U14665 (N_14665,N_14503,N_14455);
nor U14666 (N_14666,N_14476,N_14519);
xnor U14667 (N_14667,N_14450,N_14487);
and U14668 (N_14668,N_14486,N_14502);
or U14669 (N_14669,N_14479,N_14545);
or U14670 (N_14670,N_14476,N_14410);
or U14671 (N_14671,N_14558,N_14432);
or U14672 (N_14672,N_14432,N_14460);
nand U14673 (N_14673,N_14518,N_14429);
or U14674 (N_14674,N_14489,N_14407);
nand U14675 (N_14675,N_14448,N_14462);
and U14676 (N_14676,N_14518,N_14413);
xor U14677 (N_14677,N_14540,N_14529);
nor U14678 (N_14678,N_14431,N_14553);
nand U14679 (N_14679,N_14472,N_14445);
nor U14680 (N_14680,N_14521,N_14513);
and U14681 (N_14681,N_14535,N_14481);
or U14682 (N_14682,N_14483,N_14464);
and U14683 (N_14683,N_14454,N_14410);
and U14684 (N_14684,N_14412,N_14428);
and U14685 (N_14685,N_14528,N_14500);
and U14686 (N_14686,N_14442,N_14458);
nand U14687 (N_14687,N_14427,N_14444);
or U14688 (N_14688,N_14443,N_14551);
xnor U14689 (N_14689,N_14475,N_14481);
nand U14690 (N_14690,N_14415,N_14524);
or U14691 (N_14691,N_14412,N_14558);
nor U14692 (N_14692,N_14427,N_14516);
or U14693 (N_14693,N_14528,N_14513);
or U14694 (N_14694,N_14501,N_14481);
nand U14695 (N_14695,N_14473,N_14472);
or U14696 (N_14696,N_14442,N_14410);
xnor U14697 (N_14697,N_14488,N_14426);
or U14698 (N_14698,N_14432,N_14446);
or U14699 (N_14699,N_14471,N_14548);
and U14700 (N_14700,N_14535,N_14530);
nor U14701 (N_14701,N_14513,N_14482);
nand U14702 (N_14702,N_14490,N_14545);
and U14703 (N_14703,N_14497,N_14528);
and U14704 (N_14704,N_14527,N_14550);
nand U14705 (N_14705,N_14507,N_14555);
nor U14706 (N_14706,N_14433,N_14540);
and U14707 (N_14707,N_14447,N_14517);
or U14708 (N_14708,N_14536,N_14538);
or U14709 (N_14709,N_14522,N_14426);
and U14710 (N_14710,N_14553,N_14441);
and U14711 (N_14711,N_14495,N_14550);
nand U14712 (N_14712,N_14548,N_14441);
and U14713 (N_14713,N_14548,N_14434);
and U14714 (N_14714,N_14499,N_14453);
nor U14715 (N_14715,N_14521,N_14402);
nor U14716 (N_14716,N_14457,N_14498);
nand U14717 (N_14717,N_14550,N_14429);
nor U14718 (N_14718,N_14419,N_14417);
or U14719 (N_14719,N_14469,N_14487);
and U14720 (N_14720,N_14584,N_14586);
or U14721 (N_14721,N_14615,N_14689);
or U14722 (N_14722,N_14626,N_14648);
or U14723 (N_14723,N_14631,N_14657);
xor U14724 (N_14724,N_14653,N_14684);
and U14725 (N_14725,N_14578,N_14610);
nand U14726 (N_14726,N_14617,N_14681);
nand U14727 (N_14727,N_14569,N_14683);
nand U14728 (N_14728,N_14704,N_14718);
or U14729 (N_14729,N_14716,N_14589);
xnor U14730 (N_14730,N_14658,N_14613);
nor U14731 (N_14731,N_14674,N_14564);
nand U14732 (N_14732,N_14655,N_14579);
and U14733 (N_14733,N_14625,N_14652);
and U14734 (N_14734,N_14662,N_14701);
or U14735 (N_14735,N_14565,N_14686);
or U14736 (N_14736,N_14560,N_14709);
or U14737 (N_14737,N_14566,N_14611);
or U14738 (N_14738,N_14712,N_14666);
xnor U14739 (N_14739,N_14628,N_14574);
nor U14740 (N_14740,N_14719,N_14677);
nor U14741 (N_14741,N_14580,N_14619);
nand U14742 (N_14742,N_14680,N_14606);
nor U14743 (N_14743,N_14607,N_14563);
or U14744 (N_14744,N_14585,N_14668);
xnor U14745 (N_14745,N_14632,N_14711);
or U14746 (N_14746,N_14561,N_14685);
and U14747 (N_14747,N_14616,N_14576);
nand U14748 (N_14748,N_14661,N_14637);
or U14749 (N_14749,N_14670,N_14660);
or U14750 (N_14750,N_14663,N_14699);
nor U14751 (N_14751,N_14595,N_14717);
nand U14752 (N_14752,N_14697,N_14624);
nor U14753 (N_14753,N_14633,N_14641);
nand U14754 (N_14754,N_14588,N_14667);
or U14755 (N_14755,N_14639,N_14593);
and U14756 (N_14756,N_14654,N_14571);
nor U14757 (N_14757,N_14702,N_14651);
or U14758 (N_14758,N_14592,N_14630);
xnor U14759 (N_14759,N_14706,N_14669);
nor U14760 (N_14760,N_14694,N_14696);
nand U14761 (N_14761,N_14691,N_14679);
or U14762 (N_14762,N_14597,N_14567);
nand U14763 (N_14763,N_14603,N_14713);
and U14764 (N_14764,N_14605,N_14682);
nand U14765 (N_14765,N_14714,N_14659);
nor U14766 (N_14766,N_14700,N_14664);
nand U14767 (N_14767,N_14703,N_14708);
or U14768 (N_14768,N_14687,N_14656);
or U14769 (N_14769,N_14635,N_14614);
nand U14770 (N_14770,N_14582,N_14693);
and U14771 (N_14771,N_14705,N_14665);
and U14772 (N_14772,N_14638,N_14644);
and U14773 (N_14773,N_14591,N_14570);
or U14774 (N_14774,N_14572,N_14604);
or U14775 (N_14775,N_14715,N_14643);
or U14776 (N_14776,N_14690,N_14678);
or U14777 (N_14777,N_14609,N_14562);
nand U14778 (N_14778,N_14627,N_14636);
or U14779 (N_14779,N_14675,N_14710);
nand U14780 (N_14780,N_14623,N_14618);
nand U14781 (N_14781,N_14642,N_14649);
nor U14782 (N_14782,N_14612,N_14583);
nor U14783 (N_14783,N_14575,N_14692);
nand U14784 (N_14784,N_14672,N_14647);
nor U14785 (N_14785,N_14601,N_14707);
nand U14786 (N_14786,N_14621,N_14568);
nand U14787 (N_14787,N_14673,N_14698);
or U14788 (N_14788,N_14596,N_14646);
and U14789 (N_14789,N_14594,N_14600);
and U14790 (N_14790,N_14650,N_14671);
xnor U14791 (N_14791,N_14622,N_14676);
nor U14792 (N_14792,N_14620,N_14645);
nand U14793 (N_14793,N_14587,N_14598);
and U14794 (N_14794,N_14695,N_14577);
and U14795 (N_14795,N_14634,N_14640);
and U14796 (N_14796,N_14602,N_14573);
nand U14797 (N_14797,N_14629,N_14581);
and U14798 (N_14798,N_14608,N_14590);
and U14799 (N_14799,N_14599,N_14688);
and U14800 (N_14800,N_14592,N_14572);
nor U14801 (N_14801,N_14674,N_14709);
nand U14802 (N_14802,N_14701,N_14596);
or U14803 (N_14803,N_14667,N_14578);
and U14804 (N_14804,N_14672,N_14708);
and U14805 (N_14805,N_14662,N_14698);
and U14806 (N_14806,N_14705,N_14560);
nand U14807 (N_14807,N_14640,N_14671);
xnor U14808 (N_14808,N_14647,N_14597);
nand U14809 (N_14809,N_14654,N_14710);
or U14810 (N_14810,N_14566,N_14692);
and U14811 (N_14811,N_14589,N_14689);
nand U14812 (N_14812,N_14606,N_14587);
xor U14813 (N_14813,N_14633,N_14699);
nand U14814 (N_14814,N_14574,N_14673);
nor U14815 (N_14815,N_14584,N_14670);
and U14816 (N_14816,N_14573,N_14620);
xnor U14817 (N_14817,N_14658,N_14607);
nand U14818 (N_14818,N_14592,N_14616);
or U14819 (N_14819,N_14679,N_14639);
or U14820 (N_14820,N_14710,N_14639);
xor U14821 (N_14821,N_14571,N_14701);
nand U14822 (N_14822,N_14630,N_14638);
nor U14823 (N_14823,N_14680,N_14589);
nor U14824 (N_14824,N_14594,N_14630);
nor U14825 (N_14825,N_14591,N_14608);
nand U14826 (N_14826,N_14638,N_14565);
or U14827 (N_14827,N_14574,N_14701);
or U14828 (N_14828,N_14695,N_14652);
nor U14829 (N_14829,N_14589,N_14666);
nand U14830 (N_14830,N_14638,N_14625);
nand U14831 (N_14831,N_14609,N_14597);
nor U14832 (N_14832,N_14619,N_14633);
nor U14833 (N_14833,N_14697,N_14682);
and U14834 (N_14834,N_14648,N_14588);
nand U14835 (N_14835,N_14562,N_14587);
or U14836 (N_14836,N_14617,N_14679);
nor U14837 (N_14837,N_14629,N_14614);
or U14838 (N_14838,N_14601,N_14704);
or U14839 (N_14839,N_14680,N_14563);
or U14840 (N_14840,N_14643,N_14659);
and U14841 (N_14841,N_14639,N_14568);
and U14842 (N_14842,N_14685,N_14674);
or U14843 (N_14843,N_14618,N_14694);
nor U14844 (N_14844,N_14615,N_14599);
nand U14845 (N_14845,N_14603,N_14718);
and U14846 (N_14846,N_14626,N_14665);
and U14847 (N_14847,N_14578,N_14634);
and U14848 (N_14848,N_14591,N_14710);
nor U14849 (N_14849,N_14688,N_14665);
and U14850 (N_14850,N_14699,N_14585);
nor U14851 (N_14851,N_14569,N_14714);
or U14852 (N_14852,N_14602,N_14670);
and U14853 (N_14853,N_14637,N_14593);
and U14854 (N_14854,N_14583,N_14592);
nor U14855 (N_14855,N_14719,N_14663);
nor U14856 (N_14856,N_14666,N_14607);
xnor U14857 (N_14857,N_14628,N_14678);
or U14858 (N_14858,N_14616,N_14618);
and U14859 (N_14859,N_14582,N_14666);
nor U14860 (N_14860,N_14639,N_14718);
or U14861 (N_14861,N_14611,N_14638);
nand U14862 (N_14862,N_14616,N_14627);
or U14863 (N_14863,N_14662,N_14637);
nand U14864 (N_14864,N_14676,N_14710);
or U14865 (N_14865,N_14673,N_14596);
and U14866 (N_14866,N_14636,N_14660);
or U14867 (N_14867,N_14638,N_14663);
nand U14868 (N_14868,N_14629,N_14583);
nor U14869 (N_14869,N_14705,N_14717);
and U14870 (N_14870,N_14689,N_14639);
nand U14871 (N_14871,N_14561,N_14642);
nand U14872 (N_14872,N_14675,N_14575);
or U14873 (N_14873,N_14607,N_14620);
and U14874 (N_14874,N_14623,N_14611);
xnor U14875 (N_14875,N_14590,N_14631);
xnor U14876 (N_14876,N_14600,N_14696);
nor U14877 (N_14877,N_14589,N_14650);
nand U14878 (N_14878,N_14704,N_14638);
and U14879 (N_14879,N_14669,N_14674);
or U14880 (N_14880,N_14848,N_14768);
nor U14881 (N_14881,N_14875,N_14832);
nand U14882 (N_14882,N_14861,N_14845);
xnor U14883 (N_14883,N_14759,N_14846);
or U14884 (N_14884,N_14830,N_14826);
and U14885 (N_14885,N_14720,N_14751);
nor U14886 (N_14886,N_14860,N_14753);
nand U14887 (N_14887,N_14785,N_14781);
and U14888 (N_14888,N_14735,N_14827);
and U14889 (N_14889,N_14786,N_14758);
or U14890 (N_14890,N_14764,N_14800);
nand U14891 (N_14891,N_14793,N_14856);
nand U14892 (N_14892,N_14765,N_14774);
nor U14893 (N_14893,N_14797,N_14796);
xnor U14894 (N_14894,N_14798,N_14844);
or U14895 (N_14895,N_14835,N_14825);
and U14896 (N_14896,N_14857,N_14839);
or U14897 (N_14897,N_14740,N_14782);
or U14898 (N_14898,N_14849,N_14779);
nor U14899 (N_14899,N_14778,N_14867);
nand U14900 (N_14900,N_14772,N_14806);
or U14901 (N_14901,N_14794,N_14819);
nor U14902 (N_14902,N_14811,N_14842);
or U14903 (N_14903,N_14721,N_14731);
nand U14904 (N_14904,N_14757,N_14807);
and U14905 (N_14905,N_14855,N_14726);
and U14906 (N_14906,N_14725,N_14852);
or U14907 (N_14907,N_14854,N_14780);
or U14908 (N_14908,N_14822,N_14730);
nand U14909 (N_14909,N_14791,N_14850);
or U14910 (N_14910,N_14727,N_14804);
nand U14911 (N_14911,N_14790,N_14802);
or U14912 (N_14912,N_14733,N_14808);
nand U14913 (N_14913,N_14870,N_14868);
nor U14914 (N_14914,N_14879,N_14776);
or U14915 (N_14915,N_14801,N_14738);
xor U14916 (N_14916,N_14744,N_14723);
nand U14917 (N_14917,N_14770,N_14828);
or U14918 (N_14918,N_14817,N_14872);
nor U14919 (N_14919,N_14836,N_14766);
nor U14920 (N_14920,N_14853,N_14820);
nor U14921 (N_14921,N_14787,N_14821);
and U14922 (N_14922,N_14877,N_14812);
or U14923 (N_14923,N_14810,N_14871);
or U14924 (N_14924,N_14763,N_14754);
nor U14925 (N_14925,N_14829,N_14750);
nand U14926 (N_14926,N_14737,N_14874);
nand U14927 (N_14927,N_14784,N_14783);
and U14928 (N_14928,N_14818,N_14729);
or U14929 (N_14929,N_14809,N_14876);
nand U14930 (N_14930,N_14805,N_14851);
nand U14931 (N_14931,N_14732,N_14789);
nor U14932 (N_14932,N_14878,N_14777);
or U14933 (N_14933,N_14724,N_14815);
nor U14934 (N_14934,N_14756,N_14739);
nand U14935 (N_14935,N_14761,N_14859);
nor U14936 (N_14936,N_14773,N_14746);
nor U14937 (N_14937,N_14858,N_14803);
xnor U14938 (N_14938,N_14741,N_14834);
nand U14939 (N_14939,N_14749,N_14748);
nand U14940 (N_14940,N_14873,N_14823);
and U14941 (N_14941,N_14838,N_14767);
and U14942 (N_14942,N_14866,N_14745);
or U14943 (N_14943,N_14865,N_14752);
or U14944 (N_14944,N_14769,N_14722);
nand U14945 (N_14945,N_14742,N_14862);
nand U14946 (N_14946,N_14771,N_14792);
nand U14947 (N_14947,N_14788,N_14837);
and U14948 (N_14948,N_14831,N_14824);
or U14949 (N_14949,N_14841,N_14816);
and U14950 (N_14950,N_14734,N_14755);
nor U14951 (N_14951,N_14869,N_14863);
nor U14952 (N_14952,N_14762,N_14743);
nor U14953 (N_14953,N_14736,N_14728);
or U14954 (N_14954,N_14833,N_14814);
or U14955 (N_14955,N_14775,N_14799);
nor U14956 (N_14956,N_14760,N_14864);
xor U14957 (N_14957,N_14813,N_14795);
or U14958 (N_14958,N_14840,N_14747);
nand U14959 (N_14959,N_14847,N_14843);
nor U14960 (N_14960,N_14792,N_14738);
nand U14961 (N_14961,N_14770,N_14810);
and U14962 (N_14962,N_14749,N_14762);
or U14963 (N_14963,N_14737,N_14763);
xor U14964 (N_14964,N_14842,N_14780);
or U14965 (N_14965,N_14833,N_14732);
and U14966 (N_14966,N_14758,N_14863);
nand U14967 (N_14967,N_14804,N_14803);
and U14968 (N_14968,N_14856,N_14732);
or U14969 (N_14969,N_14760,N_14823);
and U14970 (N_14970,N_14732,N_14849);
xnor U14971 (N_14971,N_14865,N_14847);
and U14972 (N_14972,N_14763,N_14820);
and U14973 (N_14973,N_14846,N_14812);
nand U14974 (N_14974,N_14736,N_14836);
xor U14975 (N_14975,N_14846,N_14765);
nand U14976 (N_14976,N_14720,N_14738);
nor U14977 (N_14977,N_14783,N_14829);
nand U14978 (N_14978,N_14829,N_14839);
and U14979 (N_14979,N_14843,N_14776);
or U14980 (N_14980,N_14853,N_14877);
and U14981 (N_14981,N_14835,N_14828);
nor U14982 (N_14982,N_14803,N_14761);
nand U14983 (N_14983,N_14868,N_14730);
or U14984 (N_14984,N_14743,N_14752);
and U14985 (N_14985,N_14844,N_14809);
and U14986 (N_14986,N_14834,N_14813);
and U14987 (N_14987,N_14728,N_14853);
or U14988 (N_14988,N_14768,N_14761);
and U14989 (N_14989,N_14757,N_14734);
nor U14990 (N_14990,N_14760,N_14773);
or U14991 (N_14991,N_14859,N_14720);
and U14992 (N_14992,N_14837,N_14750);
nand U14993 (N_14993,N_14819,N_14789);
or U14994 (N_14994,N_14760,N_14862);
nand U14995 (N_14995,N_14739,N_14728);
and U14996 (N_14996,N_14874,N_14859);
nand U14997 (N_14997,N_14768,N_14748);
or U14998 (N_14998,N_14833,N_14753);
or U14999 (N_14999,N_14854,N_14750);
xnor U15000 (N_15000,N_14867,N_14828);
and U15001 (N_15001,N_14770,N_14790);
nor U15002 (N_15002,N_14811,N_14760);
or U15003 (N_15003,N_14747,N_14835);
nor U15004 (N_15004,N_14844,N_14786);
nand U15005 (N_15005,N_14870,N_14767);
nor U15006 (N_15006,N_14759,N_14842);
nor U15007 (N_15007,N_14779,N_14802);
and U15008 (N_15008,N_14723,N_14796);
or U15009 (N_15009,N_14816,N_14743);
nand U15010 (N_15010,N_14820,N_14860);
and U15011 (N_15011,N_14803,N_14785);
nand U15012 (N_15012,N_14809,N_14838);
xor U15013 (N_15013,N_14824,N_14720);
nor U15014 (N_15014,N_14810,N_14879);
and U15015 (N_15015,N_14801,N_14752);
xnor U15016 (N_15016,N_14731,N_14750);
and U15017 (N_15017,N_14811,N_14852);
or U15018 (N_15018,N_14826,N_14822);
and U15019 (N_15019,N_14796,N_14748);
nand U15020 (N_15020,N_14759,N_14744);
xor U15021 (N_15021,N_14776,N_14846);
or U15022 (N_15022,N_14816,N_14771);
nand U15023 (N_15023,N_14752,N_14744);
xor U15024 (N_15024,N_14737,N_14825);
nand U15025 (N_15025,N_14803,N_14826);
nand U15026 (N_15026,N_14878,N_14810);
and U15027 (N_15027,N_14755,N_14839);
nor U15028 (N_15028,N_14762,N_14878);
xor U15029 (N_15029,N_14816,N_14761);
nor U15030 (N_15030,N_14833,N_14829);
xnor U15031 (N_15031,N_14797,N_14721);
and U15032 (N_15032,N_14857,N_14816);
nor U15033 (N_15033,N_14745,N_14773);
nor U15034 (N_15034,N_14872,N_14850);
nor U15035 (N_15035,N_14721,N_14767);
nand U15036 (N_15036,N_14835,N_14866);
and U15037 (N_15037,N_14839,N_14805);
and U15038 (N_15038,N_14825,N_14876);
nor U15039 (N_15039,N_14779,N_14788);
and U15040 (N_15040,N_14992,N_14962);
or U15041 (N_15041,N_15005,N_15013);
and U15042 (N_15042,N_14976,N_14950);
or U15043 (N_15043,N_14902,N_14898);
xor U15044 (N_15044,N_15018,N_14941);
and U15045 (N_15045,N_15028,N_14978);
and U15046 (N_15046,N_14980,N_14972);
and U15047 (N_15047,N_15021,N_14964);
and U15048 (N_15048,N_14905,N_14921);
nor U15049 (N_15049,N_15027,N_15020);
or U15050 (N_15050,N_15034,N_14987);
or U15051 (N_15051,N_15009,N_14938);
and U15052 (N_15052,N_14940,N_15016);
nand U15053 (N_15053,N_14882,N_14925);
nor U15054 (N_15054,N_14883,N_14995);
and U15055 (N_15055,N_14909,N_14954);
nor U15056 (N_15056,N_14977,N_14997);
nand U15057 (N_15057,N_14931,N_14918);
nor U15058 (N_15058,N_15014,N_15002);
and U15059 (N_15059,N_14919,N_15029);
or U15060 (N_15060,N_14924,N_14994);
xnor U15061 (N_15061,N_14990,N_14979);
and U15062 (N_15062,N_14891,N_14965);
and U15063 (N_15063,N_14900,N_14966);
nand U15064 (N_15064,N_15017,N_14959);
or U15065 (N_15065,N_14951,N_14906);
nand U15066 (N_15066,N_14970,N_14910);
and U15067 (N_15067,N_14963,N_14881);
and U15068 (N_15068,N_14920,N_14880);
nand U15069 (N_15069,N_14958,N_15024);
nand U15070 (N_15070,N_14989,N_14968);
nand U15071 (N_15071,N_14934,N_14932);
nand U15072 (N_15072,N_15019,N_14985);
or U15073 (N_15073,N_14939,N_14929);
nand U15074 (N_15074,N_14991,N_14969);
nor U15075 (N_15075,N_14901,N_14897);
or U15076 (N_15076,N_15003,N_14890);
and U15077 (N_15077,N_14894,N_14911);
xnor U15078 (N_15078,N_14993,N_15023);
nor U15079 (N_15079,N_14904,N_15038);
nor U15080 (N_15080,N_14998,N_14949);
xor U15081 (N_15081,N_14935,N_14927);
xor U15082 (N_15082,N_14999,N_15035);
or U15083 (N_15083,N_14884,N_14996);
nor U15084 (N_15084,N_14899,N_14915);
nand U15085 (N_15085,N_14937,N_14895);
nand U15086 (N_15086,N_14946,N_14988);
nor U15087 (N_15087,N_14907,N_14892);
nand U15088 (N_15088,N_15006,N_15037);
nand U15089 (N_15089,N_14914,N_14916);
or U15090 (N_15090,N_14912,N_15036);
and U15091 (N_15091,N_14888,N_14971);
nor U15092 (N_15092,N_14984,N_14922);
nor U15093 (N_15093,N_15001,N_14967);
nand U15094 (N_15094,N_14948,N_15033);
xnor U15095 (N_15095,N_14947,N_14983);
nor U15096 (N_15096,N_14893,N_15025);
and U15097 (N_15097,N_14981,N_14942);
or U15098 (N_15098,N_14933,N_14975);
nor U15099 (N_15099,N_15030,N_14956);
or U15100 (N_15100,N_15000,N_14974);
xor U15101 (N_15101,N_14903,N_15012);
or U15102 (N_15102,N_15011,N_14928);
xnor U15103 (N_15103,N_15015,N_15022);
or U15104 (N_15104,N_15010,N_14896);
or U15105 (N_15105,N_14952,N_14930);
and U15106 (N_15106,N_14960,N_14986);
xor U15107 (N_15107,N_14923,N_15007);
and U15108 (N_15108,N_14885,N_14926);
xnor U15109 (N_15109,N_14943,N_14982);
or U15110 (N_15110,N_14944,N_14913);
nand U15111 (N_15111,N_15026,N_14889);
nand U15112 (N_15112,N_15032,N_14908);
and U15113 (N_15113,N_15039,N_14953);
nor U15114 (N_15114,N_14955,N_14961);
xnor U15115 (N_15115,N_14917,N_14936);
nor U15116 (N_15116,N_14957,N_15031);
or U15117 (N_15117,N_15008,N_14886);
nand U15118 (N_15118,N_14945,N_14973);
nand U15119 (N_15119,N_15004,N_14887);
and U15120 (N_15120,N_14934,N_14888);
and U15121 (N_15121,N_14930,N_14936);
nor U15122 (N_15122,N_14985,N_14943);
or U15123 (N_15123,N_14920,N_14959);
xnor U15124 (N_15124,N_14981,N_14957);
and U15125 (N_15125,N_14961,N_14974);
or U15126 (N_15126,N_14951,N_15010);
xor U15127 (N_15127,N_14931,N_14985);
and U15128 (N_15128,N_14901,N_15029);
and U15129 (N_15129,N_14914,N_14932);
and U15130 (N_15130,N_14880,N_15038);
nand U15131 (N_15131,N_14921,N_15039);
and U15132 (N_15132,N_14885,N_15011);
nor U15133 (N_15133,N_15029,N_14897);
or U15134 (N_15134,N_15017,N_14977);
and U15135 (N_15135,N_14993,N_14968);
nand U15136 (N_15136,N_15011,N_14883);
or U15137 (N_15137,N_15037,N_14907);
or U15138 (N_15138,N_14917,N_14940);
nand U15139 (N_15139,N_14902,N_14949);
and U15140 (N_15140,N_14945,N_14917);
nand U15141 (N_15141,N_14978,N_15034);
nor U15142 (N_15142,N_14909,N_14887);
or U15143 (N_15143,N_14952,N_14982);
nor U15144 (N_15144,N_14939,N_15024);
and U15145 (N_15145,N_14902,N_14906);
or U15146 (N_15146,N_15039,N_14896);
xnor U15147 (N_15147,N_14942,N_15009);
and U15148 (N_15148,N_14905,N_14937);
and U15149 (N_15149,N_14919,N_15030);
xnor U15150 (N_15150,N_14988,N_15038);
and U15151 (N_15151,N_14919,N_14971);
nor U15152 (N_15152,N_14986,N_14945);
or U15153 (N_15153,N_14952,N_14953);
nand U15154 (N_15154,N_14969,N_14933);
nand U15155 (N_15155,N_15036,N_14906);
nand U15156 (N_15156,N_15015,N_14880);
nand U15157 (N_15157,N_14909,N_15003);
xnor U15158 (N_15158,N_14939,N_14916);
and U15159 (N_15159,N_14899,N_14945);
nand U15160 (N_15160,N_14950,N_15024);
and U15161 (N_15161,N_15011,N_14963);
and U15162 (N_15162,N_14978,N_14916);
xor U15163 (N_15163,N_14987,N_14927);
nand U15164 (N_15164,N_14912,N_14882);
and U15165 (N_15165,N_14974,N_15011);
and U15166 (N_15166,N_14937,N_14915);
and U15167 (N_15167,N_14969,N_14884);
nor U15168 (N_15168,N_15012,N_14965);
and U15169 (N_15169,N_15010,N_15017);
or U15170 (N_15170,N_14979,N_15028);
nor U15171 (N_15171,N_14974,N_15029);
and U15172 (N_15172,N_14971,N_14994);
xnor U15173 (N_15173,N_14915,N_15003);
and U15174 (N_15174,N_14912,N_14899);
nand U15175 (N_15175,N_15027,N_14985);
and U15176 (N_15176,N_15029,N_14954);
nand U15177 (N_15177,N_15020,N_15009);
nor U15178 (N_15178,N_15020,N_14942);
xnor U15179 (N_15179,N_14994,N_14983);
xnor U15180 (N_15180,N_15000,N_15017);
xor U15181 (N_15181,N_14945,N_14908);
nor U15182 (N_15182,N_14997,N_14950);
nor U15183 (N_15183,N_14892,N_14964);
and U15184 (N_15184,N_15037,N_15007);
nand U15185 (N_15185,N_14904,N_14973);
and U15186 (N_15186,N_14921,N_15035);
nor U15187 (N_15187,N_14994,N_14913);
xnor U15188 (N_15188,N_14881,N_15011);
or U15189 (N_15189,N_14928,N_15002);
or U15190 (N_15190,N_14988,N_15024);
and U15191 (N_15191,N_14931,N_14946);
xor U15192 (N_15192,N_14967,N_14882);
nand U15193 (N_15193,N_14964,N_14903);
nand U15194 (N_15194,N_14899,N_14931);
nor U15195 (N_15195,N_14977,N_14961);
xor U15196 (N_15196,N_14894,N_14925);
nand U15197 (N_15197,N_15024,N_14965);
nor U15198 (N_15198,N_14991,N_14931);
nor U15199 (N_15199,N_14949,N_14945);
and U15200 (N_15200,N_15119,N_15145);
or U15201 (N_15201,N_15064,N_15084);
or U15202 (N_15202,N_15089,N_15163);
xnor U15203 (N_15203,N_15093,N_15161);
nor U15204 (N_15204,N_15047,N_15196);
nor U15205 (N_15205,N_15056,N_15147);
nor U15206 (N_15206,N_15199,N_15104);
nor U15207 (N_15207,N_15054,N_15085);
xnor U15208 (N_15208,N_15045,N_15137);
and U15209 (N_15209,N_15197,N_15059);
and U15210 (N_15210,N_15156,N_15158);
nand U15211 (N_15211,N_15080,N_15055);
and U15212 (N_15212,N_15051,N_15164);
xor U15213 (N_15213,N_15072,N_15166);
nand U15214 (N_15214,N_15063,N_15133);
and U15215 (N_15215,N_15125,N_15132);
or U15216 (N_15216,N_15136,N_15173);
nand U15217 (N_15217,N_15171,N_15139);
nand U15218 (N_15218,N_15094,N_15127);
nand U15219 (N_15219,N_15135,N_15068);
nor U15220 (N_15220,N_15131,N_15146);
nor U15221 (N_15221,N_15151,N_15193);
nand U15222 (N_15222,N_15101,N_15073);
xnor U15223 (N_15223,N_15046,N_15062);
nand U15224 (N_15224,N_15181,N_15184);
xor U15225 (N_15225,N_15042,N_15120);
nand U15226 (N_15226,N_15088,N_15191);
or U15227 (N_15227,N_15187,N_15178);
and U15228 (N_15228,N_15162,N_15070);
nand U15229 (N_15229,N_15061,N_15076);
xnor U15230 (N_15230,N_15109,N_15040);
nor U15231 (N_15231,N_15179,N_15103);
nor U15232 (N_15232,N_15149,N_15078);
xor U15233 (N_15233,N_15044,N_15105);
and U15234 (N_15234,N_15067,N_15150);
nor U15235 (N_15235,N_15160,N_15107);
nand U15236 (N_15236,N_15053,N_15118);
and U15237 (N_15237,N_15092,N_15071);
nand U15238 (N_15238,N_15129,N_15140);
nand U15239 (N_15239,N_15102,N_15192);
xnor U15240 (N_15240,N_15087,N_15077);
nor U15241 (N_15241,N_15195,N_15048);
and U15242 (N_15242,N_15153,N_15113);
nor U15243 (N_15243,N_15110,N_15096);
nand U15244 (N_15244,N_15086,N_15126);
and U15245 (N_15245,N_15112,N_15177);
nand U15246 (N_15246,N_15095,N_15041);
nor U15247 (N_15247,N_15052,N_15081);
or U15248 (N_15248,N_15188,N_15189);
nand U15249 (N_15249,N_15194,N_15098);
nand U15250 (N_15250,N_15058,N_15182);
nor U15251 (N_15251,N_15090,N_15183);
xor U15252 (N_15252,N_15123,N_15043);
or U15253 (N_15253,N_15114,N_15190);
xnor U15254 (N_15254,N_15165,N_15116);
and U15255 (N_15255,N_15176,N_15091);
nand U15256 (N_15256,N_15154,N_15124);
and U15257 (N_15257,N_15134,N_15185);
xor U15258 (N_15258,N_15128,N_15172);
nand U15259 (N_15259,N_15168,N_15141);
and U15260 (N_15260,N_15144,N_15097);
nand U15261 (N_15261,N_15075,N_15175);
nor U15262 (N_15262,N_15167,N_15115);
or U15263 (N_15263,N_15198,N_15130);
nor U15264 (N_15264,N_15108,N_15074);
or U15265 (N_15265,N_15148,N_15111);
and U15266 (N_15266,N_15138,N_15155);
or U15267 (N_15267,N_15117,N_15186);
and U15268 (N_15268,N_15057,N_15157);
nand U15269 (N_15269,N_15082,N_15100);
nand U15270 (N_15270,N_15069,N_15050);
nand U15271 (N_15271,N_15121,N_15083);
nor U15272 (N_15272,N_15180,N_15159);
and U15273 (N_15273,N_15142,N_15066);
and U15274 (N_15274,N_15099,N_15122);
and U15275 (N_15275,N_15174,N_15169);
and U15276 (N_15276,N_15152,N_15060);
or U15277 (N_15277,N_15065,N_15106);
nor U15278 (N_15278,N_15049,N_15079);
nand U15279 (N_15279,N_15143,N_15170);
nor U15280 (N_15280,N_15062,N_15086);
or U15281 (N_15281,N_15166,N_15182);
nor U15282 (N_15282,N_15064,N_15087);
nor U15283 (N_15283,N_15044,N_15184);
xor U15284 (N_15284,N_15040,N_15175);
nor U15285 (N_15285,N_15126,N_15057);
nand U15286 (N_15286,N_15105,N_15046);
xor U15287 (N_15287,N_15179,N_15048);
xor U15288 (N_15288,N_15057,N_15146);
nor U15289 (N_15289,N_15096,N_15081);
xor U15290 (N_15290,N_15059,N_15071);
xor U15291 (N_15291,N_15096,N_15056);
nand U15292 (N_15292,N_15062,N_15166);
and U15293 (N_15293,N_15187,N_15193);
nand U15294 (N_15294,N_15069,N_15163);
nor U15295 (N_15295,N_15118,N_15074);
and U15296 (N_15296,N_15075,N_15156);
nand U15297 (N_15297,N_15197,N_15068);
and U15298 (N_15298,N_15171,N_15059);
nand U15299 (N_15299,N_15106,N_15140);
nand U15300 (N_15300,N_15196,N_15139);
xnor U15301 (N_15301,N_15055,N_15154);
nand U15302 (N_15302,N_15120,N_15165);
and U15303 (N_15303,N_15133,N_15155);
nand U15304 (N_15304,N_15150,N_15186);
or U15305 (N_15305,N_15123,N_15102);
nand U15306 (N_15306,N_15194,N_15145);
or U15307 (N_15307,N_15164,N_15198);
and U15308 (N_15308,N_15084,N_15139);
and U15309 (N_15309,N_15164,N_15146);
nor U15310 (N_15310,N_15189,N_15045);
nand U15311 (N_15311,N_15067,N_15180);
xor U15312 (N_15312,N_15138,N_15183);
or U15313 (N_15313,N_15064,N_15184);
or U15314 (N_15314,N_15135,N_15054);
nor U15315 (N_15315,N_15154,N_15159);
nand U15316 (N_15316,N_15148,N_15089);
nand U15317 (N_15317,N_15166,N_15145);
or U15318 (N_15318,N_15159,N_15140);
or U15319 (N_15319,N_15116,N_15153);
nor U15320 (N_15320,N_15122,N_15050);
nor U15321 (N_15321,N_15080,N_15186);
nand U15322 (N_15322,N_15087,N_15150);
nor U15323 (N_15323,N_15059,N_15040);
or U15324 (N_15324,N_15148,N_15068);
and U15325 (N_15325,N_15128,N_15081);
nor U15326 (N_15326,N_15072,N_15074);
and U15327 (N_15327,N_15059,N_15198);
nand U15328 (N_15328,N_15166,N_15084);
nor U15329 (N_15329,N_15171,N_15149);
and U15330 (N_15330,N_15046,N_15132);
nand U15331 (N_15331,N_15115,N_15161);
and U15332 (N_15332,N_15157,N_15125);
or U15333 (N_15333,N_15080,N_15177);
xnor U15334 (N_15334,N_15111,N_15166);
and U15335 (N_15335,N_15051,N_15170);
nor U15336 (N_15336,N_15078,N_15161);
nor U15337 (N_15337,N_15074,N_15137);
xnor U15338 (N_15338,N_15195,N_15100);
nand U15339 (N_15339,N_15049,N_15151);
and U15340 (N_15340,N_15181,N_15195);
xnor U15341 (N_15341,N_15050,N_15100);
and U15342 (N_15342,N_15135,N_15108);
and U15343 (N_15343,N_15107,N_15051);
nor U15344 (N_15344,N_15062,N_15095);
and U15345 (N_15345,N_15132,N_15154);
nor U15346 (N_15346,N_15150,N_15069);
xor U15347 (N_15347,N_15146,N_15094);
nand U15348 (N_15348,N_15171,N_15165);
or U15349 (N_15349,N_15184,N_15177);
or U15350 (N_15350,N_15131,N_15040);
nand U15351 (N_15351,N_15150,N_15118);
nor U15352 (N_15352,N_15198,N_15107);
or U15353 (N_15353,N_15196,N_15046);
nand U15354 (N_15354,N_15167,N_15053);
nor U15355 (N_15355,N_15097,N_15089);
or U15356 (N_15356,N_15154,N_15187);
or U15357 (N_15357,N_15191,N_15150);
or U15358 (N_15358,N_15105,N_15086);
and U15359 (N_15359,N_15087,N_15103);
and U15360 (N_15360,N_15352,N_15233);
or U15361 (N_15361,N_15282,N_15227);
and U15362 (N_15362,N_15247,N_15260);
nor U15363 (N_15363,N_15236,N_15310);
nand U15364 (N_15364,N_15250,N_15205);
or U15365 (N_15365,N_15294,N_15289);
and U15366 (N_15366,N_15330,N_15311);
and U15367 (N_15367,N_15223,N_15312);
or U15368 (N_15368,N_15217,N_15219);
and U15369 (N_15369,N_15345,N_15305);
and U15370 (N_15370,N_15254,N_15208);
nor U15371 (N_15371,N_15256,N_15241);
nor U15372 (N_15372,N_15317,N_15277);
nor U15373 (N_15373,N_15339,N_15350);
nor U15374 (N_15374,N_15213,N_15320);
nor U15375 (N_15375,N_15235,N_15270);
and U15376 (N_15376,N_15334,N_15251);
and U15377 (N_15377,N_15353,N_15264);
or U15378 (N_15378,N_15321,N_15257);
or U15379 (N_15379,N_15287,N_15207);
nor U15380 (N_15380,N_15234,N_15304);
or U15381 (N_15381,N_15252,N_15301);
nor U15382 (N_15382,N_15333,N_15303);
and U15383 (N_15383,N_15245,N_15242);
nand U15384 (N_15384,N_15232,N_15324);
xnor U15385 (N_15385,N_15238,N_15275);
nor U15386 (N_15386,N_15284,N_15265);
and U15387 (N_15387,N_15271,N_15300);
nor U15388 (N_15388,N_15239,N_15231);
nor U15389 (N_15389,N_15206,N_15212);
nand U15390 (N_15390,N_15273,N_15209);
and U15391 (N_15391,N_15210,N_15279);
or U15392 (N_15392,N_15225,N_15296);
and U15393 (N_15393,N_15261,N_15344);
nand U15394 (N_15394,N_15295,N_15338);
nor U15395 (N_15395,N_15288,N_15268);
nand U15396 (N_15396,N_15307,N_15244);
nor U15397 (N_15397,N_15337,N_15259);
nand U15398 (N_15398,N_15281,N_15220);
nor U15399 (N_15399,N_15258,N_15297);
nand U15400 (N_15400,N_15349,N_15328);
nand U15401 (N_15401,N_15286,N_15354);
nor U15402 (N_15402,N_15292,N_15359);
nor U15403 (N_15403,N_15229,N_15329);
nand U15404 (N_15404,N_15331,N_15322);
nand U15405 (N_15405,N_15230,N_15298);
nand U15406 (N_15406,N_15218,N_15318);
nand U15407 (N_15407,N_15224,N_15336);
nor U15408 (N_15408,N_15342,N_15262);
nand U15409 (N_15409,N_15348,N_15306);
xnor U15410 (N_15410,N_15203,N_15202);
and U15411 (N_15411,N_15278,N_15243);
or U15412 (N_15412,N_15248,N_15316);
nor U15413 (N_15413,N_15253,N_15274);
or U15414 (N_15414,N_15263,N_15214);
or U15415 (N_15415,N_15276,N_15269);
nand U15416 (N_15416,N_15343,N_15285);
nor U15417 (N_15417,N_15200,N_15335);
and U15418 (N_15418,N_15246,N_15308);
nand U15419 (N_15419,N_15358,N_15249);
or U15420 (N_15420,N_15290,N_15346);
nor U15421 (N_15421,N_15326,N_15267);
or U15422 (N_15422,N_15299,N_15216);
nor U15423 (N_15423,N_15215,N_15266);
or U15424 (N_15424,N_15315,N_15237);
and U15425 (N_15425,N_15293,N_15341);
nand U15426 (N_15426,N_15291,N_15325);
nor U15427 (N_15427,N_15355,N_15211);
nand U15428 (N_15428,N_15280,N_15240);
nor U15429 (N_15429,N_15204,N_15302);
nand U15430 (N_15430,N_15309,N_15283);
or U15431 (N_15431,N_15347,N_15222);
nand U15432 (N_15432,N_15340,N_15332);
or U15433 (N_15433,N_15313,N_15272);
or U15434 (N_15434,N_15255,N_15323);
or U15435 (N_15435,N_15201,N_15351);
nand U15436 (N_15436,N_15327,N_15314);
and U15437 (N_15437,N_15221,N_15319);
nor U15438 (N_15438,N_15228,N_15356);
or U15439 (N_15439,N_15357,N_15226);
nand U15440 (N_15440,N_15330,N_15285);
or U15441 (N_15441,N_15341,N_15236);
nor U15442 (N_15442,N_15202,N_15217);
or U15443 (N_15443,N_15310,N_15265);
nor U15444 (N_15444,N_15319,N_15310);
and U15445 (N_15445,N_15234,N_15312);
nor U15446 (N_15446,N_15223,N_15221);
nor U15447 (N_15447,N_15204,N_15255);
nand U15448 (N_15448,N_15269,N_15334);
nand U15449 (N_15449,N_15275,N_15265);
and U15450 (N_15450,N_15342,N_15211);
nor U15451 (N_15451,N_15333,N_15218);
nor U15452 (N_15452,N_15266,N_15324);
and U15453 (N_15453,N_15315,N_15303);
xnor U15454 (N_15454,N_15211,N_15265);
nand U15455 (N_15455,N_15200,N_15329);
nand U15456 (N_15456,N_15246,N_15271);
nand U15457 (N_15457,N_15226,N_15209);
xor U15458 (N_15458,N_15260,N_15259);
xor U15459 (N_15459,N_15338,N_15349);
nand U15460 (N_15460,N_15263,N_15255);
xnor U15461 (N_15461,N_15339,N_15359);
or U15462 (N_15462,N_15346,N_15245);
nor U15463 (N_15463,N_15328,N_15342);
or U15464 (N_15464,N_15217,N_15300);
nor U15465 (N_15465,N_15200,N_15253);
nand U15466 (N_15466,N_15279,N_15308);
nor U15467 (N_15467,N_15230,N_15338);
nand U15468 (N_15468,N_15290,N_15241);
xor U15469 (N_15469,N_15210,N_15339);
nand U15470 (N_15470,N_15242,N_15322);
nand U15471 (N_15471,N_15294,N_15297);
nand U15472 (N_15472,N_15311,N_15357);
and U15473 (N_15473,N_15312,N_15294);
and U15474 (N_15474,N_15240,N_15281);
xor U15475 (N_15475,N_15202,N_15292);
and U15476 (N_15476,N_15345,N_15227);
xnor U15477 (N_15477,N_15330,N_15243);
nor U15478 (N_15478,N_15209,N_15298);
nand U15479 (N_15479,N_15316,N_15209);
or U15480 (N_15480,N_15266,N_15297);
or U15481 (N_15481,N_15327,N_15343);
nor U15482 (N_15482,N_15258,N_15307);
or U15483 (N_15483,N_15338,N_15200);
nor U15484 (N_15484,N_15341,N_15309);
or U15485 (N_15485,N_15291,N_15295);
nand U15486 (N_15486,N_15307,N_15339);
nor U15487 (N_15487,N_15338,N_15352);
or U15488 (N_15488,N_15232,N_15280);
nor U15489 (N_15489,N_15306,N_15291);
nand U15490 (N_15490,N_15351,N_15358);
nand U15491 (N_15491,N_15353,N_15222);
or U15492 (N_15492,N_15231,N_15298);
or U15493 (N_15493,N_15337,N_15246);
nor U15494 (N_15494,N_15202,N_15333);
nand U15495 (N_15495,N_15315,N_15277);
nand U15496 (N_15496,N_15200,N_15315);
nand U15497 (N_15497,N_15205,N_15255);
nand U15498 (N_15498,N_15202,N_15229);
and U15499 (N_15499,N_15287,N_15229);
nor U15500 (N_15500,N_15203,N_15283);
or U15501 (N_15501,N_15282,N_15252);
or U15502 (N_15502,N_15227,N_15290);
or U15503 (N_15503,N_15267,N_15353);
nand U15504 (N_15504,N_15335,N_15207);
xor U15505 (N_15505,N_15235,N_15254);
or U15506 (N_15506,N_15269,N_15343);
and U15507 (N_15507,N_15221,N_15354);
or U15508 (N_15508,N_15304,N_15322);
and U15509 (N_15509,N_15322,N_15334);
xor U15510 (N_15510,N_15262,N_15239);
and U15511 (N_15511,N_15212,N_15296);
or U15512 (N_15512,N_15336,N_15201);
and U15513 (N_15513,N_15319,N_15290);
or U15514 (N_15514,N_15255,N_15209);
and U15515 (N_15515,N_15263,N_15355);
or U15516 (N_15516,N_15204,N_15288);
or U15517 (N_15517,N_15220,N_15307);
or U15518 (N_15518,N_15302,N_15268);
and U15519 (N_15519,N_15213,N_15276);
nand U15520 (N_15520,N_15392,N_15395);
nor U15521 (N_15521,N_15504,N_15390);
or U15522 (N_15522,N_15447,N_15427);
and U15523 (N_15523,N_15462,N_15443);
or U15524 (N_15524,N_15380,N_15430);
nand U15525 (N_15525,N_15498,N_15436);
xor U15526 (N_15526,N_15481,N_15410);
and U15527 (N_15527,N_15367,N_15373);
nor U15528 (N_15528,N_15490,N_15381);
or U15529 (N_15529,N_15433,N_15508);
or U15530 (N_15530,N_15453,N_15489);
nor U15531 (N_15531,N_15362,N_15467);
xor U15532 (N_15532,N_15431,N_15484);
or U15533 (N_15533,N_15474,N_15421);
nand U15534 (N_15534,N_15406,N_15376);
and U15535 (N_15535,N_15411,N_15510);
nor U15536 (N_15536,N_15385,N_15459);
or U15537 (N_15537,N_15448,N_15505);
nand U15538 (N_15538,N_15394,N_15440);
or U15539 (N_15539,N_15519,N_15438);
or U15540 (N_15540,N_15400,N_15384);
xnor U15541 (N_15541,N_15449,N_15457);
and U15542 (N_15542,N_15401,N_15425);
nand U15543 (N_15543,N_15468,N_15458);
nor U15544 (N_15544,N_15399,N_15383);
nand U15545 (N_15545,N_15428,N_15461);
nor U15546 (N_15546,N_15407,N_15469);
and U15547 (N_15547,N_15471,N_15413);
nand U15548 (N_15548,N_15497,N_15450);
and U15549 (N_15549,N_15402,N_15493);
or U15550 (N_15550,N_15404,N_15432);
or U15551 (N_15551,N_15398,N_15397);
nor U15552 (N_15552,N_15364,N_15517);
nand U15553 (N_15553,N_15420,N_15502);
nand U15554 (N_15554,N_15518,N_15415);
or U15555 (N_15555,N_15513,N_15377);
nand U15556 (N_15556,N_15492,N_15422);
nor U15557 (N_15557,N_15374,N_15516);
nand U15558 (N_15558,N_15500,N_15485);
nand U15559 (N_15559,N_15366,N_15414);
nand U15560 (N_15560,N_15465,N_15408);
xor U15561 (N_15561,N_15509,N_15506);
xor U15562 (N_15562,N_15491,N_15486);
nor U15563 (N_15563,N_15463,N_15393);
xnor U15564 (N_15564,N_15451,N_15507);
nand U15565 (N_15565,N_15429,N_15455);
and U15566 (N_15566,N_15379,N_15499);
xnor U15567 (N_15567,N_15442,N_15405);
or U15568 (N_15568,N_15487,N_15419);
nor U15569 (N_15569,N_15488,N_15389);
and U15570 (N_15570,N_15424,N_15360);
or U15571 (N_15571,N_15483,N_15470);
and U15572 (N_15572,N_15512,N_15386);
nor U15573 (N_15573,N_15372,N_15466);
nand U15574 (N_15574,N_15444,N_15480);
nand U15575 (N_15575,N_15472,N_15479);
and U15576 (N_15576,N_15503,N_15454);
or U15577 (N_15577,N_15426,N_15370);
nor U15578 (N_15578,N_15417,N_15371);
xor U15579 (N_15579,N_15476,N_15473);
nor U15580 (N_15580,N_15435,N_15501);
nor U15581 (N_15581,N_15494,N_15478);
nor U15582 (N_15582,N_15495,N_15446);
nor U15583 (N_15583,N_15456,N_15396);
nor U15584 (N_15584,N_15368,N_15416);
or U15585 (N_15585,N_15378,N_15482);
or U15586 (N_15586,N_15412,N_15445);
nand U15587 (N_15587,N_15460,N_15418);
and U15588 (N_15588,N_15514,N_15496);
and U15589 (N_15589,N_15403,N_15511);
and U15590 (N_15590,N_15369,N_15437);
nor U15591 (N_15591,N_15387,N_15382);
or U15592 (N_15592,N_15441,N_15452);
and U15593 (N_15593,N_15434,N_15388);
nor U15594 (N_15594,N_15439,N_15477);
and U15595 (N_15595,N_15375,N_15475);
and U15596 (N_15596,N_15423,N_15365);
xnor U15597 (N_15597,N_15363,N_15464);
nor U15598 (N_15598,N_15409,N_15391);
nand U15599 (N_15599,N_15515,N_15361);
and U15600 (N_15600,N_15476,N_15414);
nor U15601 (N_15601,N_15466,N_15399);
or U15602 (N_15602,N_15397,N_15515);
and U15603 (N_15603,N_15381,N_15382);
nor U15604 (N_15604,N_15439,N_15442);
or U15605 (N_15605,N_15364,N_15476);
nor U15606 (N_15606,N_15392,N_15444);
or U15607 (N_15607,N_15509,N_15505);
nand U15608 (N_15608,N_15435,N_15461);
nor U15609 (N_15609,N_15471,N_15477);
xor U15610 (N_15610,N_15421,N_15437);
or U15611 (N_15611,N_15515,N_15432);
or U15612 (N_15612,N_15394,N_15424);
nand U15613 (N_15613,N_15489,N_15447);
or U15614 (N_15614,N_15468,N_15446);
or U15615 (N_15615,N_15423,N_15411);
nand U15616 (N_15616,N_15427,N_15519);
nor U15617 (N_15617,N_15445,N_15417);
nor U15618 (N_15618,N_15467,N_15494);
nor U15619 (N_15619,N_15440,N_15511);
or U15620 (N_15620,N_15472,N_15414);
or U15621 (N_15621,N_15457,N_15463);
nand U15622 (N_15622,N_15510,N_15404);
or U15623 (N_15623,N_15415,N_15464);
nand U15624 (N_15624,N_15376,N_15369);
or U15625 (N_15625,N_15502,N_15468);
or U15626 (N_15626,N_15507,N_15361);
nor U15627 (N_15627,N_15472,N_15415);
or U15628 (N_15628,N_15435,N_15471);
nor U15629 (N_15629,N_15473,N_15462);
nand U15630 (N_15630,N_15379,N_15391);
nor U15631 (N_15631,N_15483,N_15412);
nor U15632 (N_15632,N_15449,N_15463);
nor U15633 (N_15633,N_15400,N_15415);
or U15634 (N_15634,N_15503,N_15452);
nor U15635 (N_15635,N_15417,N_15387);
nor U15636 (N_15636,N_15418,N_15402);
xor U15637 (N_15637,N_15433,N_15487);
xnor U15638 (N_15638,N_15415,N_15513);
xnor U15639 (N_15639,N_15406,N_15400);
xnor U15640 (N_15640,N_15428,N_15394);
nor U15641 (N_15641,N_15401,N_15478);
and U15642 (N_15642,N_15377,N_15501);
nand U15643 (N_15643,N_15455,N_15423);
and U15644 (N_15644,N_15380,N_15460);
nand U15645 (N_15645,N_15393,N_15412);
or U15646 (N_15646,N_15395,N_15418);
xor U15647 (N_15647,N_15422,N_15395);
or U15648 (N_15648,N_15511,N_15414);
and U15649 (N_15649,N_15404,N_15455);
nand U15650 (N_15650,N_15442,N_15512);
nor U15651 (N_15651,N_15429,N_15487);
nor U15652 (N_15652,N_15431,N_15425);
nand U15653 (N_15653,N_15365,N_15394);
or U15654 (N_15654,N_15457,N_15393);
nor U15655 (N_15655,N_15451,N_15508);
or U15656 (N_15656,N_15493,N_15407);
nand U15657 (N_15657,N_15456,N_15369);
nor U15658 (N_15658,N_15447,N_15511);
and U15659 (N_15659,N_15454,N_15439);
nor U15660 (N_15660,N_15470,N_15412);
or U15661 (N_15661,N_15459,N_15452);
xor U15662 (N_15662,N_15374,N_15368);
nor U15663 (N_15663,N_15458,N_15364);
xor U15664 (N_15664,N_15369,N_15471);
or U15665 (N_15665,N_15482,N_15418);
xor U15666 (N_15666,N_15494,N_15516);
nand U15667 (N_15667,N_15420,N_15373);
nor U15668 (N_15668,N_15423,N_15471);
xor U15669 (N_15669,N_15506,N_15430);
nor U15670 (N_15670,N_15387,N_15451);
or U15671 (N_15671,N_15407,N_15390);
and U15672 (N_15672,N_15410,N_15360);
nand U15673 (N_15673,N_15381,N_15372);
nand U15674 (N_15674,N_15430,N_15478);
xor U15675 (N_15675,N_15474,N_15388);
nor U15676 (N_15676,N_15373,N_15511);
nor U15677 (N_15677,N_15459,N_15431);
nor U15678 (N_15678,N_15505,N_15378);
xnor U15679 (N_15679,N_15474,N_15473);
or U15680 (N_15680,N_15575,N_15648);
or U15681 (N_15681,N_15586,N_15538);
nor U15682 (N_15682,N_15617,N_15626);
nor U15683 (N_15683,N_15633,N_15590);
nor U15684 (N_15684,N_15663,N_15523);
nor U15685 (N_15685,N_15536,N_15566);
xor U15686 (N_15686,N_15591,N_15585);
and U15687 (N_15687,N_15602,N_15580);
nor U15688 (N_15688,N_15544,N_15641);
nand U15689 (N_15689,N_15659,N_15646);
xor U15690 (N_15690,N_15561,N_15645);
nand U15691 (N_15691,N_15603,N_15587);
and U15692 (N_15692,N_15653,N_15522);
or U15693 (N_15693,N_15627,N_15572);
nor U15694 (N_15694,N_15540,N_15598);
nand U15695 (N_15695,N_15573,N_15657);
nor U15696 (N_15696,N_15570,N_15640);
and U15697 (N_15697,N_15619,N_15562);
nor U15698 (N_15698,N_15565,N_15604);
and U15699 (N_15699,N_15616,N_15678);
nor U15700 (N_15700,N_15609,N_15525);
nand U15701 (N_15701,N_15545,N_15599);
nor U15702 (N_15702,N_15569,N_15661);
nor U15703 (N_15703,N_15652,N_15531);
xor U15704 (N_15704,N_15529,N_15608);
nor U15705 (N_15705,N_15625,N_15632);
xor U15706 (N_15706,N_15669,N_15611);
and U15707 (N_15707,N_15672,N_15556);
nor U15708 (N_15708,N_15612,N_15601);
nand U15709 (N_15709,N_15621,N_15624);
and U15710 (N_15710,N_15660,N_15597);
or U15711 (N_15711,N_15647,N_15635);
or U15712 (N_15712,N_15539,N_15614);
or U15713 (N_15713,N_15662,N_15579);
or U15714 (N_15714,N_15592,N_15606);
or U15715 (N_15715,N_15642,N_15637);
and U15716 (N_15716,N_15552,N_15639);
nor U15717 (N_15717,N_15634,N_15673);
nand U15718 (N_15718,N_15548,N_15607);
and U15719 (N_15719,N_15558,N_15533);
nand U15720 (N_15720,N_15583,N_15527);
and U15721 (N_15721,N_15571,N_15521);
xor U15722 (N_15722,N_15589,N_15650);
xor U15723 (N_15723,N_15594,N_15555);
nor U15724 (N_15724,N_15574,N_15644);
and U15725 (N_15725,N_15674,N_15553);
nand U15726 (N_15726,N_15567,N_15542);
or U15727 (N_15727,N_15551,N_15643);
nand U15728 (N_15728,N_15547,N_15655);
xor U15729 (N_15729,N_15671,N_15581);
nand U15730 (N_15730,N_15557,N_15620);
nor U15731 (N_15731,N_15622,N_15630);
nand U15732 (N_15732,N_15537,N_15568);
and U15733 (N_15733,N_15615,N_15543);
nor U15734 (N_15734,N_15679,N_15550);
xor U15735 (N_15735,N_15677,N_15520);
or U15736 (N_15736,N_15593,N_15596);
or U15737 (N_15737,N_15667,N_15605);
xnor U15738 (N_15738,N_15546,N_15549);
or U15739 (N_15739,N_15576,N_15563);
xor U15740 (N_15740,N_15541,N_15675);
and U15741 (N_15741,N_15524,N_15535);
xor U15742 (N_15742,N_15560,N_15613);
nor U15743 (N_15743,N_15528,N_15564);
or U15744 (N_15744,N_15654,N_15582);
nor U15745 (N_15745,N_15658,N_15623);
and U15746 (N_15746,N_15584,N_15526);
or U15747 (N_15747,N_15651,N_15665);
and U15748 (N_15748,N_15595,N_15588);
and U15749 (N_15749,N_15628,N_15656);
nand U15750 (N_15750,N_15668,N_15554);
and U15751 (N_15751,N_15666,N_15638);
nor U15752 (N_15752,N_15530,N_15618);
nor U15753 (N_15753,N_15532,N_15534);
nor U15754 (N_15754,N_15636,N_15577);
and U15755 (N_15755,N_15649,N_15670);
nor U15756 (N_15756,N_15676,N_15631);
or U15757 (N_15757,N_15664,N_15578);
and U15758 (N_15758,N_15559,N_15600);
nand U15759 (N_15759,N_15629,N_15610);
xnor U15760 (N_15760,N_15564,N_15672);
nand U15761 (N_15761,N_15537,N_15625);
xor U15762 (N_15762,N_15637,N_15524);
nand U15763 (N_15763,N_15587,N_15606);
or U15764 (N_15764,N_15658,N_15589);
xor U15765 (N_15765,N_15569,N_15524);
nand U15766 (N_15766,N_15541,N_15645);
nand U15767 (N_15767,N_15672,N_15664);
nand U15768 (N_15768,N_15589,N_15601);
nor U15769 (N_15769,N_15575,N_15638);
or U15770 (N_15770,N_15571,N_15639);
nand U15771 (N_15771,N_15579,N_15619);
or U15772 (N_15772,N_15638,N_15546);
nor U15773 (N_15773,N_15644,N_15537);
nor U15774 (N_15774,N_15593,N_15660);
or U15775 (N_15775,N_15602,N_15567);
nand U15776 (N_15776,N_15660,N_15588);
or U15777 (N_15777,N_15569,N_15530);
nand U15778 (N_15778,N_15599,N_15528);
and U15779 (N_15779,N_15562,N_15651);
or U15780 (N_15780,N_15605,N_15581);
nand U15781 (N_15781,N_15614,N_15576);
nor U15782 (N_15782,N_15638,N_15528);
or U15783 (N_15783,N_15554,N_15535);
xor U15784 (N_15784,N_15653,N_15546);
or U15785 (N_15785,N_15584,N_15547);
and U15786 (N_15786,N_15575,N_15533);
or U15787 (N_15787,N_15540,N_15523);
or U15788 (N_15788,N_15586,N_15532);
xnor U15789 (N_15789,N_15550,N_15528);
nand U15790 (N_15790,N_15666,N_15560);
or U15791 (N_15791,N_15578,N_15537);
nand U15792 (N_15792,N_15610,N_15521);
or U15793 (N_15793,N_15594,N_15608);
or U15794 (N_15794,N_15526,N_15656);
nor U15795 (N_15795,N_15527,N_15565);
or U15796 (N_15796,N_15594,N_15601);
xnor U15797 (N_15797,N_15641,N_15573);
nor U15798 (N_15798,N_15678,N_15594);
and U15799 (N_15799,N_15595,N_15622);
nand U15800 (N_15800,N_15571,N_15592);
or U15801 (N_15801,N_15606,N_15621);
or U15802 (N_15802,N_15577,N_15606);
and U15803 (N_15803,N_15678,N_15541);
nand U15804 (N_15804,N_15522,N_15675);
nand U15805 (N_15805,N_15557,N_15532);
or U15806 (N_15806,N_15549,N_15593);
nand U15807 (N_15807,N_15556,N_15596);
xnor U15808 (N_15808,N_15568,N_15604);
and U15809 (N_15809,N_15555,N_15565);
nor U15810 (N_15810,N_15564,N_15545);
or U15811 (N_15811,N_15628,N_15590);
nor U15812 (N_15812,N_15645,N_15589);
or U15813 (N_15813,N_15630,N_15592);
and U15814 (N_15814,N_15641,N_15577);
and U15815 (N_15815,N_15563,N_15679);
or U15816 (N_15816,N_15607,N_15577);
nor U15817 (N_15817,N_15621,N_15639);
and U15818 (N_15818,N_15628,N_15556);
nand U15819 (N_15819,N_15644,N_15552);
nor U15820 (N_15820,N_15671,N_15578);
nor U15821 (N_15821,N_15666,N_15544);
nand U15822 (N_15822,N_15578,N_15539);
nor U15823 (N_15823,N_15521,N_15625);
nor U15824 (N_15824,N_15653,N_15647);
and U15825 (N_15825,N_15562,N_15567);
and U15826 (N_15826,N_15670,N_15658);
or U15827 (N_15827,N_15532,N_15533);
or U15828 (N_15828,N_15679,N_15636);
nor U15829 (N_15829,N_15602,N_15612);
nand U15830 (N_15830,N_15628,N_15521);
and U15831 (N_15831,N_15553,N_15602);
or U15832 (N_15832,N_15561,N_15676);
nor U15833 (N_15833,N_15609,N_15624);
and U15834 (N_15834,N_15562,N_15630);
or U15835 (N_15835,N_15591,N_15570);
nor U15836 (N_15836,N_15651,N_15568);
and U15837 (N_15837,N_15678,N_15521);
nand U15838 (N_15838,N_15550,N_15603);
or U15839 (N_15839,N_15549,N_15671);
nand U15840 (N_15840,N_15705,N_15762);
xor U15841 (N_15841,N_15813,N_15795);
and U15842 (N_15842,N_15799,N_15839);
and U15843 (N_15843,N_15684,N_15786);
nand U15844 (N_15844,N_15708,N_15713);
and U15845 (N_15845,N_15814,N_15732);
or U15846 (N_15846,N_15822,N_15827);
nor U15847 (N_15847,N_15737,N_15817);
or U15848 (N_15848,N_15826,N_15836);
nor U15849 (N_15849,N_15793,N_15735);
nand U15850 (N_15850,N_15729,N_15719);
and U15851 (N_15851,N_15750,N_15728);
or U15852 (N_15852,N_15821,N_15801);
nand U15853 (N_15853,N_15781,N_15830);
or U15854 (N_15854,N_15716,N_15797);
and U15855 (N_15855,N_15753,N_15774);
nand U15856 (N_15856,N_15697,N_15760);
nand U15857 (N_15857,N_15761,N_15816);
nor U15858 (N_15858,N_15711,N_15806);
nor U15859 (N_15859,N_15752,N_15741);
and U15860 (N_15860,N_15833,N_15775);
nor U15861 (N_15861,N_15740,N_15754);
or U15862 (N_15862,N_15743,N_15755);
and U15863 (N_15863,N_15688,N_15773);
xnor U15864 (N_15864,N_15691,N_15784);
xor U15865 (N_15865,N_15772,N_15710);
xor U15866 (N_15866,N_15718,N_15748);
and U15867 (N_15867,N_15702,N_15776);
nand U15868 (N_15868,N_15681,N_15824);
and U15869 (N_15869,N_15837,N_15777);
nor U15870 (N_15870,N_15690,N_15689);
nand U15871 (N_15871,N_15739,N_15707);
nor U15872 (N_15872,N_15742,N_15693);
or U15873 (N_15873,N_15831,N_15721);
xnor U15874 (N_15874,N_15763,N_15696);
or U15875 (N_15875,N_15727,N_15828);
nor U15876 (N_15876,N_15787,N_15745);
and U15877 (N_15877,N_15800,N_15723);
nand U15878 (N_15878,N_15744,N_15794);
and U15879 (N_15879,N_15686,N_15766);
nand U15880 (N_15880,N_15714,N_15695);
xnor U15881 (N_15881,N_15717,N_15796);
nor U15882 (N_15882,N_15730,N_15791);
xnor U15883 (N_15883,N_15804,N_15764);
nor U15884 (N_15884,N_15738,N_15699);
or U15885 (N_15885,N_15692,N_15835);
or U15886 (N_15886,N_15768,N_15724);
or U15887 (N_15887,N_15683,N_15703);
nand U15888 (N_15888,N_15782,N_15734);
and U15889 (N_15889,N_15685,N_15789);
nor U15890 (N_15890,N_15798,N_15694);
nand U15891 (N_15891,N_15747,N_15709);
or U15892 (N_15892,N_15811,N_15785);
and U15893 (N_15893,N_15812,N_15759);
nor U15894 (N_15894,N_15725,N_15825);
and U15895 (N_15895,N_15832,N_15819);
or U15896 (N_15896,N_15720,N_15682);
or U15897 (N_15897,N_15749,N_15770);
or U15898 (N_15898,N_15790,N_15783);
nand U15899 (N_15899,N_15736,N_15767);
nor U15900 (N_15900,N_15731,N_15704);
nor U15901 (N_15901,N_15805,N_15829);
xor U15902 (N_15902,N_15765,N_15838);
or U15903 (N_15903,N_15815,N_15698);
nand U15904 (N_15904,N_15808,N_15779);
nor U15905 (N_15905,N_15700,N_15809);
and U15906 (N_15906,N_15756,N_15803);
nor U15907 (N_15907,N_15820,N_15778);
or U15908 (N_15908,N_15722,N_15758);
nor U15909 (N_15909,N_15701,N_15733);
or U15910 (N_15910,N_15769,N_15810);
and U15911 (N_15911,N_15680,N_15802);
nand U15912 (N_15912,N_15726,N_15757);
nand U15913 (N_15913,N_15771,N_15706);
or U15914 (N_15914,N_15746,N_15807);
nand U15915 (N_15915,N_15687,N_15751);
nand U15916 (N_15916,N_15823,N_15792);
nor U15917 (N_15917,N_15780,N_15788);
or U15918 (N_15918,N_15818,N_15834);
xor U15919 (N_15919,N_15715,N_15712);
nor U15920 (N_15920,N_15768,N_15831);
nand U15921 (N_15921,N_15796,N_15794);
xor U15922 (N_15922,N_15837,N_15731);
nand U15923 (N_15923,N_15801,N_15771);
nor U15924 (N_15924,N_15752,N_15734);
nor U15925 (N_15925,N_15759,N_15682);
or U15926 (N_15926,N_15707,N_15728);
nor U15927 (N_15927,N_15739,N_15736);
nor U15928 (N_15928,N_15688,N_15771);
or U15929 (N_15929,N_15699,N_15833);
and U15930 (N_15930,N_15799,N_15736);
nor U15931 (N_15931,N_15682,N_15767);
nor U15932 (N_15932,N_15812,N_15713);
nor U15933 (N_15933,N_15727,N_15710);
nand U15934 (N_15934,N_15696,N_15764);
nand U15935 (N_15935,N_15784,N_15778);
nand U15936 (N_15936,N_15680,N_15828);
nor U15937 (N_15937,N_15695,N_15745);
and U15938 (N_15938,N_15737,N_15725);
and U15939 (N_15939,N_15760,N_15762);
or U15940 (N_15940,N_15826,N_15685);
nor U15941 (N_15941,N_15716,N_15807);
nor U15942 (N_15942,N_15705,N_15697);
or U15943 (N_15943,N_15819,N_15797);
nor U15944 (N_15944,N_15803,N_15693);
nand U15945 (N_15945,N_15830,N_15695);
and U15946 (N_15946,N_15733,N_15763);
and U15947 (N_15947,N_15837,N_15793);
or U15948 (N_15948,N_15705,N_15803);
or U15949 (N_15949,N_15838,N_15740);
or U15950 (N_15950,N_15753,N_15785);
or U15951 (N_15951,N_15839,N_15762);
and U15952 (N_15952,N_15805,N_15837);
or U15953 (N_15953,N_15794,N_15816);
and U15954 (N_15954,N_15772,N_15721);
and U15955 (N_15955,N_15769,N_15795);
nand U15956 (N_15956,N_15691,N_15797);
nand U15957 (N_15957,N_15730,N_15703);
nor U15958 (N_15958,N_15817,N_15830);
or U15959 (N_15959,N_15839,N_15703);
nor U15960 (N_15960,N_15705,N_15773);
or U15961 (N_15961,N_15786,N_15694);
xnor U15962 (N_15962,N_15688,N_15762);
or U15963 (N_15963,N_15816,N_15817);
nor U15964 (N_15964,N_15772,N_15737);
nor U15965 (N_15965,N_15704,N_15790);
or U15966 (N_15966,N_15692,N_15697);
or U15967 (N_15967,N_15696,N_15780);
and U15968 (N_15968,N_15760,N_15714);
or U15969 (N_15969,N_15741,N_15682);
nor U15970 (N_15970,N_15816,N_15745);
or U15971 (N_15971,N_15784,N_15726);
nand U15972 (N_15972,N_15815,N_15689);
nand U15973 (N_15973,N_15835,N_15682);
and U15974 (N_15974,N_15726,N_15747);
nand U15975 (N_15975,N_15804,N_15800);
nor U15976 (N_15976,N_15813,N_15784);
nand U15977 (N_15977,N_15716,N_15766);
nand U15978 (N_15978,N_15795,N_15784);
nand U15979 (N_15979,N_15714,N_15715);
xor U15980 (N_15980,N_15775,N_15683);
and U15981 (N_15981,N_15704,N_15764);
and U15982 (N_15982,N_15793,N_15792);
and U15983 (N_15983,N_15760,N_15758);
xor U15984 (N_15984,N_15826,N_15749);
and U15985 (N_15985,N_15722,N_15705);
nor U15986 (N_15986,N_15752,N_15832);
nand U15987 (N_15987,N_15699,N_15753);
nor U15988 (N_15988,N_15697,N_15704);
or U15989 (N_15989,N_15799,N_15722);
or U15990 (N_15990,N_15694,N_15791);
xnor U15991 (N_15991,N_15758,N_15790);
xnor U15992 (N_15992,N_15702,N_15685);
and U15993 (N_15993,N_15729,N_15698);
nor U15994 (N_15994,N_15806,N_15828);
and U15995 (N_15995,N_15809,N_15748);
nand U15996 (N_15996,N_15753,N_15728);
or U15997 (N_15997,N_15811,N_15690);
or U15998 (N_15998,N_15837,N_15830);
or U15999 (N_15999,N_15745,N_15741);
and U16000 (N_16000,N_15994,N_15891);
nor U16001 (N_16001,N_15974,N_15884);
or U16002 (N_16002,N_15933,N_15943);
or U16003 (N_16003,N_15944,N_15968);
nor U16004 (N_16004,N_15865,N_15907);
nand U16005 (N_16005,N_15980,N_15864);
xor U16006 (N_16006,N_15956,N_15961);
or U16007 (N_16007,N_15924,N_15991);
nor U16008 (N_16008,N_15958,N_15881);
or U16009 (N_16009,N_15918,N_15925);
nor U16010 (N_16010,N_15928,N_15885);
nand U16011 (N_16011,N_15841,N_15901);
or U16012 (N_16012,N_15967,N_15935);
or U16013 (N_16013,N_15983,N_15923);
and U16014 (N_16014,N_15982,N_15846);
and U16015 (N_16015,N_15979,N_15986);
nand U16016 (N_16016,N_15963,N_15894);
nand U16017 (N_16017,N_15888,N_15949);
nor U16018 (N_16018,N_15992,N_15987);
nand U16019 (N_16019,N_15904,N_15849);
nand U16020 (N_16020,N_15851,N_15882);
xor U16021 (N_16021,N_15927,N_15939);
nor U16022 (N_16022,N_15984,N_15930);
or U16023 (N_16023,N_15970,N_15937);
nand U16024 (N_16024,N_15916,N_15975);
or U16025 (N_16025,N_15879,N_15945);
xnor U16026 (N_16026,N_15899,N_15951);
or U16027 (N_16027,N_15912,N_15840);
nor U16028 (N_16028,N_15997,N_15900);
nand U16029 (N_16029,N_15856,N_15981);
nand U16030 (N_16030,N_15914,N_15898);
or U16031 (N_16031,N_15957,N_15875);
nand U16032 (N_16032,N_15929,N_15932);
or U16033 (N_16033,N_15852,N_15878);
or U16034 (N_16034,N_15964,N_15947);
and U16035 (N_16035,N_15938,N_15863);
and U16036 (N_16036,N_15883,N_15965);
nor U16037 (N_16037,N_15880,N_15859);
xnor U16038 (N_16038,N_15969,N_15936);
nor U16039 (N_16039,N_15843,N_15940);
nand U16040 (N_16040,N_15948,N_15893);
nor U16041 (N_16041,N_15911,N_15960);
nor U16042 (N_16042,N_15931,N_15996);
nor U16043 (N_16043,N_15871,N_15934);
xor U16044 (N_16044,N_15972,N_15946);
nand U16045 (N_16045,N_15860,N_15917);
or U16046 (N_16046,N_15853,N_15913);
xnor U16047 (N_16047,N_15942,N_15877);
and U16048 (N_16048,N_15941,N_15897);
nor U16049 (N_16049,N_15874,N_15887);
and U16050 (N_16050,N_15858,N_15903);
nor U16051 (N_16051,N_15902,N_15985);
nand U16052 (N_16052,N_15890,N_15872);
and U16053 (N_16053,N_15869,N_15868);
and U16054 (N_16054,N_15976,N_15862);
and U16055 (N_16055,N_15962,N_15906);
and U16056 (N_16056,N_15988,N_15850);
xor U16057 (N_16057,N_15966,N_15895);
or U16058 (N_16058,N_15861,N_15995);
xnor U16059 (N_16059,N_15848,N_15855);
and U16060 (N_16060,N_15892,N_15919);
nand U16061 (N_16061,N_15978,N_15908);
nand U16062 (N_16062,N_15870,N_15905);
nand U16063 (N_16063,N_15909,N_15873);
xor U16064 (N_16064,N_15866,N_15977);
nand U16065 (N_16065,N_15845,N_15886);
and U16066 (N_16066,N_15959,N_15954);
nor U16067 (N_16067,N_15973,N_15998);
or U16068 (N_16068,N_15953,N_15922);
and U16069 (N_16069,N_15842,N_15990);
nor U16070 (N_16070,N_15889,N_15876);
or U16071 (N_16071,N_15854,N_15971);
xor U16072 (N_16072,N_15857,N_15847);
nand U16073 (N_16073,N_15999,N_15915);
and U16074 (N_16074,N_15955,N_15993);
nand U16075 (N_16075,N_15926,N_15989);
nor U16076 (N_16076,N_15950,N_15896);
xor U16077 (N_16077,N_15910,N_15867);
nand U16078 (N_16078,N_15921,N_15844);
nor U16079 (N_16079,N_15920,N_15952);
nor U16080 (N_16080,N_15893,N_15993);
or U16081 (N_16081,N_15948,N_15864);
and U16082 (N_16082,N_15974,N_15998);
and U16083 (N_16083,N_15928,N_15910);
xor U16084 (N_16084,N_15985,N_15981);
and U16085 (N_16085,N_15902,N_15919);
and U16086 (N_16086,N_15926,N_15941);
and U16087 (N_16087,N_15857,N_15871);
nor U16088 (N_16088,N_15895,N_15925);
nor U16089 (N_16089,N_15863,N_15843);
xnor U16090 (N_16090,N_15868,N_15845);
nand U16091 (N_16091,N_15853,N_15942);
nor U16092 (N_16092,N_15845,N_15975);
nand U16093 (N_16093,N_15872,N_15841);
nand U16094 (N_16094,N_15911,N_15897);
or U16095 (N_16095,N_15877,N_15999);
nand U16096 (N_16096,N_15864,N_15876);
and U16097 (N_16097,N_15847,N_15985);
and U16098 (N_16098,N_15942,N_15963);
nor U16099 (N_16099,N_15970,N_15913);
or U16100 (N_16100,N_15850,N_15915);
nor U16101 (N_16101,N_15940,N_15939);
and U16102 (N_16102,N_15905,N_15853);
xor U16103 (N_16103,N_15995,N_15955);
nor U16104 (N_16104,N_15861,N_15878);
nor U16105 (N_16105,N_15983,N_15921);
xor U16106 (N_16106,N_15938,N_15998);
or U16107 (N_16107,N_15906,N_15961);
nand U16108 (N_16108,N_15893,N_15979);
and U16109 (N_16109,N_15934,N_15982);
nand U16110 (N_16110,N_15886,N_15855);
and U16111 (N_16111,N_15946,N_15957);
or U16112 (N_16112,N_15971,N_15881);
and U16113 (N_16113,N_15949,N_15891);
nand U16114 (N_16114,N_15873,N_15901);
and U16115 (N_16115,N_15905,N_15910);
nor U16116 (N_16116,N_15875,N_15984);
nor U16117 (N_16117,N_15961,N_15895);
nand U16118 (N_16118,N_15967,N_15862);
nor U16119 (N_16119,N_15921,N_15966);
or U16120 (N_16120,N_15963,N_15997);
nand U16121 (N_16121,N_15875,N_15987);
or U16122 (N_16122,N_15870,N_15943);
nand U16123 (N_16123,N_15917,N_15899);
nor U16124 (N_16124,N_15960,N_15865);
xnor U16125 (N_16125,N_15908,N_15867);
nand U16126 (N_16126,N_15863,N_15928);
xnor U16127 (N_16127,N_15997,N_15898);
or U16128 (N_16128,N_15987,N_15994);
or U16129 (N_16129,N_15864,N_15853);
or U16130 (N_16130,N_15929,N_15930);
and U16131 (N_16131,N_15874,N_15897);
or U16132 (N_16132,N_15883,N_15850);
nor U16133 (N_16133,N_15994,N_15940);
or U16134 (N_16134,N_15852,N_15972);
or U16135 (N_16135,N_15852,N_15922);
xnor U16136 (N_16136,N_15963,N_15961);
nand U16137 (N_16137,N_15947,N_15987);
or U16138 (N_16138,N_15931,N_15874);
xor U16139 (N_16139,N_15873,N_15896);
and U16140 (N_16140,N_15944,N_15953);
or U16141 (N_16141,N_15995,N_15922);
nor U16142 (N_16142,N_15978,N_15884);
or U16143 (N_16143,N_15989,N_15999);
xor U16144 (N_16144,N_15871,N_15906);
nand U16145 (N_16145,N_15928,N_15950);
xor U16146 (N_16146,N_15857,N_15936);
xnor U16147 (N_16147,N_15955,N_15944);
and U16148 (N_16148,N_15990,N_15939);
and U16149 (N_16149,N_15919,N_15967);
xor U16150 (N_16150,N_15911,N_15928);
or U16151 (N_16151,N_15972,N_15954);
xor U16152 (N_16152,N_15860,N_15878);
xnor U16153 (N_16153,N_15949,N_15845);
or U16154 (N_16154,N_15983,N_15859);
and U16155 (N_16155,N_15847,N_15912);
nor U16156 (N_16156,N_15882,N_15966);
nor U16157 (N_16157,N_15961,N_15994);
xnor U16158 (N_16158,N_15922,N_15923);
nor U16159 (N_16159,N_15902,N_15888);
xor U16160 (N_16160,N_16031,N_16156);
xnor U16161 (N_16161,N_16056,N_16116);
nor U16162 (N_16162,N_16118,N_16067);
or U16163 (N_16163,N_16136,N_16090);
xnor U16164 (N_16164,N_16150,N_16131);
xnor U16165 (N_16165,N_16024,N_16078);
nor U16166 (N_16166,N_16140,N_16020);
nor U16167 (N_16167,N_16127,N_16138);
and U16168 (N_16168,N_16085,N_16076);
nor U16169 (N_16169,N_16135,N_16004);
and U16170 (N_16170,N_16007,N_16089);
xor U16171 (N_16171,N_16117,N_16110);
nor U16172 (N_16172,N_16036,N_16055);
xor U16173 (N_16173,N_16032,N_16010);
and U16174 (N_16174,N_16096,N_16021);
or U16175 (N_16175,N_16072,N_16148);
or U16176 (N_16176,N_16122,N_16120);
nor U16177 (N_16177,N_16023,N_16083);
and U16178 (N_16178,N_16026,N_16153);
or U16179 (N_16179,N_16124,N_16054);
or U16180 (N_16180,N_16144,N_16149);
nand U16181 (N_16181,N_16104,N_16079);
nor U16182 (N_16182,N_16129,N_16048);
and U16183 (N_16183,N_16147,N_16111);
xnor U16184 (N_16184,N_16015,N_16014);
xor U16185 (N_16185,N_16029,N_16134);
or U16186 (N_16186,N_16109,N_16086);
and U16187 (N_16187,N_16001,N_16106);
xor U16188 (N_16188,N_16042,N_16017);
xor U16189 (N_16189,N_16061,N_16057);
nor U16190 (N_16190,N_16082,N_16145);
nor U16191 (N_16191,N_16098,N_16088);
nand U16192 (N_16192,N_16094,N_16113);
or U16193 (N_16193,N_16070,N_16003);
nand U16194 (N_16194,N_16151,N_16022);
or U16195 (N_16195,N_16158,N_16073);
nor U16196 (N_16196,N_16006,N_16033);
or U16197 (N_16197,N_16099,N_16039);
nor U16198 (N_16198,N_16027,N_16050);
and U16199 (N_16199,N_16066,N_16077);
xnor U16200 (N_16200,N_16005,N_16051);
nor U16201 (N_16201,N_16108,N_16125);
or U16202 (N_16202,N_16016,N_16084);
or U16203 (N_16203,N_16097,N_16081);
nand U16204 (N_16204,N_16064,N_16040);
nand U16205 (N_16205,N_16000,N_16107);
nand U16206 (N_16206,N_16009,N_16154);
nand U16207 (N_16207,N_16071,N_16063);
or U16208 (N_16208,N_16047,N_16102);
or U16209 (N_16209,N_16019,N_16065);
or U16210 (N_16210,N_16159,N_16105);
or U16211 (N_16211,N_16041,N_16052);
nor U16212 (N_16212,N_16152,N_16049);
and U16213 (N_16213,N_16062,N_16037);
nor U16214 (N_16214,N_16139,N_16074);
or U16215 (N_16215,N_16087,N_16128);
and U16216 (N_16216,N_16034,N_16095);
or U16217 (N_16217,N_16011,N_16112);
or U16218 (N_16218,N_16101,N_16146);
nand U16219 (N_16219,N_16038,N_16114);
nor U16220 (N_16220,N_16093,N_16028);
nor U16221 (N_16221,N_16103,N_16013);
or U16222 (N_16222,N_16126,N_16045);
nand U16223 (N_16223,N_16141,N_16143);
and U16224 (N_16224,N_16018,N_16068);
and U16225 (N_16225,N_16157,N_16142);
nand U16226 (N_16226,N_16008,N_16043);
or U16227 (N_16227,N_16092,N_16058);
nor U16228 (N_16228,N_16121,N_16133);
and U16229 (N_16229,N_16123,N_16080);
nor U16230 (N_16230,N_16002,N_16030);
or U16231 (N_16231,N_16044,N_16059);
nand U16232 (N_16232,N_16075,N_16137);
nor U16233 (N_16233,N_16025,N_16132);
or U16234 (N_16234,N_16069,N_16053);
nor U16235 (N_16235,N_16046,N_16155);
or U16236 (N_16236,N_16130,N_16035);
xor U16237 (N_16237,N_16060,N_16091);
nand U16238 (N_16238,N_16100,N_16012);
or U16239 (N_16239,N_16115,N_16119);
or U16240 (N_16240,N_16009,N_16116);
or U16241 (N_16241,N_16088,N_16027);
and U16242 (N_16242,N_16019,N_16017);
or U16243 (N_16243,N_16002,N_16140);
and U16244 (N_16244,N_16039,N_16097);
and U16245 (N_16245,N_16154,N_16019);
nor U16246 (N_16246,N_16101,N_16130);
or U16247 (N_16247,N_16112,N_16088);
and U16248 (N_16248,N_16050,N_16066);
and U16249 (N_16249,N_16047,N_16130);
nand U16250 (N_16250,N_16086,N_16049);
or U16251 (N_16251,N_16004,N_16069);
nor U16252 (N_16252,N_16117,N_16025);
xnor U16253 (N_16253,N_16100,N_16056);
nand U16254 (N_16254,N_16058,N_16043);
nor U16255 (N_16255,N_16056,N_16079);
nor U16256 (N_16256,N_16010,N_16140);
nor U16257 (N_16257,N_16041,N_16104);
or U16258 (N_16258,N_16158,N_16021);
or U16259 (N_16259,N_16036,N_16085);
and U16260 (N_16260,N_16008,N_16010);
xnor U16261 (N_16261,N_16150,N_16106);
or U16262 (N_16262,N_16058,N_16085);
xnor U16263 (N_16263,N_16086,N_16021);
nand U16264 (N_16264,N_16027,N_16152);
or U16265 (N_16265,N_16074,N_16147);
nor U16266 (N_16266,N_16028,N_16125);
or U16267 (N_16267,N_16101,N_16002);
nand U16268 (N_16268,N_16001,N_16073);
and U16269 (N_16269,N_16062,N_16019);
or U16270 (N_16270,N_16106,N_16121);
nor U16271 (N_16271,N_16150,N_16076);
nor U16272 (N_16272,N_16059,N_16054);
or U16273 (N_16273,N_16031,N_16119);
nor U16274 (N_16274,N_16105,N_16129);
and U16275 (N_16275,N_16100,N_16047);
and U16276 (N_16276,N_16093,N_16035);
nor U16277 (N_16277,N_16077,N_16138);
nand U16278 (N_16278,N_16039,N_16142);
and U16279 (N_16279,N_16100,N_16105);
nor U16280 (N_16280,N_16024,N_16117);
and U16281 (N_16281,N_16031,N_16093);
and U16282 (N_16282,N_16125,N_16029);
nand U16283 (N_16283,N_16045,N_16124);
nor U16284 (N_16284,N_16021,N_16055);
and U16285 (N_16285,N_16149,N_16135);
and U16286 (N_16286,N_16116,N_16052);
nor U16287 (N_16287,N_16078,N_16080);
or U16288 (N_16288,N_16054,N_16073);
nand U16289 (N_16289,N_16114,N_16108);
or U16290 (N_16290,N_16030,N_16067);
and U16291 (N_16291,N_16035,N_16041);
and U16292 (N_16292,N_16068,N_16029);
nand U16293 (N_16293,N_16136,N_16055);
xnor U16294 (N_16294,N_16023,N_16097);
nor U16295 (N_16295,N_16078,N_16097);
and U16296 (N_16296,N_16009,N_16043);
or U16297 (N_16297,N_16098,N_16008);
xnor U16298 (N_16298,N_16148,N_16145);
nor U16299 (N_16299,N_16151,N_16130);
nand U16300 (N_16300,N_16052,N_16077);
and U16301 (N_16301,N_16151,N_16066);
xor U16302 (N_16302,N_16094,N_16103);
or U16303 (N_16303,N_16063,N_16043);
or U16304 (N_16304,N_16113,N_16006);
nand U16305 (N_16305,N_16109,N_16084);
nor U16306 (N_16306,N_16077,N_16071);
and U16307 (N_16307,N_16135,N_16013);
nand U16308 (N_16308,N_16017,N_16026);
nor U16309 (N_16309,N_16092,N_16114);
nand U16310 (N_16310,N_16105,N_16022);
and U16311 (N_16311,N_16041,N_16157);
xor U16312 (N_16312,N_16035,N_16148);
xnor U16313 (N_16313,N_16070,N_16044);
nand U16314 (N_16314,N_16089,N_16111);
or U16315 (N_16315,N_16071,N_16093);
nor U16316 (N_16316,N_16020,N_16036);
and U16317 (N_16317,N_16027,N_16091);
and U16318 (N_16318,N_16097,N_16004);
nor U16319 (N_16319,N_16043,N_16011);
and U16320 (N_16320,N_16310,N_16245);
and U16321 (N_16321,N_16193,N_16185);
and U16322 (N_16322,N_16229,N_16212);
nor U16323 (N_16323,N_16241,N_16225);
nor U16324 (N_16324,N_16163,N_16300);
and U16325 (N_16325,N_16227,N_16248);
nor U16326 (N_16326,N_16306,N_16194);
or U16327 (N_16327,N_16219,N_16224);
nand U16328 (N_16328,N_16258,N_16287);
and U16329 (N_16329,N_16246,N_16221);
xor U16330 (N_16330,N_16308,N_16206);
or U16331 (N_16331,N_16284,N_16292);
and U16332 (N_16332,N_16257,N_16214);
nor U16333 (N_16333,N_16278,N_16189);
nand U16334 (N_16334,N_16176,N_16238);
nand U16335 (N_16335,N_16199,N_16253);
or U16336 (N_16336,N_16209,N_16303);
nand U16337 (N_16337,N_16311,N_16205);
nor U16338 (N_16338,N_16228,N_16313);
nand U16339 (N_16339,N_16309,N_16234);
nor U16340 (N_16340,N_16236,N_16235);
and U16341 (N_16341,N_16289,N_16290);
or U16342 (N_16342,N_16315,N_16262);
nand U16343 (N_16343,N_16216,N_16307);
nor U16344 (N_16344,N_16318,N_16218);
and U16345 (N_16345,N_16291,N_16252);
nor U16346 (N_16346,N_16197,N_16312);
nand U16347 (N_16347,N_16317,N_16196);
and U16348 (N_16348,N_16222,N_16179);
nand U16349 (N_16349,N_16200,N_16204);
and U16350 (N_16350,N_16302,N_16255);
nor U16351 (N_16351,N_16170,N_16319);
and U16352 (N_16352,N_16295,N_16277);
nand U16353 (N_16353,N_16191,N_16180);
nor U16354 (N_16354,N_16296,N_16161);
xor U16355 (N_16355,N_16215,N_16243);
nor U16356 (N_16356,N_16169,N_16210);
nor U16357 (N_16357,N_16165,N_16249);
xor U16358 (N_16358,N_16247,N_16174);
or U16359 (N_16359,N_16175,N_16226);
nor U16360 (N_16360,N_16260,N_16251);
nor U16361 (N_16361,N_16263,N_16183);
nand U16362 (N_16362,N_16301,N_16181);
and U16363 (N_16363,N_16250,N_16265);
or U16364 (N_16364,N_16294,N_16207);
xnor U16365 (N_16365,N_16195,N_16232);
xnor U16366 (N_16366,N_16259,N_16242);
and U16367 (N_16367,N_16217,N_16266);
nand U16368 (N_16368,N_16173,N_16283);
nor U16369 (N_16369,N_16187,N_16280);
or U16370 (N_16370,N_16167,N_16293);
and U16371 (N_16371,N_16288,N_16201);
and U16372 (N_16372,N_16244,N_16186);
nor U16373 (N_16373,N_16168,N_16192);
nor U16374 (N_16374,N_16268,N_16281);
and U16375 (N_16375,N_16177,N_16254);
nor U16376 (N_16376,N_16272,N_16286);
or U16377 (N_16377,N_16298,N_16267);
nand U16378 (N_16378,N_16273,N_16198);
and U16379 (N_16379,N_16237,N_16160);
nand U16380 (N_16380,N_16213,N_16240);
and U16381 (N_16381,N_16271,N_16279);
and U16382 (N_16382,N_16256,N_16233);
nand U16383 (N_16383,N_16202,N_16172);
nand U16384 (N_16384,N_16230,N_16269);
nand U16385 (N_16385,N_16316,N_16261);
nand U16386 (N_16386,N_16239,N_16231);
and U16387 (N_16387,N_16285,N_16264);
or U16388 (N_16388,N_16276,N_16282);
nand U16389 (N_16389,N_16162,N_16275);
xnor U16390 (N_16390,N_16208,N_16274);
nand U16391 (N_16391,N_16171,N_16297);
or U16392 (N_16392,N_16314,N_16184);
nor U16393 (N_16393,N_16203,N_16220);
nor U16394 (N_16394,N_16299,N_16178);
nor U16395 (N_16395,N_16164,N_16305);
or U16396 (N_16396,N_16304,N_16182);
nand U16397 (N_16397,N_16223,N_16190);
and U16398 (N_16398,N_16270,N_16188);
and U16399 (N_16399,N_16211,N_16166);
nor U16400 (N_16400,N_16305,N_16285);
or U16401 (N_16401,N_16213,N_16279);
or U16402 (N_16402,N_16266,N_16219);
nand U16403 (N_16403,N_16248,N_16234);
nor U16404 (N_16404,N_16160,N_16180);
nand U16405 (N_16405,N_16290,N_16176);
or U16406 (N_16406,N_16282,N_16296);
nor U16407 (N_16407,N_16318,N_16186);
and U16408 (N_16408,N_16188,N_16195);
nand U16409 (N_16409,N_16208,N_16185);
and U16410 (N_16410,N_16259,N_16196);
nand U16411 (N_16411,N_16230,N_16253);
or U16412 (N_16412,N_16257,N_16280);
xor U16413 (N_16413,N_16254,N_16193);
or U16414 (N_16414,N_16304,N_16195);
nand U16415 (N_16415,N_16238,N_16297);
nor U16416 (N_16416,N_16206,N_16306);
and U16417 (N_16417,N_16208,N_16160);
and U16418 (N_16418,N_16257,N_16255);
nor U16419 (N_16419,N_16182,N_16277);
or U16420 (N_16420,N_16201,N_16174);
nor U16421 (N_16421,N_16218,N_16315);
and U16422 (N_16422,N_16241,N_16221);
nand U16423 (N_16423,N_16269,N_16243);
nand U16424 (N_16424,N_16197,N_16228);
nand U16425 (N_16425,N_16318,N_16263);
nor U16426 (N_16426,N_16265,N_16200);
and U16427 (N_16427,N_16319,N_16233);
and U16428 (N_16428,N_16280,N_16182);
and U16429 (N_16429,N_16170,N_16257);
or U16430 (N_16430,N_16222,N_16209);
and U16431 (N_16431,N_16312,N_16238);
or U16432 (N_16432,N_16277,N_16275);
xor U16433 (N_16433,N_16246,N_16258);
or U16434 (N_16434,N_16176,N_16222);
or U16435 (N_16435,N_16292,N_16290);
nor U16436 (N_16436,N_16171,N_16314);
xor U16437 (N_16437,N_16162,N_16265);
nand U16438 (N_16438,N_16245,N_16281);
nor U16439 (N_16439,N_16228,N_16226);
and U16440 (N_16440,N_16219,N_16274);
nand U16441 (N_16441,N_16231,N_16192);
and U16442 (N_16442,N_16310,N_16318);
or U16443 (N_16443,N_16244,N_16272);
and U16444 (N_16444,N_16275,N_16229);
or U16445 (N_16445,N_16251,N_16313);
or U16446 (N_16446,N_16246,N_16280);
nand U16447 (N_16447,N_16299,N_16163);
nor U16448 (N_16448,N_16194,N_16191);
nor U16449 (N_16449,N_16176,N_16204);
xor U16450 (N_16450,N_16243,N_16196);
nand U16451 (N_16451,N_16197,N_16318);
nor U16452 (N_16452,N_16248,N_16217);
nand U16453 (N_16453,N_16300,N_16286);
nand U16454 (N_16454,N_16283,N_16175);
nor U16455 (N_16455,N_16313,N_16211);
nor U16456 (N_16456,N_16230,N_16314);
or U16457 (N_16457,N_16180,N_16212);
xor U16458 (N_16458,N_16303,N_16223);
nor U16459 (N_16459,N_16161,N_16178);
or U16460 (N_16460,N_16263,N_16206);
or U16461 (N_16461,N_16186,N_16223);
nand U16462 (N_16462,N_16243,N_16232);
nand U16463 (N_16463,N_16274,N_16304);
nand U16464 (N_16464,N_16185,N_16267);
or U16465 (N_16465,N_16314,N_16317);
xnor U16466 (N_16466,N_16287,N_16309);
or U16467 (N_16467,N_16200,N_16297);
or U16468 (N_16468,N_16310,N_16265);
nor U16469 (N_16469,N_16287,N_16248);
nor U16470 (N_16470,N_16271,N_16304);
or U16471 (N_16471,N_16165,N_16297);
nor U16472 (N_16472,N_16311,N_16294);
and U16473 (N_16473,N_16192,N_16198);
and U16474 (N_16474,N_16234,N_16168);
or U16475 (N_16475,N_16232,N_16312);
xor U16476 (N_16476,N_16239,N_16160);
or U16477 (N_16477,N_16304,N_16319);
nor U16478 (N_16478,N_16221,N_16236);
nor U16479 (N_16479,N_16161,N_16198);
nand U16480 (N_16480,N_16405,N_16378);
nand U16481 (N_16481,N_16446,N_16431);
nor U16482 (N_16482,N_16354,N_16384);
or U16483 (N_16483,N_16420,N_16403);
xnor U16484 (N_16484,N_16453,N_16357);
nand U16485 (N_16485,N_16460,N_16339);
nor U16486 (N_16486,N_16424,N_16331);
xor U16487 (N_16487,N_16335,N_16418);
or U16488 (N_16488,N_16345,N_16465);
nand U16489 (N_16489,N_16346,N_16373);
nor U16490 (N_16490,N_16321,N_16474);
nor U16491 (N_16491,N_16472,N_16391);
or U16492 (N_16492,N_16351,N_16401);
nand U16493 (N_16493,N_16320,N_16459);
or U16494 (N_16494,N_16364,N_16374);
and U16495 (N_16495,N_16417,N_16477);
or U16496 (N_16496,N_16326,N_16443);
nor U16497 (N_16497,N_16438,N_16385);
nand U16498 (N_16498,N_16455,N_16323);
nor U16499 (N_16499,N_16444,N_16437);
nand U16500 (N_16500,N_16458,N_16402);
xor U16501 (N_16501,N_16383,N_16361);
nor U16502 (N_16502,N_16473,N_16333);
xnor U16503 (N_16503,N_16362,N_16451);
and U16504 (N_16504,N_16434,N_16435);
or U16505 (N_16505,N_16375,N_16344);
nand U16506 (N_16506,N_16440,N_16388);
and U16507 (N_16507,N_16421,N_16408);
and U16508 (N_16508,N_16468,N_16399);
or U16509 (N_16509,N_16347,N_16426);
or U16510 (N_16510,N_16476,N_16380);
and U16511 (N_16511,N_16366,N_16400);
nor U16512 (N_16512,N_16479,N_16450);
nand U16513 (N_16513,N_16348,N_16397);
nand U16514 (N_16514,N_16360,N_16423);
and U16515 (N_16515,N_16356,N_16461);
xnor U16516 (N_16516,N_16328,N_16419);
nor U16517 (N_16517,N_16432,N_16466);
xnor U16518 (N_16518,N_16343,N_16336);
nand U16519 (N_16519,N_16386,N_16324);
nand U16520 (N_16520,N_16454,N_16330);
or U16521 (N_16521,N_16463,N_16379);
nand U16522 (N_16522,N_16377,N_16342);
and U16523 (N_16523,N_16387,N_16422);
nand U16524 (N_16524,N_16327,N_16449);
and U16525 (N_16525,N_16412,N_16365);
nand U16526 (N_16526,N_16329,N_16398);
or U16527 (N_16527,N_16441,N_16395);
nor U16528 (N_16528,N_16334,N_16475);
nor U16529 (N_16529,N_16325,N_16368);
nor U16530 (N_16530,N_16478,N_16404);
nand U16531 (N_16531,N_16358,N_16322);
or U16532 (N_16532,N_16390,N_16470);
nand U16533 (N_16533,N_16467,N_16427);
nand U16534 (N_16534,N_16382,N_16353);
xnor U16535 (N_16535,N_16436,N_16359);
nor U16536 (N_16536,N_16447,N_16363);
nor U16537 (N_16537,N_16337,N_16462);
nand U16538 (N_16538,N_16414,N_16396);
nand U16539 (N_16539,N_16376,N_16371);
or U16540 (N_16540,N_16350,N_16448);
nor U16541 (N_16541,N_16439,N_16457);
nand U16542 (N_16542,N_16433,N_16429);
nor U16543 (N_16543,N_16349,N_16392);
nor U16544 (N_16544,N_16411,N_16340);
or U16545 (N_16545,N_16416,N_16471);
nand U16546 (N_16546,N_16430,N_16367);
nand U16547 (N_16547,N_16389,N_16464);
nand U16548 (N_16548,N_16452,N_16445);
or U16549 (N_16549,N_16381,N_16332);
or U16550 (N_16550,N_16413,N_16456);
nor U16551 (N_16551,N_16442,N_16415);
nand U16552 (N_16552,N_16469,N_16355);
nor U16553 (N_16553,N_16394,N_16370);
nand U16554 (N_16554,N_16393,N_16428);
or U16555 (N_16555,N_16407,N_16341);
and U16556 (N_16556,N_16409,N_16425);
nor U16557 (N_16557,N_16406,N_16410);
nand U16558 (N_16558,N_16338,N_16369);
and U16559 (N_16559,N_16352,N_16372);
nand U16560 (N_16560,N_16353,N_16445);
or U16561 (N_16561,N_16364,N_16337);
xor U16562 (N_16562,N_16447,N_16344);
nor U16563 (N_16563,N_16449,N_16450);
and U16564 (N_16564,N_16360,N_16422);
nor U16565 (N_16565,N_16461,N_16478);
or U16566 (N_16566,N_16392,N_16405);
or U16567 (N_16567,N_16446,N_16429);
or U16568 (N_16568,N_16356,N_16329);
nor U16569 (N_16569,N_16460,N_16447);
nand U16570 (N_16570,N_16436,N_16333);
or U16571 (N_16571,N_16441,N_16431);
nand U16572 (N_16572,N_16454,N_16476);
nand U16573 (N_16573,N_16426,N_16429);
nand U16574 (N_16574,N_16374,N_16467);
nor U16575 (N_16575,N_16354,N_16349);
and U16576 (N_16576,N_16349,N_16430);
and U16577 (N_16577,N_16336,N_16361);
and U16578 (N_16578,N_16430,N_16399);
and U16579 (N_16579,N_16425,N_16350);
or U16580 (N_16580,N_16334,N_16370);
and U16581 (N_16581,N_16357,N_16380);
xnor U16582 (N_16582,N_16451,N_16406);
nand U16583 (N_16583,N_16437,N_16336);
nor U16584 (N_16584,N_16324,N_16340);
nand U16585 (N_16585,N_16479,N_16419);
or U16586 (N_16586,N_16383,N_16393);
xnor U16587 (N_16587,N_16333,N_16361);
nor U16588 (N_16588,N_16412,N_16469);
or U16589 (N_16589,N_16354,N_16379);
nor U16590 (N_16590,N_16387,N_16363);
or U16591 (N_16591,N_16338,N_16423);
nor U16592 (N_16592,N_16403,N_16321);
or U16593 (N_16593,N_16453,N_16432);
xor U16594 (N_16594,N_16439,N_16467);
or U16595 (N_16595,N_16468,N_16466);
or U16596 (N_16596,N_16447,N_16422);
or U16597 (N_16597,N_16392,N_16325);
and U16598 (N_16598,N_16436,N_16395);
or U16599 (N_16599,N_16478,N_16402);
nand U16600 (N_16600,N_16364,N_16454);
or U16601 (N_16601,N_16324,N_16362);
or U16602 (N_16602,N_16363,N_16384);
nand U16603 (N_16603,N_16367,N_16383);
nor U16604 (N_16604,N_16386,N_16462);
nor U16605 (N_16605,N_16320,N_16455);
or U16606 (N_16606,N_16445,N_16396);
nor U16607 (N_16607,N_16381,N_16457);
nor U16608 (N_16608,N_16344,N_16429);
nor U16609 (N_16609,N_16458,N_16449);
or U16610 (N_16610,N_16354,N_16364);
and U16611 (N_16611,N_16421,N_16459);
or U16612 (N_16612,N_16453,N_16379);
or U16613 (N_16613,N_16422,N_16373);
nor U16614 (N_16614,N_16433,N_16477);
nor U16615 (N_16615,N_16410,N_16478);
nor U16616 (N_16616,N_16356,N_16369);
nor U16617 (N_16617,N_16467,N_16428);
nand U16618 (N_16618,N_16359,N_16402);
or U16619 (N_16619,N_16408,N_16356);
and U16620 (N_16620,N_16475,N_16414);
and U16621 (N_16621,N_16391,N_16413);
nand U16622 (N_16622,N_16320,N_16371);
and U16623 (N_16623,N_16357,N_16370);
xor U16624 (N_16624,N_16419,N_16382);
and U16625 (N_16625,N_16399,N_16337);
nand U16626 (N_16626,N_16446,N_16456);
nand U16627 (N_16627,N_16411,N_16373);
nand U16628 (N_16628,N_16320,N_16372);
xor U16629 (N_16629,N_16394,N_16472);
nand U16630 (N_16630,N_16417,N_16381);
and U16631 (N_16631,N_16403,N_16356);
or U16632 (N_16632,N_16382,N_16437);
and U16633 (N_16633,N_16346,N_16412);
or U16634 (N_16634,N_16373,N_16471);
and U16635 (N_16635,N_16469,N_16327);
nand U16636 (N_16636,N_16343,N_16405);
and U16637 (N_16637,N_16454,N_16409);
nand U16638 (N_16638,N_16415,N_16432);
nand U16639 (N_16639,N_16335,N_16450);
nand U16640 (N_16640,N_16540,N_16607);
or U16641 (N_16641,N_16549,N_16508);
nand U16642 (N_16642,N_16569,N_16585);
xnor U16643 (N_16643,N_16589,N_16502);
nor U16644 (N_16644,N_16586,N_16595);
nor U16645 (N_16645,N_16612,N_16521);
and U16646 (N_16646,N_16551,N_16587);
xor U16647 (N_16647,N_16544,N_16517);
nor U16648 (N_16648,N_16611,N_16615);
and U16649 (N_16649,N_16494,N_16532);
nand U16650 (N_16650,N_16594,N_16571);
and U16651 (N_16651,N_16510,N_16545);
nand U16652 (N_16652,N_16499,N_16602);
or U16653 (N_16653,N_16489,N_16610);
and U16654 (N_16654,N_16538,N_16542);
nand U16655 (N_16655,N_16634,N_16503);
xnor U16656 (N_16656,N_16482,N_16627);
nand U16657 (N_16657,N_16591,N_16516);
nand U16658 (N_16658,N_16636,N_16509);
nor U16659 (N_16659,N_16547,N_16534);
or U16660 (N_16660,N_16605,N_16531);
xor U16661 (N_16661,N_16632,N_16548);
nand U16662 (N_16662,N_16487,N_16576);
or U16663 (N_16663,N_16480,N_16581);
nor U16664 (N_16664,N_16635,N_16565);
and U16665 (N_16665,N_16512,N_16578);
nand U16666 (N_16666,N_16572,N_16579);
and U16667 (N_16667,N_16570,N_16600);
and U16668 (N_16668,N_16630,N_16619);
or U16669 (N_16669,N_16527,N_16501);
and U16670 (N_16670,N_16568,N_16598);
and U16671 (N_16671,N_16537,N_16513);
nor U16672 (N_16672,N_16564,N_16523);
nor U16673 (N_16673,N_16546,N_16608);
nand U16674 (N_16674,N_16574,N_16530);
nand U16675 (N_16675,N_16535,N_16628);
or U16676 (N_16676,N_16604,N_16582);
or U16677 (N_16677,N_16563,N_16567);
and U16678 (N_16678,N_16518,N_16488);
or U16679 (N_16679,N_16614,N_16484);
xnor U16680 (N_16680,N_16491,N_16631);
and U16681 (N_16681,N_16486,N_16507);
and U16682 (N_16682,N_16533,N_16638);
nor U16683 (N_16683,N_16637,N_16560);
and U16684 (N_16684,N_16511,N_16596);
nand U16685 (N_16685,N_16559,N_16520);
and U16686 (N_16686,N_16492,N_16577);
or U16687 (N_16687,N_16500,N_16555);
nor U16688 (N_16688,N_16493,N_16498);
and U16689 (N_16689,N_16504,N_16519);
or U16690 (N_16690,N_16528,N_16485);
or U16691 (N_16691,N_16506,N_16624);
nand U16692 (N_16692,N_16603,N_16495);
nor U16693 (N_16693,N_16622,N_16558);
nand U16694 (N_16694,N_16522,N_16556);
or U16695 (N_16695,N_16590,N_16633);
and U16696 (N_16696,N_16609,N_16514);
nand U16697 (N_16697,N_16621,N_16561);
or U16698 (N_16698,N_16639,N_16490);
and U16699 (N_16699,N_16562,N_16606);
and U16700 (N_16700,N_16526,N_16557);
nor U16701 (N_16701,N_16505,N_16515);
nor U16702 (N_16702,N_16573,N_16481);
nor U16703 (N_16703,N_16583,N_16613);
nor U16704 (N_16704,N_16601,N_16541);
nor U16705 (N_16705,N_16543,N_16552);
and U16706 (N_16706,N_16616,N_16626);
and U16707 (N_16707,N_16625,N_16497);
nand U16708 (N_16708,N_16588,N_16496);
xor U16709 (N_16709,N_16584,N_16550);
nand U16710 (N_16710,N_16599,N_16593);
nand U16711 (N_16711,N_16529,N_16592);
and U16712 (N_16712,N_16566,N_16597);
and U16713 (N_16713,N_16539,N_16623);
or U16714 (N_16714,N_16553,N_16525);
or U16715 (N_16715,N_16620,N_16524);
or U16716 (N_16716,N_16536,N_16575);
nand U16717 (N_16717,N_16629,N_16617);
xor U16718 (N_16718,N_16580,N_16483);
and U16719 (N_16719,N_16554,N_16618);
nand U16720 (N_16720,N_16596,N_16585);
nand U16721 (N_16721,N_16620,N_16568);
nand U16722 (N_16722,N_16532,N_16495);
or U16723 (N_16723,N_16526,N_16513);
nor U16724 (N_16724,N_16622,N_16481);
or U16725 (N_16725,N_16490,N_16526);
and U16726 (N_16726,N_16573,N_16489);
nand U16727 (N_16727,N_16595,N_16532);
or U16728 (N_16728,N_16533,N_16579);
nand U16729 (N_16729,N_16559,N_16544);
and U16730 (N_16730,N_16564,N_16524);
xor U16731 (N_16731,N_16569,N_16578);
or U16732 (N_16732,N_16505,N_16527);
nor U16733 (N_16733,N_16626,N_16588);
and U16734 (N_16734,N_16562,N_16573);
nor U16735 (N_16735,N_16512,N_16584);
xnor U16736 (N_16736,N_16575,N_16577);
nand U16737 (N_16737,N_16581,N_16529);
or U16738 (N_16738,N_16558,N_16528);
nor U16739 (N_16739,N_16618,N_16481);
nand U16740 (N_16740,N_16607,N_16508);
nor U16741 (N_16741,N_16587,N_16495);
nand U16742 (N_16742,N_16556,N_16568);
nor U16743 (N_16743,N_16505,N_16522);
nor U16744 (N_16744,N_16586,N_16514);
xor U16745 (N_16745,N_16564,N_16485);
nand U16746 (N_16746,N_16569,N_16633);
nand U16747 (N_16747,N_16548,N_16588);
or U16748 (N_16748,N_16637,N_16601);
and U16749 (N_16749,N_16516,N_16582);
or U16750 (N_16750,N_16586,N_16503);
nand U16751 (N_16751,N_16575,N_16637);
and U16752 (N_16752,N_16603,N_16549);
xor U16753 (N_16753,N_16525,N_16558);
xnor U16754 (N_16754,N_16535,N_16514);
and U16755 (N_16755,N_16510,N_16594);
or U16756 (N_16756,N_16520,N_16502);
and U16757 (N_16757,N_16592,N_16535);
and U16758 (N_16758,N_16535,N_16529);
or U16759 (N_16759,N_16570,N_16582);
and U16760 (N_16760,N_16544,N_16534);
or U16761 (N_16761,N_16577,N_16485);
or U16762 (N_16762,N_16585,N_16605);
or U16763 (N_16763,N_16552,N_16503);
nor U16764 (N_16764,N_16505,N_16592);
or U16765 (N_16765,N_16580,N_16513);
and U16766 (N_16766,N_16523,N_16639);
nand U16767 (N_16767,N_16599,N_16614);
or U16768 (N_16768,N_16498,N_16593);
nand U16769 (N_16769,N_16544,N_16556);
nor U16770 (N_16770,N_16622,N_16525);
and U16771 (N_16771,N_16558,N_16617);
and U16772 (N_16772,N_16574,N_16583);
nor U16773 (N_16773,N_16506,N_16562);
and U16774 (N_16774,N_16521,N_16569);
or U16775 (N_16775,N_16571,N_16557);
or U16776 (N_16776,N_16511,N_16551);
nand U16777 (N_16777,N_16483,N_16614);
or U16778 (N_16778,N_16561,N_16515);
nand U16779 (N_16779,N_16536,N_16497);
or U16780 (N_16780,N_16515,N_16630);
nand U16781 (N_16781,N_16585,N_16608);
and U16782 (N_16782,N_16533,N_16535);
nand U16783 (N_16783,N_16580,N_16556);
nand U16784 (N_16784,N_16531,N_16513);
nor U16785 (N_16785,N_16602,N_16590);
nand U16786 (N_16786,N_16503,N_16532);
nor U16787 (N_16787,N_16491,N_16589);
nand U16788 (N_16788,N_16629,N_16602);
or U16789 (N_16789,N_16501,N_16609);
and U16790 (N_16790,N_16482,N_16580);
and U16791 (N_16791,N_16631,N_16619);
or U16792 (N_16792,N_16514,N_16599);
nand U16793 (N_16793,N_16497,N_16540);
nor U16794 (N_16794,N_16540,N_16581);
xnor U16795 (N_16795,N_16525,N_16604);
xor U16796 (N_16796,N_16630,N_16561);
or U16797 (N_16797,N_16531,N_16627);
xnor U16798 (N_16798,N_16546,N_16585);
and U16799 (N_16799,N_16507,N_16617);
or U16800 (N_16800,N_16724,N_16728);
nor U16801 (N_16801,N_16697,N_16718);
or U16802 (N_16802,N_16752,N_16745);
nand U16803 (N_16803,N_16787,N_16750);
nor U16804 (N_16804,N_16759,N_16783);
and U16805 (N_16805,N_16690,N_16756);
xnor U16806 (N_16806,N_16712,N_16676);
and U16807 (N_16807,N_16656,N_16658);
or U16808 (N_16808,N_16673,N_16738);
or U16809 (N_16809,N_16777,N_16726);
and U16810 (N_16810,N_16688,N_16735);
and U16811 (N_16811,N_16746,N_16739);
xnor U16812 (N_16812,N_16786,N_16730);
nor U16813 (N_16813,N_16644,N_16749);
nor U16814 (N_16814,N_16751,N_16797);
nand U16815 (N_16815,N_16766,N_16655);
and U16816 (N_16816,N_16686,N_16702);
or U16817 (N_16817,N_16679,N_16651);
xor U16818 (N_16818,N_16737,N_16683);
and U16819 (N_16819,N_16691,N_16727);
nand U16820 (N_16820,N_16641,N_16785);
and U16821 (N_16821,N_16663,N_16687);
nor U16822 (N_16822,N_16769,N_16798);
nand U16823 (N_16823,N_16707,N_16703);
nand U16824 (N_16824,N_16720,N_16781);
and U16825 (N_16825,N_16761,N_16714);
or U16826 (N_16826,N_16770,N_16700);
nor U16827 (N_16827,N_16732,N_16747);
nor U16828 (N_16828,N_16701,N_16775);
and U16829 (N_16829,N_16689,N_16742);
or U16830 (N_16830,N_16657,N_16760);
nand U16831 (N_16831,N_16767,N_16706);
nand U16832 (N_16832,N_16744,N_16722);
xnor U16833 (N_16833,N_16698,N_16672);
and U16834 (N_16834,N_16741,N_16662);
nand U16835 (N_16835,N_16771,N_16729);
nand U16836 (N_16836,N_16674,N_16725);
nand U16837 (N_16837,N_16757,N_16647);
nor U16838 (N_16838,N_16649,N_16723);
and U16839 (N_16839,N_16758,N_16789);
xnor U16840 (N_16840,N_16792,N_16665);
xnor U16841 (N_16841,N_16740,N_16659);
nor U16842 (N_16842,N_16768,N_16710);
xnor U16843 (N_16843,N_16645,N_16779);
or U16844 (N_16844,N_16754,N_16772);
nor U16845 (N_16845,N_16793,N_16668);
and U16846 (N_16846,N_16640,N_16708);
or U16847 (N_16847,N_16704,N_16650);
or U16848 (N_16848,N_16762,N_16646);
nand U16849 (N_16849,N_16664,N_16682);
nand U16850 (N_16850,N_16755,N_16764);
and U16851 (N_16851,N_16675,N_16719);
and U16852 (N_16852,N_16660,N_16780);
or U16853 (N_16853,N_16795,N_16791);
nand U16854 (N_16854,N_16654,N_16694);
and U16855 (N_16855,N_16788,N_16670);
or U16856 (N_16856,N_16695,N_16774);
and U16857 (N_16857,N_16748,N_16684);
nor U16858 (N_16858,N_16705,N_16782);
xnor U16859 (N_16859,N_16677,N_16716);
nand U16860 (N_16860,N_16661,N_16696);
xnor U16861 (N_16861,N_16715,N_16681);
and U16862 (N_16862,N_16709,N_16667);
or U16863 (N_16863,N_16776,N_16643);
nor U16864 (N_16864,N_16666,N_16733);
or U16865 (N_16865,N_16799,N_16796);
or U16866 (N_16866,N_16648,N_16731);
xor U16867 (N_16867,N_16693,N_16753);
nor U16868 (N_16868,N_16736,N_16721);
and U16869 (N_16869,N_16671,N_16778);
xnor U16870 (N_16870,N_16653,N_16790);
or U16871 (N_16871,N_16734,N_16685);
or U16872 (N_16872,N_16652,N_16743);
nand U16873 (N_16873,N_16773,N_16692);
or U16874 (N_16874,N_16669,N_16713);
and U16875 (N_16875,N_16717,N_16763);
nor U16876 (N_16876,N_16678,N_16784);
xor U16877 (N_16877,N_16680,N_16765);
nand U16878 (N_16878,N_16711,N_16642);
nand U16879 (N_16879,N_16699,N_16794);
or U16880 (N_16880,N_16794,N_16679);
nand U16881 (N_16881,N_16688,N_16648);
nand U16882 (N_16882,N_16678,N_16742);
and U16883 (N_16883,N_16757,N_16709);
nor U16884 (N_16884,N_16691,N_16659);
or U16885 (N_16885,N_16731,N_16792);
or U16886 (N_16886,N_16699,N_16695);
and U16887 (N_16887,N_16772,N_16707);
nand U16888 (N_16888,N_16729,N_16698);
nand U16889 (N_16889,N_16659,N_16731);
and U16890 (N_16890,N_16788,N_16720);
nor U16891 (N_16891,N_16749,N_16761);
or U16892 (N_16892,N_16699,N_16696);
or U16893 (N_16893,N_16718,N_16746);
or U16894 (N_16894,N_16697,N_16647);
nand U16895 (N_16895,N_16782,N_16783);
nand U16896 (N_16896,N_16667,N_16653);
nand U16897 (N_16897,N_16656,N_16653);
nor U16898 (N_16898,N_16651,N_16764);
nand U16899 (N_16899,N_16728,N_16721);
nand U16900 (N_16900,N_16755,N_16681);
nor U16901 (N_16901,N_16780,N_16738);
or U16902 (N_16902,N_16767,N_16680);
nor U16903 (N_16903,N_16671,N_16683);
nand U16904 (N_16904,N_16753,N_16740);
and U16905 (N_16905,N_16689,N_16700);
nor U16906 (N_16906,N_16723,N_16697);
nor U16907 (N_16907,N_16770,N_16781);
and U16908 (N_16908,N_16671,N_16681);
and U16909 (N_16909,N_16718,N_16674);
or U16910 (N_16910,N_16679,N_16660);
nor U16911 (N_16911,N_16698,N_16655);
and U16912 (N_16912,N_16716,N_16722);
and U16913 (N_16913,N_16663,N_16692);
nor U16914 (N_16914,N_16725,N_16737);
and U16915 (N_16915,N_16799,N_16770);
nand U16916 (N_16916,N_16645,N_16744);
xnor U16917 (N_16917,N_16683,N_16744);
nand U16918 (N_16918,N_16731,N_16645);
xor U16919 (N_16919,N_16704,N_16780);
nand U16920 (N_16920,N_16789,N_16684);
xor U16921 (N_16921,N_16659,N_16736);
or U16922 (N_16922,N_16795,N_16750);
nand U16923 (N_16923,N_16795,N_16746);
and U16924 (N_16924,N_16733,N_16661);
xor U16925 (N_16925,N_16777,N_16699);
and U16926 (N_16926,N_16717,N_16664);
and U16927 (N_16927,N_16715,N_16785);
xor U16928 (N_16928,N_16688,N_16696);
nor U16929 (N_16929,N_16747,N_16661);
xor U16930 (N_16930,N_16781,N_16785);
and U16931 (N_16931,N_16706,N_16748);
or U16932 (N_16932,N_16720,N_16780);
xnor U16933 (N_16933,N_16668,N_16758);
and U16934 (N_16934,N_16725,N_16646);
nand U16935 (N_16935,N_16766,N_16661);
and U16936 (N_16936,N_16641,N_16782);
nand U16937 (N_16937,N_16794,N_16772);
nor U16938 (N_16938,N_16669,N_16678);
or U16939 (N_16939,N_16729,N_16736);
and U16940 (N_16940,N_16709,N_16766);
xnor U16941 (N_16941,N_16648,N_16658);
or U16942 (N_16942,N_16762,N_16650);
nand U16943 (N_16943,N_16732,N_16700);
nand U16944 (N_16944,N_16736,N_16698);
nand U16945 (N_16945,N_16711,N_16762);
nor U16946 (N_16946,N_16790,N_16681);
or U16947 (N_16947,N_16743,N_16760);
nor U16948 (N_16948,N_16749,N_16754);
or U16949 (N_16949,N_16707,N_16799);
nand U16950 (N_16950,N_16648,N_16762);
nor U16951 (N_16951,N_16736,N_16700);
or U16952 (N_16952,N_16670,N_16688);
and U16953 (N_16953,N_16670,N_16758);
xnor U16954 (N_16954,N_16793,N_16710);
nor U16955 (N_16955,N_16667,N_16712);
nor U16956 (N_16956,N_16776,N_16667);
nand U16957 (N_16957,N_16791,N_16713);
or U16958 (N_16958,N_16781,N_16726);
nor U16959 (N_16959,N_16780,N_16672);
or U16960 (N_16960,N_16841,N_16920);
nand U16961 (N_16961,N_16810,N_16933);
and U16962 (N_16962,N_16839,N_16906);
or U16963 (N_16963,N_16931,N_16867);
or U16964 (N_16964,N_16859,N_16806);
and U16965 (N_16965,N_16958,N_16814);
and U16966 (N_16966,N_16916,N_16942);
nand U16967 (N_16967,N_16881,N_16945);
nand U16968 (N_16968,N_16832,N_16882);
nor U16969 (N_16969,N_16913,N_16877);
nor U16970 (N_16970,N_16929,N_16890);
nand U16971 (N_16971,N_16915,N_16866);
or U16972 (N_16972,N_16807,N_16860);
and U16973 (N_16973,N_16909,N_16956);
nor U16974 (N_16974,N_16932,N_16850);
and U16975 (N_16975,N_16918,N_16887);
nor U16976 (N_16976,N_16871,N_16917);
nand U16977 (N_16977,N_16959,N_16809);
or U16978 (N_16978,N_16910,N_16886);
or U16979 (N_16979,N_16837,N_16891);
nor U16980 (N_16980,N_16828,N_16822);
and U16981 (N_16981,N_16957,N_16800);
nand U16982 (N_16982,N_16901,N_16827);
nand U16983 (N_16983,N_16897,N_16889);
nor U16984 (N_16984,N_16879,N_16878);
nor U16985 (N_16985,N_16849,N_16936);
nor U16986 (N_16986,N_16944,N_16869);
and U16987 (N_16987,N_16876,N_16904);
nor U16988 (N_16988,N_16811,N_16863);
and U16989 (N_16989,N_16820,N_16935);
and U16990 (N_16990,N_16898,N_16924);
nor U16991 (N_16991,N_16934,N_16836);
and U16992 (N_16992,N_16812,N_16834);
nor U16993 (N_16993,N_16831,N_16838);
or U16994 (N_16994,N_16941,N_16856);
nor U16995 (N_16995,N_16946,N_16953);
nor U16996 (N_16996,N_16872,N_16949);
nand U16997 (N_16997,N_16902,N_16930);
or U16998 (N_16998,N_16895,N_16847);
nor U16999 (N_16999,N_16870,N_16845);
nor U17000 (N_17000,N_16923,N_16821);
nor U17001 (N_17001,N_16926,N_16844);
nand U17002 (N_17002,N_16899,N_16907);
nand U17003 (N_17003,N_16903,N_16857);
xor U17004 (N_17004,N_16880,N_16928);
nor U17005 (N_17005,N_16817,N_16846);
or U17006 (N_17006,N_16818,N_16803);
and U17007 (N_17007,N_16852,N_16911);
xor U17008 (N_17008,N_16939,N_16833);
nand U17009 (N_17009,N_16905,N_16805);
nor U17010 (N_17010,N_16842,N_16825);
or U17011 (N_17011,N_16912,N_16854);
or U17012 (N_17012,N_16873,N_16874);
nor U17013 (N_17013,N_16851,N_16853);
nor U17014 (N_17014,N_16885,N_16921);
or U17015 (N_17015,N_16840,N_16925);
xnor U17016 (N_17016,N_16816,N_16943);
nand U17017 (N_17017,N_16819,N_16896);
nand U17018 (N_17018,N_16919,N_16829);
xor U17019 (N_17019,N_16937,N_16861);
and U17020 (N_17020,N_16855,N_16802);
and U17021 (N_17021,N_16823,N_16883);
or U17022 (N_17022,N_16952,N_16824);
nand U17023 (N_17023,N_16801,N_16938);
and U17024 (N_17024,N_16947,N_16922);
and U17025 (N_17025,N_16948,N_16927);
nor U17026 (N_17026,N_16940,N_16858);
nand U17027 (N_17027,N_16813,N_16894);
or U17028 (N_17028,N_16865,N_16862);
xnor U17029 (N_17029,N_16815,N_16830);
nor U17030 (N_17030,N_16888,N_16900);
nor U17031 (N_17031,N_16914,N_16848);
or U17032 (N_17032,N_16893,N_16826);
nor U17033 (N_17033,N_16955,N_16808);
and U17034 (N_17034,N_16951,N_16875);
nor U17035 (N_17035,N_16864,N_16884);
and U17036 (N_17036,N_16954,N_16835);
nand U17037 (N_17037,N_16868,N_16804);
or U17038 (N_17038,N_16908,N_16892);
and U17039 (N_17039,N_16843,N_16950);
nand U17040 (N_17040,N_16811,N_16827);
xnor U17041 (N_17041,N_16882,N_16941);
nand U17042 (N_17042,N_16823,N_16944);
or U17043 (N_17043,N_16926,N_16808);
nand U17044 (N_17044,N_16896,N_16862);
and U17045 (N_17045,N_16843,N_16904);
xor U17046 (N_17046,N_16894,N_16946);
nor U17047 (N_17047,N_16882,N_16916);
or U17048 (N_17048,N_16806,N_16949);
nor U17049 (N_17049,N_16807,N_16872);
or U17050 (N_17050,N_16920,N_16924);
nand U17051 (N_17051,N_16808,N_16941);
nor U17052 (N_17052,N_16817,N_16822);
xor U17053 (N_17053,N_16898,N_16950);
nand U17054 (N_17054,N_16862,N_16927);
nor U17055 (N_17055,N_16909,N_16957);
or U17056 (N_17056,N_16840,N_16959);
nand U17057 (N_17057,N_16943,N_16940);
xor U17058 (N_17058,N_16908,N_16878);
and U17059 (N_17059,N_16850,N_16846);
and U17060 (N_17060,N_16949,N_16887);
or U17061 (N_17061,N_16807,N_16914);
nand U17062 (N_17062,N_16936,N_16886);
nand U17063 (N_17063,N_16876,N_16914);
nand U17064 (N_17064,N_16949,N_16852);
or U17065 (N_17065,N_16883,N_16834);
nor U17066 (N_17066,N_16842,N_16930);
and U17067 (N_17067,N_16920,N_16898);
nand U17068 (N_17068,N_16827,N_16864);
nor U17069 (N_17069,N_16847,N_16907);
nand U17070 (N_17070,N_16819,N_16921);
or U17071 (N_17071,N_16855,N_16844);
and U17072 (N_17072,N_16817,N_16915);
and U17073 (N_17073,N_16930,N_16869);
nor U17074 (N_17074,N_16850,N_16893);
or U17075 (N_17075,N_16940,N_16957);
and U17076 (N_17076,N_16925,N_16818);
and U17077 (N_17077,N_16814,N_16930);
nand U17078 (N_17078,N_16898,N_16802);
or U17079 (N_17079,N_16945,N_16909);
nor U17080 (N_17080,N_16907,N_16908);
xor U17081 (N_17081,N_16921,N_16886);
or U17082 (N_17082,N_16846,N_16803);
nand U17083 (N_17083,N_16803,N_16899);
and U17084 (N_17084,N_16936,N_16892);
or U17085 (N_17085,N_16860,N_16871);
or U17086 (N_17086,N_16876,N_16949);
or U17087 (N_17087,N_16889,N_16902);
xor U17088 (N_17088,N_16800,N_16868);
and U17089 (N_17089,N_16856,N_16909);
nand U17090 (N_17090,N_16870,N_16843);
and U17091 (N_17091,N_16959,N_16803);
nand U17092 (N_17092,N_16849,N_16815);
and U17093 (N_17093,N_16809,N_16886);
or U17094 (N_17094,N_16830,N_16834);
and U17095 (N_17095,N_16949,N_16864);
or U17096 (N_17096,N_16872,N_16844);
and U17097 (N_17097,N_16956,N_16907);
and U17098 (N_17098,N_16860,N_16954);
and U17099 (N_17099,N_16953,N_16951);
and U17100 (N_17100,N_16945,N_16925);
nor U17101 (N_17101,N_16946,N_16803);
and U17102 (N_17102,N_16842,N_16848);
nand U17103 (N_17103,N_16903,N_16863);
nor U17104 (N_17104,N_16855,N_16938);
or U17105 (N_17105,N_16908,N_16894);
or U17106 (N_17106,N_16812,N_16850);
or U17107 (N_17107,N_16829,N_16855);
and U17108 (N_17108,N_16885,N_16872);
nor U17109 (N_17109,N_16957,N_16906);
nand U17110 (N_17110,N_16910,N_16862);
nor U17111 (N_17111,N_16845,N_16909);
or U17112 (N_17112,N_16859,N_16908);
and U17113 (N_17113,N_16942,N_16948);
or U17114 (N_17114,N_16903,N_16929);
or U17115 (N_17115,N_16843,N_16956);
nand U17116 (N_17116,N_16807,N_16908);
nor U17117 (N_17117,N_16875,N_16811);
and U17118 (N_17118,N_16929,N_16856);
xor U17119 (N_17119,N_16805,N_16811);
nor U17120 (N_17120,N_16993,N_17106);
nor U17121 (N_17121,N_17017,N_16973);
or U17122 (N_17122,N_17070,N_17095);
nand U17123 (N_17123,N_17071,N_17042);
and U17124 (N_17124,N_17029,N_16991);
and U17125 (N_17125,N_17039,N_16981);
nand U17126 (N_17126,N_17012,N_17066);
and U17127 (N_17127,N_17020,N_17015);
nand U17128 (N_17128,N_17072,N_17030);
or U17129 (N_17129,N_16960,N_16992);
or U17130 (N_17130,N_17045,N_17115);
or U17131 (N_17131,N_17024,N_17019);
nand U17132 (N_17132,N_17105,N_16977);
nand U17133 (N_17133,N_17097,N_17076);
nor U17134 (N_17134,N_17033,N_17018);
nand U17135 (N_17135,N_17078,N_17092);
nor U17136 (N_17136,N_16999,N_17084);
or U17137 (N_17137,N_17050,N_17113);
and U17138 (N_17138,N_17090,N_17001);
or U17139 (N_17139,N_17040,N_17116);
nor U17140 (N_17140,N_17041,N_17061);
and U17141 (N_17141,N_17016,N_16970);
and U17142 (N_17142,N_16963,N_17036);
and U17143 (N_17143,N_17088,N_17096);
nand U17144 (N_17144,N_17021,N_17044);
and U17145 (N_17145,N_17100,N_17002);
nand U17146 (N_17146,N_17117,N_17079);
or U17147 (N_17147,N_16980,N_17109);
nor U17148 (N_17148,N_17074,N_16974);
nor U17149 (N_17149,N_16967,N_17058);
or U17150 (N_17150,N_17101,N_16982);
and U17151 (N_17151,N_16965,N_17028);
or U17152 (N_17152,N_17091,N_16968);
nor U17153 (N_17153,N_16994,N_17006);
xor U17154 (N_17154,N_17059,N_17063);
and U17155 (N_17155,N_16979,N_17089);
nand U17156 (N_17156,N_17085,N_16966);
nor U17157 (N_17157,N_17013,N_17047);
nand U17158 (N_17158,N_16988,N_17065);
nor U17159 (N_17159,N_17077,N_17069);
nor U17160 (N_17160,N_17064,N_16976);
nor U17161 (N_17161,N_16987,N_16986);
and U17162 (N_17162,N_16989,N_17087);
nor U17163 (N_17163,N_17034,N_17111);
nand U17164 (N_17164,N_16972,N_17035);
nor U17165 (N_17165,N_17032,N_16964);
or U17166 (N_17166,N_16997,N_17062);
or U17167 (N_17167,N_17114,N_17054);
nor U17168 (N_17168,N_17043,N_16998);
xor U17169 (N_17169,N_17031,N_17060);
nand U17170 (N_17170,N_16962,N_17057);
or U17171 (N_17171,N_17112,N_16983);
nand U17172 (N_17172,N_17104,N_17086);
or U17173 (N_17173,N_17055,N_17108);
nand U17174 (N_17174,N_17037,N_17075);
nand U17175 (N_17175,N_17011,N_17093);
nor U17176 (N_17176,N_17000,N_17073);
or U17177 (N_17177,N_17102,N_17004);
nand U17178 (N_17178,N_17022,N_17007);
nand U17179 (N_17179,N_17094,N_16961);
nor U17180 (N_17180,N_17026,N_16996);
and U17181 (N_17181,N_17027,N_17008);
and U17182 (N_17182,N_17081,N_17010);
nand U17183 (N_17183,N_17005,N_17119);
and U17184 (N_17184,N_17098,N_16985);
nor U17185 (N_17185,N_16971,N_17118);
or U17186 (N_17186,N_17067,N_17014);
xor U17187 (N_17187,N_17103,N_17009);
or U17188 (N_17188,N_17038,N_17025);
or U17189 (N_17189,N_17080,N_17110);
and U17190 (N_17190,N_16978,N_17068);
or U17191 (N_17191,N_17053,N_17049);
nand U17192 (N_17192,N_16984,N_17003);
nor U17193 (N_17193,N_17099,N_16969);
xnor U17194 (N_17194,N_17051,N_17107);
nor U17195 (N_17195,N_16990,N_17083);
nand U17196 (N_17196,N_17046,N_17082);
xor U17197 (N_17197,N_16995,N_17048);
nor U17198 (N_17198,N_17023,N_16975);
or U17199 (N_17199,N_17052,N_17056);
xnor U17200 (N_17200,N_17067,N_17002);
or U17201 (N_17201,N_17007,N_17080);
nand U17202 (N_17202,N_17001,N_17081);
and U17203 (N_17203,N_17100,N_17114);
nand U17204 (N_17204,N_17079,N_17007);
or U17205 (N_17205,N_17091,N_16979);
or U17206 (N_17206,N_17033,N_17091);
and U17207 (N_17207,N_17030,N_16972);
nand U17208 (N_17208,N_17065,N_17068);
xnor U17209 (N_17209,N_16966,N_17036);
nor U17210 (N_17210,N_17085,N_17029);
nand U17211 (N_17211,N_17014,N_17088);
xnor U17212 (N_17212,N_17083,N_17004);
or U17213 (N_17213,N_17034,N_17024);
nand U17214 (N_17214,N_17007,N_17031);
and U17215 (N_17215,N_16999,N_17107);
and U17216 (N_17216,N_17065,N_17054);
or U17217 (N_17217,N_17118,N_17103);
or U17218 (N_17218,N_16972,N_17102);
and U17219 (N_17219,N_16970,N_17047);
xor U17220 (N_17220,N_17005,N_17096);
nand U17221 (N_17221,N_17056,N_17046);
or U17222 (N_17222,N_16963,N_17015);
nand U17223 (N_17223,N_16986,N_16963);
and U17224 (N_17224,N_17057,N_17075);
nand U17225 (N_17225,N_17012,N_17118);
nor U17226 (N_17226,N_17100,N_17050);
and U17227 (N_17227,N_16987,N_17114);
and U17228 (N_17228,N_17001,N_16988);
xor U17229 (N_17229,N_17012,N_17011);
and U17230 (N_17230,N_17004,N_17089);
nor U17231 (N_17231,N_16960,N_17041);
nor U17232 (N_17232,N_17088,N_17059);
and U17233 (N_17233,N_17087,N_17062);
nor U17234 (N_17234,N_16993,N_17052);
and U17235 (N_17235,N_17020,N_17055);
nand U17236 (N_17236,N_17059,N_16965);
nand U17237 (N_17237,N_17103,N_17067);
and U17238 (N_17238,N_17072,N_17091);
and U17239 (N_17239,N_17012,N_16990);
and U17240 (N_17240,N_16996,N_17097);
nand U17241 (N_17241,N_16972,N_17092);
nor U17242 (N_17242,N_17117,N_17029);
and U17243 (N_17243,N_17034,N_17022);
or U17244 (N_17244,N_17063,N_17092);
or U17245 (N_17245,N_17052,N_17068);
nor U17246 (N_17246,N_17064,N_16980);
and U17247 (N_17247,N_17034,N_17054);
nor U17248 (N_17248,N_17008,N_16991);
nor U17249 (N_17249,N_17041,N_17038);
nand U17250 (N_17250,N_17077,N_17046);
nor U17251 (N_17251,N_16995,N_17040);
or U17252 (N_17252,N_17085,N_17038);
nor U17253 (N_17253,N_17041,N_17021);
or U17254 (N_17254,N_17071,N_16981);
or U17255 (N_17255,N_17112,N_17057);
nor U17256 (N_17256,N_17015,N_16983);
and U17257 (N_17257,N_17027,N_16983);
xor U17258 (N_17258,N_17061,N_17004);
nand U17259 (N_17259,N_17048,N_17105);
or U17260 (N_17260,N_17118,N_17108);
and U17261 (N_17261,N_17025,N_17111);
nand U17262 (N_17262,N_17018,N_17079);
or U17263 (N_17263,N_16975,N_16997);
and U17264 (N_17264,N_17099,N_17052);
nand U17265 (N_17265,N_17113,N_16975);
and U17266 (N_17266,N_17024,N_16989);
nor U17267 (N_17267,N_17050,N_16979);
and U17268 (N_17268,N_17049,N_16980);
and U17269 (N_17269,N_16976,N_17049);
or U17270 (N_17270,N_17081,N_17068);
xnor U17271 (N_17271,N_17092,N_17005);
and U17272 (N_17272,N_17010,N_16988);
nor U17273 (N_17273,N_17012,N_17001);
or U17274 (N_17274,N_17119,N_16983);
nor U17275 (N_17275,N_17013,N_17034);
nor U17276 (N_17276,N_17053,N_17067);
xor U17277 (N_17277,N_17017,N_17096);
nand U17278 (N_17278,N_17073,N_17025);
and U17279 (N_17279,N_17030,N_16997);
or U17280 (N_17280,N_17248,N_17246);
nand U17281 (N_17281,N_17237,N_17195);
nor U17282 (N_17282,N_17247,N_17129);
xnor U17283 (N_17283,N_17260,N_17267);
nand U17284 (N_17284,N_17207,N_17158);
nor U17285 (N_17285,N_17160,N_17176);
nor U17286 (N_17286,N_17212,N_17251);
nand U17287 (N_17287,N_17208,N_17189);
xnor U17288 (N_17288,N_17214,N_17133);
nor U17289 (N_17289,N_17161,N_17229);
nand U17290 (N_17290,N_17183,N_17187);
and U17291 (N_17291,N_17264,N_17139);
nand U17292 (N_17292,N_17234,N_17249);
or U17293 (N_17293,N_17209,N_17140);
nand U17294 (N_17294,N_17204,N_17170);
xor U17295 (N_17295,N_17174,N_17220);
or U17296 (N_17296,N_17159,N_17203);
nor U17297 (N_17297,N_17223,N_17134);
nor U17298 (N_17298,N_17157,N_17132);
nor U17299 (N_17299,N_17205,N_17142);
xnor U17300 (N_17300,N_17269,N_17181);
nor U17301 (N_17301,N_17263,N_17166);
nand U17302 (N_17302,N_17256,N_17135);
nand U17303 (N_17303,N_17252,N_17184);
and U17304 (N_17304,N_17198,N_17180);
and U17305 (N_17305,N_17255,N_17165);
xor U17306 (N_17306,N_17143,N_17227);
and U17307 (N_17307,N_17153,N_17210);
nand U17308 (N_17308,N_17137,N_17240);
or U17309 (N_17309,N_17164,N_17231);
or U17310 (N_17310,N_17215,N_17224);
xor U17311 (N_17311,N_17202,N_17141);
or U17312 (N_17312,N_17156,N_17125);
nor U17313 (N_17313,N_17197,N_17236);
nand U17314 (N_17314,N_17254,N_17276);
or U17315 (N_17315,N_17238,N_17225);
nor U17316 (N_17316,N_17122,N_17257);
or U17317 (N_17317,N_17121,N_17173);
or U17318 (N_17318,N_17235,N_17162);
and U17319 (N_17319,N_17178,N_17128);
nor U17320 (N_17320,N_17278,N_17154);
nand U17321 (N_17321,N_17136,N_17192);
and U17322 (N_17322,N_17279,N_17138);
nor U17323 (N_17323,N_17123,N_17222);
nor U17324 (N_17324,N_17230,N_17241);
xor U17325 (N_17325,N_17262,N_17185);
nand U17326 (N_17326,N_17270,N_17219);
nand U17327 (N_17327,N_17146,N_17145);
nand U17328 (N_17328,N_17211,N_17179);
nand U17329 (N_17329,N_17194,N_17206);
nor U17330 (N_17330,N_17274,N_17167);
nand U17331 (N_17331,N_17131,N_17265);
nand U17332 (N_17332,N_17243,N_17268);
nand U17333 (N_17333,N_17186,N_17193);
or U17334 (N_17334,N_17196,N_17188);
and U17335 (N_17335,N_17150,N_17199);
nor U17336 (N_17336,N_17261,N_17259);
nor U17337 (N_17337,N_17266,N_17201);
nor U17338 (N_17338,N_17163,N_17120);
and U17339 (N_17339,N_17124,N_17126);
and U17340 (N_17340,N_17168,N_17169);
or U17341 (N_17341,N_17277,N_17190);
nand U17342 (N_17342,N_17244,N_17144);
nand U17343 (N_17343,N_17271,N_17242);
nand U17344 (N_17344,N_17149,N_17232);
nor U17345 (N_17345,N_17172,N_17273);
xor U17346 (N_17346,N_17250,N_17275);
or U17347 (N_17347,N_17151,N_17148);
and U17348 (N_17348,N_17175,N_17272);
nor U17349 (N_17349,N_17221,N_17217);
nor U17350 (N_17350,N_17228,N_17233);
or U17351 (N_17351,N_17171,N_17258);
nand U17352 (N_17352,N_17253,N_17177);
nand U17353 (N_17353,N_17155,N_17127);
and U17354 (N_17354,N_17245,N_17147);
nor U17355 (N_17355,N_17130,N_17213);
nand U17356 (N_17356,N_17200,N_17239);
and U17357 (N_17357,N_17218,N_17216);
nor U17358 (N_17358,N_17191,N_17226);
nand U17359 (N_17359,N_17182,N_17152);
nand U17360 (N_17360,N_17253,N_17213);
nand U17361 (N_17361,N_17130,N_17206);
or U17362 (N_17362,N_17122,N_17235);
and U17363 (N_17363,N_17229,N_17140);
xnor U17364 (N_17364,N_17144,N_17235);
and U17365 (N_17365,N_17236,N_17277);
nand U17366 (N_17366,N_17165,N_17214);
or U17367 (N_17367,N_17234,N_17225);
xor U17368 (N_17368,N_17144,N_17136);
nand U17369 (N_17369,N_17138,N_17135);
nor U17370 (N_17370,N_17262,N_17251);
nand U17371 (N_17371,N_17187,N_17211);
or U17372 (N_17372,N_17124,N_17257);
and U17373 (N_17373,N_17132,N_17215);
nor U17374 (N_17374,N_17178,N_17160);
and U17375 (N_17375,N_17127,N_17187);
nor U17376 (N_17376,N_17155,N_17184);
nor U17377 (N_17377,N_17205,N_17274);
or U17378 (N_17378,N_17125,N_17266);
nor U17379 (N_17379,N_17253,N_17279);
and U17380 (N_17380,N_17228,N_17238);
and U17381 (N_17381,N_17225,N_17149);
or U17382 (N_17382,N_17139,N_17237);
nor U17383 (N_17383,N_17137,N_17195);
and U17384 (N_17384,N_17184,N_17168);
nand U17385 (N_17385,N_17130,N_17214);
nand U17386 (N_17386,N_17256,N_17272);
or U17387 (N_17387,N_17271,N_17272);
and U17388 (N_17388,N_17259,N_17210);
and U17389 (N_17389,N_17156,N_17145);
nand U17390 (N_17390,N_17121,N_17136);
xor U17391 (N_17391,N_17172,N_17239);
and U17392 (N_17392,N_17124,N_17142);
and U17393 (N_17393,N_17149,N_17154);
nor U17394 (N_17394,N_17141,N_17236);
and U17395 (N_17395,N_17176,N_17245);
or U17396 (N_17396,N_17154,N_17258);
nor U17397 (N_17397,N_17184,N_17195);
and U17398 (N_17398,N_17261,N_17144);
nand U17399 (N_17399,N_17128,N_17157);
xor U17400 (N_17400,N_17211,N_17151);
or U17401 (N_17401,N_17274,N_17149);
and U17402 (N_17402,N_17250,N_17149);
nand U17403 (N_17403,N_17172,N_17205);
nor U17404 (N_17404,N_17221,N_17176);
nand U17405 (N_17405,N_17274,N_17248);
or U17406 (N_17406,N_17189,N_17194);
or U17407 (N_17407,N_17148,N_17209);
and U17408 (N_17408,N_17265,N_17178);
or U17409 (N_17409,N_17243,N_17173);
xnor U17410 (N_17410,N_17210,N_17277);
or U17411 (N_17411,N_17279,N_17185);
or U17412 (N_17412,N_17212,N_17229);
nor U17413 (N_17413,N_17208,N_17222);
nor U17414 (N_17414,N_17154,N_17174);
or U17415 (N_17415,N_17197,N_17256);
nand U17416 (N_17416,N_17235,N_17188);
nor U17417 (N_17417,N_17183,N_17124);
or U17418 (N_17418,N_17128,N_17255);
and U17419 (N_17419,N_17158,N_17137);
nor U17420 (N_17420,N_17226,N_17127);
xor U17421 (N_17421,N_17263,N_17279);
nand U17422 (N_17422,N_17161,N_17268);
nand U17423 (N_17423,N_17147,N_17161);
and U17424 (N_17424,N_17145,N_17253);
and U17425 (N_17425,N_17233,N_17168);
nor U17426 (N_17426,N_17214,N_17168);
nand U17427 (N_17427,N_17244,N_17122);
nand U17428 (N_17428,N_17215,N_17155);
nand U17429 (N_17429,N_17194,N_17276);
xor U17430 (N_17430,N_17122,N_17194);
and U17431 (N_17431,N_17160,N_17142);
nor U17432 (N_17432,N_17147,N_17158);
nand U17433 (N_17433,N_17245,N_17138);
nor U17434 (N_17434,N_17182,N_17149);
xnor U17435 (N_17435,N_17263,N_17221);
nand U17436 (N_17436,N_17278,N_17140);
nand U17437 (N_17437,N_17252,N_17179);
and U17438 (N_17438,N_17160,N_17174);
nand U17439 (N_17439,N_17194,N_17211);
nor U17440 (N_17440,N_17289,N_17330);
nand U17441 (N_17441,N_17290,N_17389);
nand U17442 (N_17442,N_17419,N_17365);
or U17443 (N_17443,N_17380,N_17418);
xnor U17444 (N_17444,N_17333,N_17358);
and U17445 (N_17445,N_17406,N_17430);
or U17446 (N_17446,N_17382,N_17308);
or U17447 (N_17447,N_17386,N_17310);
nor U17448 (N_17448,N_17309,N_17295);
nand U17449 (N_17449,N_17307,N_17306);
and U17450 (N_17450,N_17345,N_17428);
xnor U17451 (N_17451,N_17313,N_17281);
nor U17452 (N_17452,N_17392,N_17320);
nor U17453 (N_17453,N_17400,N_17401);
nand U17454 (N_17454,N_17364,N_17414);
nand U17455 (N_17455,N_17360,N_17394);
nor U17456 (N_17456,N_17293,N_17422);
nand U17457 (N_17457,N_17356,N_17311);
xnor U17458 (N_17458,N_17397,N_17416);
or U17459 (N_17459,N_17425,N_17421);
or U17460 (N_17460,N_17375,N_17336);
and U17461 (N_17461,N_17322,N_17390);
or U17462 (N_17462,N_17357,N_17434);
or U17463 (N_17463,N_17427,N_17341);
nor U17464 (N_17464,N_17298,N_17362);
and U17465 (N_17465,N_17292,N_17299);
nor U17466 (N_17466,N_17324,N_17370);
nor U17467 (N_17467,N_17346,N_17319);
nor U17468 (N_17468,N_17305,N_17438);
nor U17469 (N_17469,N_17371,N_17355);
nand U17470 (N_17470,N_17409,N_17353);
or U17471 (N_17471,N_17300,N_17368);
nor U17472 (N_17472,N_17399,N_17412);
or U17473 (N_17473,N_17315,N_17294);
or U17474 (N_17474,N_17435,N_17436);
nor U17475 (N_17475,N_17391,N_17420);
nand U17476 (N_17476,N_17326,N_17302);
or U17477 (N_17477,N_17407,N_17429);
nand U17478 (N_17478,N_17351,N_17282);
xor U17479 (N_17479,N_17384,N_17331);
nand U17480 (N_17480,N_17378,N_17348);
nor U17481 (N_17481,N_17361,N_17334);
nor U17482 (N_17482,N_17318,N_17424);
nor U17483 (N_17483,N_17321,N_17372);
or U17484 (N_17484,N_17343,N_17433);
nor U17485 (N_17485,N_17297,N_17437);
nor U17486 (N_17486,N_17410,N_17342);
and U17487 (N_17487,N_17396,N_17325);
nand U17488 (N_17488,N_17393,N_17347);
nand U17489 (N_17489,N_17340,N_17439);
nand U17490 (N_17490,N_17363,N_17316);
and U17491 (N_17491,N_17423,N_17344);
and U17492 (N_17492,N_17312,N_17402);
xor U17493 (N_17493,N_17323,N_17349);
and U17494 (N_17494,N_17359,N_17301);
or U17495 (N_17495,N_17350,N_17432);
xnor U17496 (N_17496,N_17303,N_17403);
and U17497 (N_17497,N_17404,N_17426);
or U17498 (N_17498,N_17337,N_17338);
nand U17499 (N_17499,N_17374,N_17398);
nand U17500 (N_17500,N_17369,N_17376);
and U17501 (N_17501,N_17385,N_17328);
or U17502 (N_17502,N_17317,N_17408);
nand U17503 (N_17503,N_17383,N_17286);
or U17504 (N_17504,N_17379,N_17431);
or U17505 (N_17505,N_17377,N_17327);
nand U17506 (N_17506,N_17288,N_17332);
or U17507 (N_17507,N_17413,N_17387);
nand U17508 (N_17508,N_17283,N_17417);
or U17509 (N_17509,N_17352,N_17366);
xnor U17510 (N_17510,N_17388,N_17304);
xnor U17511 (N_17511,N_17411,N_17291);
or U17512 (N_17512,N_17296,N_17280);
nand U17513 (N_17513,N_17314,N_17329);
or U17514 (N_17514,N_17415,N_17373);
nor U17515 (N_17515,N_17354,N_17287);
or U17516 (N_17516,N_17339,N_17367);
or U17517 (N_17517,N_17381,N_17405);
nand U17518 (N_17518,N_17395,N_17284);
and U17519 (N_17519,N_17285,N_17335);
and U17520 (N_17520,N_17376,N_17330);
and U17521 (N_17521,N_17354,N_17296);
and U17522 (N_17522,N_17370,N_17404);
nand U17523 (N_17523,N_17431,N_17313);
nor U17524 (N_17524,N_17308,N_17372);
or U17525 (N_17525,N_17330,N_17410);
or U17526 (N_17526,N_17410,N_17338);
and U17527 (N_17527,N_17304,N_17337);
or U17528 (N_17528,N_17360,N_17426);
nand U17529 (N_17529,N_17389,N_17340);
nand U17530 (N_17530,N_17303,N_17337);
nand U17531 (N_17531,N_17310,N_17416);
and U17532 (N_17532,N_17388,N_17381);
or U17533 (N_17533,N_17356,N_17401);
or U17534 (N_17534,N_17305,N_17422);
nor U17535 (N_17535,N_17366,N_17315);
or U17536 (N_17536,N_17329,N_17308);
nor U17537 (N_17537,N_17345,N_17364);
nor U17538 (N_17538,N_17384,N_17338);
or U17539 (N_17539,N_17389,N_17368);
xnor U17540 (N_17540,N_17405,N_17346);
nand U17541 (N_17541,N_17302,N_17340);
or U17542 (N_17542,N_17373,N_17362);
and U17543 (N_17543,N_17422,N_17394);
or U17544 (N_17544,N_17313,N_17331);
xnor U17545 (N_17545,N_17384,N_17376);
or U17546 (N_17546,N_17334,N_17436);
nand U17547 (N_17547,N_17287,N_17418);
or U17548 (N_17548,N_17346,N_17419);
and U17549 (N_17549,N_17406,N_17434);
or U17550 (N_17550,N_17433,N_17356);
nor U17551 (N_17551,N_17347,N_17329);
nor U17552 (N_17552,N_17307,N_17302);
nand U17553 (N_17553,N_17415,N_17425);
nand U17554 (N_17554,N_17426,N_17399);
nand U17555 (N_17555,N_17401,N_17342);
or U17556 (N_17556,N_17307,N_17351);
or U17557 (N_17557,N_17351,N_17418);
nor U17558 (N_17558,N_17397,N_17324);
nor U17559 (N_17559,N_17333,N_17345);
nor U17560 (N_17560,N_17283,N_17294);
nand U17561 (N_17561,N_17432,N_17284);
or U17562 (N_17562,N_17370,N_17428);
nand U17563 (N_17563,N_17419,N_17434);
nor U17564 (N_17564,N_17420,N_17396);
and U17565 (N_17565,N_17416,N_17302);
nand U17566 (N_17566,N_17373,N_17355);
nand U17567 (N_17567,N_17310,N_17292);
and U17568 (N_17568,N_17439,N_17330);
nand U17569 (N_17569,N_17286,N_17365);
or U17570 (N_17570,N_17386,N_17362);
and U17571 (N_17571,N_17314,N_17319);
nand U17572 (N_17572,N_17333,N_17352);
nor U17573 (N_17573,N_17404,N_17355);
nand U17574 (N_17574,N_17377,N_17362);
and U17575 (N_17575,N_17342,N_17396);
nand U17576 (N_17576,N_17325,N_17376);
and U17577 (N_17577,N_17413,N_17349);
nor U17578 (N_17578,N_17375,N_17321);
nor U17579 (N_17579,N_17396,N_17353);
and U17580 (N_17580,N_17310,N_17345);
and U17581 (N_17581,N_17359,N_17307);
and U17582 (N_17582,N_17311,N_17370);
or U17583 (N_17583,N_17378,N_17436);
nand U17584 (N_17584,N_17321,N_17297);
or U17585 (N_17585,N_17329,N_17352);
nor U17586 (N_17586,N_17416,N_17280);
or U17587 (N_17587,N_17299,N_17420);
and U17588 (N_17588,N_17334,N_17390);
nand U17589 (N_17589,N_17396,N_17354);
and U17590 (N_17590,N_17285,N_17283);
nand U17591 (N_17591,N_17284,N_17307);
xor U17592 (N_17592,N_17422,N_17386);
and U17593 (N_17593,N_17417,N_17287);
xor U17594 (N_17594,N_17366,N_17429);
nor U17595 (N_17595,N_17350,N_17286);
nor U17596 (N_17596,N_17280,N_17331);
or U17597 (N_17597,N_17412,N_17401);
nor U17598 (N_17598,N_17361,N_17287);
and U17599 (N_17599,N_17396,N_17361);
nand U17600 (N_17600,N_17522,N_17504);
xnor U17601 (N_17601,N_17448,N_17546);
or U17602 (N_17602,N_17581,N_17515);
nand U17603 (N_17603,N_17517,N_17529);
and U17604 (N_17604,N_17580,N_17582);
and U17605 (N_17605,N_17458,N_17533);
nand U17606 (N_17606,N_17579,N_17550);
nand U17607 (N_17607,N_17551,N_17568);
nand U17608 (N_17608,N_17564,N_17468);
and U17609 (N_17609,N_17501,N_17594);
nand U17610 (N_17610,N_17491,N_17526);
nor U17611 (N_17611,N_17471,N_17454);
or U17612 (N_17612,N_17498,N_17575);
or U17613 (N_17613,N_17478,N_17475);
and U17614 (N_17614,N_17554,N_17542);
or U17615 (N_17615,N_17500,N_17518);
nand U17616 (N_17616,N_17560,N_17510);
or U17617 (N_17617,N_17490,N_17495);
xor U17618 (N_17618,N_17527,N_17577);
nor U17619 (N_17619,N_17512,N_17553);
and U17620 (N_17620,N_17535,N_17484);
xnor U17621 (N_17621,N_17480,N_17441);
or U17622 (N_17622,N_17442,N_17597);
nor U17623 (N_17623,N_17492,N_17552);
nor U17624 (N_17624,N_17584,N_17509);
nand U17625 (N_17625,N_17549,N_17483);
or U17626 (N_17626,N_17534,N_17567);
xnor U17627 (N_17627,N_17489,N_17595);
or U17628 (N_17628,N_17596,N_17592);
and U17629 (N_17629,N_17545,N_17470);
and U17630 (N_17630,N_17586,N_17443);
xor U17631 (N_17631,N_17457,N_17486);
nand U17632 (N_17632,N_17599,N_17530);
nor U17633 (N_17633,N_17467,N_17520);
or U17634 (N_17634,N_17485,N_17481);
xnor U17635 (N_17635,N_17569,N_17466);
nor U17636 (N_17636,N_17449,N_17456);
nor U17637 (N_17637,N_17591,N_17519);
and U17638 (N_17638,N_17557,N_17462);
and U17639 (N_17639,N_17487,N_17506);
xor U17640 (N_17640,N_17562,N_17465);
and U17641 (N_17641,N_17548,N_17573);
nand U17642 (N_17642,N_17514,N_17461);
and U17643 (N_17643,N_17440,N_17587);
xnor U17644 (N_17644,N_17521,N_17479);
nor U17645 (N_17645,N_17588,N_17539);
nand U17646 (N_17646,N_17544,N_17532);
and U17647 (N_17647,N_17531,N_17473);
nand U17648 (N_17648,N_17541,N_17507);
nor U17649 (N_17649,N_17476,N_17516);
and U17650 (N_17650,N_17472,N_17574);
or U17651 (N_17651,N_17555,N_17499);
and U17652 (N_17652,N_17488,N_17477);
or U17653 (N_17653,N_17558,N_17525);
nor U17654 (N_17654,N_17508,N_17452);
and U17655 (N_17655,N_17445,N_17559);
or U17656 (N_17656,N_17474,N_17523);
nand U17657 (N_17657,N_17453,N_17511);
nor U17658 (N_17658,N_17589,N_17444);
nand U17659 (N_17659,N_17446,N_17578);
or U17660 (N_17660,N_17447,N_17543);
or U17661 (N_17661,N_17566,N_17540);
xnor U17662 (N_17662,N_17547,N_17469);
nor U17663 (N_17663,N_17463,N_17536);
and U17664 (N_17664,N_17593,N_17503);
nor U17665 (N_17665,N_17571,N_17537);
nor U17666 (N_17666,N_17502,N_17524);
nand U17667 (N_17667,N_17572,N_17561);
nor U17668 (N_17668,N_17459,N_17451);
or U17669 (N_17669,N_17576,N_17493);
nor U17670 (N_17670,N_17565,N_17464);
or U17671 (N_17671,N_17482,N_17496);
or U17672 (N_17672,N_17590,N_17494);
nor U17673 (N_17673,N_17538,N_17505);
nand U17674 (N_17674,N_17583,N_17455);
nand U17675 (N_17675,N_17570,N_17460);
xor U17676 (N_17676,N_17513,N_17585);
nand U17677 (N_17677,N_17450,N_17556);
and U17678 (N_17678,N_17598,N_17528);
and U17679 (N_17679,N_17563,N_17497);
and U17680 (N_17680,N_17541,N_17540);
or U17681 (N_17681,N_17481,N_17473);
nor U17682 (N_17682,N_17538,N_17561);
nor U17683 (N_17683,N_17454,N_17527);
and U17684 (N_17684,N_17509,N_17596);
nor U17685 (N_17685,N_17520,N_17491);
nor U17686 (N_17686,N_17552,N_17545);
nor U17687 (N_17687,N_17518,N_17495);
or U17688 (N_17688,N_17534,N_17452);
or U17689 (N_17689,N_17551,N_17596);
xnor U17690 (N_17690,N_17534,N_17597);
xor U17691 (N_17691,N_17515,N_17523);
nand U17692 (N_17692,N_17465,N_17522);
and U17693 (N_17693,N_17577,N_17568);
nand U17694 (N_17694,N_17508,N_17454);
nor U17695 (N_17695,N_17462,N_17598);
and U17696 (N_17696,N_17542,N_17508);
nor U17697 (N_17697,N_17476,N_17490);
or U17698 (N_17698,N_17552,N_17587);
and U17699 (N_17699,N_17507,N_17504);
nand U17700 (N_17700,N_17456,N_17513);
nand U17701 (N_17701,N_17484,N_17584);
nor U17702 (N_17702,N_17552,N_17535);
nand U17703 (N_17703,N_17510,N_17499);
and U17704 (N_17704,N_17527,N_17570);
and U17705 (N_17705,N_17541,N_17498);
and U17706 (N_17706,N_17444,N_17551);
and U17707 (N_17707,N_17467,N_17443);
xor U17708 (N_17708,N_17447,N_17550);
or U17709 (N_17709,N_17450,N_17589);
or U17710 (N_17710,N_17450,N_17596);
and U17711 (N_17711,N_17500,N_17503);
nand U17712 (N_17712,N_17476,N_17474);
nand U17713 (N_17713,N_17503,N_17455);
and U17714 (N_17714,N_17526,N_17484);
or U17715 (N_17715,N_17589,N_17510);
nand U17716 (N_17716,N_17444,N_17597);
nand U17717 (N_17717,N_17506,N_17455);
xor U17718 (N_17718,N_17550,N_17455);
or U17719 (N_17719,N_17451,N_17464);
xor U17720 (N_17720,N_17484,N_17527);
and U17721 (N_17721,N_17502,N_17478);
nor U17722 (N_17722,N_17569,N_17586);
nor U17723 (N_17723,N_17599,N_17548);
or U17724 (N_17724,N_17580,N_17555);
nand U17725 (N_17725,N_17496,N_17468);
and U17726 (N_17726,N_17456,N_17448);
or U17727 (N_17727,N_17512,N_17454);
and U17728 (N_17728,N_17493,N_17537);
nor U17729 (N_17729,N_17531,N_17499);
nor U17730 (N_17730,N_17592,N_17480);
or U17731 (N_17731,N_17454,N_17583);
nand U17732 (N_17732,N_17444,N_17494);
nor U17733 (N_17733,N_17440,N_17466);
and U17734 (N_17734,N_17451,N_17448);
or U17735 (N_17735,N_17565,N_17476);
xnor U17736 (N_17736,N_17507,N_17499);
or U17737 (N_17737,N_17575,N_17584);
or U17738 (N_17738,N_17521,N_17465);
or U17739 (N_17739,N_17466,N_17448);
or U17740 (N_17740,N_17522,N_17590);
nor U17741 (N_17741,N_17579,N_17446);
nor U17742 (N_17742,N_17528,N_17578);
or U17743 (N_17743,N_17464,N_17556);
and U17744 (N_17744,N_17461,N_17478);
nor U17745 (N_17745,N_17541,N_17564);
nand U17746 (N_17746,N_17499,N_17473);
nor U17747 (N_17747,N_17504,N_17584);
or U17748 (N_17748,N_17531,N_17528);
and U17749 (N_17749,N_17483,N_17523);
nor U17750 (N_17750,N_17585,N_17485);
and U17751 (N_17751,N_17551,N_17469);
nor U17752 (N_17752,N_17565,N_17590);
nor U17753 (N_17753,N_17551,N_17518);
or U17754 (N_17754,N_17584,N_17581);
xnor U17755 (N_17755,N_17509,N_17580);
nand U17756 (N_17756,N_17595,N_17565);
nor U17757 (N_17757,N_17481,N_17451);
and U17758 (N_17758,N_17448,N_17446);
or U17759 (N_17759,N_17502,N_17595);
and U17760 (N_17760,N_17604,N_17616);
nand U17761 (N_17761,N_17655,N_17685);
and U17762 (N_17762,N_17610,N_17658);
or U17763 (N_17763,N_17715,N_17719);
or U17764 (N_17764,N_17710,N_17723);
or U17765 (N_17765,N_17619,N_17670);
nand U17766 (N_17766,N_17759,N_17611);
and U17767 (N_17767,N_17735,N_17635);
xor U17768 (N_17768,N_17712,N_17628);
nor U17769 (N_17769,N_17743,N_17681);
nor U17770 (N_17770,N_17623,N_17713);
nand U17771 (N_17771,N_17736,N_17705);
and U17772 (N_17772,N_17640,N_17684);
nor U17773 (N_17773,N_17674,N_17652);
nor U17774 (N_17774,N_17607,N_17672);
xnor U17775 (N_17775,N_17663,N_17608);
and U17776 (N_17776,N_17660,N_17673);
or U17777 (N_17777,N_17682,N_17615);
or U17778 (N_17778,N_17744,N_17679);
nor U17779 (N_17779,N_17707,N_17637);
nor U17780 (N_17780,N_17742,N_17677);
nand U17781 (N_17781,N_17714,N_17751);
nand U17782 (N_17782,N_17621,N_17692);
nor U17783 (N_17783,N_17702,N_17749);
nand U17784 (N_17784,N_17666,N_17727);
or U17785 (N_17785,N_17728,N_17624);
nand U17786 (N_17786,N_17617,N_17643);
nand U17787 (N_17787,N_17746,N_17739);
nor U17788 (N_17788,N_17647,N_17694);
or U17789 (N_17789,N_17745,N_17734);
or U17790 (N_17790,N_17696,N_17612);
nand U17791 (N_17791,N_17693,N_17691);
nand U17792 (N_17792,N_17717,N_17718);
nand U17793 (N_17793,N_17758,N_17730);
and U17794 (N_17794,N_17689,N_17667);
and U17795 (N_17795,N_17625,N_17644);
xnor U17796 (N_17796,N_17669,N_17676);
nor U17797 (N_17797,N_17731,N_17662);
nand U17798 (N_17798,N_17645,N_17722);
and U17799 (N_17799,N_17729,N_17750);
or U17800 (N_17800,N_17600,N_17650);
or U17801 (N_17801,N_17738,N_17683);
nand U17802 (N_17802,N_17701,N_17602);
nand U17803 (N_17803,N_17695,N_17726);
xnor U17804 (N_17804,N_17630,N_17627);
nor U17805 (N_17805,N_17639,N_17646);
nor U17806 (N_17806,N_17747,N_17706);
or U17807 (N_17807,N_17724,N_17687);
xnor U17808 (N_17808,N_17649,N_17641);
nor U17809 (N_17809,N_17620,N_17653);
and U17810 (N_17810,N_17698,N_17757);
and U17811 (N_17811,N_17680,N_17725);
nand U17812 (N_17812,N_17618,N_17675);
nand U17813 (N_17813,N_17638,N_17711);
nor U17814 (N_17814,N_17664,N_17697);
xnor U17815 (N_17815,N_17678,N_17651);
or U17816 (N_17816,N_17752,N_17632);
nor U17817 (N_17817,N_17606,N_17631);
nand U17818 (N_17818,N_17659,N_17657);
nor U17819 (N_17819,N_17613,N_17690);
and U17820 (N_17820,N_17629,N_17648);
or U17821 (N_17821,N_17634,N_17756);
or U17822 (N_17822,N_17733,N_17741);
nand U17823 (N_17823,N_17703,N_17626);
nor U17824 (N_17824,N_17665,N_17753);
nand U17825 (N_17825,N_17688,N_17614);
nand U17826 (N_17826,N_17636,N_17603);
and U17827 (N_17827,N_17700,N_17686);
or U17828 (N_17828,N_17609,N_17754);
and U17829 (N_17829,N_17668,N_17661);
or U17830 (N_17830,N_17748,N_17732);
nor U17831 (N_17831,N_17601,N_17740);
or U17832 (N_17832,N_17671,N_17605);
and U17833 (N_17833,N_17755,N_17654);
nor U17834 (N_17834,N_17721,N_17699);
xnor U17835 (N_17835,N_17709,N_17622);
nand U17836 (N_17836,N_17737,N_17704);
and U17837 (N_17837,N_17716,N_17708);
nor U17838 (N_17838,N_17633,N_17656);
nand U17839 (N_17839,N_17720,N_17642);
or U17840 (N_17840,N_17717,N_17641);
xnor U17841 (N_17841,N_17728,N_17745);
nand U17842 (N_17842,N_17740,N_17673);
and U17843 (N_17843,N_17716,N_17713);
or U17844 (N_17844,N_17754,N_17630);
nor U17845 (N_17845,N_17669,N_17705);
nand U17846 (N_17846,N_17602,N_17695);
nor U17847 (N_17847,N_17697,N_17731);
nand U17848 (N_17848,N_17625,N_17650);
nand U17849 (N_17849,N_17718,N_17699);
nor U17850 (N_17850,N_17715,N_17658);
and U17851 (N_17851,N_17621,N_17699);
nand U17852 (N_17852,N_17602,N_17757);
nand U17853 (N_17853,N_17628,N_17684);
nor U17854 (N_17854,N_17749,N_17708);
or U17855 (N_17855,N_17705,N_17602);
nand U17856 (N_17856,N_17719,N_17757);
and U17857 (N_17857,N_17601,N_17703);
and U17858 (N_17858,N_17658,N_17698);
xor U17859 (N_17859,N_17701,N_17754);
and U17860 (N_17860,N_17637,N_17737);
nand U17861 (N_17861,N_17620,N_17688);
xor U17862 (N_17862,N_17677,N_17702);
or U17863 (N_17863,N_17649,N_17655);
xnor U17864 (N_17864,N_17721,N_17684);
or U17865 (N_17865,N_17650,N_17736);
and U17866 (N_17866,N_17701,N_17756);
or U17867 (N_17867,N_17677,N_17657);
or U17868 (N_17868,N_17755,N_17615);
and U17869 (N_17869,N_17638,N_17673);
nand U17870 (N_17870,N_17603,N_17704);
or U17871 (N_17871,N_17630,N_17667);
nor U17872 (N_17872,N_17725,N_17654);
nand U17873 (N_17873,N_17638,N_17728);
nand U17874 (N_17874,N_17755,N_17736);
nor U17875 (N_17875,N_17639,N_17608);
nand U17876 (N_17876,N_17731,N_17644);
nand U17877 (N_17877,N_17692,N_17607);
nor U17878 (N_17878,N_17653,N_17742);
nor U17879 (N_17879,N_17683,N_17724);
nand U17880 (N_17880,N_17614,N_17674);
or U17881 (N_17881,N_17613,N_17758);
nand U17882 (N_17882,N_17639,N_17604);
or U17883 (N_17883,N_17669,N_17636);
and U17884 (N_17884,N_17661,N_17731);
or U17885 (N_17885,N_17718,N_17643);
nor U17886 (N_17886,N_17703,N_17753);
xnor U17887 (N_17887,N_17699,N_17636);
nor U17888 (N_17888,N_17644,N_17752);
nor U17889 (N_17889,N_17628,N_17743);
nand U17890 (N_17890,N_17680,N_17676);
or U17891 (N_17891,N_17670,N_17631);
nand U17892 (N_17892,N_17649,N_17746);
and U17893 (N_17893,N_17725,N_17753);
nand U17894 (N_17894,N_17690,N_17650);
or U17895 (N_17895,N_17624,N_17646);
xor U17896 (N_17896,N_17717,N_17614);
or U17897 (N_17897,N_17638,N_17717);
or U17898 (N_17898,N_17736,N_17753);
and U17899 (N_17899,N_17736,N_17751);
and U17900 (N_17900,N_17678,N_17693);
nand U17901 (N_17901,N_17617,N_17685);
nor U17902 (N_17902,N_17724,N_17643);
nand U17903 (N_17903,N_17719,N_17667);
nor U17904 (N_17904,N_17682,N_17621);
and U17905 (N_17905,N_17645,N_17735);
nor U17906 (N_17906,N_17649,N_17627);
nand U17907 (N_17907,N_17640,N_17697);
nor U17908 (N_17908,N_17710,N_17717);
or U17909 (N_17909,N_17693,N_17719);
or U17910 (N_17910,N_17727,N_17614);
nor U17911 (N_17911,N_17695,N_17733);
nand U17912 (N_17912,N_17714,N_17644);
nor U17913 (N_17913,N_17613,N_17673);
nor U17914 (N_17914,N_17627,N_17736);
nor U17915 (N_17915,N_17703,N_17693);
nand U17916 (N_17916,N_17751,N_17631);
nor U17917 (N_17917,N_17737,N_17735);
or U17918 (N_17918,N_17756,N_17711);
nand U17919 (N_17919,N_17674,N_17703);
xor U17920 (N_17920,N_17871,N_17803);
xnor U17921 (N_17921,N_17900,N_17858);
xor U17922 (N_17922,N_17830,N_17798);
xnor U17923 (N_17923,N_17856,N_17776);
nor U17924 (N_17924,N_17885,N_17851);
nand U17925 (N_17925,N_17883,N_17904);
and U17926 (N_17926,N_17810,N_17905);
nand U17927 (N_17927,N_17818,N_17799);
or U17928 (N_17928,N_17865,N_17783);
and U17929 (N_17929,N_17822,N_17850);
nor U17930 (N_17930,N_17910,N_17895);
xor U17931 (N_17931,N_17886,N_17864);
or U17932 (N_17932,N_17764,N_17857);
nand U17933 (N_17933,N_17828,N_17877);
nand U17934 (N_17934,N_17805,N_17890);
nand U17935 (N_17935,N_17908,N_17911);
nor U17936 (N_17936,N_17785,N_17863);
and U17937 (N_17937,N_17898,N_17846);
nor U17938 (N_17938,N_17889,N_17887);
and U17939 (N_17939,N_17913,N_17762);
or U17940 (N_17940,N_17795,N_17876);
xor U17941 (N_17941,N_17859,N_17845);
nor U17942 (N_17942,N_17832,N_17809);
nand U17943 (N_17943,N_17769,N_17834);
nand U17944 (N_17944,N_17773,N_17820);
nand U17945 (N_17945,N_17881,N_17804);
xnor U17946 (N_17946,N_17918,N_17782);
nor U17947 (N_17947,N_17796,N_17853);
and U17948 (N_17948,N_17878,N_17872);
nand U17949 (N_17949,N_17867,N_17766);
nor U17950 (N_17950,N_17844,N_17812);
nor U17951 (N_17951,N_17774,N_17793);
nor U17952 (N_17952,N_17847,N_17914);
nand U17953 (N_17953,N_17888,N_17906);
or U17954 (N_17954,N_17891,N_17816);
nor U17955 (N_17955,N_17879,N_17814);
or U17956 (N_17956,N_17824,N_17896);
nor U17957 (N_17957,N_17835,N_17842);
or U17958 (N_17958,N_17868,N_17790);
and U17959 (N_17959,N_17817,N_17841);
nor U17960 (N_17960,N_17772,N_17915);
and U17961 (N_17961,N_17806,N_17848);
or U17962 (N_17962,N_17843,N_17909);
nand U17963 (N_17963,N_17781,N_17839);
or U17964 (N_17964,N_17778,N_17775);
and U17965 (N_17965,N_17899,N_17849);
nor U17966 (N_17966,N_17760,N_17791);
and U17967 (N_17967,N_17784,N_17902);
nand U17968 (N_17968,N_17855,N_17852);
nand U17969 (N_17969,N_17768,N_17763);
nor U17970 (N_17970,N_17894,N_17837);
and U17971 (N_17971,N_17815,N_17821);
nand U17972 (N_17972,N_17771,N_17780);
nor U17973 (N_17973,N_17819,N_17892);
or U17974 (N_17974,N_17912,N_17807);
nor U17975 (N_17975,N_17767,N_17802);
or U17976 (N_17976,N_17823,N_17875);
nand U17977 (N_17977,N_17840,N_17893);
or U17978 (N_17978,N_17811,N_17861);
or U17979 (N_17979,N_17869,N_17825);
nand U17980 (N_17980,N_17903,N_17789);
nor U17981 (N_17981,N_17833,N_17882);
and U17982 (N_17982,N_17860,N_17800);
and U17983 (N_17983,N_17916,N_17813);
nand U17984 (N_17984,N_17907,N_17770);
or U17985 (N_17985,N_17777,N_17884);
and U17986 (N_17986,N_17779,N_17901);
and U17987 (N_17987,N_17797,N_17794);
and U17988 (N_17988,N_17854,N_17788);
nor U17989 (N_17989,N_17831,N_17826);
nor U17990 (N_17990,N_17870,N_17786);
nand U17991 (N_17991,N_17880,N_17836);
and U17992 (N_17992,N_17765,N_17874);
and U17993 (N_17993,N_17897,N_17919);
or U17994 (N_17994,N_17792,N_17808);
and U17995 (N_17995,N_17761,N_17787);
nand U17996 (N_17996,N_17873,N_17829);
nor U17997 (N_17997,N_17917,N_17866);
nor U17998 (N_17998,N_17801,N_17838);
nor U17999 (N_17999,N_17827,N_17862);
or U18000 (N_18000,N_17871,N_17834);
xnor U18001 (N_18001,N_17814,N_17843);
or U18002 (N_18002,N_17829,N_17882);
xor U18003 (N_18003,N_17792,N_17844);
nor U18004 (N_18004,N_17809,N_17893);
xnor U18005 (N_18005,N_17916,N_17891);
xor U18006 (N_18006,N_17864,N_17846);
or U18007 (N_18007,N_17862,N_17845);
nand U18008 (N_18008,N_17778,N_17804);
nor U18009 (N_18009,N_17852,N_17829);
xnor U18010 (N_18010,N_17877,N_17762);
and U18011 (N_18011,N_17796,N_17919);
nor U18012 (N_18012,N_17912,N_17800);
and U18013 (N_18013,N_17851,N_17879);
nor U18014 (N_18014,N_17898,N_17800);
and U18015 (N_18015,N_17833,N_17878);
nor U18016 (N_18016,N_17863,N_17901);
and U18017 (N_18017,N_17833,N_17781);
nor U18018 (N_18018,N_17817,N_17847);
nor U18019 (N_18019,N_17864,N_17904);
nand U18020 (N_18020,N_17789,N_17763);
nor U18021 (N_18021,N_17815,N_17767);
nor U18022 (N_18022,N_17909,N_17905);
nor U18023 (N_18023,N_17771,N_17821);
xor U18024 (N_18024,N_17787,N_17807);
nor U18025 (N_18025,N_17807,N_17917);
nor U18026 (N_18026,N_17912,N_17762);
and U18027 (N_18027,N_17814,N_17825);
nor U18028 (N_18028,N_17809,N_17879);
nand U18029 (N_18029,N_17811,N_17806);
or U18030 (N_18030,N_17813,N_17840);
nand U18031 (N_18031,N_17826,N_17852);
nor U18032 (N_18032,N_17897,N_17827);
xnor U18033 (N_18033,N_17837,N_17826);
xor U18034 (N_18034,N_17788,N_17777);
nand U18035 (N_18035,N_17863,N_17797);
nand U18036 (N_18036,N_17826,N_17788);
or U18037 (N_18037,N_17902,N_17907);
nor U18038 (N_18038,N_17857,N_17782);
and U18039 (N_18039,N_17775,N_17912);
or U18040 (N_18040,N_17763,N_17782);
or U18041 (N_18041,N_17770,N_17894);
nor U18042 (N_18042,N_17881,N_17791);
or U18043 (N_18043,N_17869,N_17891);
nor U18044 (N_18044,N_17788,N_17909);
xnor U18045 (N_18045,N_17776,N_17891);
nand U18046 (N_18046,N_17762,N_17894);
or U18047 (N_18047,N_17856,N_17783);
nor U18048 (N_18048,N_17848,N_17882);
or U18049 (N_18049,N_17849,N_17812);
or U18050 (N_18050,N_17782,N_17787);
xor U18051 (N_18051,N_17826,N_17778);
and U18052 (N_18052,N_17760,N_17847);
nand U18053 (N_18053,N_17848,N_17837);
and U18054 (N_18054,N_17892,N_17813);
nand U18055 (N_18055,N_17917,N_17908);
nand U18056 (N_18056,N_17771,N_17896);
or U18057 (N_18057,N_17881,N_17872);
nor U18058 (N_18058,N_17777,N_17766);
and U18059 (N_18059,N_17877,N_17862);
or U18060 (N_18060,N_17908,N_17877);
xor U18061 (N_18061,N_17765,N_17845);
and U18062 (N_18062,N_17870,N_17783);
or U18063 (N_18063,N_17874,N_17776);
or U18064 (N_18064,N_17793,N_17762);
xor U18065 (N_18065,N_17760,N_17813);
or U18066 (N_18066,N_17830,N_17895);
nor U18067 (N_18067,N_17869,N_17892);
xnor U18068 (N_18068,N_17918,N_17786);
or U18069 (N_18069,N_17830,N_17880);
nor U18070 (N_18070,N_17803,N_17867);
and U18071 (N_18071,N_17865,N_17785);
nand U18072 (N_18072,N_17844,N_17834);
nor U18073 (N_18073,N_17830,N_17858);
and U18074 (N_18074,N_17762,N_17841);
nor U18075 (N_18075,N_17795,N_17822);
nand U18076 (N_18076,N_17822,N_17788);
and U18077 (N_18077,N_17891,N_17770);
or U18078 (N_18078,N_17858,N_17904);
nor U18079 (N_18079,N_17852,N_17878);
xnor U18080 (N_18080,N_18049,N_18027);
nor U18081 (N_18081,N_17922,N_17989);
and U18082 (N_18082,N_18003,N_18059);
and U18083 (N_18083,N_18021,N_18035);
and U18084 (N_18084,N_17943,N_17968);
and U18085 (N_18085,N_18053,N_17938);
nor U18086 (N_18086,N_18078,N_17973);
or U18087 (N_18087,N_18055,N_18045);
nor U18088 (N_18088,N_18013,N_17987);
and U18089 (N_18089,N_17928,N_18073);
or U18090 (N_18090,N_18034,N_18040);
or U18091 (N_18091,N_18006,N_17983);
or U18092 (N_18092,N_18041,N_18039);
nor U18093 (N_18093,N_17966,N_17942);
or U18094 (N_18094,N_17986,N_18075);
and U18095 (N_18095,N_17945,N_18016);
and U18096 (N_18096,N_18033,N_18029);
or U18097 (N_18097,N_18015,N_17949);
and U18098 (N_18098,N_17971,N_18010);
or U18099 (N_18099,N_17932,N_18077);
xor U18100 (N_18100,N_17990,N_17994);
or U18101 (N_18101,N_17924,N_18048);
xor U18102 (N_18102,N_17936,N_17930);
and U18103 (N_18103,N_18028,N_18000);
or U18104 (N_18104,N_18023,N_17927);
and U18105 (N_18105,N_18038,N_17929);
or U18106 (N_18106,N_17925,N_18019);
and U18107 (N_18107,N_17933,N_18012);
nand U18108 (N_18108,N_17955,N_18071);
nor U18109 (N_18109,N_17962,N_18067);
nor U18110 (N_18110,N_18069,N_17976);
or U18111 (N_18111,N_18056,N_17965);
nor U18112 (N_18112,N_18072,N_17982);
and U18113 (N_18113,N_18026,N_17940);
nor U18114 (N_18114,N_17985,N_17920);
nand U18115 (N_18115,N_17984,N_17934);
or U18116 (N_18116,N_18024,N_17923);
or U18117 (N_18117,N_18042,N_17958);
nor U18118 (N_18118,N_17997,N_18009);
and U18119 (N_18119,N_17956,N_17993);
nor U18120 (N_18120,N_18068,N_18002);
or U18121 (N_18121,N_18007,N_18062);
or U18122 (N_18122,N_18001,N_18052);
nand U18123 (N_18123,N_17939,N_17941);
nor U18124 (N_18124,N_18011,N_17954);
and U18125 (N_18125,N_17950,N_17946);
nor U18126 (N_18126,N_17964,N_18022);
nand U18127 (N_18127,N_18044,N_17944);
xnor U18128 (N_18128,N_17935,N_17975);
and U18129 (N_18129,N_17988,N_18058);
or U18130 (N_18130,N_17948,N_18008);
or U18131 (N_18131,N_17951,N_18061);
or U18132 (N_18132,N_17992,N_17967);
nand U18133 (N_18133,N_18025,N_18066);
and U18134 (N_18134,N_17981,N_17998);
and U18135 (N_18135,N_18031,N_18064);
xor U18136 (N_18136,N_18004,N_17974);
or U18137 (N_18137,N_17996,N_17957);
xor U18138 (N_18138,N_17972,N_17979);
or U18139 (N_18139,N_18020,N_18036);
xor U18140 (N_18140,N_17995,N_17947);
nand U18141 (N_18141,N_17959,N_18030);
nor U18142 (N_18142,N_17952,N_17980);
nor U18143 (N_18143,N_17999,N_18046);
or U18144 (N_18144,N_18054,N_18063);
xnor U18145 (N_18145,N_18079,N_18065);
or U18146 (N_18146,N_17960,N_17963);
or U18147 (N_18147,N_17970,N_18060);
nor U18148 (N_18148,N_18037,N_17977);
or U18149 (N_18149,N_17969,N_18057);
or U18150 (N_18150,N_17953,N_18076);
and U18151 (N_18151,N_18017,N_18043);
nand U18152 (N_18152,N_18047,N_17921);
xnor U18153 (N_18153,N_18070,N_17931);
nand U18154 (N_18154,N_17937,N_18074);
xor U18155 (N_18155,N_17926,N_18005);
and U18156 (N_18156,N_18050,N_17991);
nor U18157 (N_18157,N_18051,N_18032);
nand U18158 (N_18158,N_17978,N_18014);
and U18159 (N_18159,N_17961,N_18018);
and U18160 (N_18160,N_17981,N_18044);
or U18161 (N_18161,N_18003,N_18041);
nand U18162 (N_18162,N_18009,N_17944);
xnor U18163 (N_18163,N_18077,N_18063);
and U18164 (N_18164,N_17999,N_18029);
nor U18165 (N_18165,N_17974,N_17922);
nand U18166 (N_18166,N_17942,N_18017);
xnor U18167 (N_18167,N_17928,N_17974);
nand U18168 (N_18168,N_18046,N_17922);
or U18169 (N_18169,N_18036,N_18040);
nand U18170 (N_18170,N_18052,N_18064);
and U18171 (N_18171,N_17993,N_17947);
or U18172 (N_18172,N_18014,N_18052);
and U18173 (N_18173,N_17969,N_18050);
nor U18174 (N_18174,N_17975,N_17921);
nor U18175 (N_18175,N_18041,N_17995);
and U18176 (N_18176,N_17976,N_17996);
or U18177 (N_18177,N_17970,N_17949);
nand U18178 (N_18178,N_17966,N_18033);
nand U18179 (N_18179,N_17975,N_18066);
xor U18180 (N_18180,N_17956,N_18020);
and U18181 (N_18181,N_18054,N_18078);
xnor U18182 (N_18182,N_18062,N_17967);
or U18183 (N_18183,N_17968,N_18007);
nand U18184 (N_18184,N_18049,N_17926);
or U18185 (N_18185,N_17933,N_18046);
xor U18186 (N_18186,N_18052,N_18063);
or U18187 (N_18187,N_17950,N_17981);
or U18188 (N_18188,N_18000,N_18002);
and U18189 (N_18189,N_18055,N_17971);
nand U18190 (N_18190,N_18050,N_17974);
and U18191 (N_18191,N_17935,N_17939);
or U18192 (N_18192,N_18071,N_18051);
xnor U18193 (N_18193,N_17990,N_18070);
nor U18194 (N_18194,N_18054,N_18016);
and U18195 (N_18195,N_17954,N_17950);
nor U18196 (N_18196,N_18028,N_17977);
and U18197 (N_18197,N_17979,N_17934);
nor U18198 (N_18198,N_17951,N_17959);
or U18199 (N_18199,N_17946,N_18003);
and U18200 (N_18200,N_18026,N_17932);
xnor U18201 (N_18201,N_17966,N_18073);
nand U18202 (N_18202,N_17994,N_17921);
and U18203 (N_18203,N_18071,N_17947);
and U18204 (N_18204,N_17955,N_18063);
and U18205 (N_18205,N_17926,N_18010);
xor U18206 (N_18206,N_18057,N_17945);
and U18207 (N_18207,N_18026,N_17924);
nor U18208 (N_18208,N_17965,N_17940);
or U18209 (N_18209,N_17934,N_17975);
nand U18210 (N_18210,N_18021,N_17971);
and U18211 (N_18211,N_18073,N_18003);
and U18212 (N_18212,N_18025,N_17983);
nand U18213 (N_18213,N_17940,N_17968);
nor U18214 (N_18214,N_18035,N_17993);
nand U18215 (N_18215,N_18037,N_17973);
xnor U18216 (N_18216,N_17984,N_18032);
nor U18217 (N_18217,N_17927,N_18072);
and U18218 (N_18218,N_17934,N_17976);
nor U18219 (N_18219,N_18040,N_17950);
nor U18220 (N_18220,N_18060,N_17929);
and U18221 (N_18221,N_18025,N_18078);
nor U18222 (N_18222,N_17994,N_18056);
nor U18223 (N_18223,N_17953,N_17965);
nor U18224 (N_18224,N_17999,N_18023);
and U18225 (N_18225,N_17992,N_17996);
nor U18226 (N_18226,N_17943,N_18009);
and U18227 (N_18227,N_17961,N_17921);
nor U18228 (N_18228,N_18055,N_18002);
and U18229 (N_18229,N_18071,N_17954);
nand U18230 (N_18230,N_17967,N_17978);
and U18231 (N_18231,N_17995,N_17966);
nand U18232 (N_18232,N_17988,N_18059);
nor U18233 (N_18233,N_18040,N_18064);
or U18234 (N_18234,N_17923,N_18050);
nand U18235 (N_18235,N_17997,N_18017);
and U18236 (N_18236,N_17931,N_18014);
nor U18237 (N_18237,N_18025,N_18002);
nand U18238 (N_18238,N_17987,N_18068);
nand U18239 (N_18239,N_18069,N_18060);
or U18240 (N_18240,N_18178,N_18173);
xnor U18241 (N_18241,N_18146,N_18193);
nand U18242 (N_18242,N_18150,N_18199);
and U18243 (N_18243,N_18155,N_18153);
or U18244 (N_18244,N_18096,N_18165);
or U18245 (N_18245,N_18128,N_18167);
nand U18246 (N_18246,N_18124,N_18100);
xor U18247 (N_18247,N_18162,N_18123);
and U18248 (N_18248,N_18111,N_18149);
nor U18249 (N_18249,N_18105,N_18235);
and U18250 (N_18250,N_18122,N_18188);
or U18251 (N_18251,N_18103,N_18210);
and U18252 (N_18252,N_18177,N_18216);
nor U18253 (N_18253,N_18197,N_18098);
xor U18254 (N_18254,N_18211,N_18109);
nand U18255 (N_18255,N_18179,N_18175);
and U18256 (N_18256,N_18104,N_18114);
nor U18257 (N_18257,N_18182,N_18130);
and U18258 (N_18258,N_18201,N_18190);
or U18259 (N_18259,N_18081,N_18170);
nand U18260 (N_18260,N_18160,N_18168);
nand U18261 (N_18261,N_18234,N_18184);
xor U18262 (N_18262,N_18126,N_18135);
nand U18263 (N_18263,N_18140,N_18231);
nand U18264 (N_18264,N_18089,N_18110);
nand U18265 (N_18265,N_18106,N_18120);
nand U18266 (N_18266,N_18176,N_18091);
or U18267 (N_18267,N_18136,N_18181);
nand U18268 (N_18268,N_18218,N_18097);
nand U18269 (N_18269,N_18239,N_18185);
nor U18270 (N_18270,N_18230,N_18151);
nor U18271 (N_18271,N_18093,N_18205);
or U18272 (N_18272,N_18137,N_18186);
or U18273 (N_18273,N_18159,N_18166);
or U18274 (N_18274,N_18192,N_18119);
and U18275 (N_18275,N_18116,N_18219);
nand U18276 (N_18276,N_18198,N_18132);
or U18277 (N_18277,N_18236,N_18115);
or U18278 (N_18278,N_18131,N_18206);
nor U18279 (N_18279,N_18129,N_18221);
or U18280 (N_18280,N_18214,N_18134);
xor U18281 (N_18281,N_18156,N_18112);
nor U18282 (N_18282,N_18090,N_18147);
xor U18283 (N_18283,N_18215,N_18092);
or U18284 (N_18284,N_18208,N_18087);
or U18285 (N_18285,N_18187,N_18200);
xor U18286 (N_18286,N_18095,N_18172);
or U18287 (N_18287,N_18083,N_18174);
nor U18288 (N_18288,N_18225,N_18094);
and U18289 (N_18289,N_18194,N_18113);
nand U18290 (N_18290,N_18191,N_18080);
or U18291 (N_18291,N_18227,N_18161);
or U18292 (N_18292,N_18169,N_18144);
nor U18293 (N_18293,N_18145,N_18183);
or U18294 (N_18294,N_18127,N_18139);
nand U18295 (N_18295,N_18148,N_18118);
nand U18296 (N_18296,N_18088,N_18202);
nand U18297 (N_18297,N_18099,N_18158);
or U18298 (N_18298,N_18082,N_18143);
or U18299 (N_18299,N_18180,N_18222);
or U18300 (N_18300,N_18121,N_18203);
and U18301 (N_18301,N_18212,N_18085);
or U18302 (N_18302,N_18195,N_18224);
nand U18303 (N_18303,N_18107,N_18141);
nor U18304 (N_18304,N_18152,N_18209);
nand U18305 (N_18305,N_18217,N_18220);
xnor U18306 (N_18306,N_18226,N_18204);
or U18307 (N_18307,N_18142,N_18228);
nand U18308 (N_18308,N_18086,N_18102);
xor U18309 (N_18309,N_18084,N_18163);
nand U18310 (N_18310,N_18229,N_18233);
and U18311 (N_18311,N_18223,N_18138);
nor U18312 (N_18312,N_18154,N_18125);
and U18313 (N_18313,N_18108,N_18133);
nor U18314 (N_18314,N_18237,N_18232);
or U18315 (N_18315,N_18213,N_18189);
nand U18316 (N_18316,N_18238,N_18164);
and U18317 (N_18317,N_18101,N_18171);
xor U18318 (N_18318,N_18157,N_18196);
and U18319 (N_18319,N_18117,N_18207);
nand U18320 (N_18320,N_18204,N_18152);
nand U18321 (N_18321,N_18221,N_18227);
nor U18322 (N_18322,N_18092,N_18134);
or U18323 (N_18323,N_18113,N_18158);
nor U18324 (N_18324,N_18219,N_18181);
xor U18325 (N_18325,N_18182,N_18186);
or U18326 (N_18326,N_18099,N_18081);
or U18327 (N_18327,N_18199,N_18113);
nand U18328 (N_18328,N_18119,N_18209);
xnor U18329 (N_18329,N_18214,N_18199);
or U18330 (N_18330,N_18205,N_18145);
xnor U18331 (N_18331,N_18123,N_18125);
xor U18332 (N_18332,N_18199,N_18188);
and U18333 (N_18333,N_18172,N_18132);
nand U18334 (N_18334,N_18210,N_18117);
or U18335 (N_18335,N_18150,N_18093);
and U18336 (N_18336,N_18095,N_18194);
or U18337 (N_18337,N_18160,N_18115);
and U18338 (N_18338,N_18160,N_18109);
nor U18339 (N_18339,N_18112,N_18096);
or U18340 (N_18340,N_18178,N_18097);
and U18341 (N_18341,N_18185,N_18197);
and U18342 (N_18342,N_18118,N_18125);
nand U18343 (N_18343,N_18191,N_18116);
and U18344 (N_18344,N_18230,N_18092);
nor U18345 (N_18345,N_18228,N_18081);
or U18346 (N_18346,N_18222,N_18201);
xnor U18347 (N_18347,N_18131,N_18151);
xnor U18348 (N_18348,N_18174,N_18140);
or U18349 (N_18349,N_18119,N_18140);
and U18350 (N_18350,N_18119,N_18236);
nor U18351 (N_18351,N_18165,N_18159);
xor U18352 (N_18352,N_18102,N_18221);
or U18353 (N_18353,N_18117,N_18121);
nand U18354 (N_18354,N_18238,N_18113);
nor U18355 (N_18355,N_18239,N_18140);
and U18356 (N_18356,N_18131,N_18162);
or U18357 (N_18357,N_18182,N_18232);
and U18358 (N_18358,N_18143,N_18170);
and U18359 (N_18359,N_18235,N_18215);
xnor U18360 (N_18360,N_18124,N_18175);
or U18361 (N_18361,N_18134,N_18202);
nor U18362 (N_18362,N_18170,N_18121);
or U18363 (N_18363,N_18156,N_18202);
nand U18364 (N_18364,N_18112,N_18154);
or U18365 (N_18365,N_18143,N_18146);
or U18366 (N_18366,N_18187,N_18198);
and U18367 (N_18367,N_18120,N_18082);
and U18368 (N_18368,N_18208,N_18145);
nor U18369 (N_18369,N_18093,N_18158);
or U18370 (N_18370,N_18186,N_18189);
nand U18371 (N_18371,N_18175,N_18188);
nor U18372 (N_18372,N_18239,N_18166);
or U18373 (N_18373,N_18231,N_18236);
nand U18374 (N_18374,N_18173,N_18116);
or U18375 (N_18375,N_18165,N_18195);
nand U18376 (N_18376,N_18216,N_18126);
xnor U18377 (N_18377,N_18119,N_18080);
nand U18378 (N_18378,N_18200,N_18111);
nand U18379 (N_18379,N_18086,N_18207);
nand U18380 (N_18380,N_18136,N_18125);
and U18381 (N_18381,N_18181,N_18097);
xor U18382 (N_18382,N_18152,N_18234);
nor U18383 (N_18383,N_18132,N_18185);
or U18384 (N_18384,N_18159,N_18202);
nor U18385 (N_18385,N_18130,N_18097);
nor U18386 (N_18386,N_18195,N_18132);
nand U18387 (N_18387,N_18211,N_18210);
nand U18388 (N_18388,N_18216,N_18167);
and U18389 (N_18389,N_18104,N_18221);
nor U18390 (N_18390,N_18197,N_18128);
and U18391 (N_18391,N_18226,N_18083);
xor U18392 (N_18392,N_18222,N_18152);
nor U18393 (N_18393,N_18172,N_18199);
and U18394 (N_18394,N_18137,N_18173);
or U18395 (N_18395,N_18119,N_18155);
and U18396 (N_18396,N_18164,N_18223);
and U18397 (N_18397,N_18203,N_18188);
nor U18398 (N_18398,N_18136,N_18174);
xnor U18399 (N_18399,N_18087,N_18102);
or U18400 (N_18400,N_18248,N_18268);
and U18401 (N_18401,N_18254,N_18335);
nand U18402 (N_18402,N_18368,N_18247);
or U18403 (N_18403,N_18243,N_18296);
nor U18404 (N_18404,N_18287,N_18285);
and U18405 (N_18405,N_18306,N_18379);
nor U18406 (N_18406,N_18371,N_18342);
and U18407 (N_18407,N_18338,N_18341);
nor U18408 (N_18408,N_18277,N_18264);
and U18409 (N_18409,N_18383,N_18299);
nor U18410 (N_18410,N_18259,N_18369);
and U18411 (N_18411,N_18298,N_18331);
nor U18412 (N_18412,N_18286,N_18290);
nor U18413 (N_18413,N_18289,N_18275);
nor U18414 (N_18414,N_18387,N_18326);
xor U18415 (N_18415,N_18263,N_18359);
nor U18416 (N_18416,N_18318,N_18303);
or U18417 (N_18417,N_18399,N_18271);
nand U18418 (N_18418,N_18283,N_18255);
and U18419 (N_18419,N_18280,N_18385);
nor U18420 (N_18420,N_18324,N_18334);
nor U18421 (N_18421,N_18391,N_18281);
or U18422 (N_18422,N_18282,N_18313);
and U18423 (N_18423,N_18328,N_18362);
nand U18424 (N_18424,N_18396,N_18310);
xnor U18425 (N_18425,N_18261,N_18312);
nor U18426 (N_18426,N_18376,N_18392);
nand U18427 (N_18427,N_18244,N_18314);
nand U18428 (N_18428,N_18241,N_18357);
or U18429 (N_18429,N_18294,N_18355);
and U18430 (N_18430,N_18364,N_18257);
nand U18431 (N_18431,N_18378,N_18323);
and U18432 (N_18432,N_18301,N_18339);
nor U18433 (N_18433,N_18384,N_18363);
xnor U18434 (N_18434,N_18380,N_18388);
and U18435 (N_18435,N_18272,N_18386);
or U18436 (N_18436,N_18278,N_18373);
and U18437 (N_18437,N_18375,N_18381);
nor U18438 (N_18438,N_18293,N_18353);
nor U18439 (N_18439,N_18309,N_18398);
and U18440 (N_18440,N_18350,N_18333);
or U18441 (N_18441,N_18307,N_18395);
or U18442 (N_18442,N_18343,N_18377);
nor U18443 (N_18443,N_18358,N_18394);
nor U18444 (N_18444,N_18240,N_18300);
and U18445 (N_18445,N_18346,N_18332);
xor U18446 (N_18446,N_18251,N_18365);
nor U18447 (N_18447,N_18345,N_18258);
or U18448 (N_18448,N_18325,N_18361);
xor U18449 (N_18449,N_18337,N_18389);
and U18450 (N_18450,N_18279,N_18252);
or U18451 (N_18451,N_18246,N_18321);
or U18452 (N_18452,N_18265,N_18266);
or U18453 (N_18453,N_18356,N_18330);
nand U18454 (N_18454,N_18260,N_18382);
and U18455 (N_18455,N_18311,N_18308);
nand U18456 (N_18456,N_18320,N_18245);
nor U18457 (N_18457,N_18322,N_18370);
or U18458 (N_18458,N_18295,N_18319);
nor U18459 (N_18459,N_18276,N_18249);
xnor U18460 (N_18460,N_18253,N_18367);
nor U18461 (N_18461,N_18256,N_18354);
nor U18462 (N_18462,N_18336,N_18262);
or U18463 (N_18463,N_18352,N_18344);
and U18464 (N_18464,N_18273,N_18242);
or U18465 (N_18465,N_18347,N_18270);
nand U18466 (N_18466,N_18302,N_18267);
xnor U18467 (N_18467,N_18340,N_18393);
xnor U18468 (N_18468,N_18397,N_18250);
xor U18469 (N_18469,N_18374,N_18351);
xor U18470 (N_18470,N_18390,N_18349);
xnor U18471 (N_18471,N_18304,N_18372);
nand U18472 (N_18472,N_18284,N_18288);
or U18473 (N_18473,N_18291,N_18366);
and U18474 (N_18474,N_18348,N_18292);
nor U18475 (N_18475,N_18329,N_18269);
or U18476 (N_18476,N_18327,N_18316);
and U18477 (N_18477,N_18297,N_18315);
and U18478 (N_18478,N_18305,N_18360);
nor U18479 (N_18479,N_18317,N_18274);
or U18480 (N_18480,N_18357,N_18260);
or U18481 (N_18481,N_18247,N_18337);
nand U18482 (N_18482,N_18290,N_18382);
and U18483 (N_18483,N_18352,N_18283);
or U18484 (N_18484,N_18307,N_18262);
and U18485 (N_18485,N_18281,N_18362);
nor U18486 (N_18486,N_18300,N_18315);
nor U18487 (N_18487,N_18287,N_18329);
or U18488 (N_18488,N_18368,N_18388);
and U18489 (N_18489,N_18379,N_18346);
and U18490 (N_18490,N_18243,N_18277);
xnor U18491 (N_18491,N_18244,N_18388);
nor U18492 (N_18492,N_18384,N_18308);
nor U18493 (N_18493,N_18304,N_18344);
and U18494 (N_18494,N_18377,N_18328);
or U18495 (N_18495,N_18308,N_18294);
nor U18496 (N_18496,N_18367,N_18290);
or U18497 (N_18497,N_18381,N_18285);
or U18498 (N_18498,N_18276,N_18366);
nor U18499 (N_18499,N_18341,N_18244);
nor U18500 (N_18500,N_18278,N_18308);
and U18501 (N_18501,N_18376,N_18310);
or U18502 (N_18502,N_18328,N_18295);
nor U18503 (N_18503,N_18295,N_18340);
or U18504 (N_18504,N_18367,N_18300);
nor U18505 (N_18505,N_18333,N_18373);
and U18506 (N_18506,N_18335,N_18390);
nand U18507 (N_18507,N_18379,N_18359);
or U18508 (N_18508,N_18262,N_18399);
nor U18509 (N_18509,N_18303,N_18263);
nor U18510 (N_18510,N_18292,N_18253);
nand U18511 (N_18511,N_18393,N_18269);
nand U18512 (N_18512,N_18368,N_18271);
and U18513 (N_18513,N_18342,N_18289);
nand U18514 (N_18514,N_18390,N_18317);
nor U18515 (N_18515,N_18352,N_18286);
or U18516 (N_18516,N_18297,N_18388);
and U18517 (N_18517,N_18312,N_18300);
and U18518 (N_18518,N_18317,N_18369);
and U18519 (N_18519,N_18305,N_18281);
and U18520 (N_18520,N_18316,N_18301);
or U18521 (N_18521,N_18320,N_18342);
nor U18522 (N_18522,N_18300,N_18279);
nor U18523 (N_18523,N_18249,N_18323);
nor U18524 (N_18524,N_18368,N_18326);
and U18525 (N_18525,N_18286,N_18348);
nor U18526 (N_18526,N_18291,N_18240);
or U18527 (N_18527,N_18359,N_18399);
nand U18528 (N_18528,N_18265,N_18393);
nor U18529 (N_18529,N_18313,N_18319);
and U18530 (N_18530,N_18310,N_18248);
nand U18531 (N_18531,N_18330,N_18361);
nor U18532 (N_18532,N_18317,N_18318);
and U18533 (N_18533,N_18283,N_18324);
nand U18534 (N_18534,N_18359,N_18256);
and U18535 (N_18535,N_18379,N_18391);
nor U18536 (N_18536,N_18383,N_18354);
or U18537 (N_18537,N_18313,N_18293);
nor U18538 (N_18538,N_18247,N_18374);
nand U18539 (N_18539,N_18291,N_18360);
nand U18540 (N_18540,N_18380,N_18320);
nor U18541 (N_18541,N_18273,N_18243);
nand U18542 (N_18542,N_18396,N_18254);
or U18543 (N_18543,N_18364,N_18320);
nand U18544 (N_18544,N_18312,N_18245);
nor U18545 (N_18545,N_18339,N_18324);
nand U18546 (N_18546,N_18313,N_18362);
nor U18547 (N_18547,N_18295,N_18275);
nor U18548 (N_18548,N_18390,N_18313);
nand U18549 (N_18549,N_18261,N_18314);
and U18550 (N_18550,N_18393,N_18245);
or U18551 (N_18551,N_18338,N_18395);
or U18552 (N_18552,N_18289,N_18361);
nand U18553 (N_18553,N_18329,N_18393);
nor U18554 (N_18554,N_18283,N_18350);
xnor U18555 (N_18555,N_18274,N_18393);
xnor U18556 (N_18556,N_18298,N_18360);
nor U18557 (N_18557,N_18308,N_18319);
nor U18558 (N_18558,N_18373,N_18302);
and U18559 (N_18559,N_18389,N_18318);
or U18560 (N_18560,N_18496,N_18511);
nor U18561 (N_18561,N_18558,N_18536);
xnor U18562 (N_18562,N_18482,N_18432);
and U18563 (N_18563,N_18530,N_18437);
nor U18564 (N_18564,N_18551,N_18448);
nor U18565 (N_18565,N_18419,N_18460);
xnor U18566 (N_18566,N_18475,N_18520);
and U18567 (N_18567,N_18410,N_18523);
nor U18568 (N_18568,N_18453,N_18540);
nor U18569 (N_18569,N_18491,N_18461);
nand U18570 (N_18570,N_18462,N_18521);
xnor U18571 (N_18571,N_18423,N_18512);
nor U18572 (N_18572,N_18472,N_18554);
nand U18573 (N_18573,N_18470,N_18443);
or U18574 (N_18574,N_18426,N_18434);
nor U18575 (N_18575,N_18487,N_18539);
nor U18576 (N_18576,N_18495,N_18514);
and U18577 (N_18577,N_18502,N_18499);
and U18578 (N_18578,N_18446,N_18485);
and U18579 (N_18579,N_18494,N_18500);
nor U18580 (N_18580,N_18459,N_18455);
nor U18581 (N_18581,N_18430,N_18477);
nor U18582 (N_18582,N_18409,N_18552);
or U18583 (N_18583,N_18549,N_18450);
or U18584 (N_18584,N_18407,N_18454);
nor U18585 (N_18585,N_18479,N_18559);
or U18586 (N_18586,N_18489,N_18517);
and U18587 (N_18587,N_18403,N_18401);
xor U18588 (N_18588,N_18555,N_18515);
xor U18589 (N_18589,N_18445,N_18405);
nand U18590 (N_18590,N_18447,N_18421);
nor U18591 (N_18591,N_18550,N_18457);
nand U18592 (N_18592,N_18424,N_18490);
xnor U18593 (N_18593,N_18546,N_18404);
xor U18594 (N_18594,N_18509,N_18506);
or U18595 (N_18595,N_18422,N_18471);
or U18596 (N_18596,N_18541,N_18441);
and U18597 (N_18597,N_18547,N_18466);
or U18598 (N_18598,N_18412,N_18469);
and U18599 (N_18599,N_18537,N_18474);
nand U18600 (N_18600,N_18526,N_18435);
nor U18601 (N_18601,N_18400,N_18483);
nor U18602 (N_18602,N_18532,N_18436);
or U18603 (N_18603,N_18473,N_18516);
nor U18604 (N_18604,N_18535,N_18519);
nand U18605 (N_18605,N_18406,N_18420);
nand U18606 (N_18606,N_18463,N_18525);
nor U18607 (N_18607,N_18465,N_18504);
and U18608 (N_18608,N_18542,N_18431);
nand U18609 (N_18609,N_18553,N_18497);
nand U18610 (N_18610,N_18458,N_18414);
or U18611 (N_18611,N_18545,N_18418);
nor U18612 (N_18612,N_18524,N_18478);
or U18613 (N_18613,N_18451,N_18534);
nor U18614 (N_18614,N_18501,N_18518);
nor U18615 (N_18615,N_18408,N_18527);
and U18616 (N_18616,N_18508,N_18492);
nand U18617 (N_18617,N_18510,N_18480);
nor U18618 (N_18618,N_18402,N_18449);
or U18619 (N_18619,N_18544,N_18456);
and U18620 (N_18620,N_18522,N_18415);
xnor U18621 (N_18621,N_18548,N_18425);
nand U18622 (N_18622,N_18433,N_18486);
nor U18623 (N_18623,N_18513,N_18444);
and U18624 (N_18624,N_18416,N_18543);
or U18625 (N_18625,N_18503,N_18464);
nor U18626 (N_18626,N_18531,N_18528);
and U18627 (N_18627,N_18452,N_18556);
and U18628 (N_18628,N_18429,N_18529);
nand U18629 (N_18629,N_18505,N_18440);
nand U18630 (N_18630,N_18439,N_18538);
nand U18631 (N_18631,N_18428,N_18493);
or U18632 (N_18632,N_18557,N_18488);
nand U18633 (N_18633,N_18411,N_18438);
nor U18634 (N_18634,N_18442,N_18413);
and U18635 (N_18635,N_18533,N_18427);
xnor U18636 (N_18636,N_18481,N_18417);
nand U18637 (N_18637,N_18467,N_18498);
and U18638 (N_18638,N_18507,N_18476);
or U18639 (N_18639,N_18468,N_18484);
and U18640 (N_18640,N_18516,N_18493);
and U18641 (N_18641,N_18401,N_18417);
or U18642 (N_18642,N_18403,N_18525);
or U18643 (N_18643,N_18472,N_18460);
or U18644 (N_18644,N_18465,N_18509);
xnor U18645 (N_18645,N_18400,N_18414);
or U18646 (N_18646,N_18443,N_18452);
nand U18647 (N_18647,N_18496,N_18526);
and U18648 (N_18648,N_18436,N_18484);
nand U18649 (N_18649,N_18445,N_18478);
nor U18650 (N_18650,N_18406,N_18493);
nand U18651 (N_18651,N_18427,N_18475);
and U18652 (N_18652,N_18505,N_18475);
nand U18653 (N_18653,N_18475,N_18541);
or U18654 (N_18654,N_18422,N_18405);
nand U18655 (N_18655,N_18516,N_18456);
and U18656 (N_18656,N_18504,N_18461);
or U18657 (N_18657,N_18447,N_18448);
or U18658 (N_18658,N_18466,N_18405);
xor U18659 (N_18659,N_18443,N_18481);
nand U18660 (N_18660,N_18516,N_18497);
or U18661 (N_18661,N_18521,N_18490);
nand U18662 (N_18662,N_18433,N_18536);
nor U18663 (N_18663,N_18466,N_18514);
nand U18664 (N_18664,N_18444,N_18517);
or U18665 (N_18665,N_18426,N_18454);
xor U18666 (N_18666,N_18416,N_18421);
nand U18667 (N_18667,N_18509,N_18543);
nor U18668 (N_18668,N_18421,N_18530);
nand U18669 (N_18669,N_18546,N_18490);
nor U18670 (N_18670,N_18514,N_18510);
and U18671 (N_18671,N_18430,N_18411);
and U18672 (N_18672,N_18429,N_18534);
or U18673 (N_18673,N_18532,N_18527);
nand U18674 (N_18674,N_18463,N_18501);
nand U18675 (N_18675,N_18499,N_18456);
or U18676 (N_18676,N_18429,N_18443);
nand U18677 (N_18677,N_18543,N_18469);
and U18678 (N_18678,N_18551,N_18438);
and U18679 (N_18679,N_18494,N_18444);
or U18680 (N_18680,N_18403,N_18480);
and U18681 (N_18681,N_18499,N_18442);
nand U18682 (N_18682,N_18472,N_18474);
or U18683 (N_18683,N_18415,N_18555);
nand U18684 (N_18684,N_18477,N_18439);
and U18685 (N_18685,N_18459,N_18474);
and U18686 (N_18686,N_18433,N_18483);
nand U18687 (N_18687,N_18493,N_18453);
and U18688 (N_18688,N_18545,N_18462);
nand U18689 (N_18689,N_18419,N_18544);
nor U18690 (N_18690,N_18471,N_18473);
and U18691 (N_18691,N_18472,N_18498);
xnor U18692 (N_18692,N_18454,N_18556);
or U18693 (N_18693,N_18477,N_18446);
nand U18694 (N_18694,N_18556,N_18558);
and U18695 (N_18695,N_18437,N_18554);
nor U18696 (N_18696,N_18497,N_18506);
and U18697 (N_18697,N_18479,N_18495);
xnor U18698 (N_18698,N_18499,N_18423);
nand U18699 (N_18699,N_18524,N_18423);
nor U18700 (N_18700,N_18431,N_18453);
or U18701 (N_18701,N_18470,N_18541);
nand U18702 (N_18702,N_18551,N_18541);
and U18703 (N_18703,N_18503,N_18510);
nor U18704 (N_18704,N_18524,N_18409);
nand U18705 (N_18705,N_18412,N_18510);
nor U18706 (N_18706,N_18519,N_18518);
and U18707 (N_18707,N_18538,N_18470);
nand U18708 (N_18708,N_18512,N_18470);
xor U18709 (N_18709,N_18487,N_18462);
nand U18710 (N_18710,N_18471,N_18508);
nand U18711 (N_18711,N_18458,N_18467);
and U18712 (N_18712,N_18494,N_18473);
and U18713 (N_18713,N_18436,N_18455);
or U18714 (N_18714,N_18422,N_18480);
nand U18715 (N_18715,N_18433,N_18442);
and U18716 (N_18716,N_18450,N_18497);
xnor U18717 (N_18717,N_18510,N_18482);
xnor U18718 (N_18718,N_18510,N_18465);
or U18719 (N_18719,N_18464,N_18467);
or U18720 (N_18720,N_18624,N_18665);
nor U18721 (N_18721,N_18688,N_18617);
and U18722 (N_18722,N_18631,N_18644);
nand U18723 (N_18723,N_18663,N_18671);
or U18724 (N_18724,N_18706,N_18641);
xor U18725 (N_18725,N_18656,N_18608);
nor U18726 (N_18726,N_18694,N_18611);
nand U18727 (N_18727,N_18570,N_18669);
and U18728 (N_18728,N_18576,N_18610);
and U18729 (N_18729,N_18604,N_18680);
and U18730 (N_18730,N_18698,N_18686);
xnor U18731 (N_18731,N_18649,N_18590);
or U18732 (N_18732,N_18705,N_18661);
xnor U18733 (N_18733,N_18677,N_18690);
and U18734 (N_18734,N_18629,N_18660);
and U18735 (N_18735,N_18579,N_18710);
or U18736 (N_18736,N_18685,N_18613);
xnor U18737 (N_18737,N_18683,N_18603);
nand U18738 (N_18738,N_18572,N_18560);
or U18739 (N_18739,N_18569,N_18634);
xor U18740 (N_18740,N_18582,N_18676);
or U18741 (N_18741,N_18668,N_18702);
or U18742 (N_18742,N_18609,N_18696);
or U18743 (N_18743,N_18673,N_18638);
and U18744 (N_18744,N_18714,N_18701);
nand U18745 (N_18745,N_18635,N_18692);
and U18746 (N_18746,N_18562,N_18639);
nand U18747 (N_18747,N_18623,N_18614);
nor U18748 (N_18748,N_18650,N_18647);
or U18749 (N_18749,N_18670,N_18715);
nor U18750 (N_18750,N_18672,N_18718);
or U18751 (N_18751,N_18612,N_18620);
nor U18752 (N_18752,N_18648,N_18598);
nor U18753 (N_18753,N_18607,N_18667);
nor U18754 (N_18754,N_18574,N_18713);
nor U18755 (N_18755,N_18693,N_18678);
and U18756 (N_18756,N_18584,N_18566);
nor U18757 (N_18757,N_18703,N_18616);
nand U18758 (N_18758,N_18657,N_18711);
nor U18759 (N_18759,N_18666,N_18632);
nand U18760 (N_18760,N_18597,N_18708);
nor U18761 (N_18761,N_18691,N_18712);
nor U18762 (N_18762,N_18640,N_18674);
and U18763 (N_18763,N_18687,N_18592);
nor U18764 (N_18764,N_18575,N_18605);
nor U18765 (N_18765,N_18675,N_18568);
and U18766 (N_18766,N_18580,N_18646);
nand U18767 (N_18767,N_18571,N_18626);
and U18768 (N_18768,N_18561,N_18630);
nand U18769 (N_18769,N_18606,N_18618);
nor U18770 (N_18770,N_18600,N_18636);
or U18771 (N_18771,N_18601,N_18642);
and U18772 (N_18772,N_18596,N_18587);
nand U18773 (N_18773,N_18679,N_18622);
xor U18774 (N_18774,N_18586,N_18684);
and U18775 (N_18775,N_18615,N_18578);
nand U18776 (N_18776,N_18682,N_18573);
nor U18777 (N_18777,N_18643,N_18564);
or U18778 (N_18778,N_18704,N_18577);
and U18779 (N_18779,N_18565,N_18567);
and U18780 (N_18780,N_18653,N_18581);
and U18781 (N_18781,N_18602,N_18595);
and U18782 (N_18782,N_18700,N_18716);
nand U18783 (N_18783,N_18719,N_18628);
and U18784 (N_18784,N_18697,N_18651);
nand U18785 (N_18785,N_18681,N_18619);
nor U18786 (N_18786,N_18563,N_18625);
or U18787 (N_18787,N_18621,N_18662);
and U18788 (N_18788,N_18633,N_18589);
or U18789 (N_18789,N_18717,N_18695);
and U18790 (N_18790,N_18699,N_18654);
and U18791 (N_18791,N_18594,N_18652);
and U18792 (N_18792,N_18659,N_18591);
and U18793 (N_18793,N_18583,N_18664);
or U18794 (N_18794,N_18637,N_18588);
or U18795 (N_18795,N_18627,N_18658);
or U18796 (N_18796,N_18585,N_18655);
nand U18797 (N_18797,N_18599,N_18707);
nor U18798 (N_18798,N_18709,N_18689);
or U18799 (N_18799,N_18593,N_18645);
or U18800 (N_18800,N_18684,N_18596);
and U18801 (N_18801,N_18632,N_18706);
or U18802 (N_18802,N_18570,N_18702);
nand U18803 (N_18803,N_18612,N_18689);
or U18804 (N_18804,N_18625,N_18628);
nand U18805 (N_18805,N_18694,N_18585);
nor U18806 (N_18806,N_18573,N_18697);
nor U18807 (N_18807,N_18600,N_18625);
or U18808 (N_18808,N_18560,N_18710);
nor U18809 (N_18809,N_18697,N_18564);
and U18810 (N_18810,N_18596,N_18563);
or U18811 (N_18811,N_18657,N_18599);
nor U18812 (N_18812,N_18666,N_18694);
nand U18813 (N_18813,N_18657,N_18646);
nor U18814 (N_18814,N_18568,N_18676);
nor U18815 (N_18815,N_18582,N_18572);
nor U18816 (N_18816,N_18658,N_18697);
nor U18817 (N_18817,N_18637,N_18635);
and U18818 (N_18818,N_18694,N_18628);
nand U18819 (N_18819,N_18691,N_18573);
and U18820 (N_18820,N_18602,N_18678);
nor U18821 (N_18821,N_18614,N_18682);
or U18822 (N_18822,N_18585,N_18688);
nand U18823 (N_18823,N_18718,N_18657);
nand U18824 (N_18824,N_18623,N_18595);
and U18825 (N_18825,N_18638,N_18600);
nand U18826 (N_18826,N_18706,N_18704);
or U18827 (N_18827,N_18612,N_18638);
nand U18828 (N_18828,N_18626,N_18587);
nand U18829 (N_18829,N_18579,N_18609);
nand U18830 (N_18830,N_18645,N_18585);
xnor U18831 (N_18831,N_18593,N_18717);
nor U18832 (N_18832,N_18691,N_18710);
nor U18833 (N_18833,N_18712,N_18563);
or U18834 (N_18834,N_18567,N_18679);
nor U18835 (N_18835,N_18571,N_18692);
or U18836 (N_18836,N_18578,N_18586);
nor U18837 (N_18837,N_18568,N_18663);
nor U18838 (N_18838,N_18655,N_18649);
or U18839 (N_18839,N_18658,N_18612);
and U18840 (N_18840,N_18654,N_18617);
nor U18841 (N_18841,N_18619,N_18668);
or U18842 (N_18842,N_18704,N_18591);
nor U18843 (N_18843,N_18681,N_18581);
and U18844 (N_18844,N_18672,N_18627);
and U18845 (N_18845,N_18659,N_18716);
and U18846 (N_18846,N_18668,N_18676);
and U18847 (N_18847,N_18705,N_18712);
nor U18848 (N_18848,N_18691,N_18668);
or U18849 (N_18849,N_18705,N_18568);
nor U18850 (N_18850,N_18719,N_18615);
nor U18851 (N_18851,N_18610,N_18715);
and U18852 (N_18852,N_18673,N_18672);
nand U18853 (N_18853,N_18660,N_18573);
or U18854 (N_18854,N_18621,N_18597);
or U18855 (N_18855,N_18668,N_18682);
nor U18856 (N_18856,N_18658,N_18585);
nand U18857 (N_18857,N_18631,N_18626);
and U18858 (N_18858,N_18576,N_18587);
nand U18859 (N_18859,N_18677,N_18567);
or U18860 (N_18860,N_18624,N_18671);
and U18861 (N_18861,N_18605,N_18715);
nand U18862 (N_18862,N_18670,N_18622);
or U18863 (N_18863,N_18639,N_18569);
nand U18864 (N_18864,N_18674,N_18688);
xnor U18865 (N_18865,N_18606,N_18702);
and U18866 (N_18866,N_18620,N_18591);
nor U18867 (N_18867,N_18691,N_18688);
xnor U18868 (N_18868,N_18666,N_18679);
xnor U18869 (N_18869,N_18582,N_18565);
or U18870 (N_18870,N_18633,N_18605);
nand U18871 (N_18871,N_18718,N_18646);
nor U18872 (N_18872,N_18677,N_18675);
nand U18873 (N_18873,N_18712,N_18661);
and U18874 (N_18874,N_18648,N_18694);
or U18875 (N_18875,N_18660,N_18685);
and U18876 (N_18876,N_18706,N_18719);
and U18877 (N_18877,N_18692,N_18641);
nor U18878 (N_18878,N_18700,N_18616);
nor U18879 (N_18879,N_18715,N_18620);
or U18880 (N_18880,N_18856,N_18747);
nor U18881 (N_18881,N_18777,N_18857);
nand U18882 (N_18882,N_18741,N_18764);
nor U18883 (N_18883,N_18726,N_18773);
nor U18884 (N_18884,N_18838,N_18758);
xor U18885 (N_18885,N_18854,N_18834);
or U18886 (N_18886,N_18735,N_18815);
and U18887 (N_18887,N_18754,N_18829);
nand U18888 (N_18888,N_18745,N_18774);
or U18889 (N_18889,N_18751,N_18844);
xnor U18890 (N_18890,N_18819,N_18836);
nor U18891 (N_18891,N_18811,N_18721);
and U18892 (N_18892,N_18753,N_18866);
or U18893 (N_18893,N_18782,N_18862);
and U18894 (N_18894,N_18845,N_18865);
or U18895 (N_18895,N_18869,N_18732);
nand U18896 (N_18896,N_18822,N_18796);
and U18897 (N_18897,N_18816,N_18737);
nor U18898 (N_18898,N_18757,N_18722);
nor U18899 (N_18899,N_18874,N_18739);
xnor U18900 (N_18900,N_18775,N_18763);
nand U18901 (N_18901,N_18784,N_18791);
and U18902 (N_18902,N_18772,N_18848);
and U18903 (N_18903,N_18795,N_18876);
nand U18904 (N_18904,N_18787,N_18759);
nand U18905 (N_18905,N_18805,N_18841);
or U18906 (N_18906,N_18790,N_18851);
and U18907 (N_18907,N_18867,N_18756);
nor U18908 (N_18908,N_18750,N_18767);
and U18909 (N_18909,N_18794,N_18785);
nand U18910 (N_18910,N_18868,N_18800);
nor U18911 (N_18911,N_18799,N_18731);
nand U18912 (N_18912,N_18870,N_18810);
xnor U18913 (N_18913,N_18780,N_18814);
or U18914 (N_18914,N_18840,N_18727);
or U18915 (N_18915,N_18778,N_18723);
and U18916 (N_18916,N_18744,N_18812);
or U18917 (N_18917,N_18797,N_18783);
or U18918 (N_18918,N_18789,N_18835);
and U18919 (N_18919,N_18755,N_18831);
or U18920 (N_18920,N_18742,N_18821);
nor U18921 (N_18921,N_18740,N_18761);
and U18922 (N_18922,N_18738,N_18864);
and U18923 (N_18923,N_18769,N_18839);
or U18924 (N_18924,N_18765,N_18825);
and U18925 (N_18925,N_18752,N_18771);
or U18926 (N_18926,N_18875,N_18720);
and U18927 (N_18927,N_18804,N_18733);
nand U18928 (N_18928,N_18760,N_18847);
and U18929 (N_18929,N_18817,N_18846);
nor U18930 (N_18930,N_18850,N_18872);
nor U18931 (N_18931,N_18749,N_18746);
xnor U18932 (N_18932,N_18748,N_18826);
and U18933 (N_18933,N_18861,N_18853);
xor U18934 (N_18934,N_18824,N_18852);
nor U18935 (N_18935,N_18779,N_18770);
xor U18936 (N_18936,N_18828,N_18792);
or U18937 (N_18937,N_18798,N_18837);
nand U18938 (N_18938,N_18729,N_18823);
xnor U18939 (N_18939,N_18807,N_18736);
xnor U18940 (N_18940,N_18730,N_18808);
or U18941 (N_18941,N_18743,N_18842);
nor U18942 (N_18942,N_18768,N_18818);
xor U18943 (N_18943,N_18813,N_18849);
or U18944 (N_18944,N_18806,N_18833);
or U18945 (N_18945,N_18877,N_18860);
nor U18946 (N_18946,N_18873,N_18809);
nor U18947 (N_18947,N_18802,N_18871);
and U18948 (N_18948,N_18820,N_18878);
or U18949 (N_18949,N_18855,N_18776);
or U18950 (N_18950,N_18725,N_18781);
nand U18951 (N_18951,N_18830,N_18766);
or U18952 (N_18952,N_18859,N_18734);
or U18953 (N_18953,N_18728,N_18724);
and U18954 (N_18954,N_18801,N_18863);
and U18955 (N_18955,N_18832,N_18788);
and U18956 (N_18956,N_18803,N_18843);
nand U18957 (N_18957,N_18762,N_18879);
nand U18958 (N_18958,N_18827,N_18786);
or U18959 (N_18959,N_18793,N_18858);
or U18960 (N_18960,N_18773,N_18805);
and U18961 (N_18961,N_18736,N_18801);
nand U18962 (N_18962,N_18733,N_18762);
or U18963 (N_18963,N_18870,N_18854);
nor U18964 (N_18964,N_18851,N_18744);
nand U18965 (N_18965,N_18837,N_18791);
nand U18966 (N_18966,N_18847,N_18768);
nor U18967 (N_18967,N_18721,N_18774);
or U18968 (N_18968,N_18834,N_18774);
and U18969 (N_18969,N_18848,N_18869);
xnor U18970 (N_18970,N_18785,N_18781);
nor U18971 (N_18971,N_18872,N_18812);
nand U18972 (N_18972,N_18834,N_18874);
and U18973 (N_18973,N_18775,N_18722);
nand U18974 (N_18974,N_18794,N_18776);
nor U18975 (N_18975,N_18735,N_18778);
and U18976 (N_18976,N_18850,N_18727);
nor U18977 (N_18977,N_18726,N_18747);
nor U18978 (N_18978,N_18795,N_18728);
and U18979 (N_18979,N_18780,N_18859);
or U18980 (N_18980,N_18800,N_18751);
nand U18981 (N_18981,N_18792,N_18771);
or U18982 (N_18982,N_18835,N_18763);
xor U18983 (N_18983,N_18849,N_18801);
nor U18984 (N_18984,N_18831,N_18866);
nor U18985 (N_18985,N_18862,N_18817);
xor U18986 (N_18986,N_18822,N_18792);
or U18987 (N_18987,N_18775,N_18729);
xnor U18988 (N_18988,N_18866,N_18867);
or U18989 (N_18989,N_18785,N_18743);
or U18990 (N_18990,N_18851,N_18868);
nand U18991 (N_18991,N_18756,N_18798);
nand U18992 (N_18992,N_18771,N_18818);
nand U18993 (N_18993,N_18827,N_18846);
xnor U18994 (N_18994,N_18757,N_18850);
nor U18995 (N_18995,N_18768,N_18837);
nand U18996 (N_18996,N_18742,N_18806);
and U18997 (N_18997,N_18771,N_18728);
xor U18998 (N_18998,N_18720,N_18874);
nand U18999 (N_18999,N_18787,N_18801);
nand U19000 (N_19000,N_18765,N_18807);
nor U19001 (N_19001,N_18732,N_18759);
and U19002 (N_19002,N_18789,N_18767);
nor U19003 (N_19003,N_18802,N_18866);
and U19004 (N_19004,N_18841,N_18810);
and U19005 (N_19005,N_18730,N_18810);
nand U19006 (N_19006,N_18731,N_18785);
or U19007 (N_19007,N_18808,N_18733);
or U19008 (N_19008,N_18743,N_18808);
and U19009 (N_19009,N_18782,N_18849);
or U19010 (N_19010,N_18805,N_18760);
and U19011 (N_19011,N_18815,N_18786);
and U19012 (N_19012,N_18727,N_18795);
nand U19013 (N_19013,N_18726,N_18877);
nand U19014 (N_19014,N_18812,N_18845);
nor U19015 (N_19015,N_18795,N_18788);
nor U19016 (N_19016,N_18804,N_18854);
nand U19017 (N_19017,N_18870,N_18844);
and U19018 (N_19018,N_18841,N_18739);
nand U19019 (N_19019,N_18829,N_18865);
and U19020 (N_19020,N_18809,N_18722);
nor U19021 (N_19021,N_18873,N_18739);
and U19022 (N_19022,N_18842,N_18798);
and U19023 (N_19023,N_18866,N_18765);
xor U19024 (N_19024,N_18837,N_18743);
nand U19025 (N_19025,N_18821,N_18723);
or U19026 (N_19026,N_18722,N_18732);
nand U19027 (N_19027,N_18848,N_18741);
and U19028 (N_19028,N_18847,N_18798);
nor U19029 (N_19029,N_18760,N_18871);
or U19030 (N_19030,N_18830,N_18786);
and U19031 (N_19031,N_18732,N_18868);
and U19032 (N_19032,N_18765,N_18756);
nor U19033 (N_19033,N_18787,N_18849);
nor U19034 (N_19034,N_18744,N_18825);
nor U19035 (N_19035,N_18838,N_18755);
nor U19036 (N_19036,N_18838,N_18745);
nand U19037 (N_19037,N_18827,N_18861);
and U19038 (N_19038,N_18794,N_18803);
and U19039 (N_19039,N_18763,N_18838);
and U19040 (N_19040,N_18976,N_19037);
nand U19041 (N_19041,N_18972,N_18964);
nor U19042 (N_19042,N_19039,N_18888);
nand U19043 (N_19043,N_18902,N_18961);
xor U19044 (N_19044,N_18928,N_18971);
nand U19045 (N_19045,N_19019,N_18952);
or U19046 (N_19046,N_18892,N_19031);
and U19047 (N_19047,N_18917,N_18975);
and U19048 (N_19048,N_18897,N_19015);
and U19049 (N_19049,N_18939,N_19023);
xnor U19050 (N_19050,N_18989,N_18957);
nor U19051 (N_19051,N_19001,N_18881);
nand U19052 (N_19052,N_18950,N_18967);
nor U19053 (N_19053,N_18966,N_18981);
and U19054 (N_19054,N_18915,N_19030);
nor U19055 (N_19055,N_18908,N_19006);
nand U19056 (N_19056,N_19036,N_18986);
or U19057 (N_19057,N_19007,N_18940);
or U19058 (N_19058,N_18980,N_18987);
xor U19059 (N_19059,N_18899,N_18895);
nand U19060 (N_19060,N_18962,N_19022);
nor U19061 (N_19061,N_18909,N_18911);
or U19062 (N_19062,N_18935,N_19021);
nand U19063 (N_19063,N_18919,N_18951);
nand U19064 (N_19064,N_18930,N_18936);
or U19065 (N_19065,N_19003,N_18913);
nand U19066 (N_19066,N_18990,N_18898);
or U19067 (N_19067,N_18973,N_19017);
nor U19068 (N_19068,N_18901,N_18883);
nand U19069 (N_19069,N_19033,N_18927);
xor U19070 (N_19070,N_19014,N_18983);
and U19071 (N_19071,N_18922,N_19000);
or U19072 (N_19072,N_18894,N_18947);
and U19073 (N_19073,N_18923,N_18906);
nor U19074 (N_19074,N_18905,N_19034);
and U19075 (N_19075,N_18925,N_19038);
or U19076 (N_19076,N_18933,N_18988);
and U19077 (N_19077,N_18904,N_19020);
or U19078 (N_19078,N_19002,N_18996);
nor U19079 (N_19079,N_18889,N_18924);
or U19080 (N_19080,N_18912,N_18968);
nor U19081 (N_19081,N_18982,N_18965);
or U19082 (N_19082,N_18963,N_19024);
nor U19083 (N_19083,N_18970,N_18960);
xnor U19084 (N_19084,N_18920,N_19011);
nand U19085 (N_19085,N_18934,N_18999);
nand U19086 (N_19086,N_19004,N_18900);
nor U19087 (N_19087,N_19027,N_18921);
or U19088 (N_19088,N_18954,N_18938);
xnor U19089 (N_19089,N_19032,N_18943);
or U19090 (N_19090,N_18979,N_18880);
and U19091 (N_19091,N_18931,N_18885);
nor U19092 (N_19092,N_19018,N_18944);
and U19093 (N_19093,N_19025,N_18942);
nand U19094 (N_19094,N_18992,N_18903);
or U19095 (N_19095,N_18969,N_19035);
nor U19096 (N_19096,N_19029,N_18998);
xnor U19097 (N_19097,N_18945,N_18887);
or U19098 (N_19098,N_18958,N_18907);
and U19099 (N_19099,N_18959,N_18948);
nor U19100 (N_19100,N_19026,N_18918);
or U19101 (N_19101,N_18956,N_18891);
nand U19102 (N_19102,N_19005,N_18946);
or U19103 (N_19103,N_19013,N_18910);
or U19104 (N_19104,N_18890,N_18978);
or U19105 (N_19105,N_18886,N_19028);
nand U19106 (N_19106,N_18941,N_18985);
or U19107 (N_19107,N_18994,N_18977);
nor U19108 (N_19108,N_18896,N_18916);
nand U19109 (N_19109,N_18955,N_18995);
or U19110 (N_19110,N_18974,N_18884);
nor U19111 (N_19111,N_18914,N_18953);
nand U19112 (N_19112,N_18937,N_18882);
and U19113 (N_19113,N_18926,N_18993);
nand U19114 (N_19114,N_19010,N_18991);
or U19115 (N_19115,N_19016,N_18932);
nand U19116 (N_19116,N_19008,N_18997);
or U19117 (N_19117,N_18893,N_18949);
or U19118 (N_19118,N_18929,N_19012);
xor U19119 (N_19119,N_18984,N_19009);
or U19120 (N_19120,N_18917,N_18949);
or U19121 (N_19121,N_18886,N_18887);
and U19122 (N_19122,N_18961,N_19005);
and U19123 (N_19123,N_19024,N_18954);
and U19124 (N_19124,N_18979,N_18903);
nand U19125 (N_19125,N_18993,N_19025);
nand U19126 (N_19126,N_19007,N_18957);
and U19127 (N_19127,N_19020,N_19016);
nor U19128 (N_19128,N_18993,N_18940);
and U19129 (N_19129,N_18904,N_18958);
xor U19130 (N_19130,N_18981,N_18937);
nor U19131 (N_19131,N_18952,N_18967);
and U19132 (N_19132,N_19023,N_18999);
or U19133 (N_19133,N_18881,N_19026);
or U19134 (N_19134,N_18959,N_18919);
nand U19135 (N_19135,N_18897,N_19003);
nand U19136 (N_19136,N_19005,N_19020);
xnor U19137 (N_19137,N_18882,N_18905);
and U19138 (N_19138,N_18969,N_19032);
or U19139 (N_19139,N_19028,N_19001);
or U19140 (N_19140,N_19033,N_18906);
or U19141 (N_19141,N_18937,N_19025);
nand U19142 (N_19142,N_18989,N_18967);
and U19143 (N_19143,N_18969,N_18996);
xnor U19144 (N_19144,N_18930,N_18907);
or U19145 (N_19145,N_18917,N_18984);
or U19146 (N_19146,N_18997,N_18896);
xnor U19147 (N_19147,N_18918,N_19024);
xor U19148 (N_19148,N_19007,N_18936);
and U19149 (N_19149,N_18911,N_18987);
and U19150 (N_19150,N_18894,N_19035);
nor U19151 (N_19151,N_19020,N_18890);
nor U19152 (N_19152,N_18945,N_18938);
nor U19153 (N_19153,N_18945,N_18965);
nand U19154 (N_19154,N_18947,N_19005);
xnor U19155 (N_19155,N_18966,N_18933);
or U19156 (N_19156,N_19038,N_19028);
nor U19157 (N_19157,N_18974,N_19034);
nand U19158 (N_19158,N_18946,N_18966);
nand U19159 (N_19159,N_18947,N_18939);
nand U19160 (N_19160,N_18894,N_18930);
nor U19161 (N_19161,N_18914,N_18916);
nor U19162 (N_19162,N_18998,N_19012);
nand U19163 (N_19163,N_18967,N_18974);
and U19164 (N_19164,N_18899,N_18892);
or U19165 (N_19165,N_19014,N_18934);
nor U19166 (N_19166,N_18955,N_18957);
nor U19167 (N_19167,N_19019,N_18903);
xor U19168 (N_19168,N_18985,N_18900);
or U19169 (N_19169,N_18916,N_18983);
nor U19170 (N_19170,N_18997,N_18950);
nand U19171 (N_19171,N_18960,N_18980);
and U19172 (N_19172,N_18889,N_18901);
or U19173 (N_19173,N_19014,N_18974);
nand U19174 (N_19174,N_18943,N_18897);
nand U19175 (N_19175,N_18883,N_18993);
nor U19176 (N_19176,N_18969,N_18946);
nor U19177 (N_19177,N_18990,N_19012);
or U19178 (N_19178,N_19018,N_18907);
or U19179 (N_19179,N_18886,N_19021);
or U19180 (N_19180,N_18909,N_18966);
nand U19181 (N_19181,N_18997,N_18934);
or U19182 (N_19182,N_18895,N_18967);
nand U19183 (N_19183,N_18966,N_18885);
nand U19184 (N_19184,N_18921,N_18911);
and U19185 (N_19185,N_18885,N_18954);
or U19186 (N_19186,N_18907,N_18906);
and U19187 (N_19187,N_19017,N_18974);
nor U19188 (N_19188,N_18936,N_18887);
and U19189 (N_19189,N_18987,N_18891);
nand U19190 (N_19190,N_18906,N_19037);
nor U19191 (N_19191,N_18951,N_18904);
or U19192 (N_19192,N_18891,N_18998);
and U19193 (N_19193,N_18902,N_18972);
xnor U19194 (N_19194,N_18930,N_18906);
xor U19195 (N_19195,N_18913,N_18971);
nor U19196 (N_19196,N_19014,N_18924);
nand U19197 (N_19197,N_18927,N_18901);
nand U19198 (N_19198,N_18979,N_19037);
or U19199 (N_19199,N_18963,N_18942);
nor U19200 (N_19200,N_19199,N_19057);
nand U19201 (N_19201,N_19146,N_19130);
and U19202 (N_19202,N_19095,N_19060);
or U19203 (N_19203,N_19118,N_19087);
and U19204 (N_19204,N_19140,N_19068);
nand U19205 (N_19205,N_19188,N_19101);
and U19206 (N_19206,N_19189,N_19108);
nor U19207 (N_19207,N_19184,N_19195);
nand U19208 (N_19208,N_19114,N_19181);
nor U19209 (N_19209,N_19104,N_19136);
and U19210 (N_19210,N_19058,N_19128);
or U19211 (N_19211,N_19059,N_19049);
nor U19212 (N_19212,N_19077,N_19169);
xnor U19213 (N_19213,N_19124,N_19078);
nand U19214 (N_19214,N_19134,N_19066);
nand U19215 (N_19215,N_19121,N_19089);
and U19216 (N_19216,N_19129,N_19145);
nand U19217 (N_19217,N_19086,N_19067);
nand U19218 (N_19218,N_19081,N_19163);
and U19219 (N_19219,N_19174,N_19138);
nand U19220 (N_19220,N_19069,N_19045);
or U19221 (N_19221,N_19074,N_19061);
and U19222 (N_19222,N_19097,N_19105);
nand U19223 (N_19223,N_19092,N_19178);
xnor U19224 (N_19224,N_19191,N_19151);
nand U19225 (N_19225,N_19041,N_19051);
xor U19226 (N_19226,N_19177,N_19091);
xor U19227 (N_19227,N_19112,N_19122);
nor U19228 (N_19228,N_19168,N_19107);
nor U19229 (N_19229,N_19125,N_19166);
nor U19230 (N_19230,N_19090,N_19182);
or U19231 (N_19231,N_19126,N_19096);
xnor U19232 (N_19232,N_19161,N_19042);
xnor U19233 (N_19233,N_19071,N_19047);
xnor U19234 (N_19234,N_19186,N_19153);
or U19235 (N_19235,N_19149,N_19076);
nand U19236 (N_19236,N_19070,N_19080);
nor U19237 (N_19237,N_19131,N_19043);
or U19238 (N_19238,N_19053,N_19185);
or U19239 (N_19239,N_19046,N_19198);
or U19240 (N_19240,N_19175,N_19119);
or U19241 (N_19241,N_19102,N_19159);
and U19242 (N_19242,N_19082,N_19179);
or U19243 (N_19243,N_19157,N_19137);
or U19244 (N_19244,N_19075,N_19065);
xnor U19245 (N_19245,N_19120,N_19064);
nand U19246 (N_19246,N_19147,N_19143);
and U19247 (N_19247,N_19088,N_19099);
nor U19248 (N_19248,N_19063,N_19176);
or U19249 (N_19249,N_19073,N_19117);
xor U19250 (N_19250,N_19154,N_19072);
and U19251 (N_19251,N_19167,N_19100);
and U19252 (N_19252,N_19098,N_19079);
or U19253 (N_19253,N_19183,N_19103);
or U19254 (N_19254,N_19194,N_19160);
or U19255 (N_19255,N_19109,N_19052);
xor U19256 (N_19256,N_19196,N_19171);
and U19257 (N_19257,N_19192,N_19110);
nand U19258 (N_19258,N_19141,N_19085);
nand U19259 (N_19259,N_19116,N_19135);
nand U19260 (N_19260,N_19148,N_19093);
or U19261 (N_19261,N_19164,N_19170);
nor U19262 (N_19262,N_19150,N_19113);
nand U19263 (N_19263,N_19193,N_19173);
nand U19264 (N_19264,N_19162,N_19172);
xor U19265 (N_19265,N_19084,N_19055);
nand U19266 (N_19266,N_19165,N_19156);
or U19267 (N_19267,N_19180,N_19127);
xnor U19268 (N_19268,N_19048,N_19190);
nand U19269 (N_19269,N_19115,N_19139);
nand U19270 (N_19270,N_19094,N_19044);
or U19271 (N_19271,N_19106,N_19111);
nand U19272 (N_19272,N_19144,N_19050);
nor U19273 (N_19273,N_19187,N_19083);
and U19274 (N_19274,N_19133,N_19054);
xor U19275 (N_19275,N_19062,N_19158);
or U19276 (N_19276,N_19152,N_19155);
nand U19277 (N_19277,N_19142,N_19040);
or U19278 (N_19278,N_19123,N_19056);
xnor U19279 (N_19279,N_19197,N_19132);
nor U19280 (N_19280,N_19107,N_19166);
nand U19281 (N_19281,N_19189,N_19067);
xor U19282 (N_19282,N_19188,N_19180);
nor U19283 (N_19283,N_19176,N_19141);
and U19284 (N_19284,N_19114,N_19047);
or U19285 (N_19285,N_19179,N_19196);
and U19286 (N_19286,N_19196,N_19091);
and U19287 (N_19287,N_19181,N_19083);
or U19288 (N_19288,N_19138,N_19127);
nor U19289 (N_19289,N_19133,N_19067);
nand U19290 (N_19290,N_19161,N_19157);
nand U19291 (N_19291,N_19059,N_19051);
or U19292 (N_19292,N_19120,N_19158);
nor U19293 (N_19293,N_19153,N_19135);
nor U19294 (N_19294,N_19153,N_19144);
nor U19295 (N_19295,N_19062,N_19069);
and U19296 (N_19296,N_19061,N_19192);
xnor U19297 (N_19297,N_19158,N_19086);
nand U19298 (N_19298,N_19111,N_19135);
nand U19299 (N_19299,N_19154,N_19152);
nor U19300 (N_19300,N_19153,N_19149);
nor U19301 (N_19301,N_19123,N_19106);
or U19302 (N_19302,N_19152,N_19066);
and U19303 (N_19303,N_19089,N_19052);
and U19304 (N_19304,N_19102,N_19084);
or U19305 (N_19305,N_19045,N_19088);
nor U19306 (N_19306,N_19148,N_19193);
and U19307 (N_19307,N_19047,N_19158);
nand U19308 (N_19308,N_19140,N_19176);
nand U19309 (N_19309,N_19132,N_19199);
nor U19310 (N_19310,N_19138,N_19170);
or U19311 (N_19311,N_19158,N_19181);
and U19312 (N_19312,N_19155,N_19169);
nand U19313 (N_19313,N_19045,N_19100);
nand U19314 (N_19314,N_19102,N_19168);
xor U19315 (N_19315,N_19076,N_19073);
and U19316 (N_19316,N_19069,N_19180);
nor U19317 (N_19317,N_19041,N_19169);
nor U19318 (N_19318,N_19177,N_19182);
nor U19319 (N_19319,N_19098,N_19105);
and U19320 (N_19320,N_19043,N_19154);
or U19321 (N_19321,N_19083,N_19186);
nor U19322 (N_19322,N_19106,N_19085);
nor U19323 (N_19323,N_19043,N_19100);
and U19324 (N_19324,N_19188,N_19115);
and U19325 (N_19325,N_19175,N_19137);
xor U19326 (N_19326,N_19188,N_19079);
or U19327 (N_19327,N_19107,N_19136);
nor U19328 (N_19328,N_19101,N_19086);
nand U19329 (N_19329,N_19054,N_19063);
xor U19330 (N_19330,N_19096,N_19065);
nand U19331 (N_19331,N_19197,N_19151);
and U19332 (N_19332,N_19166,N_19087);
nand U19333 (N_19333,N_19190,N_19129);
nand U19334 (N_19334,N_19079,N_19109);
or U19335 (N_19335,N_19181,N_19156);
xor U19336 (N_19336,N_19186,N_19096);
and U19337 (N_19337,N_19097,N_19100);
nor U19338 (N_19338,N_19110,N_19184);
and U19339 (N_19339,N_19094,N_19174);
or U19340 (N_19340,N_19049,N_19134);
xnor U19341 (N_19341,N_19109,N_19151);
nand U19342 (N_19342,N_19146,N_19116);
nand U19343 (N_19343,N_19068,N_19073);
and U19344 (N_19344,N_19107,N_19082);
xnor U19345 (N_19345,N_19085,N_19077);
or U19346 (N_19346,N_19117,N_19088);
or U19347 (N_19347,N_19195,N_19177);
nor U19348 (N_19348,N_19053,N_19073);
or U19349 (N_19349,N_19059,N_19092);
xnor U19350 (N_19350,N_19147,N_19100);
or U19351 (N_19351,N_19074,N_19057);
nor U19352 (N_19352,N_19137,N_19142);
or U19353 (N_19353,N_19140,N_19149);
or U19354 (N_19354,N_19180,N_19192);
and U19355 (N_19355,N_19131,N_19144);
nor U19356 (N_19356,N_19040,N_19071);
or U19357 (N_19357,N_19177,N_19115);
and U19358 (N_19358,N_19171,N_19154);
nor U19359 (N_19359,N_19158,N_19199);
nor U19360 (N_19360,N_19207,N_19225);
or U19361 (N_19361,N_19306,N_19357);
and U19362 (N_19362,N_19243,N_19309);
nor U19363 (N_19363,N_19214,N_19329);
or U19364 (N_19364,N_19343,N_19319);
and U19365 (N_19365,N_19253,N_19301);
xnor U19366 (N_19366,N_19236,N_19336);
nand U19367 (N_19367,N_19347,N_19328);
nor U19368 (N_19368,N_19317,N_19304);
and U19369 (N_19369,N_19266,N_19292);
nor U19370 (N_19370,N_19258,N_19332);
nor U19371 (N_19371,N_19335,N_19259);
nor U19372 (N_19372,N_19264,N_19260);
nor U19373 (N_19373,N_19269,N_19284);
nand U19374 (N_19374,N_19256,N_19263);
nor U19375 (N_19375,N_19272,N_19281);
and U19376 (N_19376,N_19303,N_19356);
or U19377 (N_19377,N_19300,N_19315);
nor U19378 (N_19378,N_19215,N_19311);
and U19379 (N_19379,N_19277,N_19331);
nor U19380 (N_19380,N_19341,N_19358);
xnor U19381 (N_19381,N_19238,N_19349);
nor U19382 (N_19382,N_19313,N_19282);
and U19383 (N_19383,N_19250,N_19254);
xnor U19384 (N_19384,N_19279,N_19200);
or U19385 (N_19385,N_19345,N_19247);
and U19386 (N_19386,N_19299,N_19296);
nand U19387 (N_19387,N_19219,N_19323);
nand U19388 (N_19388,N_19233,N_19257);
or U19389 (N_19389,N_19204,N_19226);
nor U19390 (N_19390,N_19230,N_19223);
and U19391 (N_19391,N_19235,N_19248);
xnor U19392 (N_19392,N_19244,N_19213);
nand U19393 (N_19393,N_19337,N_19320);
nor U19394 (N_19394,N_19327,N_19294);
nor U19395 (N_19395,N_19308,N_19261);
or U19396 (N_19396,N_19339,N_19350);
xnor U19397 (N_19397,N_19271,N_19237);
nand U19398 (N_19398,N_19203,N_19216);
nor U19399 (N_19399,N_19346,N_19275);
or U19400 (N_19400,N_19289,N_19338);
or U19401 (N_19401,N_19228,N_19352);
nor U19402 (N_19402,N_19217,N_19344);
nor U19403 (N_19403,N_19334,N_19297);
and U19404 (N_19404,N_19286,N_19262);
nand U19405 (N_19405,N_19206,N_19288);
nand U19406 (N_19406,N_19325,N_19240);
or U19407 (N_19407,N_19295,N_19274);
xor U19408 (N_19408,N_19229,N_19324);
or U19409 (N_19409,N_19333,N_19273);
or U19410 (N_19410,N_19267,N_19314);
and U19411 (N_19411,N_19330,N_19340);
nand U19412 (N_19412,N_19252,N_19307);
and U19413 (N_19413,N_19321,N_19224);
and U19414 (N_19414,N_19316,N_19302);
nand U19415 (N_19415,N_19231,N_19268);
nand U19416 (N_19416,N_19239,N_19241);
nand U19417 (N_19417,N_19342,N_19234);
nor U19418 (N_19418,N_19351,N_19348);
nand U19419 (N_19419,N_19287,N_19285);
or U19420 (N_19420,N_19305,N_19291);
or U19421 (N_19421,N_19353,N_19202);
and U19422 (N_19422,N_19276,N_19355);
nand U19423 (N_19423,N_19265,N_19354);
xnor U19424 (N_19424,N_19318,N_19210);
xnor U19425 (N_19425,N_19312,N_19249);
nand U19426 (N_19426,N_19242,N_19245);
nand U19427 (N_19427,N_19293,N_19283);
or U19428 (N_19428,N_19298,N_19310);
nor U19429 (N_19429,N_19278,N_19222);
xnor U19430 (N_19430,N_19211,N_19280);
or U19431 (N_19431,N_19208,N_19227);
and U19432 (N_19432,N_19232,N_19251);
or U19433 (N_19433,N_19212,N_19220);
nor U19434 (N_19434,N_19209,N_19290);
nor U19435 (N_19435,N_19218,N_19270);
and U19436 (N_19436,N_19221,N_19359);
and U19437 (N_19437,N_19322,N_19201);
nand U19438 (N_19438,N_19255,N_19205);
and U19439 (N_19439,N_19326,N_19246);
nand U19440 (N_19440,N_19226,N_19217);
nand U19441 (N_19441,N_19255,N_19262);
xnor U19442 (N_19442,N_19249,N_19234);
and U19443 (N_19443,N_19324,N_19235);
nor U19444 (N_19444,N_19223,N_19242);
and U19445 (N_19445,N_19207,N_19300);
or U19446 (N_19446,N_19201,N_19346);
or U19447 (N_19447,N_19294,N_19337);
xor U19448 (N_19448,N_19206,N_19327);
and U19449 (N_19449,N_19300,N_19311);
xnor U19450 (N_19450,N_19252,N_19339);
or U19451 (N_19451,N_19243,N_19338);
nand U19452 (N_19452,N_19228,N_19301);
nand U19453 (N_19453,N_19210,N_19245);
xor U19454 (N_19454,N_19241,N_19319);
and U19455 (N_19455,N_19349,N_19212);
nand U19456 (N_19456,N_19348,N_19321);
and U19457 (N_19457,N_19316,N_19257);
or U19458 (N_19458,N_19254,N_19203);
nor U19459 (N_19459,N_19266,N_19278);
nor U19460 (N_19460,N_19208,N_19260);
and U19461 (N_19461,N_19257,N_19276);
nor U19462 (N_19462,N_19353,N_19281);
and U19463 (N_19463,N_19227,N_19260);
nand U19464 (N_19464,N_19309,N_19245);
nand U19465 (N_19465,N_19283,N_19280);
nand U19466 (N_19466,N_19255,N_19279);
xor U19467 (N_19467,N_19217,N_19310);
or U19468 (N_19468,N_19200,N_19234);
and U19469 (N_19469,N_19344,N_19295);
or U19470 (N_19470,N_19247,N_19306);
xor U19471 (N_19471,N_19348,N_19208);
nand U19472 (N_19472,N_19294,N_19295);
nor U19473 (N_19473,N_19226,N_19301);
nand U19474 (N_19474,N_19274,N_19336);
or U19475 (N_19475,N_19206,N_19347);
nand U19476 (N_19476,N_19273,N_19234);
or U19477 (N_19477,N_19210,N_19320);
and U19478 (N_19478,N_19219,N_19254);
nand U19479 (N_19479,N_19325,N_19208);
nor U19480 (N_19480,N_19239,N_19230);
nor U19481 (N_19481,N_19317,N_19275);
or U19482 (N_19482,N_19244,N_19287);
or U19483 (N_19483,N_19352,N_19203);
or U19484 (N_19484,N_19249,N_19320);
or U19485 (N_19485,N_19307,N_19266);
nand U19486 (N_19486,N_19279,N_19302);
xor U19487 (N_19487,N_19350,N_19306);
or U19488 (N_19488,N_19358,N_19271);
nand U19489 (N_19489,N_19291,N_19232);
nor U19490 (N_19490,N_19241,N_19253);
or U19491 (N_19491,N_19326,N_19254);
and U19492 (N_19492,N_19310,N_19355);
or U19493 (N_19493,N_19289,N_19230);
or U19494 (N_19494,N_19239,N_19234);
xor U19495 (N_19495,N_19219,N_19230);
or U19496 (N_19496,N_19319,N_19253);
xor U19497 (N_19497,N_19292,N_19345);
and U19498 (N_19498,N_19226,N_19225);
or U19499 (N_19499,N_19219,N_19313);
xor U19500 (N_19500,N_19327,N_19248);
and U19501 (N_19501,N_19253,N_19283);
nor U19502 (N_19502,N_19266,N_19210);
nor U19503 (N_19503,N_19258,N_19289);
xnor U19504 (N_19504,N_19315,N_19328);
nor U19505 (N_19505,N_19225,N_19202);
or U19506 (N_19506,N_19221,N_19234);
and U19507 (N_19507,N_19216,N_19230);
nand U19508 (N_19508,N_19207,N_19244);
and U19509 (N_19509,N_19271,N_19270);
xor U19510 (N_19510,N_19322,N_19288);
nor U19511 (N_19511,N_19201,N_19267);
nand U19512 (N_19512,N_19229,N_19216);
nor U19513 (N_19513,N_19258,N_19351);
nor U19514 (N_19514,N_19273,N_19295);
or U19515 (N_19515,N_19339,N_19306);
nor U19516 (N_19516,N_19327,N_19217);
or U19517 (N_19517,N_19332,N_19273);
nand U19518 (N_19518,N_19351,N_19317);
nor U19519 (N_19519,N_19352,N_19252);
and U19520 (N_19520,N_19429,N_19430);
nor U19521 (N_19521,N_19464,N_19452);
xnor U19522 (N_19522,N_19489,N_19494);
nand U19523 (N_19523,N_19419,N_19365);
or U19524 (N_19524,N_19425,N_19479);
or U19525 (N_19525,N_19373,N_19367);
nor U19526 (N_19526,N_19423,N_19441);
and U19527 (N_19527,N_19453,N_19444);
and U19528 (N_19528,N_19360,N_19438);
nor U19529 (N_19529,N_19379,N_19462);
or U19530 (N_19530,N_19390,N_19370);
nand U19531 (N_19531,N_19488,N_19381);
nand U19532 (N_19532,N_19407,N_19431);
and U19533 (N_19533,N_19509,N_19363);
nor U19534 (N_19534,N_19426,N_19480);
or U19535 (N_19535,N_19457,N_19391);
and U19536 (N_19536,N_19507,N_19369);
or U19537 (N_19537,N_19411,N_19513);
and U19538 (N_19538,N_19404,N_19465);
nand U19539 (N_19539,N_19415,N_19421);
or U19540 (N_19540,N_19382,N_19493);
or U19541 (N_19541,N_19477,N_19417);
and U19542 (N_19542,N_19422,N_19472);
or U19543 (N_19543,N_19362,N_19420);
nand U19544 (N_19544,N_19481,N_19449);
or U19545 (N_19545,N_19458,N_19502);
nor U19546 (N_19546,N_19505,N_19424);
xnor U19547 (N_19547,N_19374,N_19482);
xnor U19548 (N_19548,N_19361,N_19518);
or U19549 (N_19549,N_19447,N_19440);
or U19550 (N_19550,N_19508,N_19403);
and U19551 (N_19551,N_19484,N_19434);
nand U19552 (N_19552,N_19433,N_19387);
or U19553 (N_19553,N_19517,N_19446);
nand U19554 (N_19554,N_19519,N_19485);
nor U19555 (N_19555,N_19497,N_19451);
nor U19556 (N_19556,N_19468,N_19386);
xor U19557 (N_19557,N_19375,N_19510);
and U19558 (N_19558,N_19377,N_19475);
nand U19559 (N_19559,N_19435,N_19490);
or U19560 (N_19560,N_19445,N_19439);
or U19561 (N_19561,N_19392,N_19413);
and U19562 (N_19562,N_19496,N_19474);
and U19563 (N_19563,N_19463,N_19514);
or U19564 (N_19564,N_19408,N_19380);
or U19565 (N_19565,N_19414,N_19478);
nor U19566 (N_19566,N_19383,N_19402);
and U19567 (N_19567,N_19476,N_19506);
and U19568 (N_19568,N_19409,N_19492);
nand U19569 (N_19569,N_19371,N_19372);
and U19570 (N_19570,N_19459,N_19384);
nand U19571 (N_19571,N_19460,N_19442);
xnor U19572 (N_19572,N_19388,N_19418);
or U19573 (N_19573,N_19397,N_19394);
and U19574 (N_19574,N_19503,N_19455);
or U19575 (N_19575,N_19406,N_19491);
nor U19576 (N_19576,N_19461,N_19471);
and U19577 (N_19577,N_19443,N_19399);
nand U19578 (N_19578,N_19450,N_19454);
or U19579 (N_19579,N_19412,N_19395);
or U19580 (N_19580,N_19393,N_19436);
nor U19581 (N_19581,N_19511,N_19378);
xnor U19582 (N_19582,N_19486,N_19466);
nor U19583 (N_19583,N_19398,N_19401);
nand U19584 (N_19584,N_19368,N_19499);
and U19585 (N_19585,N_19500,N_19515);
or U19586 (N_19586,N_19473,N_19469);
nor U19587 (N_19587,N_19456,N_19448);
nor U19588 (N_19588,N_19432,N_19467);
and U19589 (N_19589,N_19376,N_19364);
and U19590 (N_19590,N_19428,N_19501);
nor U19591 (N_19591,N_19437,N_19498);
nand U19592 (N_19592,N_19495,N_19405);
nor U19593 (N_19593,N_19483,N_19416);
nor U19594 (N_19594,N_19396,N_19385);
nor U19595 (N_19595,N_19512,N_19389);
nand U19596 (N_19596,N_19400,N_19504);
nor U19597 (N_19597,N_19487,N_19427);
and U19598 (N_19598,N_19410,N_19470);
or U19599 (N_19599,N_19516,N_19366);
nor U19600 (N_19600,N_19382,N_19486);
and U19601 (N_19601,N_19370,N_19438);
nor U19602 (N_19602,N_19477,N_19443);
or U19603 (N_19603,N_19388,N_19441);
and U19604 (N_19604,N_19364,N_19422);
nor U19605 (N_19605,N_19386,N_19483);
nor U19606 (N_19606,N_19455,N_19514);
and U19607 (N_19607,N_19380,N_19386);
or U19608 (N_19608,N_19517,N_19403);
nand U19609 (N_19609,N_19468,N_19443);
and U19610 (N_19610,N_19380,N_19477);
nand U19611 (N_19611,N_19463,N_19444);
and U19612 (N_19612,N_19472,N_19447);
and U19613 (N_19613,N_19471,N_19506);
nor U19614 (N_19614,N_19488,N_19506);
or U19615 (N_19615,N_19474,N_19382);
xor U19616 (N_19616,N_19489,N_19458);
nor U19617 (N_19617,N_19373,N_19477);
nand U19618 (N_19618,N_19437,N_19370);
nand U19619 (N_19619,N_19485,N_19456);
or U19620 (N_19620,N_19470,N_19431);
xor U19621 (N_19621,N_19461,N_19519);
and U19622 (N_19622,N_19422,N_19421);
nand U19623 (N_19623,N_19511,N_19461);
or U19624 (N_19624,N_19369,N_19437);
xnor U19625 (N_19625,N_19459,N_19509);
or U19626 (N_19626,N_19413,N_19367);
nor U19627 (N_19627,N_19446,N_19411);
xnor U19628 (N_19628,N_19519,N_19438);
or U19629 (N_19629,N_19435,N_19394);
or U19630 (N_19630,N_19472,N_19483);
xor U19631 (N_19631,N_19473,N_19495);
or U19632 (N_19632,N_19468,N_19374);
nor U19633 (N_19633,N_19402,N_19372);
or U19634 (N_19634,N_19487,N_19458);
or U19635 (N_19635,N_19367,N_19510);
nor U19636 (N_19636,N_19415,N_19491);
xnor U19637 (N_19637,N_19454,N_19387);
or U19638 (N_19638,N_19360,N_19475);
nand U19639 (N_19639,N_19498,N_19422);
and U19640 (N_19640,N_19378,N_19482);
xnor U19641 (N_19641,N_19389,N_19414);
nand U19642 (N_19642,N_19517,N_19383);
nand U19643 (N_19643,N_19426,N_19392);
xnor U19644 (N_19644,N_19364,N_19457);
nor U19645 (N_19645,N_19371,N_19374);
or U19646 (N_19646,N_19382,N_19479);
nand U19647 (N_19647,N_19383,N_19448);
and U19648 (N_19648,N_19459,N_19363);
nor U19649 (N_19649,N_19413,N_19489);
and U19650 (N_19650,N_19451,N_19492);
or U19651 (N_19651,N_19500,N_19390);
or U19652 (N_19652,N_19421,N_19375);
nor U19653 (N_19653,N_19417,N_19392);
xnor U19654 (N_19654,N_19413,N_19437);
xnor U19655 (N_19655,N_19414,N_19509);
nand U19656 (N_19656,N_19387,N_19421);
nand U19657 (N_19657,N_19470,N_19389);
nand U19658 (N_19658,N_19369,N_19407);
nand U19659 (N_19659,N_19380,N_19475);
or U19660 (N_19660,N_19370,N_19429);
nor U19661 (N_19661,N_19384,N_19440);
or U19662 (N_19662,N_19418,N_19449);
nand U19663 (N_19663,N_19507,N_19483);
nand U19664 (N_19664,N_19491,N_19515);
and U19665 (N_19665,N_19436,N_19503);
nand U19666 (N_19666,N_19472,N_19377);
xor U19667 (N_19667,N_19502,N_19372);
nand U19668 (N_19668,N_19460,N_19417);
nand U19669 (N_19669,N_19419,N_19477);
and U19670 (N_19670,N_19397,N_19513);
or U19671 (N_19671,N_19432,N_19415);
nor U19672 (N_19672,N_19452,N_19389);
nand U19673 (N_19673,N_19511,N_19371);
nor U19674 (N_19674,N_19380,N_19416);
or U19675 (N_19675,N_19470,N_19379);
and U19676 (N_19676,N_19516,N_19422);
nor U19677 (N_19677,N_19421,N_19519);
or U19678 (N_19678,N_19513,N_19406);
nor U19679 (N_19679,N_19484,N_19371);
nor U19680 (N_19680,N_19610,N_19580);
nand U19681 (N_19681,N_19531,N_19623);
nor U19682 (N_19682,N_19555,N_19678);
or U19683 (N_19683,N_19553,N_19664);
or U19684 (N_19684,N_19629,N_19535);
or U19685 (N_19685,N_19603,N_19599);
nor U19686 (N_19686,N_19671,N_19591);
or U19687 (N_19687,N_19594,N_19608);
and U19688 (N_19688,N_19666,N_19564);
nor U19689 (N_19689,N_19578,N_19676);
nor U19690 (N_19690,N_19614,N_19543);
xor U19691 (N_19691,N_19650,N_19538);
nor U19692 (N_19692,N_19572,N_19657);
nor U19693 (N_19693,N_19654,N_19616);
and U19694 (N_19694,N_19540,N_19659);
and U19695 (N_19695,N_19662,N_19596);
or U19696 (N_19696,N_19552,N_19669);
nor U19697 (N_19697,N_19658,N_19645);
or U19698 (N_19698,N_19571,N_19632);
and U19699 (N_19699,N_19670,N_19611);
xor U19700 (N_19700,N_19667,N_19620);
nand U19701 (N_19701,N_19529,N_19576);
and U19702 (N_19702,N_19642,N_19637);
nor U19703 (N_19703,N_19646,N_19534);
and U19704 (N_19704,N_19618,N_19612);
xor U19705 (N_19705,N_19522,N_19565);
nor U19706 (N_19706,N_19528,N_19537);
or U19707 (N_19707,N_19624,N_19527);
or U19708 (N_19708,N_19556,N_19668);
nor U19709 (N_19709,N_19619,N_19577);
nor U19710 (N_19710,N_19652,N_19597);
nor U19711 (N_19711,N_19649,N_19633);
or U19712 (N_19712,N_19651,N_19585);
nand U19713 (N_19713,N_19536,N_19566);
or U19714 (N_19714,N_19533,N_19648);
nor U19715 (N_19715,N_19550,N_19638);
nand U19716 (N_19716,N_19575,N_19656);
nand U19717 (N_19717,N_19627,N_19523);
and U19718 (N_19718,N_19586,N_19588);
nand U19719 (N_19719,N_19615,N_19568);
nand U19720 (N_19720,N_19634,N_19567);
xor U19721 (N_19721,N_19547,N_19545);
nand U19722 (N_19722,N_19622,N_19605);
nor U19723 (N_19723,N_19600,N_19582);
or U19724 (N_19724,N_19581,N_19675);
or U19725 (N_19725,N_19607,N_19631);
or U19726 (N_19726,N_19539,N_19551);
and U19727 (N_19727,N_19625,N_19593);
nand U19728 (N_19728,N_19640,N_19592);
and U19729 (N_19729,N_19617,N_19587);
and U19730 (N_19730,N_19604,N_19644);
nor U19731 (N_19731,N_19554,N_19679);
nor U19732 (N_19732,N_19639,N_19655);
or U19733 (N_19733,N_19590,N_19674);
and U19734 (N_19734,N_19559,N_19601);
and U19735 (N_19735,N_19525,N_19665);
nor U19736 (N_19736,N_19560,N_19641);
nand U19737 (N_19737,N_19548,N_19549);
or U19738 (N_19738,N_19613,N_19595);
nor U19739 (N_19739,N_19541,N_19609);
nand U19740 (N_19740,N_19574,N_19544);
or U19741 (N_19741,N_19569,N_19561);
xnor U19742 (N_19742,N_19598,N_19546);
and U19743 (N_19743,N_19653,N_19628);
or U19744 (N_19744,N_19530,N_19672);
or U19745 (N_19745,N_19636,N_19621);
nand U19746 (N_19746,N_19635,N_19626);
and U19747 (N_19747,N_19661,N_19520);
and U19748 (N_19748,N_19557,N_19532);
nand U19749 (N_19749,N_19606,N_19647);
or U19750 (N_19750,N_19660,N_19558);
xor U19751 (N_19751,N_19583,N_19589);
and U19752 (N_19752,N_19643,N_19584);
and U19753 (N_19753,N_19602,N_19673);
nor U19754 (N_19754,N_19524,N_19663);
or U19755 (N_19755,N_19562,N_19521);
xor U19756 (N_19756,N_19579,N_19677);
nand U19757 (N_19757,N_19563,N_19542);
nor U19758 (N_19758,N_19570,N_19526);
and U19759 (N_19759,N_19630,N_19573);
nor U19760 (N_19760,N_19663,N_19552);
and U19761 (N_19761,N_19606,N_19617);
and U19762 (N_19762,N_19625,N_19572);
nand U19763 (N_19763,N_19597,N_19566);
and U19764 (N_19764,N_19538,N_19559);
or U19765 (N_19765,N_19637,N_19533);
nand U19766 (N_19766,N_19564,N_19654);
or U19767 (N_19767,N_19529,N_19628);
and U19768 (N_19768,N_19594,N_19575);
or U19769 (N_19769,N_19535,N_19635);
or U19770 (N_19770,N_19666,N_19544);
or U19771 (N_19771,N_19627,N_19645);
nor U19772 (N_19772,N_19583,N_19556);
nand U19773 (N_19773,N_19523,N_19613);
and U19774 (N_19774,N_19660,N_19616);
nand U19775 (N_19775,N_19673,N_19635);
nor U19776 (N_19776,N_19525,N_19632);
and U19777 (N_19777,N_19546,N_19655);
and U19778 (N_19778,N_19672,N_19633);
xnor U19779 (N_19779,N_19561,N_19615);
nand U19780 (N_19780,N_19553,N_19559);
or U19781 (N_19781,N_19617,N_19553);
or U19782 (N_19782,N_19534,N_19600);
xnor U19783 (N_19783,N_19630,N_19618);
nor U19784 (N_19784,N_19650,N_19652);
nor U19785 (N_19785,N_19609,N_19524);
nand U19786 (N_19786,N_19576,N_19561);
or U19787 (N_19787,N_19600,N_19658);
or U19788 (N_19788,N_19580,N_19668);
and U19789 (N_19789,N_19610,N_19576);
and U19790 (N_19790,N_19522,N_19553);
or U19791 (N_19791,N_19627,N_19543);
and U19792 (N_19792,N_19612,N_19538);
or U19793 (N_19793,N_19579,N_19621);
nor U19794 (N_19794,N_19544,N_19614);
nand U19795 (N_19795,N_19613,N_19678);
and U19796 (N_19796,N_19677,N_19535);
xor U19797 (N_19797,N_19520,N_19612);
nand U19798 (N_19798,N_19634,N_19583);
or U19799 (N_19799,N_19656,N_19592);
or U19800 (N_19800,N_19671,N_19645);
xnor U19801 (N_19801,N_19596,N_19668);
xor U19802 (N_19802,N_19556,N_19566);
or U19803 (N_19803,N_19574,N_19662);
and U19804 (N_19804,N_19570,N_19525);
xnor U19805 (N_19805,N_19625,N_19541);
or U19806 (N_19806,N_19540,N_19555);
nand U19807 (N_19807,N_19648,N_19545);
and U19808 (N_19808,N_19660,N_19586);
and U19809 (N_19809,N_19547,N_19619);
and U19810 (N_19810,N_19649,N_19637);
nor U19811 (N_19811,N_19626,N_19671);
nand U19812 (N_19812,N_19624,N_19561);
and U19813 (N_19813,N_19634,N_19564);
or U19814 (N_19814,N_19673,N_19562);
nor U19815 (N_19815,N_19579,N_19555);
nor U19816 (N_19816,N_19553,N_19667);
xnor U19817 (N_19817,N_19650,N_19545);
or U19818 (N_19818,N_19545,N_19645);
nor U19819 (N_19819,N_19557,N_19649);
or U19820 (N_19820,N_19642,N_19677);
nand U19821 (N_19821,N_19546,N_19526);
nor U19822 (N_19822,N_19616,N_19596);
xnor U19823 (N_19823,N_19565,N_19570);
nor U19824 (N_19824,N_19531,N_19670);
and U19825 (N_19825,N_19640,N_19534);
or U19826 (N_19826,N_19599,N_19547);
nor U19827 (N_19827,N_19524,N_19593);
nor U19828 (N_19828,N_19551,N_19644);
nand U19829 (N_19829,N_19538,N_19613);
nor U19830 (N_19830,N_19568,N_19526);
xor U19831 (N_19831,N_19525,N_19636);
and U19832 (N_19832,N_19552,N_19520);
or U19833 (N_19833,N_19679,N_19558);
or U19834 (N_19834,N_19619,N_19587);
nor U19835 (N_19835,N_19599,N_19678);
nor U19836 (N_19836,N_19526,N_19533);
and U19837 (N_19837,N_19600,N_19616);
nor U19838 (N_19838,N_19607,N_19568);
or U19839 (N_19839,N_19675,N_19622);
and U19840 (N_19840,N_19739,N_19778);
or U19841 (N_19841,N_19683,N_19764);
or U19842 (N_19842,N_19809,N_19745);
nor U19843 (N_19843,N_19751,N_19796);
xor U19844 (N_19844,N_19718,N_19743);
and U19845 (N_19845,N_19763,N_19775);
nand U19846 (N_19846,N_19756,N_19771);
nor U19847 (N_19847,N_19702,N_19754);
nor U19848 (N_19848,N_19768,N_19783);
nand U19849 (N_19849,N_19733,N_19760);
or U19850 (N_19850,N_19715,N_19772);
nor U19851 (N_19851,N_19681,N_19803);
and U19852 (N_19852,N_19738,N_19806);
and U19853 (N_19853,N_19832,N_19680);
nor U19854 (N_19854,N_19747,N_19822);
or U19855 (N_19855,N_19692,N_19740);
or U19856 (N_19856,N_19696,N_19838);
or U19857 (N_19857,N_19825,N_19789);
and U19858 (N_19858,N_19730,N_19716);
nand U19859 (N_19859,N_19812,N_19773);
and U19860 (N_19860,N_19779,N_19807);
nor U19861 (N_19861,N_19792,N_19688);
and U19862 (N_19862,N_19707,N_19826);
nor U19863 (N_19863,N_19788,N_19695);
or U19864 (N_19864,N_19828,N_19719);
or U19865 (N_19865,N_19837,N_19804);
or U19866 (N_19866,N_19801,N_19777);
nand U19867 (N_19867,N_19752,N_19782);
and U19868 (N_19868,N_19709,N_19731);
nand U19869 (N_19869,N_19713,N_19781);
or U19870 (N_19870,N_19735,N_19706);
or U19871 (N_19871,N_19817,N_19831);
and U19872 (N_19872,N_19805,N_19700);
nor U19873 (N_19873,N_19682,N_19794);
or U19874 (N_19874,N_19830,N_19711);
nand U19875 (N_19875,N_19699,N_19793);
or U19876 (N_19876,N_19684,N_19802);
xor U19877 (N_19877,N_19834,N_19734);
nand U19878 (N_19878,N_19780,N_19710);
and U19879 (N_19879,N_19755,N_19712);
nor U19880 (N_19880,N_19686,N_19767);
nand U19881 (N_19881,N_19704,N_19705);
nand U19882 (N_19882,N_19758,N_19766);
nand U19883 (N_19883,N_19721,N_19818);
and U19884 (N_19884,N_19725,N_19714);
and U19885 (N_19885,N_19765,N_19827);
nor U19886 (N_19886,N_19697,N_19757);
and U19887 (N_19887,N_19720,N_19741);
and U19888 (N_19888,N_19691,N_19811);
nor U19889 (N_19889,N_19823,N_19759);
or U19890 (N_19890,N_19819,N_19798);
xor U19891 (N_19891,N_19698,N_19816);
nor U19892 (N_19892,N_19748,N_19808);
nand U19893 (N_19893,N_19753,N_19749);
and U19894 (N_19894,N_19728,N_19685);
nor U19895 (N_19895,N_19726,N_19839);
nand U19896 (N_19896,N_19761,N_19708);
nor U19897 (N_19897,N_19737,N_19791);
and U19898 (N_19898,N_19814,N_19703);
nor U19899 (N_19899,N_19821,N_19746);
nand U19900 (N_19900,N_19769,N_19787);
nand U19901 (N_19901,N_19723,N_19776);
nand U19902 (N_19902,N_19732,N_19687);
nor U19903 (N_19903,N_19810,N_19770);
or U19904 (N_19904,N_19784,N_19833);
nand U19905 (N_19905,N_19736,N_19820);
or U19906 (N_19906,N_19795,N_19722);
nand U19907 (N_19907,N_19701,N_19790);
nor U19908 (N_19908,N_19750,N_19724);
or U19909 (N_19909,N_19762,N_19829);
or U19910 (N_19910,N_19689,N_19800);
and U19911 (N_19911,N_19742,N_19774);
and U19912 (N_19912,N_19694,N_19797);
nor U19913 (N_19913,N_19824,N_19690);
nor U19914 (N_19914,N_19785,N_19727);
xnor U19915 (N_19915,N_19815,N_19835);
or U19916 (N_19916,N_19744,N_19729);
nor U19917 (N_19917,N_19693,N_19717);
xnor U19918 (N_19918,N_19799,N_19813);
or U19919 (N_19919,N_19786,N_19836);
or U19920 (N_19920,N_19742,N_19779);
and U19921 (N_19921,N_19711,N_19724);
nand U19922 (N_19922,N_19784,N_19752);
xnor U19923 (N_19923,N_19837,N_19686);
and U19924 (N_19924,N_19838,N_19834);
or U19925 (N_19925,N_19771,N_19722);
or U19926 (N_19926,N_19831,N_19803);
nand U19927 (N_19927,N_19815,N_19740);
nand U19928 (N_19928,N_19808,N_19817);
nand U19929 (N_19929,N_19782,N_19770);
xnor U19930 (N_19930,N_19701,N_19815);
or U19931 (N_19931,N_19769,N_19763);
nor U19932 (N_19932,N_19747,N_19682);
nor U19933 (N_19933,N_19789,N_19820);
or U19934 (N_19934,N_19817,N_19746);
nor U19935 (N_19935,N_19696,N_19786);
nor U19936 (N_19936,N_19725,N_19813);
or U19937 (N_19937,N_19774,N_19798);
nor U19938 (N_19938,N_19810,N_19802);
or U19939 (N_19939,N_19749,N_19706);
and U19940 (N_19940,N_19784,N_19689);
nand U19941 (N_19941,N_19689,N_19745);
or U19942 (N_19942,N_19831,N_19829);
or U19943 (N_19943,N_19769,N_19794);
or U19944 (N_19944,N_19722,N_19755);
nor U19945 (N_19945,N_19732,N_19756);
nor U19946 (N_19946,N_19834,N_19805);
nor U19947 (N_19947,N_19776,N_19706);
and U19948 (N_19948,N_19690,N_19770);
nor U19949 (N_19949,N_19725,N_19711);
nor U19950 (N_19950,N_19823,N_19694);
xor U19951 (N_19951,N_19767,N_19711);
nor U19952 (N_19952,N_19783,N_19696);
nor U19953 (N_19953,N_19760,N_19763);
or U19954 (N_19954,N_19715,N_19820);
nand U19955 (N_19955,N_19712,N_19822);
or U19956 (N_19956,N_19702,N_19741);
nand U19957 (N_19957,N_19724,N_19734);
and U19958 (N_19958,N_19814,N_19732);
xnor U19959 (N_19959,N_19731,N_19693);
or U19960 (N_19960,N_19719,N_19684);
or U19961 (N_19961,N_19772,N_19696);
and U19962 (N_19962,N_19825,N_19739);
and U19963 (N_19963,N_19747,N_19708);
and U19964 (N_19964,N_19702,N_19829);
xnor U19965 (N_19965,N_19839,N_19763);
or U19966 (N_19966,N_19696,N_19768);
and U19967 (N_19967,N_19828,N_19744);
nand U19968 (N_19968,N_19812,N_19756);
or U19969 (N_19969,N_19703,N_19711);
and U19970 (N_19970,N_19771,N_19729);
nand U19971 (N_19971,N_19802,N_19826);
or U19972 (N_19972,N_19809,N_19747);
nor U19973 (N_19973,N_19737,N_19754);
and U19974 (N_19974,N_19817,N_19814);
and U19975 (N_19975,N_19685,N_19832);
and U19976 (N_19976,N_19833,N_19811);
nand U19977 (N_19977,N_19694,N_19698);
and U19978 (N_19978,N_19810,N_19789);
nor U19979 (N_19979,N_19723,N_19819);
or U19980 (N_19980,N_19763,N_19796);
and U19981 (N_19981,N_19801,N_19768);
or U19982 (N_19982,N_19803,N_19817);
or U19983 (N_19983,N_19754,N_19685);
nand U19984 (N_19984,N_19720,N_19709);
nand U19985 (N_19985,N_19778,N_19839);
nor U19986 (N_19986,N_19717,N_19798);
or U19987 (N_19987,N_19777,N_19813);
and U19988 (N_19988,N_19704,N_19778);
nor U19989 (N_19989,N_19705,N_19723);
nor U19990 (N_19990,N_19825,N_19711);
nand U19991 (N_19991,N_19709,N_19746);
or U19992 (N_19992,N_19703,N_19682);
nor U19993 (N_19993,N_19710,N_19727);
and U19994 (N_19994,N_19797,N_19702);
nor U19995 (N_19995,N_19839,N_19814);
nor U19996 (N_19996,N_19697,N_19770);
and U19997 (N_19997,N_19713,N_19718);
and U19998 (N_19998,N_19739,N_19696);
nand U19999 (N_19999,N_19684,N_19787);
nand UO_0 (O_0,N_19964,N_19979);
and UO_1 (O_1,N_19956,N_19845);
or UO_2 (O_2,N_19885,N_19933);
nor UO_3 (O_3,N_19993,N_19897);
nor UO_4 (O_4,N_19983,N_19977);
or UO_5 (O_5,N_19867,N_19930);
nor UO_6 (O_6,N_19940,N_19972);
xnor UO_7 (O_7,N_19973,N_19911);
and UO_8 (O_8,N_19880,N_19939);
and UO_9 (O_9,N_19941,N_19970);
and UO_10 (O_10,N_19944,N_19948);
or UO_11 (O_11,N_19987,N_19986);
nand UO_12 (O_12,N_19869,N_19998);
nand UO_13 (O_13,N_19886,N_19932);
xor UO_14 (O_14,N_19990,N_19892);
and UO_15 (O_15,N_19859,N_19848);
nor UO_16 (O_16,N_19863,N_19954);
nor UO_17 (O_17,N_19900,N_19996);
nand UO_18 (O_18,N_19898,N_19934);
xor UO_19 (O_19,N_19881,N_19883);
xnor UO_20 (O_20,N_19920,N_19899);
nand UO_21 (O_21,N_19908,N_19893);
nor UO_22 (O_22,N_19874,N_19955);
nor UO_23 (O_23,N_19976,N_19852);
and UO_24 (O_24,N_19957,N_19992);
or UO_25 (O_25,N_19936,N_19914);
nand UO_26 (O_26,N_19887,N_19884);
and UO_27 (O_27,N_19862,N_19858);
or UO_28 (O_28,N_19844,N_19966);
or UO_29 (O_29,N_19925,N_19907);
nor UO_30 (O_30,N_19906,N_19951);
nand UO_31 (O_31,N_19994,N_19963);
xnor UO_32 (O_32,N_19988,N_19856);
nor UO_33 (O_33,N_19913,N_19849);
nand UO_34 (O_34,N_19919,N_19857);
and UO_35 (O_35,N_19952,N_19995);
nor UO_36 (O_36,N_19937,N_19922);
and UO_37 (O_37,N_19926,N_19910);
nor UO_38 (O_38,N_19864,N_19962);
nor UO_39 (O_39,N_19890,N_19905);
or UO_40 (O_40,N_19841,N_19980);
and UO_41 (O_41,N_19846,N_19982);
and UO_42 (O_42,N_19974,N_19969);
nor UO_43 (O_43,N_19959,N_19923);
nand UO_44 (O_44,N_19921,N_19953);
and UO_45 (O_45,N_19927,N_19918);
nor UO_46 (O_46,N_19978,N_19968);
nand UO_47 (O_47,N_19871,N_19855);
or UO_48 (O_48,N_19938,N_19868);
nand UO_49 (O_49,N_19958,N_19928);
nor UO_50 (O_50,N_19971,N_19967);
or UO_51 (O_51,N_19985,N_19960);
and UO_52 (O_52,N_19997,N_19989);
nand UO_53 (O_53,N_19894,N_19861);
and UO_54 (O_54,N_19877,N_19931);
xnor UO_55 (O_55,N_19870,N_19854);
nor UO_56 (O_56,N_19895,N_19999);
or UO_57 (O_57,N_19949,N_19909);
or UO_58 (O_58,N_19860,N_19946);
and UO_59 (O_59,N_19902,N_19842);
and UO_60 (O_60,N_19876,N_19984);
nand UO_61 (O_61,N_19942,N_19850);
or UO_62 (O_62,N_19853,N_19903);
xnor UO_63 (O_63,N_19879,N_19961);
and UO_64 (O_64,N_19929,N_19847);
and UO_65 (O_65,N_19891,N_19947);
nand UO_66 (O_66,N_19896,N_19917);
and UO_67 (O_67,N_19873,N_19866);
nor UO_68 (O_68,N_19865,N_19935);
nor UO_69 (O_69,N_19889,N_19912);
or UO_70 (O_70,N_19904,N_19975);
and UO_71 (O_71,N_19916,N_19840);
nand UO_72 (O_72,N_19872,N_19950);
and UO_73 (O_73,N_19915,N_19991);
nor UO_74 (O_74,N_19878,N_19981);
xnor UO_75 (O_75,N_19965,N_19924);
nor UO_76 (O_76,N_19851,N_19875);
nand UO_77 (O_77,N_19882,N_19901);
xor UO_78 (O_78,N_19945,N_19888);
xnor UO_79 (O_79,N_19843,N_19943);
or UO_80 (O_80,N_19948,N_19884);
or UO_81 (O_81,N_19946,N_19935);
or UO_82 (O_82,N_19990,N_19844);
or UO_83 (O_83,N_19963,N_19908);
nor UO_84 (O_84,N_19975,N_19985);
and UO_85 (O_85,N_19937,N_19872);
nand UO_86 (O_86,N_19846,N_19988);
and UO_87 (O_87,N_19903,N_19851);
nand UO_88 (O_88,N_19909,N_19900);
nor UO_89 (O_89,N_19985,N_19895);
nand UO_90 (O_90,N_19938,N_19880);
or UO_91 (O_91,N_19971,N_19865);
nand UO_92 (O_92,N_19880,N_19840);
or UO_93 (O_93,N_19926,N_19990);
nor UO_94 (O_94,N_19852,N_19956);
or UO_95 (O_95,N_19925,N_19887);
nand UO_96 (O_96,N_19935,N_19949);
nor UO_97 (O_97,N_19879,N_19972);
and UO_98 (O_98,N_19932,N_19896);
or UO_99 (O_99,N_19866,N_19841);
nand UO_100 (O_100,N_19866,N_19994);
nor UO_101 (O_101,N_19951,N_19991);
xor UO_102 (O_102,N_19921,N_19930);
and UO_103 (O_103,N_19968,N_19973);
xnor UO_104 (O_104,N_19871,N_19919);
nand UO_105 (O_105,N_19879,N_19951);
xnor UO_106 (O_106,N_19970,N_19962);
and UO_107 (O_107,N_19862,N_19926);
nand UO_108 (O_108,N_19971,N_19895);
nor UO_109 (O_109,N_19994,N_19957);
nand UO_110 (O_110,N_19960,N_19945);
xor UO_111 (O_111,N_19997,N_19874);
or UO_112 (O_112,N_19883,N_19970);
nor UO_113 (O_113,N_19987,N_19984);
xnor UO_114 (O_114,N_19941,N_19995);
nand UO_115 (O_115,N_19911,N_19855);
and UO_116 (O_116,N_19918,N_19867);
and UO_117 (O_117,N_19872,N_19885);
nor UO_118 (O_118,N_19969,N_19932);
nor UO_119 (O_119,N_19898,N_19866);
or UO_120 (O_120,N_19926,N_19971);
or UO_121 (O_121,N_19945,N_19998);
nand UO_122 (O_122,N_19958,N_19892);
nand UO_123 (O_123,N_19884,N_19917);
or UO_124 (O_124,N_19912,N_19894);
or UO_125 (O_125,N_19972,N_19868);
nand UO_126 (O_126,N_19918,N_19933);
nor UO_127 (O_127,N_19899,N_19984);
nor UO_128 (O_128,N_19997,N_19852);
nor UO_129 (O_129,N_19874,N_19870);
xnor UO_130 (O_130,N_19912,N_19865);
nand UO_131 (O_131,N_19860,N_19901);
nand UO_132 (O_132,N_19980,N_19870);
xnor UO_133 (O_133,N_19841,N_19888);
nand UO_134 (O_134,N_19955,N_19884);
nor UO_135 (O_135,N_19947,N_19942);
and UO_136 (O_136,N_19908,N_19890);
and UO_137 (O_137,N_19962,N_19997);
nand UO_138 (O_138,N_19992,N_19987);
and UO_139 (O_139,N_19914,N_19876);
nand UO_140 (O_140,N_19928,N_19966);
nand UO_141 (O_141,N_19917,N_19943);
nand UO_142 (O_142,N_19924,N_19969);
nor UO_143 (O_143,N_19866,N_19964);
or UO_144 (O_144,N_19945,N_19972);
or UO_145 (O_145,N_19944,N_19971);
xor UO_146 (O_146,N_19993,N_19926);
nand UO_147 (O_147,N_19841,N_19851);
nor UO_148 (O_148,N_19973,N_19984);
nor UO_149 (O_149,N_19941,N_19987);
or UO_150 (O_150,N_19871,N_19870);
nor UO_151 (O_151,N_19916,N_19867);
nand UO_152 (O_152,N_19968,N_19921);
xor UO_153 (O_153,N_19933,N_19943);
or UO_154 (O_154,N_19939,N_19910);
nand UO_155 (O_155,N_19948,N_19974);
nand UO_156 (O_156,N_19937,N_19911);
or UO_157 (O_157,N_19885,N_19928);
nor UO_158 (O_158,N_19938,N_19890);
nand UO_159 (O_159,N_19871,N_19888);
or UO_160 (O_160,N_19870,N_19924);
and UO_161 (O_161,N_19936,N_19980);
and UO_162 (O_162,N_19961,N_19906);
and UO_163 (O_163,N_19883,N_19865);
xnor UO_164 (O_164,N_19919,N_19897);
nor UO_165 (O_165,N_19924,N_19981);
or UO_166 (O_166,N_19958,N_19967);
nand UO_167 (O_167,N_19938,N_19865);
or UO_168 (O_168,N_19914,N_19958);
and UO_169 (O_169,N_19937,N_19962);
and UO_170 (O_170,N_19990,N_19940);
and UO_171 (O_171,N_19949,N_19960);
or UO_172 (O_172,N_19875,N_19886);
and UO_173 (O_173,N_19992,N_19934);
nand UO_174 (O_174,N_19979,N_19857);
nor UO_175 (O_175,N_19854,N_19883);
or UO_176 (O_176,N_19928,N_19888);
nor UO_177 (O_177,N_19917,N_19904);
xnor UO_178 (O_178,N_19876,N_19927);
nand UO_179 (O_179,N_19912,N_19994);
nor UO_180 (O_180,N_19966,N_19879);
nand UO_181 (O_181,N_19919,N_19950);
nand UO_182 (O_182,N_19869,N_19896);
nand UO_183 (O_183,N_19890,N_19868);
and UO_184 (O_184,N_19938,N_19877);
and UO_185 (O_185,N_19947,N_19934);
and UO_186 (O_186,N_19948,N_19859);
nor UO_187 (O_187,N_19848,N_19994);
and UO_188 (O_188,N_19891,N_19911);
xor UO_189 (O_189,N_19940,N_19912);
nand UO_190 (O_190,N_19914,N_19886);
nor UO_191 (O_191,N_19957,N_19951);
nor UO_192 (O_192,N_19878,N_19873);
nand UO_193 (O_193,N_19907,N_19971);
nand UO_194 (O_194,N_19985,N_19855);
or UO_195 (O_195,N_19893,N_19970);
xor UO_196 (O_196,N_19992,N_19883);
or UO_197 (O_197,N_19955,N_19927);
nor UO_198 (O_198,N_19984,N_19925);
xor UO_199 (O_199,N_19955,N_19982);
and UO_200 (O_200,N_19923,N_19997);
or UO_201 (O_201,N_19983,N_19864);
nand UO_202 (O_202,N_19949,N_19871);
nor UO_203 (O_203,N_19975,N_19979);
or UO_204 (O_204,N_19942,N_19885);
nor UO_205 (O_205,N_19854,N_19855);
nor UO_206 (O_206,N_19875,N_19868);
or UO_207 (O_207,N_19949,N_19941);
and UO_208 (O_208,N_19939,N_19996);
or UO_209 (O_209,N_19960,N_19990);
nor UO_210 (O_210,N_19934,N_19935);
and UO_211 (O_211,N_19908,N_19935);
or UO_212 (O_212,N_19993,N_19950);
or UO_213 (O_213,N_19934,N_19872);
or UO_214 (O_214,N_19923,N_19949);
xnor UO_215 (O_215,N_19869,N_19864);
or UO_216 (O_216,N_19863,N_19930);
xnor UO_217 (O_217,N_19988,N_19857);
and UO_218 (O_218,N_19977,N_19857);
nor UO_219 (O_219,N_19851,N_19840);
or UO_220 (O_220,N_19999,N_19952);
nor UO_221 (O_221,N_19921,N_19854);
nand UO_222 (O_222,N_19854,N_19842);
nand UO_223 (O_223,N_19975,N_19880);
and UO_224 (O_224,N_19883,N_19922);
nor UO_225 (O_225,N_19851,N_19935);
nand UO_226 (O_226,N_19938,N_19914);
xnor UO_227 (O_227,N_19946,N_19888);
nand UO_228 (O_228,N_19951,N_19869);
nand UO_229 (O_229,N_19957,N_19974);
nand UO_230 (O_230,N_19994,N_19862);
xor UO_231 (O_231,N_19934,N_19962);
nand UO_232 (O_232,N_19989,N_19898);
nor UO_233 (O_233,N_19851,N_19905);
nand UO_234 (O_234,N_19850,N_19981);
or UO_235 (O_235,N_19980,N_19966);
nand UO_236 (O_236,N_19850,N_19857);
nor UO_237 (O_237,N_19975,N_19988);
and UO_238 (O_238,N_19844,N_19943);
nand UO_239 (O_239,N_19966,N_19964);
nand UO_240 (O_240,N_19893,N_19848);
nand UO_241 (O_241,N_19889,N_19958);
nor UO_242 (O_242,N_19924,N_19987);
and UO_243 (O_243,N_19938,N_19874);
or UO_244 (O_244,N_19915,N_19855);
nand UO_245 (O_245,N_19917,N_19955);
and UO_246 (O_246,N_19859,N_19886);
nor UO_247 (O_247,N_19876,N_19870);
nand UO_248 (O_248,N_19951,N_19999);
nor UO_249 (O_249,N_19973,N_19920);
nor UO_250 (O_250,N_19862,N_19988);
or UO_251 (O_251,N_19947,N_19908);
nand UO_252 (O_252,N_19853,N_19848);
nand UO_253 (O_253,N_19862,N_19889);
nand UO_254 (O_254,N_19964,N_19858);
or UO_255 (O_255,N_19982,N_19916);
xnor UO_256 (O_256,N_19867,N_19847);
nand UO_257 (O_257,N_19888,N_19913);
nand UO_258 (O_258,N_19942,N_19888);
or UO_259 (O_259,N_19954,N_19930);
or UO_260 (O_260,N_19880,N_19943);
and UO_261 (O_261,N_19997,N_19987);
and UO_262 (O_262,N_19931,N_19922);
nand UO_263 (O_263,N_19849,N_19868);
nor UO_264 (O_264,N_19923,N_19940);
nand UO_265 (O_265,N_19934,N_19919);
or UO_266 (O_266,N_19893,N_19954);
and UO_267 (O_267,N_19874,N_19859);
and UO_268 (O_268,N_19997,N_19847);
and UO_269 (O_269,N_19897,N_19922);
nor UO_270 (O_270,N_19848,N_19914);
or UO_271 (O_271,N_19932,N_19946);
nor UO_272 (O_272,N_19887,N_19943);
nand UO_273 (O_273,N_19960,N_19964);
and UO_274 (O_274,N_19846,N_19881);
and UO_275 (O_275,N_19844,N_19952);
nor UO_276 (O_276,N_19984,N_19957);
nand UO_277 (O_277,N_19916,N_19899);
and UO_278 (O_278,N_19886,N_19840);
and UO_279 (O_279,N_19844,N_19956);
and UO_280 (O_280,N_19999,N_19918);
nand UO_281 (O_281,N_19865,N_19929);
and UO_282 (O_282,N_19908,N_19927);
or UO_283 (O_283,N_19966,N_19881);
or UO_284 (O_284,N_19909,N_19857);
nand UO_285 (O_285,N_19985,N_19882);
nor UO_286 (O_286,N_19929,N_19902);
and UO_287 (O_287,N_19884,N_19848);
xnor UO_288 (O_288,N_19904,N_19919);
or UO_289 (O_289,N_19974,N_19890);
nor UO_290 (O_290,N_19959,N_19844);
xnor UO_291 (O_291,N_19875,N_19959);
xnor UO_292 (O_292,N_19894,N_19921);
or UO_293 (O_293,N_19979,N_19961);
nor UO_294 (O_294,N_19972,N_19861);
and UO_295 (O_295,N_19935,N_19996);
or UO_296 (O_296,N_19910,N_19890);
or UO_297 (O_297,N_19842,N_19933);
or UO_298 (O_298,N_19880,N_19903);
and UO_299 (O_299,N_19929,N_19924);
and UO_300 (O_300,N_19968,N_19993);
or UO_301 (O_301,N_19937,N_19975);
nor UO_302 (O_302,N_19911,N_19933);
and UO_303 (O_303,N_19880,N_19922);
or UO_304 (O_304,N_19952,N_19875);
nand UO_305 (O_305,N_19993,N_19997);
nand UO_306 (O_306,N_19969,N_19964);
nand UO_307 (O_307,N_19896,N_19944);
and UO_308 (O_308,N_19865,N_19994);
nand UO_309 (O_309,N_19994,N_19943);
or UO_310 (O_310,N_19866,N_19850);
nand UO_311 (O_311,N_19860,N_19847);
and UO_312 (O_312,N_19979,N_19887);
or UO_313 (O_313,N_19937,N_19898);
and UO_314 (O_314,N_19932,N_19963);
nor UO_315 (O_315,N_19932,N_19928);
xnor UO_316 (O_316,N_19939,N_19893);
nand UO_317 (O_317,N_19921,N_19966);
or UO_318 (O_318,N_19932,N_19877);
or UO_319 (O_319,N_19920,N_19881);
or UO_320 (O_320,N_19919,N_19844);
nor UO_321 (O_321,N_19845,N_19935);
nand UO_322 (O_322,N_19869,N_19994);
nand UO_323 (O_323,N_19884,N_19842);
and UO_324 (O_324,N_19991,N_19874);
or UO_325 (O_325,N_19951,N_19915);
or UO_326 (O_326,N_19847,N_19973);
or UO_327 (O_327,N_19964,N_19953);
and UO_328 (O_328,N_19961,N_19919);
or UO_329 (O_329,N_19880,N_19876);
and UO_330 (O_330,N_19964,N_19973);
and UO_331 (O_331,N_19840,N_19948);
nor UO_332 (O_332,N_19932,N_19878);
and UO_333 (O_333,N_19860,N_19984);
nor UO_334 (O_334,N_19895,N_19916);
or UO_335 (O_335,N_19973,N_19965);
or UO_336 (O_336,N_19849,N_19949);
nand UO_337 (O_337,N_19841,N_19970);
and UO_338 (O_338,N_19937,N_19848);
nand UO_339 (O_339,N_19998,N_19975);
nand UO_340 (O_340,N_19882,N_19989);
or UO_341 (O_341,N_19944,N_19881);
xnor UO_342 (O_342,N_19897,N_19958);
or UO_343 (O_343,N_19957,N_19887);
nand UO_344 (O_344,N_19989,N_19904);
nor UO_345 (O_345,N_19884,N_19924);
nand UO_346 (O_346,N_19946,N_19973);
and UO_347 (O_347,N_19994,N_19845);
nor UO_348 (O_348,N_19852,N_19874);
nor UO_349 (O_349,N_19870,N_19855);
and UO_350 (O_350,N_19943,N_19860);
and UO_351 (O_351,N_19982,N_19993);
nor UO_352 (O_352,N_19852,N_19856);
or UO_353 (O_353,N_19981,N_19906);
nand UO_354 (O_354,N_19932,N_19964);
and UO_355 (O_355,N_19890,N_19986);
nand UO_356 (O_356,N_19943,N_19850);
nor UO_357 (O_357,N_19865,N_19966);
nand UO_358 (O_358,N_19903,N_19902);
nor UO_359 (O_359,N_19846,N_19909);
nor UO_360 (O_360,N_19845,N_19896);
nand UO_361 (O_361,N_19937,N_19926);
xnor UO_362 (O_362,N_19990,N_19981);
or UO_363 (O_363,N_19884,N_19984);
xor UO_364 (O_364,N_19863,N_19994);
or UO_365 (O_365,N_19948,N_19880);
and UO_366 (O_366,N_19927,N_19951);
xnor UO_367 (O_367,N_19994,N_19975);
nand UO_368 (O_368,N_19978,N_19951);
nand UO_369 (O_369,N_19951,N_19884);
nor UO_370 (O_370,N_19967,N_19987);
and UO_371 (O_371,N_19843,N_19886);
nand UO_372 (O_372,N_19980,N_19851);
nand UO_373 (O_373,N_19847,N_19879);
nor UO_374 (O_374,N_19962,N_19942);
and UO_375 (O_375,N_19956,N_19926);
nor UO_376 (O_376,N_19996,N_19948);
or UO_377 (O_377,N_19934,N_19983);
or UO_378 (O_378,N_19927,N_19989);
or UO_379 (O_379,N_19874,N_19971);
nand UO_380 (O_380,N_19860,N_19867);
nor UO_381 (O_381,N_19843,N_19847);
and UO_382 (O_382,N_19974,N_19909);
nand UO_383 (O_383,N_19980,N_19862);
nor UO_384 (O_384,N_19844,N_19982);
or UO_385 (O_385,N_19840,N_19876);
or UO_386 (O_386,N_19973,N_19954);
or UO_387 (O_387,N_19975,N_19888);
nor UO_388 (O_388,N_19847,N_19865);
or UO_389 (O_389,N_19901,N_19880);
nand UO_390 (O_390,N_19930,N_19999);
nand UO_391 (O_391,N_19873,N_19933);
or UO_392 (O_392,N_19982,N_19973);
nor UO_393 (O_393,N_19959,N_19944);
nor UO_394 (O_394,N_19979,N_19864);
or UO_395 (O_395,N_19991,N_19876);
xnor UO_396 (O_396,N_19946,N_19845);
or UO_397 (O_397,N_19893,N_19998);
nand UO_398 (O_398,N_19887,N_19971);
and UO_399 (O_399,N_19922,N_19911);
nor UO_400 (O_400,N_19870,N_19968);
nand UO_401 (O_401,N_19841,N_19862);
or UO_402 (O_402,N_19976,N_19975);
or UO_403 (O_403,N_19871,N_19849);
or UO_404 (O_404,N_19971,N_19870);
nor UO_405 (O_405,N_19944,N_19857);
nor UO_406 (O_406,N_19879,N_19984);
and UO_407 (O_407,N_19844,N_19964);
xor UO_408 (O_408,N_19993,N_19862);
nor UO_409 (O_409,N_19925,N_19961);
and UO_410 (O_410,N_19927,N_19861);
and UO_411 (O_411,N_19987,N_19970);
and UO_412 (O_412,N_19938,N_19946);
or UO_413 (O_413,N_19990,N_19967);
and UO_414 (O_414,N_19962,N_19853);
nor UO_415 (O_415,N_19920,N_19898);
or UO_416 (O_416,N_19990,N_19927);
or UO_417 (O_417,N_19919,N_19958);
nor UO_418 (O_418,N_19863,N_19998);
or UO_419 (O_419,N_19945,N_19982);
nor UO_420 (O_420,N_19884,N_19941);
and UO_421 (O_421,N_19933,N_19903);
xor UO_422 (O_422,N_19880,N_19972);
nand UO_423 (O_423,N_19991,N_19965);
nand UO_424 (O_424,N_19851,N_19995);
nand UO_425 (O_425,N_19869,N_19963);
or UO_426 (O_426,N_19914,N_19917);
or UO_427 (O_427,N_19861,N_19853);
nand UO_428 (O_428,N_19967,N_19871);
nor UO_429 (O_429,N_19859,N_19912);
or UO_430 (O_430,N_19943,N_19854);
or UO_431 (O_431,N_19875,N_19968);
nor UO_432 (O_432,N_19936,N_19869);
and UO_433 (O_433,N_19853,N_19990);
or UO_434 (O_434,N_19956,N_19919);
and UO_435 (O_435,N_19950,N_19953);
nand UO_436 (O_436,N_19925,N_19979);
and UO_437 (O_437,N_19875,N_19862);
xor UO_438 (O_438,N_19977,N_19903);
and UO_439 (O_439,N_19997,N_19891);
nand UO_440 (O_440,N_19973,N_19978);
and UO_441 (O_441,N_19929,N_19846);
nor UO_442 (O_442,N_19921,N_19856);
nor UO_443 (O_443,N_19910,N_19934);
and UO_444 (O_444,N_19906,N_19968);
nand UO_445 (O_445,N_19984,N_19983);
or UO_446 (O_446,N_19912,N_19981);
or UO_447 (O_447,N_19932,N_19913);
xor UO_448 (O_448,N_19950,N_19893);
or UO_449 (O_449,N_19844,N_19948);
xnor UO_450 (O_450,N_19942,N_19914);
xnor UO_451 (O_451,N_19980,N_19947);
and UO_452 (O_452,N_19894,N_19885);
nor UO_453 (O_453,N_19878,N_19884);
and UO_454 (O_454,N_19886,N_19861);
nor UO_455 (O_455,N_19849,N_19945);
or UO_456 (O_456,N_19893,N_19991);
or UO_457 (O_457,N_19873,N_19864);
nand UO_458 (O_458,N_19866,N_19917);
nor UO_459 (O_459,N_19970,N_19978);
nand UO_460 (O_460,N_19897,N_19990);
nor UO_461 (O_461,N_19958,N_19878);
or UO_462 (O_462,N_19882,N_19958);
or UO_463 (O_463,N_19898,N_19874);
nor UO_464 (O_464,N_19929,N_19979);
nor UO_465 (O_465,N_19883,N_19917);
nand UO_466 (O_466,N_19860,N_19925);
and UO_467 (O_467,N_19976,N_19914);
or UO_468 (O_468,N_19864,N_19981);
xnor UO_469 (O_469,N_19995,N_19973);
or UO_470 (O_470,N_19921,N_19998);
and UO_471 (O_471,N_19934,N_19858);
or UO_472 (O_472,N_19961,N_19896);
or UO_473 (O_473,N_19909,N_19887);
and UO_474 (O_474,N_19987,N_19890);
and UO_475 (O_475,N_19914,N_19918);
xnor UO_476 (O_476,N_19994,N_19936);
or UO_477 (O_477,N_19918,N_19953);
nor UO_478 (O_478,N_19959,N_19904);
nor UO_479 (O_479,N_19860,N_19921);
nor UO_480 (O_480,N_19868,N_19894);
or UO_481 (O_481,N_19868,N_19949);
nor UO_482 (O_482,N_19925,N_19974);
or UO_483 (O_483,N_19937,N_19849);
nand UO_484 (O_484,N_19988,N_19904);
and UO_485 (O_485,N_19949,N_19843);
nor UO_486 (O_486,N_19857,N_19927);
nand UO_487 (O_487,N_19929,N_19888);
nand UO_488 (O_488,N_19863,N_19969);
or UO_489 (O_489,N_19927,N_19895);
or UO_490 (O_490,N_19900,N_19954);
nand UO_491 (O_491,N_19989,N_19991);
nand UO_492 (O_492,N_19915,N_19872);
nand UO_493 (O_493,N_19950,N_19962);
xor UO_494 (O_494,N_19977,N_19937);
and UO_495 (O_495,N_19956,N_19916);
or UO_496 (O_496,N_19972,N_19984);
xor UO_497 (O_497,N_19872,N_19972);
nor UO_498 (O_498,N_19924,N_19857);
nand UO_499 (O_499,N_19879,N_19948);
nand UO_500 (O_500,N_19926,N_19934);
and UO_501 (O_501,N_19856,N_19858);
or UO_502 (O_502,N_19877,N_19888);
or UO_503 (O_503,N_19885,N_19905);
nand UO_504 (O_504,N_19929,N_19880);
xor UO_505 (O_505,N_19891,N_19869);
nand UO_506 (O_506,N_19948,N_19901);
and UO_507 (O_507,N_19921,N_19862);
and UO_508 (O_508,N_19971,N_19845);
or UO_509 (O_509,N_19865,N_19965);
nor UO_510 (O_510,N_19963,N_19943);
xnor UO_511 (O_511,N_19947,N_19922);
and UO_512 (O_512,N_19907,N_19929);
nor UO_513 (O_513,N_19902,N_19991);
nand UO_514 (O_514,N_19914,N_19850);
and UO_515 (O_515,N_19989,N_19944);
or UO_516 (O_516,N_19936,N_19897);
nand UO_517 (O_517,N_19942,N_19939);
and UO_518 (O_518,N_19983,N_19952);
or UO_519 (O_519,N_19941,N_19846);
nand UO_520 (O_520,N_19843,N_19887);
xor UO_521 (O_521,N_19917,N_19928);
and UO_522 (O_522,N_19840,N_19984);
nor UO_523 (O_523,N_19905,N_19867);
nand UO_524 (O_524,N_19898,N_19929);
nand UO_525 (O_525,N_19972,N_19858);
xor UO_526 (O_526,N_19950,N_19992);
and UO_527 (O_527,N_19876,N_19921);
nand UO_528 (O_528,N_19977,N_19861);
nand UO_529 (O_529,N_19946,N_19998);
xor UO_530 (O_530,N_19853,N_19977);
or UO_531 (O_531,N_19952,N_19882);
nand UO_532 (O_532,N_19958,N_19868);
nor UO_533 (O_533,N_19864,N_19877);
and UO_534 (O_534,N_19982,N_19964);
nand UO_535 (O_535,N_19956,N_19901);
and UO_536 (O_536,N_19927,N_19841);
xnor UO_537 (O_537,N_19904,N_19911);
nand UO_538 (O_538,N_19962,N_19846);
and UO_539 (O_539,N_19890,N_19934);
and UO_540 (O_540,N_19870,N_19900);
xnor UO_541 (O_541,N_19938,N_19983);
and UO_542 (O_542,N_19983,N_19926);
nand UO_543 (O_543,N_19942,N_19937);
nor UO_544 (O_544,N_19860,N_19955);
or UO_545 (O_545,N_19899,N_19858);
xor UO_546 (O_546,N_19860,N_19870);
nand UO_547 (O_547,N_19860,N_19923);
and UO_548 (O_548,N_19940,N_19928);
or UO_549 (O_549,N_19902,N_19871);
nor UO_550 (O_550,N_19862,N_19943);
or UO_551 (O_551,N_19895,N_19880);
nand UO_552 (O_552,N_19978,N_19843);
or UO_553 (O_553,N_19885,N_19993);
xnor UO_554 (O_554,N_19993,N_19856);
and UO_555 (O_555,N_19913,N_19851);
and UO_556 (O_556,N_19936,N_19929);
nor UO_557 (O_557,N_19901,N_19871);
xnor UO_558 (O_558,N_19996,N_19848);
nand UO_559 (O_559,N_19970,N_19953);
nand UO_560 (O_560,N_19973,N_19880);
xnor UO_561 (O_561,N_19896,N_19906);
nand UO_562 (O_562,N_19948,N_19954);
xnor UO_563 (O_563,N_19949,N_19873);
and UO_564 (O_564,N_19905,N_19949);
nor UO_565 (O_565,N_19901,N_19846);
or UO_566 (O_566,N_19907,N_19846);
and UO_567 (O_567,N_19939,N_19973);
nor UO_568 (O_568,N_19863,N_19971);
or UO_569 (O_569,N_19997,N_19870);
nor UO_570 (O_570,N_19945,N_19994);
nor UO_571 (O_571,N_19974,N_19848);
nor UO_572 (O_572,N_19857,N_19986);
xnor UO_573 (O_573,N_19920,N_19935);
nor UO_574 (O_574,N_19894,N_19985);
nand UO_575 (O_575,N_19860,N_19937);
xor UO_576 (O_576,N_19981,N_19858);
nor UO_577 (O_577,N_19846,N_19940);
xor UO_578 (O_578,N_19981,N_19982);
or UO_579 (O_579,N_19865,N_19997);
or UO_580 (O_580,N_19982,N_19948);
nand UO_581 (O_581,N_19954,N_19855);
or UO_582 (O_582,N_19939,N_19990);
and UO_583 (O_583,N_19884,N_19986);
or UO_584 (O_584,N_19930,N_19945);
nor UO_585 (O_585,N_19895,N_19963);
nor UO_586 (O_586,N_19983,N_19853);
nor UO_587 (O_587,N_19919,N_19949);
nand UO_588 (O_588,N_19901,N_19873);
nand UO_589 (O_589,N_19923,N_19908);
nor UO_590 (O_590,N_19864,N_19975);
nor UO_591 (O_591,N_19925,N_19893);
or UO_592 (O_592,N_19861,N_19918);
nand UO_593 (O_593,N_19845,N_19870);
and UO_594 (O_594,N_19868,N_19879);
or UO_595 (O_595,N_19965,N_19844);
xnor UO_596 (O_596,N_19981,N_19891);
and UO_597 (O_597,N_19868,N_19932);
nor UO_598 (O_598,N_19927,N_19867);
and UO_599 (O_599,N_19915,N_19930);
and UO_600 (O_600,N_19841,N_19936);
nand UO_601 (O_601,N_19893,N_19964);
nor UO_602 (O_602,N_19960,N_19984);
and UO_603 (O_603,N_19906,N_19917);
nand UO_604 (O_604,N_19902,N_19893);
nor UO_605 (O_605,N_19840,N_19957);
and UO_606 (O_606,N_19898,N_19888);
nand UO_607 (O_607,N_19986,N_19893);
nand UO_608 (O_608,N_19866,N_19858);
or UO_609 (O_609,N_19986,N_19935);
xor UO_610 (O_610,N_19873,N_19990);
nand UO_611 (O_611,N_19863,N_19909);
nor UO_612 (O_612,N_19995,N_19939);
and UO_613 (O_613,N_19915,N_19879);
nor UO_614 (O_614,N_19885,N_19967);
nor UO_615 (O_615,N_19916,N_19928);
nor UO_616 (O_616,N_19977,N_19944);
nand UO_617 (O_617,N_19923,N_19904);
nor UO_618 (O_618,N_19880,N_19992);
nand UO_619 (O_619,N_19979,N_19942);
nor UO_620 (O_620,N_19896,N_19855);
nor UO_621 (O_621,N_19936,N_19962);
nor UO_622 (O_622,N_19908,N_19929);
and UO_623 (O_623,N_19996,N_19954);
nor UO_624 (O_624,N_19929,N_19893);
or UO_625 (O_625,N_19947,N_19985);
nand UO_626 (O_626,N_19856,N_19867);
nand UO_627 (O_627,N_19946,N_19864);
nor UO_628 (O_628,N_19973,N_19857);
nor UO_629 (O_629,N_19985,N_19926);
or UO_630 (O_630,N_19881,N_19916);
nor UO_631 (O_631,N_19969,N_19840);
xnor UO_632 (O_632,N_19842,N_19851);
or UO_633 (O_633,N_19855,N_19992);
nor UO_634 (O_634,N_19935,N_19980);
nor UO_635 (O_635,N_19961,N_19869);
or UO_636 (O_636,N_19860,N_19889);
nand UO_637 (O_637,N_19991,N_19918);
nand UO_638 (O_638,N_19854,N_19882);
nor UO_639 (O_639,N_19886,N_19937);
nor UO_640 (O_640,N_19889,N_19971);
nand UO_641 (O_641,N_19892,N_19957);
nand UO_642 (O_642,N_19958,N_19883);
nor UO_643 (O_643,N_19962,N_19871);
nor UO_644 (O_644,N_19864,N_19851);
and UO_645 (O_645,N_19856,N_19999);
nor UO_646 (O_646,N_19921,N_19989);
or UO_647 (O_647,N_19844,N_19973);
and UO_648 (O_648,N_19969,N_19910);
nor UO_649 (O_649,N_19979,N_19852);
nor UO_650 (O_650,N_19993,N_19908);
nand UO_651 (O_651,N_19849,N_19878);
nand UO_652 (O_652,N_19877,N_19924);
or UO_653 (O_653,N_19890,N_19867);
nand UO_654 (O_654,N_19978,N_19960);
nor UO_655 (O_655,N_19943,N_19845);
nor UO_656 (O_656,N_19981,N_19992);
and UO_657 (O_657,N_19916,N_19894);
nand UO_658 (O_658,N_19861,N_19980);
xnor UO_659 (O_659,N_19882,N_19929);
nor UO_660 (O_660,N_19921,N_19883);
and UO_661 (O_661,N_19959,N_19902);
nand UO_662 (O_662,N_19991,N_19941);
nand UO_663 (O_663,N_19873,N_19982);
and UO_664 (O_664,N_19976,N_19961);
and UO_665 (O_665,N_19953,N_19956);
nor UO_666 (O_666,N_19935,N_19900);
xnor UO_667 (O_667,N_19932,N_19925);
or UO_668 (O_668,N_19841,N_19968);
and UO_669 (O_669,N_19963,N_19937);
nor UO_670 (O_670,N_19848,N_19952);
nand UO_671 (O_671,N_19897,N_19971);
and UO_672 (O_672,N_19847,N_19951);
and UO_673 (O_673,N_19872,N_19941);
xnor UO_674 (O_674,N_19900,N_19999);
or UO_675 (O_675,N_19891,N_19957);
nor UO_676 (O_676,N_19990,N_19944);
xnor UO_677 (O_677,N_19982,N_19875);
nor UO_678 (O_678,N_19866,N_19871);
nand UO_679 (O_679,N_19933,N_19946);
nor UO_680 (O_680,N_19983,N_19842);
and UO_681 (O_681,N_19990,N_19889);
nor UO_682 (O_682,N_19880,N_19867);
or UO_683 (O_683,N_19952,N_19945);
or UO_684 (O_684,N_19847,N_19924);
nand UO_685 (O_685,N_19987,N_19897);
or UO_686 (O_686,N_19931,N_19965);
nand UO_687 (O_687,N_19866,N_19929);
nor UO_688 (O_688,N_19988,N_19998);
and UO_689 (O_689,N_19954,N_19936);
nor UO_690 (O_690,N_19944,N_19865);
nor UO_691 (O_691,N_19911,N_19994);
nor UO_692 (O_692,N_19977,N_19975);
and UO_693 (O_693,N_19908,N_19856);
nor UO_694 (O_694,N_19890,N_19921);
or UO_695 (O_695,N_19974,N_19868);
nand UO_696 (O_696,N_19923,N_19883);
or UO_697 (O_697,N_19973,N_19882);
nor UO_698 (O_698,N_19844,N_19845);
and UO_699 (O_699,N_19952,N_19973);
xor UO_700 (O_700,N_19849,N_19906);
and UO_701 (O_701,N_19944,N_19983);
nor UO_702 (O_702,N_19846,N_19882);
nand UO_703 (O_703,N_19900,N_19963);
nor UO_704 (O_704,N_19852,N_19900);
and UO_705 (O_705,N_19893,N_19907);
or UO_706 (O_706,N_19971,N_19938);
nor UO_707 (O_707,N_19992,N_19997);
nand UO_708 (O_708,N_19981,N_19846);
nand UO_709 (O_709,N_19880,N_19873);
or UO_710 (O_710,N_19877,N_19972);
xnor UO_711 (O_711,N_19995,N_19852);
and UO_712 (O_712,N_19947,N_19884);
or UO_713 (O_713,N_19850,N_19995);
nand UO_714 (O_714,N_19864,N_19844);
nand UO_715 (O_715,N_19934,N_19886);
or UO_716 (O_716,N_19947,N_19902);
nand UO_717 (O_717,N_19897,N_19877);
nor UO_718 (O_718,N_19983,N_19967);
nor UO_719 (O_719,N_19936,N_19973);
xnor UO_720 (O_720,N_19943,N_19906);
nand UO_721 (O_721,N_19953,N_19995);
or UO_722 (O_722,N_19932,N_19982);
nor UO_723 (O_723,N_19989,N_19915);
nand UO_724 (O_724,N_19964,N_19987);
nor UO_725 (O_725,N_19851,N_19979);
and UO_726 (O_726,N_19941,N_19955);
nand UO_727 (O_727,N_19864,N_19924);
nand UO_728 (O_728,N_19936,N_19932);
or UO_729 (O_729,N_19843,N_19926);
nand UO_730 (O_730,N_19979,N_19971);
nor UO_731 (O_731,N_19873,N_19848);
nand UO_732 (O_732,N_19900,N_19964);
nand UO_733 (O_733,N_19884,N_19928);
or UO_734 (O_734,N_19866,N_19908);
or UO_735 (O_735,N_19900,N_19955);
nand UO_736 (O_736,N_19982,N_19956);
xnor UO_737 (O_737,N_19986,N_19901);
nand UO_738 (O_738,N_19971,N_19881);
nand UO_739 (O_739,N_19896,N_19843);
or UO_740 (O_740,N_19848,N_19862);
nor UO_741 (O_741,N_19990,N_19959);
or UO_742 (O_742,N_19852,N_19897);
nor UO_743 (O_743,N_19876,N_19900);
and UO_744 (O_744,N_19903,N_19905);
nand UO_745 (O_745,N_19851,N_19953);
xor UO_746 (O_746,N_19960,N_19994);
and UO_747 (O_747,N_19895,N_19952);
nor UO_748 (O_748,N_19909,N_19925);
and UO_749 (O_749,N_19856,N_19860);
nand UO_750 (O_750,N_19958,N_19844);
nand UO_751 (O_751,N_19895,N_19935);
nand UO_752 (O_752,N_19979,N_19968);
or UO_753 (O_753,N_19952,N_19933);
nand UO_754 (O_754,N_19970,N_19911);
and UO_755 (O_755,N_19952,N_19948);
nand UO_756 (O_756,N_19948,N_19906);
or UO_757 (O_757,N_19918,N_19983);
nor UO_758 (O_758,N_19866,N_19862);
nand UO_759 (O_759,N_19937,N_19840);
nand UO_760 (O_760,N_19889,N_19953);
nor UO_761 (O_761,N_19841,N_19996);
nand UO_762 (O_762,N_19956,N_19841);
or UO_763 (O_763,N_19844,N_19875);
nand UO_764 (O_764,N_19961,N_19897);
or UO_765 (O_765,N_19971,N_19905);
nor UO_766 (O_766,N_19842,N_19903);
and UO_767 (O_767,N_19959,N_19991);
nand UO_768 (O_768,N_19897,N_19997);
or UO_769 (O_769,N_19970,N_19857);
and UO_770 (O_770,N_19961,N_19846);
and UO_771 (O_771,N_19864,N_19910);
or UO_772 (O_772,N_19947,N_19926);
nor UO_773 (O_773,N_19896,N_19900);
and UO_774 (O_774,N_19841,N_19975);
or UO_775 (O_775,N_19881,N_19885);
or UO_776 (O_776,N_19981,N_19971);
nor UO_777 (O_777,N_19989,N_19877);
xor UO_778 (O_778,N_19911,N_19870);
and UO_779 (O_779,N_19879,N_19873);
nand UO_780 (O_780,N_19845,N_19880);
or UO_781 (O_781,N_19890,N_19882);
nand UO_782 (O_782,N_19929,N_19964);
or UO_783 (O_783,N_19981,N_19902);
and UO_784 (O_784,N_19986,N_19998);
nand UO_785 (O_785,N_19886,N_19929);
and UO_786 (O_786,N_19867,N_19865);
or UO_787 (O_787,N_19980,N_19894);
or UO_788 (O_788,N_19906,N_19924);
and UO_789 (O_789,N_19884,N_19879);
nor UO_790 (O_790,N_19948,N_19947);
and UO_791 (O_791,N_19950,N_19981);
or UO_792 (O_792,N_19911,N_19883);
and UO_793 (O_793,N_19944,N_19882);
nand UO_794 (O_794,N_19862,N_19935);
xor UO_795 (O_795,N_19938,N_19974);
or UO_796 (O_796,N_19998,N_19884);
or UO_797 (O_797,N_19921,N_19913);
xor UO_798 (O_798,N_19873,N_19845);
nor UO_799 (O_799,N_19908,N_19841);
and UO_800 (O_800,N_19856,N_19890);
xnor UO_801 (O_801,N_19940,N_19840);
xnor UO_802 (O_802,N_19954,N_19858);
or UO_803 (O_803,N_19907,N_19851);
xnor UO_804 (O_804,N_19860,N_19895);
or UO_805 (O_805,N_19900,N_19880);
nand UO_806 (O_806,N_19947,N_19916);
xor UO_807 (O_807,N_19875,N_19977);
and UO_808 (O_808,N_19994,N_19906);
nor UO_809 (O_809,N_19848,N_19876);
and UO_810 (O_810,N_19893,N_19861);
xnor UO_811 (O_811,N_19869,N_19952);
nand UO_812 (O_812,N_19998,N_19919);
nor UO_813 (O_813,N_19858,N_19871);
xor UO_814 (O_814,N_19910,N_19845);
nor UO_815 (O_815,N_19846,N_19975);
or UO_816 (O_816,N_19869,N_19907);
xnor UO_817 (O_817,N_19910,N_19918);
nand UO_818 (O_818,N_19925,N_19851);
and UO_819 (O_819,N_19962,N_19928);
and UO_820 (O_820,N_19919,N_19848);
or UO_821 (O_821,N_19921,N_19936);
nor UO_822 (O_822,N_19885,N_19859);
nand UO_823 (O_823,N_19985,N_19993);
nand UO_824 (O_824,N_19980,N_19868);
or UO_825 (O_825,N_19946,N_19974);
or UO_826 (O_826,N_19949,N_19864);
nand UO_827 (O_827,N_19993,N_19880);
or UO_828 (O_828,N_19857,N_19864);
and UO_829 (O_829,N_19905,N_19843);
and UO_830 (O_830,N_19948,N_19990);
and UO_831 (O_831,N_19896,N_19925);
nor UO_832 (O_832,N_19991,N_19945);
nor UO_833 (O_833,N_19849,N_19905);
nand UO_834 (O_834,N_19848,N_19865);
or UO_835 (O_835,N_19886,N_19865);
nor UO_836 (O_836,N_19867,N_19924);
and UO_837 (O_837,N_19911,N_19983);
or UO_838 (O_838,N_19868,N_19897);
nor UO_839 (O_839,N_19855,N_19879);
and UO_840 (O_840,N_19929,N_19961);
nand UO_841 (O_841,N_19840,N_19850);
nor UO_842 (O_842,N_19940,N_19948);
or UO_843 (O_843,N_19915,N_19905);
and UO_844 (O_844,N_19917,N_19915);
and UO_845 (O_845,N_19918,N_19841);
nor UO_846 (O_846,N_19918,N_19986);
or UO_847 (O_847,N_19844,N_19886);
and UO_848 (O_848,N_19995,N_19926);
nand UO_849 (O_849,N_19990,N_19882);
or UO_850 (O_850,N_19860,N_19979);
or UO_851 (O_851,N_19911,N_19929);
xnor UO_852 (O_852,N_19855,N_19844);
nand UO_853 (O_853,N_19949,N_19967);
nand UO_854 (O_854,N_19899,N_19948);
or UO_855 (O_855,N_19853,N_19842);
nor UO_856 (O_856,N_19906,N_19987);
nor UO_857 (O_857,N_19959,N_19852);
and UO_858 (O_858,N_19848,N_19956);
nor UO_859 (O_859,N_19941,N_19858);
nand UO_860 (O_860,N_19877,N_19911);
nand UO_861 (O_861,N_19977,N_19968);
nand UO_862 (O_862,N_19869,N_19960);
nand UO_863 (O_863,N_19846,N_19847);
nand UO_864 (O_864,N_19969,N_19975);
nand UO_865 (O_865,N_19885,N_19984);
and UO_866 (O_866,N_19901,N_19879);
nor UO_867 (O_867,N_19861,N_19898);
or UO_868 (O_868,N_19941,N_19927);
xor UO_869 (O_869,N_19851,N_19869);
xor UO_870 (O_870,N_19893,N_19870);
xnor UO_871 (O_871,N_19944,N_19874);
nand UO_872 (O_872,N_19877,N_19927);
or UO_873 (O_873,N_19949,N_19975);
nor UO_874 (O_874,N_19926,N_19931);
nand UO_875 (O_875,N_19857,N_19875);
and UO_876 (O_876,N_19940,N_19967);
and UO_877 (O_877,N_19947,N_19990);
nor UO_878 (O_878,N_19888,N_19881);
or UO_879 (O_879,N_19866,N_19869);
nand UO_880 (O_880,N_19865,N_19900);
nor UO_881 (O_881,N_19903,N_19987);
nor UO_882 (O_882,N_19992,N_19954);
and UO_883 (O_883,N_19901,N_19991);
nand UO_884 (O_884,N_19856,N_19931);
xnor UO_885 (O_885,N_19893,N_19961);
or UO_886 (O_886,N_19940,N_19857);
and UO_887 (O_887,N_19894,N_19910);
or UO_888 (O_888,N_19936,N_19842);
xor UO_889 (O_889,N_19952,N_19891);
nand UO_890 (O_890,N_19861,N_19872);
or UO_891 (O_891,N_19920,N_19863);
nor UO_892 (O_892,N_19953,N_19883);
and UO_893 (O_893,N_19952,N_19864);
or UO_894 (O_894,N_19918,N_19877);
xnor UO_895 (O_895,N_19975,N_19956);
and UO_896 (O_896,N_19991,N_19853);
nand UO_897 (O_897,N_19925,N_19993);
and UO_898 (O_898,N_19942,N_19879);
xor UO_899 (O_899,N_19976,N_19995);
nand UO_900 (O_900,N_19856,N_19952);
or UO_901 (O_901,N_19947,N_19991);
nor UO_902 (O_902,N_19878,N_19993);
nor UO_903 (O_903,N_19878,N_19841);
xnor UO_904 (O_904,N_19917,N_19902);
nand UO_905 (O_905,N_19887,N_19845);
and UO_906 (O_906,N_19875,N_19965);
xor UO_907 (O_907,N_19846,N_19928);
and UO_908 (O_908,N_19854,N_19850);
and UO_909 (O_909,N_19855,N_19936);
nand UO_910 (O_910,N_19844,N_19986);
and UO_911 (O_911,N_19894,N_19955);
or UO_912 (O_912,N_19982,N_19958);
nand UO_913 (O_913,N_19935,N_19988);
and UO_914 (O_914,N_19970,N_19982);
nand UO_915 (O_915,N_19858,N_19979);
nand UO_916 (O_916,N_19852,N_19931);
or UO_917 (O_917,N_19873,N_19974);
xnor UO_918 (O_918,N_19899,N_19913);
xnor UO_919 (O_919,N_19924,N_19872);
xor UO_920 (O_920,N_19854,N_19953);
or UO_921 (O_921,N_19977,N_19929);
nor UO_922 (O_922,N_19857,N_19881);
nand UO_923 (O_923,N_19890,N_19850);
xor UO_924 (O_924,N_19856,N_19991);
and UO_925 (O_925,N_19887,N_19965);
nand UO_926 (O_926,N_19898,N_19983);
or UO_927 (O_927,N_19990,N_19952);
xor UO_928 (O_928,N_19993,N_19976);
or UO_929 (O_929,N_19999,N_19937);
xnor UO_930 (O_930,N_19985,N_19989);
or UO_931 (O_931,N_19878,N_19842);
nand UO_932 (O_932,N_19892,N_19909);
nor UO_933 (O_933,N_19981,N_19997);
xor UO_934 (O_934,N_19880,N_19907);
nor UO_935 (O_935,N_19867,N_19923);
nor UO_936 (O_936,N_19879,N_19919);
and UO_937 (O_937,N_19856,N_19939);
or UO_938 (O_938,N_19922,N_19936);
and UO_939 (O_939,N_19874,N_19933);
nand UO_940 (O_940,N_19860,N_19875);
or UO_941 (O_941,N_19850,N_19937);
and UO_942 (O_942,N_19989,N_19941);
nor UO_943 (O_943,N_19965,N_19850);
and UO_944 (O_944,N_19996,N_19987);
nor UO_945 (O_945,N_19992,N_19971);
nor UO_946 (O_946,N_19863,N_19840);
xor UO_947 (O_947,N_19887,N_19973);
nor UO_948 (O_948,N_19966,N_19863);
and UO_949 (O_949,N_19924,N_19995);
nor UO_950 (O_950,N_19880,N_19921);
nor UO_951 (O_951,N_19969,N_19848);
nor UO_952 (O_952,N_19854,N_19975);
and UO_953 (O_953,N_19977,N_19998);
or UO_954 (O_954,N_19871,N_19937);
or UO_955 (O_955,N_19868,N_19861);
and UO_956 (O_956,N_19954,N_19972);
xnor UO_957 (O_957,N_19942,N_19895);
and UO_958 (O_958,N_19965,N_19910);
nand UO_959 (O_959,N_19944,N_19967);
nor UO_960 (O_960,N_19920,N_19988);
and UO_961 (O_961,N_19866,N_19944);
and UO_962 (O_962,N_19912,N_19918);
and UO_963 (O_963,N_19907,N_19956);
and UO_964 (O_964,N_19868,N_19874);
nand UO_965 (O_965,N_19913,N_19908);
nor UO_966 (O_966,N_19859,N_19847);
nor UO_967 (O_967,N_19977,N_19896);
and UO_968 (O_968,N_19954,N_19852);
and UO_969 (O_969,N_19878,N_19995);
nand UO_970 (O_970,N_19888,N_19978);
or UO_971 (O_971,N_19840,N_19991);
or UO_972 (O_972,N_19856,N_19963);
or UO_973 (O_973,N_19931,N_19971);
and UO_974 (O_974,N_19903,N_19983);
and UO_975 (O_975,N_19860,N_19932);
xor UO_976 (O_976,N_19905,N_19848);
nor UO_977 (O_977,N_19943,N_19871);
and UO_978 (O_978,N_19862,N_19974);
and UO_979 (O_979,N_19972,N_19893);
or UO_980 (O_980,N_19850,N_19856);
xor UO_981 (O_981,N_19975,N_19858);
nor UO_982 (O_982,N_19938,N_19867);
or UO_983 (O_983,N_19882,N_19951);
or UO_984 (O_984,N_19915,N_19893);
nor UO_985 (O_985,N_19979,N_19911);
or UO_986 (O_986,N_19960,N_19856);
nor UO_987 (O_987,N_19871,N_19875);
and UO_988 (O_988,N_19991,N_19872);
nor UO_989 (O_989,N_19893,N_19897);
nor UO_990 (O_990,N_19856,N_19943);
nor UO_991 (O_991,N_19986,N_19879);
and UO_992 (O_992,N_19935,N_19917);
xor UO_993 (O_993,N_19851,N_19951);
and UO_994 (O_994,N_19961,N_19928);
nor UO_995 (O_995,N_19924,N_19873);
nand UO_996 (O_996,N_19998,N_19864);
nand UO_997 (O_997,N_19961,N_19937);
or UO_998 (O_998,N_19846,N_19923);
nor UO_999 (O_999,N_19942,N_19970);
nor UO_1000 (O_1000,N_19894,N_19917);
and UO_1001 (O_1001,N_19956,N_19951);
and UO_1002 (O_1002,N_19972,N_19928);
nand UO_1003 (O_1003,N_19938,N_19871);
nor UO_1004 (O_1004,N_19974,N_19997);
nand UO_1005 (O_1005,N_19847,N_19884);
nor UO_1006 (O_1006,N_19896,N_19840);
or UO_1007 (O_1007,N_19993,N_19907);
and UO_1008 (O_1008,N_19843,N_19927);
nand UO_1009 (O_1009,N_19857,N_19855);
or UO_1010 (O_1010,N_19914,N_19951);
nor UO_1011 (O_1011,N_19911,N_19935);
or UO_1012 (O_1012,N_19957,N_19939);
or UO_1013 (O_1013,N_19942,N_19951);
and UO_1014 (O_1014,N_19883,N_19976);
and UO_1015 (O_1015,N_19850,N_19852);
nor UO_1016 (O_1016,N_19842,N_19855);
or UO_1017 (O_1017,N_19937,N_19925);
or UO_1018 (O_1018,N_19891,N_19879);
or UO_1019 (O_1019,N_19991,N_19907);
and UO_1020 (O_1020,N_19916,N_19975);
xnor UO_1021 (O_1021,N_19972,N_19947);
or UO_1022 (O_1022,N_19994,N_19921);
nor UO_1023 (O_1023,N_19996,N_19852);
and UO_1024 (O_1024,N_19889,N_19988);
nand UO_1025 (O_1025,N_19953,N_19929);
nand UO_1026 (O_1026,N_19965,N_19848);
and UO_1027 (O_1027,N_19971,N_19988);
nor UO_1028 (O_1028,N_19933,N_19880);
and UO_1029 (O_1029,N_19931,N_19994);
nor UO_1030 (O_1030,N_19983,N_19845);
nand UO_1031 (O_1031,N_19957,N_19846);
or UO_1032 (O_1032,N_19871,N_19980);
xor UO_1033 (O_1033,N_19871,N_19872);
or UO_1034 (O_1034,N_19970,N_19934);
nor UO_1035 (O_1035,N_19878,N_19954);
nand UO_1036 (O_1036,N_19981,N_19919);
nand UO_1037 (O_1037,N_19903,N_19899);
nor UO_1038 (O_1038,N_19945,N_19858);
xor UO_1039 (O_1039,N_19900,N_19972);
xnor UO_1040 (O_1040,N_19840,N_19852);
xor UO_1041 (O_1041,N_19840,N_19962);
and UO_1042 (O_1042,N_19891,N_19868);
nor UO_1043 (O_1043,N_19935,N_19964);
and UO_1044 (O_1044,N_19850,N_19934);
nand UO_1045 (O_1045,N_19911,N_19936);
nand UO_1046 (O_1046,N_19949,N_19914);
nand UO_1047 (O_1047,N_19897,N_19900);
nor UO_1048 (O_1048,N_19841,N_19993);
nand UO_1049 (O_1049,N_19844,N_19998);
or UO_1050 (O_1050,N_19849,N_19892);
nor UO_1051 (O_1051,N_19927,N_19865);
or UO_1052 (O_1052,N_19999,N_19925);
and UO_1053 (O_1053,N_19952,N_19920);
or UO_1054 (O_1054,N_19943,N_19913);
nand UO_1055 (O_1055,N_19928,N_19858);
nand UO_1056 (O_1056,N_19913,N_19960);
nor UO_1057 (O_1057,N_19964,N_19922);
or UO_1058 (O_1058,N_19885,N_19852);
or UO_1059 (O_1059,N_19858,N_19921);
and UO_1060 (O_1060,N_19883,N_19889);
nand UO_1061 (O_1061,N_19923,N_19892);
nand UO_1062 (O_1062,N_19924,N_19934);
nand UO_1063 (O_1063,N_19922,N_19994);
nor UO_1064 (O_1064,N_19921,N_19999);
nand UO_1065 (O_1065,N_19844,N_19979);
or UO_1066 (O_1066,N_19990,N_19987);
or UO_1067 (O_1067,N_19851,N_19901);
or UO_1068 (O_1068,N_19851,N_19950);
or UO_1069 (O_1069,N_19902,N_19861);
nand UO_1070 (O_1070,N_19854,N_19880);
nand UO_1071 (O_1071,N_19962,N_19979);
or UO_1072 (O_1072,N_19940,N_19876);
or UO_1073 (O_1073,N_19997,N_19959);
and UO_1074 (O_1074,N_19890,N_19961);
nor UO_1075 (O_1075,N_19975,N_19945);
xor UO_1076 (O_1076,N_19849,N_19995);
nand UO_1077 (O_1077,N_19845,N_19927);
nand UO_1078 (O_1078,N_19977,N_19999);
and UO_1079 (O_1079,N_19914,N_19929);
nor UO_1080 (O_1080,N_19978,N_19993);
nand UO_1081 (O_1081,N_19941,N_19983);
nor UO_1082 (O_1082,N_19902,N_19924);
nor UO_1083 (O_1083,N_19903,N_19922);
nor UO_1084 (O_1084,N_19946,N_19977);
nor UO_1085 (O_1085,N_19924,N_19882);
or UO_1086 (O_1086,N_19968,N_19853);
or UO_1087 (O_1087,N_19978,N_19907);
xnor UO_1088 (O_1088,N_19886,N_19933);
xnor UO_1089 (O_1089,N_19912,N_19879);
nor UO_1090 (O_1090,N_19942,N_19856);
xnor UO_1091 (O_1091,N_19938,N_19955);
and UO_1092 (O_1092,N_19956,N_19987);
nand UO_1093 (O_1093,N_19862,N_19950);
nor UO_1094 (O_1094,N_19901,N_19974);
nand UO_1095 (O_1095,N_19846,N_19948);
nand UO_1096 (O_1096,N_19970,N_19876);
nor UO_1097 (O_1097,N_19901,N_19848);
nor UO_1098 (O_1098,N_19847,N_19891);
or UO_1099 (O_1099,N_19964,N_19856);
xnor UO_1100 (O_1100,N_19981,N_19887);
nor UO_1101 (O_1101,N_19949,N_19888);
or UO_1102 (O_1102,N_19893,N_19992);
xnor UO_1103 (O_1103,N_19886,N_19939);
and UO_1104 (O_1104,N_19861,N_19926);
or UO_1105 (O_1105,N_19938,N_19844);
nor UO_1106 (O_1106,N_19918,N_19937);
and UO_1107 (O_1107,N_19881,N_19993);
xor UO_1108 (O_1108,N_19995,N_19894);
or UO_1109 (O_1109,N_19986,N_19967);
or UO_1110 (O_1110,N_19846,N_19874);
and UO_1111 (O_1111,N_19906,N_19989);
nor UO_1112 (O_1112,N_19868,N_19863);
and UO_1113 (O_1113,N_19871,N_19939);
or UO_1114 (O_1114,N_19956,N_19924);
and UO_1115 (O_1115,N_19878,N_19928);
or UO_1116 (O_1116,N_19854,N_19853);
nand UO_1117 (O_1117,N_19865,N_19903);
and UO_1118 (O_1118,N_19844,N_19914);
and UO_1119 (O_1119,N_19930,N_19932);
or UO_1120 (O_1120,N_19861,N_19964);
nor UO_1121 (O_1121,N_19968,N_19998);
nor UO_1122 (O_1122,N_19924,N_19930);
xnor UO_1123 (O_1123,N_19888,N_19955);
nor UO_1124 (O_1124,N_19926,N_19966);
or UO_1125 (O_1125,N_19935,N_19947);
or UO_1126 (O_1126,N_19854,N_19897);
nor UO_1127 (O_1127,N_19920,N_19964);
and UO_1128 (O_1128,N_19975,N_19876);
nor UO_1129 (O_1129,N_19995,N_19898);
nor UO_1130 (O_1130,N_19994,N_19856);
or UO_1131 (O_1131,N_19915,N_19851);
nand UO_1132 (O_1132,N_19931,N_19972);
and UO_1133 (O_1133,N_19854,N_19871);
nor UO_1134 (O_1134,N_19891,N_19855);
and UO_1135 (O_1135,N_19891,N_19963);
nand UO_1136 (O_1136,N_19852,N_19937);
and UO_1137 (O_1137,N_19962,N_19991);
xnor UO_1138 (O_1138,N_19963,N_19934);
and UO_1139 (O_1139,N_19996,N_19914);
and UO_1140 (O_1140,N_19869,N_19927);
and UO_1141 (O_1141,N_19853,N_19882);
nor UO_1142 (O_1142,N_19939,N_19971);
xor UO_1143 (O_1143,N_19998,N_19969);
nand UO_1144 (O_1144,N_19986,N_19978);
or UO_1145 (O_1145,N_19865,N_19842);
or UO_1146 (O_1146,N_19941,N_19936);
nor UO_1147 (O_1147,N_19927,N_19925);
and UO_1148 (O_1148,N_19912,N_19896);
xor UO_1149 (O_1149,N_19989,N_19993);
or UO_1150 (O_1150,N_19971,N_19982);
or UO_1151 (O_1151,N_19873,N_19905);
nor UO_1152 (O_1152,N_19886,N_19848);
and UO_1153 (O_1153,N_19994,N_19855);
or UO_1154 (O_1154,N_19919,N_19948);
xor UO_1155 (O_1155,N_19880,N_19955);
nand UO_1156 (O_1156,N_19862,N_19989);
and UO_1157 (O_1157,N_19919,N_19940);
and UO_1158 (O_1158,N_19975,N_19843);
nor UO_1159 (O_1159,N_19990,N_19914);
nand UO_1160 (O_1160,N_19947,N_19907);
or UO_1161 (O_1161,N_19917,N_19939);
nand UO_1162 (O_1162,N_19907,N_19852);
nor UO_1163 (O_1163,N_19869,N_19956);
or UO_1164 (O_1164,N_19942,N_19894);
nor UO_1165 (O_1165,N_19993,N_19961);
nor UO_1166 (O_1166,N_19976,N_19972);
and UO_1167 (O_1167,N_19931,N_19917);
xor UO_1168 (O_1168,N_19889,N_19915);
nand UO_1169 (O_1169,N_19840,N_19843);
nor UO_1170 (O_1170,N_19859,N_19993);
or UO_1171 (O_1171,N_19849,N_19867);
nand UO_1172 (O_1172,N_19985,N_19845);
and UO_1173 (O_1173,N_19936,N_19872);
or UO_1174 (O_1174,N_19919,N_19846);
or UO_1175 (O_1175,N_19887,N_19926);
and UO_1176 (O_1176,N_19879,N_19950);
and UO_1177 (O_1177,N_19905,N_19983);
xnor UO_1178 (O_1178,N_19916,N_19896);
and UO_1179 (O_1179,N_19942,N_19930);
nand UO_1180 (O_1180,N_19945,N_19901);
and UO_1181 (O_1181,N_19943,N_19916);
nor UO_1182 (O_1182,N_19962,N_19985);
nor UO_1183 (O_1183,N_19917,N_19993);
or UO_1184 (O_1184,N_19939,N_19954);
or UO_1185 (O_1185,N_19993,N_19956);
or UO_1186 (O_1186,N_19880,N_19853);
and UO_1187 (O_1187,N_19872,N_19844);
or UO_1188 (O_1188,N_19849,N_19907);
nand UO_1189 (O_1189,N_19860,N_19952);
and UO_1190 (O_1190,N_19903,N_19989);
and UO_1191 (O_1191,N_19877,N_19928);
nor UO_1192 (O_1192,N_19881,N_19904);
and UO_1193 (O_1193,N_19909,N_19962);
and UO_1194 (O_1194,N_19917,N_19927);
nor UO_1195 (O_1195,N_19902,N_19844);
nand UO_1196 (O_1196,N_19857,N_19987);
nand UO_1197 (O_1197,N_19845,N_19892);
or UO_1198 (O_1198,N_19888,N_19906);
or UO_1199 (O_1199,N_19989,N_19996);
xnor UO_1200 (O_1200,N_19992,N_19999);
xnor UO_1201 (O_1201,N_19954,N_19881);
or UO_1202 (O_1202,N_19876,N_19872);
nand UO_1203 (O_1203,N_19977,N_19992);
nor UO_1204 (O_1204,N_19864,N_19961);
nor UO_1205 (O_1205,N_19942,N_19935);
nand UO_1206 (O_1206,N_19884,N_19861);
nand UO_1207 (O_1207,N_19933,N_19930);
or UO_1208 (O_1208,N_19984,N_19847);
and UO_1209 (O_1209,N_19896,N_19889);
or UO_1210 (O_1210,N_19947,N_19878);
and UO_1211 (O_1211,N_19926,N_19854);
nor UO_1212 (O_1212,N_19972,N_19987);
or UO_1213 (O_1213,N_19979,N_19867);
nand UO_1214 (O_1214,N_19915,N_19921);
or UO_1215 (O_1215,N_19984,N_19852);
nor UO_1216 (O_1216,N_19980,N_19930);
or UO_1217 (O_1217,N_19847,N_19956);
and UO_1218 (O_1218,N_19951,N_19964);
and UO_1219 (O_1219,N_19954,N_19934);
and UO_1220 (O_1220,N_19984,N_19946);
nand UO_1221 (O_1221,N_19919,N_19969);
nor UO_1222 (O_1222,N_19908,N_19848);
nand UO_1223 (O_1223,N_19978,N_19967);
and UO_1224 (O_1224,N_19956,N_19994);
and UO_1225 (O_1225,N_19858,N_19955);
xnor UO_1226 (O_1226,N_19959,N_19951);
xor UO_1227 (O_1227,N_19999,N_19956);
and UO_1228 (O_1228,N_19863,N_19925);
and UO_1229 (O_1229,N_19954,N_19916);
xnor UO_1230 (O_1230,N_19903,N_19847);
or UO_1231 (O_1231,N_19886,N_19898);
nand UO_1232 (O_1232,N_19977,N_19867);
nor UO_1233 (O_1233,N_19900,N_19939);
nor UO_1234 (O_1234,N_19933,N_19985);
xor UO_1235 (O_1235,N_19913,N_19906);
or UO_1236 (O_1236,N_19850,N_19919);
nor UO_1237 (O_1237,N_19882,N_19957);
nand UO_1238 (O_1238,N_19994,N_19967);
nand UO_1239 (O_1239,N_19990,N_19958);
nor UO_1240 (O_1240,N_19859,N_19858);
and UO_1241 (O_1241,N_19887,N_19846);
xor UO_1242 (O_1242,N_19848,N_19915);
or UO_1243 (O_1243,N_19921,N_19992);
and UO_1244 (O_1244,N_19904,N_19991);
and UO_1245 (O_1245,N_19996,N_19953);
nand UO_1246 (O_1246,N_19982,N_19919);
and UO_1247 (O_1247,N_19910,N_19915);
nand UO_1248 (O_1248,N_19942,N_19925);
nor UO_1249 (O_1249,N_19898,N_19889);
nand UO_1250 (O_1250,N_19995,N_19980);
and UO_1251 (O_1251,N_19970,N_19886);
or UO_1252 (O_1252,N_19889,N_19967);
nor UO_1253 (O_1253,N_19936,N_19873);
or UO_1254 (O_1254,N_19942,N_19998);
xnor UO_1255 (O_1255,N_19859,N_19898);
and UO_1256 (O_1256,N_19870,N_19939);
and UO_1257 (O_1257,N_19918,N_19898);
nor UO_1258 (O_1258,N_19844,N_19921);
nand UO_1259 (O_1259,N_19859,N_19939);
and UO_1260 (O_1260,N_19903,N_19932);
xor UO_1261 (O_1261,N_19995,N_19902);
xor UO_1262 (O_1262,N_19974,N_19891);
nor UO_1263 (O_1263,N_19984,N_19974);
nor UO_1264 (O_1264,N_19850,N_19932);
nand UO_1265 (O_1265,N_19975,N_19951);
nand UO_1266 (O_1266,N_19904,N_19854);
and UO_1267 (O_1267,N_19900,N_19869);
xnor UO_1268 (O_1268,N_19858,N_19997);
or UO_1269 (O_1269,N_19968,N_19981);
nor UO_1270 (O_1270,N_19861,N_19955);
or UO_1271 (O_1271,N_19938,N_19892);
nor UO_1272 (O_1272,N_19920,N_19999);
and UO_1273 (O_1273,N_19962,N_19964);
or UO_1274 (O_1274,N_19971,N_19968);
nor UO_1275 (O_1275,N_19866,N_19936);
or UO_1276 (O_1276,N_19956,N_19932);
and UO_1277 (O_1277,N_19983,N_19919);
or UO_1278 (O_1278,N_19866,N_19877);
nor UO_1279 (O_1279,N_19865,N_19843);
nor UO_1280 (O_1280,N_19890,N_19904);
nand UO_1281 (O_1281,N_19951,N_19983);
nand UO_1282 (O_1282,N_19992,N_19844);
xor UO_1283 (O_1283,N_19908,N_19901);
or UO_1284 (O_1284,N_19863,N_19846);
and UO_1285 (O_1285,N_19924,N_19845);
or UO_1286 (O_1286,N_19905,N_19852);
and UO_1287 (O_1287,N_19884,N_19972);
nor UO_1288 (O_1288,N_19917,N_19885);
and UO_1289 (O_1289,N_19923,N_19888);
or UO_1290 (O_1290,N_19943,N_19925);
nand UO_1291 (O_1291,N_19953,N_19948);
or UO_1292 (O_1292,N_19896,N_19995);
or UO_1293 (O_1293,N_19999,N_19898);
or UO_1294 (O_1294,N_19857,N_19889);
or UO_1295 (O_1295,N_19917,N_19905);
and UO_1296 (O_1296,N_19888,N_19947);
nor UO_1297 (O_1297,N_19847,N_19870);
and UO_1298 (O_1298,N_19895,N_19918);
nand UO_1299 (O_1299,N_19996,N_19894);
nand UO_1300 (O_1300,N_19950,N_19845);
or UO_1301 (O_1301,N_19907,N_19997);
xor UO_1302 (O_1302,N_19934,N_19889);
or UO_1303 (O_1303,N_19869,N_19857);
xnor UO_1304 (O_1304,N_19904,N_19880);
xor UO_1305 (O_1305,N_19918,N_19907);
and UO_1306 (O_1306,N_19972,N_19920);
nor UO_1307 (O_1307,N_19935,N_19998);
and UO_1308 (O_1308,N_19894,N_19949);
nor UO_1309 (O_1309,N_19844,N_19975);
nor UO_1310 (O_1310,N_19976,N_19881);
and UO_1311 (O_1311,N_19960,N_19951);
nand UO_1312 (O_1312,N_19923,N_19950);
nor UO_1313 (O_1313,N_19868,N_19982);
nand UO_1314 (O_1314,N_19872,N_19903);
and UO_1315 (O_1315,N_19887,N_19922);
nor UO_1316 (O_1316,N_19987,N_19879);
and UO_1317 (O_1317,N_19912,N_19862);
xor UO_1318 (O_1318,N_19986,N_19952);
and UO_1319 (O_1319,N_19991,N_19923);
and UO_1320 (O_1320,N_19840,N_19973);
nor UO_1321 (O_1321,N_19872,N_19865);
and UO_1322 (O_1322,N_19941,N_19969);
or UO_1323 (O_1323,N_19949,N_19998);
xor UO_1324 (O_1324,N_19881,N_19866);
nand UO_1325 (O_1325,N_19899,N_19967);
and UO_1326 (O_1326,N_19949,N_19956);
and UO_1327 (O_1327,N_19944,N_19957);
or UO_1328 (O_1328,N_19946,N_19945);
nand UO_1329 (O_1329,N_19871,N_19887);
nand UO_1330 (O_1330,N_19869,N_19988);
and UO_1331 (O_1331,N_19925,N_19918);
or UO_1332 (O_1332,N_19954,N_19938);
or UO_1333 (O_1333,N_19845,N_19865);
or UO_1334 (O_1334,N_19890,N_19989);
and UO_1335 (O_1335,N_19940,N_19951);
xnor UO_1336 (O_1336,N_19956,N_19920);
xor UO_1337 (O_1337,N_19983,N_19886);
or UO_1338 (O_1338,N_19905,N_19999);
and UO_1339 (O_1339,N_19964,N_19888);
nor UO_1340 (O_1340,N_19933,N_19938);
or UO_1341 (O_1341,N_19899,N_19963);
nand UO_1342 (O_1342,N_19913,N_19894);
nor UO_1343 (O_1343,N_19978,N_19892);
and UO_1344 (O_1344,N_19889,N_19973);
nor UO_1345 (O_1345,N_19975,N_19940);
and UO_1346 (O_1346,N_19919,N_19965);
nor UO_1347 (O_1347,N_19989,N_19966);
nor UO_1348 (O_1348,N_19944,N_19984);
nor UO_1349 (O_1349,N_19919,N_19939);
nor UO_1350 (O_1350,N_19905,N_19886);
and UO_1351 (O_1351,N_19869,N_19914);
or UO_1352 (O_1352,N_19942,N_19876);
xor UO_1353 (O_1353,N_19920,N_19904);
or UO_1354 (O_1354,N_19979,N_19890);
nor UO_1355 (O_1355,N_19937,N_19941);
nand UO_1356 (O_1356,N_19939,N_19901);
and UO_1357 (O_1357,N_19949,N_19885);
and UO_1358 (O_1358,N_19965,N_19915);
or UO_1359 (O_1359,N_19976,N_19941);
and UO_1360 (O_1360,N_19857,N_19978);
and UO_1361 (O_1361,N_19913,N_19846);
or UO_1362 (O_1362,N_19972,N_19851);
nor UO_1363 (O_1363,N_19916,N_19913);
nand UO_1364 (O_1364,N_19843,N_19942);
or UO_1365 (O_1365,N_19966,N_19847);
nor UO_1366 (O_1366,N_19980,N_19944);
and UO_1367 (O_1367,N_19893,N_19856);
nor UO_1368 (O_1368,N_19890,N_19928);
and UO_1369 (O_1369,N_19884,N_19935);
and UO_1370 (O_1370,N_19993,N_19954);
or UO_1371 (O_1371,N_19953,N_19927);
and UO_1372 (O_1372,N_19953,N_19865);
nand UO_1373 (O_1373,N_19970,N_19905);
or UO_1374 (O_1374,N_19928,N_19990);
nor UO_1375 (O_1375,N_19941,N_19892);
and UO_1376 (O_1376,N_19968,N_19950);
and UO_1377 (O_1377,N_19843,N_19954);
or UO_1378 (O_1378,N_19994,N_19986);
nand UO_1379 (O_1379,N_19937,N_19841);
and UO_1380 (O_1380,N_19987,N_19902);
nor UO_1381 (O_1381,N_19931,N_19918);
and UO_1382 (O_1382,N_19862,N_19861);
xnor UO_1383 (O_1383,N_19884,N_19965);
or UO_1384 (O_1384,N_19842,N_19876);
nor UO_1385 (O_1385,N_19907,N_19916);
nor UO_1386 (O_1386,N_19925,N_19959);
and UO_1387 (O_1387,N_19892,N_19907);
or UO_1388 (O_1388,N_19996,N_19907);
nand UO_1389 (O_1389,N_19900,N_19911);
nor UO_1390 (O_1390,N_19911,N_19924);
xnor UO_1391 (O_1391,N_19869,N_19944);
xor UO_1392 (O_1392,N_19967,N_19840);
xnor UO_1393 (O_1393,N_19974,N_19886);
or UO_1394 (O_1394,N_19921,N_19869);
and UO_1395 (O_1395,N_19905,N_19874);
nor UO_1396 (O_1396,N_19971,N_19925);
nand UO_1397 (O_1397,N_19868,N_19899);
or UO_1398 (O_1398,N_19982,N_19904);
and UO_1399 (O_1399,N_19896,N_19939);
or UO_1400 (O_1400,N_19904,N_19938);
or UO_1401 (O_1401,N_19920,N_19979);
nor UO_1402 (O_1402,N_19863,N_19938);
or UO_1403 (O_1403,N_19988,N_19955);
nand UO_1404 (O_1404,N_19960,N_19936);
and UO_1405 (O_1405,N_19954,N_19841);
nor UO_1406 (O_1406,N_19916,N_19870);
or UO_1407 (O_1407,N_19915,N_19907);
nand UO_1408 (O_1408,N_19946,N_19985);
nand UO_1409 (O_1409,N_19977,N_19856);
and UO_1410 (O_1410,N_19991,N_19859);
and UO_1411 (O_1411,N_19933,N_19965);
nor UO_1412 (O_1412,N_19965,N_19842);
nor UO_1413 (O_1413,N_19886,N_19891);
nor UO_1414 (O_1414,N_19935,N_19961);
xnor UO_1415 (O_1415,N_19852,N_19883);
nor UO_1416 (O_1416,N_19956,N_19886);
or UO_1417 (O_1417,N_19923,N_19976);
nor UO_1418 (O_1418,N_19986,N_19962);
nand UO_1419 (O_1419,N_19995,N_19917);
nor UO_1420 (O_1420,N_19862,N_19961);
nand UO_1421 (O_1421,N_19950,N_19871);
and UO_1422 (O_1422,N_19888,N_19939);
nand UO_1423 (O_1423,N_19896,N_19893);
or UO_1424 (O_1424,N_19916,N_19849);
or UO_1425 (O_1425,N_19861,N_19981);
nor UO_1426 (O_1426,N_19941,N_19929);
nor UO_1427 (O_1427,N_19909,N_19984);
and UO_1428 (O_1428,N_19845,N_19934);
and UO_1429 (O_1429,N_19905,N_19954);
nand UO_1430 (O_1430,N_19859,N_19944);
xor UO_1431 (O_1431,N_19886,N_19999);
and UO_1432 (O_1432,N_19901,N_19878);
and UO_1433 (O_1433,N_19992,N_19984);
and UO_1434 (O_1434,N_19932,N_19843);
or UO_1435 (O_1435,N_19882,N_19867);
and UO_1436 (O_1436,N_19869,N_19873);
or UO_1437 (O_1437,N_19865,N_19961);
or UO_1438 (O_1438,N_19980,N_19843);
and UO_1439 (O_1439,N_19936,N_19998);
nor UO_1440 (O_1440,N_19862,N_19879);
or UO_1441 (O_1441,N_19848,N_19895);
or UO_1442 (O_1442,N_19996,N_19880);
or UO_1443 (O_1443,N_19949,N_19958);
or UO_1444 (O_1444,N_19858,N_19845);
nor UO_1445 (O_1445,N_19998,N_19934);
or UO_1446 (O_1446,N_19975,N_19885);
and UO_1447 (O_1447,N_19945,N_19933);
nand UO_1448 (O_1448,N_19912,N_19844);
xor UO_1449 (O_1449,N_19983,N_19892);
or UO_1450 (O_1450,N_19882,N_19933);
nand UO_1451 (O_1451,N_19906,N_19940);
nand UO_1452 (O_1452,N_19956,N_19968);
nand UO_1453 (O_1453,N_19896,N_19861);
nor UO_1454 (O_1454,N_19846,N_19892);
or UO_1455 (O_1455,N_19881,N_19917);
nor UO_1456 (O_1456,N_19857,N_19953);
nand UO_1457 (O_1457,N_19843,N_19979);
xnor UO_1458 (O_1458,N_19855,N_19961);
and UO_1459 (O_1459,N_19920,N_19890);
nand UO_1460 (O_1460,N_19999,N_19866);
nor UO_1461 (O_1461,N_19883,N_19938);
nand UO_1462 (O_1462,N_19892,N_19869);
nand UO_1463 (O_1463,N_19847,N_19983);
or UO_1464 (O_1464,N_19987,N_19982);
nor UO_1465 (O_1465,N_19840,N_19879);
and UO_1466 (O_1466,N_19845,N_19860);
or UO_1467 (O_1467,N_19880,N_19899);
nand UO_1468 (O_1468,N_19924,N_19860);
nor UO_1469 (O_1469,N_19977,N_19932);
nor UO_1470 (O_1470,N_19964,N_19955);
or UO_1471 (O_1471,N_19870,N_19908);
xnor UO_1472 (O_1472,N_19966,N_19848);
nand UO_1473 (O_1473,N_19881,N_19895);
nand UO_1474 (O_1474,N_19992,N_19891);
and UO_1475 (O_1475,N_19922,N_19844);
or UO_1476 (O_1476,N_19942,N_19915);
and UO_1477 (O_1477,N_19842,N_19988);
xor UO_1478 (O_1478,N_19951,N_19859);
xor UO_1479 (O_1479,N_19901,N_19916);
or UO_1480 (O_1480,N_19957,N_19945);
and UO_1481 (O_1481,N_19856,N_19967);
nand UO_1482 (O_1482,N_19993,N_19848);
xor UO_1483 (O_1483,N_19963,N_19926);
nor UO_1484 (O_1484,N_19906,N_19985);
nor UO_1485 (O_1485,N_19913,N_19861);
and UO_1486 (O_1486,N_19891,N_19958);
nand UO_1487 (O_1487,N_19902,N_19890);
or UO_1488 (O_1488,N_19955,N_19984);
nand UO_1489 (O_1489,N_19885,N_19904);
and UO_1490 (O_1490,N_19946,N_19956);
xnor UO_1491 (O_1491,N_19860,N_19951);
and UO_1492 (O_1492,N_19956,N_19934);
nor UO_1493 (O_1493,N_19846,N_19983);
nand UO_1494 (O_1494,N_19962,N_19904);
nor UO_1495 (O_1495,N_19933,N_19887);
nand UO_1496 (O_1496,N_19922,N_19908);
and UO_1497 (O_1497,N_19854,N_19846);
nor UO_1498 (O_1498,N_19914,N_19981);
or UO_1499 (O_1499,N_19934,N_19847);
xnor UO_1500 (O_1500,N_19989,N_19874);
and UO_1501 (O_1501,N_19931,N_19974);
and UO_1502 (O_1502,N_19954,N_19922);
or UO_1503 (O_1503,N_19881,N_19940);
or UO_1504 (O_1504,N_19973,N_19917);
or UO_1505 (O_1505,N_19857,N_19995);
and UO_1506 (O_1506,N_19922,N_19999);
nand UO_1507 (O_1507,N_19851,N_19917);
nand UO_1508 (O_1508,N_19983,N_19969);
nand UO_1509 (O_1509,N_19982,N_19983);
nor UO_1510 (O_1510,N_19957,N_19960);
nand UO_1511 (O_1511,N_19972,N_19981);
nor UO_1512 (O_1512,N_19891,N_19946);
or UO_1513 (O_1513,N_19964,N_19867);
and UO_1514 (O_1514,N_19847,N_19874);
and UO_1515 (O_1515,N_19862,N_19890);
and UO_1516 (O_1516,N_19969,N_19876);
nand UO_1517 (O_1517,N_19939,N_19972);
and UO_1518 (O_1518,N_19954,N_19888);
xor UO_1519 (O_1519,N_19921,N_19942);
nand UO_1520 (O_1520,N_19908,N_19992);
or UO_1521 (O_1521,N_19998,N_19910);
or UO_1522 (O_1522,N_19906,N_19946);
nand UO_1523 (O_1523,N_19873,N_19870);
or UO_1524 (O_1524,N_19874,N_19879);
nor UO_1525 (O_1525,N_19927,N_19894);
nor UO_1526 (O_1526,N_19983,N_19915);
nor UO_1527 (O_1527,N_19850,N_19933);
nor UO_1528 (O_1528,N_19990,N_19868);
or UO_1529 (O_1529,N_19904,N_19997);
nor UO_1530 (O_1530,N_19959,N_19914);
or UO_1531 (O_1531,N_19895,N_19912);
nor UO_1532 (O_1532,N_19945,N_19934);
nand UO_1533 (O_1533,N_19970,N_19866);
and UO_1534 (O_1534,N_19963,N_19903);
nand UO_1535 (O_1535,N_19915,N_19875);
nor UO_1536 (O_1536,N_19883,N_19893);
and UO_1537 (O_1537,N_19857,N_19900);
nand UO_1538 (O_1538,N_19983,N_19997);
or UO_1539 (O_1539,N_19868,N_19903);
nand UO_1540 (O_1540,N_19974,N_19859);
or UO_1541 (O_1541,N_19954,N_19877);
and UO_1542 (O_1542,N_19994,N_19899);
nand UO_1543 (O_1543,N_19923,N_19970);
xnor UO_1544 (O_1544,N_19939,N_19961);
and UO_1545 (O_1545,N_19872,N_19980);
or UO_1546 (O_1546,N_19843,N_19965);
or UO_1547 (O_1547,N_19940,N_19991);
nor UO_1548 (O_1548,N_19941,N_19922);
or UO_1549 (O_1549,N_19893,N_19928);
or UO_1550 (O_1550,N_19916,N_19929);
and UO_1551 (O_1551,N_19885,N_19858);
nor UO_1552 (O_1552,N_19888,N_19971);
and UO_1553 (O_1553,N_19867,N_19893);
or UO_1554 (O_1554,N_19974,N_19966);
and UO_1555 (O_1555,N_19921,N_19982);
nand UO_1556 (O_1556,N_19984,N_19896);
or UO_1557 (O_1557,N_19936,N_19882);
xnor UO_1558 (O_1558,N_19956,N_19883);
xnor UO_1559 (O_1559,N_19924,N_19889);
and UO_1560 (O_1560,N_19900,N_19884);
and UO_1561 (O_1561,N_19962,N_19911);
nor UO_1562 (O_1562,N_19967,N_19982);
xor UO_1563 (O_1563,N_19900,N_19945);
xnor UO_1564 (O_1564,N_19957,N_19959);
or UO_1565 (O_1565,N_19844,N_19887);
nand UO_1566 (O_1566,N_19992,N_19919);
or UO_1567 (O_1567,N_19945,N_19907);
nand UO_1568 (O_1568,N_19946,N_19869);
xor UO_1569 (O_1569,N_19906,N_19894);
xor UO_1570 (O_1570,N_19869,N_19928);
nor UO_1571 (O_1571,N_19995,N_19940);
nand UO_1572 (O_1572,N_19846,N_19855);
nor UO_1573 (O_1573,N_19898,N_19993);
and UO_1574 (O_1574,N_19865,N_19899);
nand UO_1575 (O_1575,N_19855,N_19843);
and UO_1576 (O_1576,N_19999,N_19978);
nor UO_1577 (O_1577,N_19945,N_19993);
nand UO_1578 (O_1578,N_19916,N_19967);
nor UO_1579 (O_1579,N_19972,N_19946);
and UO_1580 (O_1580,N_19946,N_19949);
and UO_1581 (O_1581,N_19972,N_19892);
and UO_1582 (O_1582,N_19925,N_19928);
or UO_1583 (O_1583,N_19894,N_19903);
nand UO_1584 (O_1584,N_19840,N_19932);
xnor UO_1585 (O_1585,N_19856,N_19863);
and UO_1586 (O_1586,N_19943,N_19973);
nor UO_1587 (O_1587,N_19922,N_19997);
nor UO_1588 (O_1588,N_19878,N_19900);
nand UO_1589 (O_1589,N_19902,N_19938);
or UO_1590 (O_1590,N_19960,N_19989);
nor UO_1591 (O_1591,N_19866,N_19948);
nor UO_1592 (O_1592,N_19996,N_19844);
or UO_1593 (O_1593,N_19914,N_19856);
and UO_1594 (O_1594,N_19982,N_19941);
nand UO_1595 (O_1595,N_19940,N_19955);
xnor UO_1596 (O_1596,N_19973,N_19879);
nand UO_1597 (O_1597,N_19933,N_19990);
nor UO_1598 (O_1598,N_19990,N_19858);
nand UO_1599 (O_1599,N_19847,N_19936);
and UO_1600 (O_1600,N_19873,N_19985);
and UO_1601 (O_1601,N_19914,N_19906);
nor UO_1602 (O_1602,N_19938,N_19920);
or UO_1603 (O_1603,N_19867,N_19941);
and UO_1604 (O_1604,N_19930,N_19970);
xnor UO_1605 (O_1605,N_19852,N_19854);
and UO_1606 (O_1606,N_19914,N_19997);
and UO_1607 (O_1607,N_19916,N_19917);
and UO_1608 (O_1608,N_19884,N_19859);
or UO_1609 (O_1609,N_19852,N_19934);
nor UO_1610 (O_1610,N_19912,N_19903);
or UO_1611 (O_1611,N_19856,N_19959);
nand UO_1612 (O_1612,N_19919,N_19988);
or UO_1613 (O_1613,N_19919,N_19953);
or UO_1614 (O_1614,N_19861,N_19965);
nor UO_1615 (O_1615,N_19921,N_19937);
nand UO_1616 (O_1616,N_19943,N_19897);
and UO_1617 (O_1617,N_19980,N_19850);
or UO_1618 (O_1618,N_19996,N_19871);
nand UO_1619 (O_1619,N_19937,N_19973);
nor UO_1620 (O_1620,N_19917,N_19859);
and UO_1621 (O_1621,N_19871,N_19934);
or UO_1622 (O_1622,N_19936,N_19920);
nand UO_1623 (O_1623,N_19881,N_19853);
and UO_1624 (O_1624,N_19842,N_19896);
and UO_1625 (O_1625,N_19989,N_19909);
nor UO_1626 (O_1626,N_19877,N_19889);
xnor UO_1627 (O_1627,N_19934,N_19913);
or UO_1628 (O_1628,N_19842,N_19919);
or UO_1629 (O_1629,N_19909,N_19880);
nand UO_1630 (O_1630,N_19860,N_19950);
nand UO_1631 (O_1631,N_19885,N_19968);
and UO_1632 (O_1632,N_19963,N_19916);
xor UO_1633 (O_1633,N_19927,N_19898);
xor UO_1634 (O_1634,N_19960,N_19973);
nand UO_1635 (O_1635,N_19864,N_19845);
or UO_1636 (O_1636,N_19900,N_19926);
xnor UO_1637 (O_1637,N_19889,N_19982);
nand UO_1638 (O_1638,N_19952,N_19943);
or UO_1639 (O_1639,N_19863,N_19923);
and UO_1640 (O_1640,N_19891,N_19973);
nand UO_1641 (O_1641,N_19907,N_19984);
or UO_1642 (O_1642,N_19927,N_19974);
and UO_1643 (O_1643,N_19866,N_19958);
xor UO_1644 (O_1644,N_19906,N_19956);
and UO_1645 (O_1645,N_19864,N_19913);
and UO_1646 (O_1646,N_19864,N_19909);
nor UO_1647 (O_1647,N_19929,N_19997);
nor UO_1648 (O_1648,N_19868,N_19954);
nand UO_1649 (O_1649,N_19960,N_19962);
xor UO_1650 (O_1650,N_19963,N_19939);
nand UO_1651 (O_1651,N_19890,N_19927);
nand UO_1652 (O_1652,N_19878,N_19906);
or UO_1653 (O_1653,N_19874,N_19950);
xor UO_1654 (O_1654,N_19884,N_19946);
nor UO_1655 (O_1655,N_19910,N_19989);
xor UO_1656 (O_1656,N_19932,N_19965);
and UO_1657 (O_1657,N_19858,N_19896);
nor UO_1658 (O_1658,N_19896,N_19918);
or UO_1659 (O_1659,N_19872,N_19922);
nor UO_1660 (O_1660,N_19905,N_19892);
xnor UO_1661 (O_1661,N_19872,N_19952);
or UO_1662 (O_1662,N_19954,N_19958);
or UO_1663 (O_1663,N_19925,N_19985);
nor UO_1664 (O_1664,N_19966,N_19985);
xor UO_1665 (O_1665,N_19940,N_19856);
or UO_1666 (O_1666,N_19971,N_19877);
nand UO_1667 (O_1667,N_19865,N_19915);
nor UO_1668 (O_1668,N_19876,N_19869);
nand UO_1669 (O_1669,N_19997,N_19850);
nand UO_1670 (O_1670,N_19862,N_19984);
xnor UO_1671 (O_1671,N_19907,N_19896);
nor UO_1672 (O_1672,N_19893,N_19886);
and UO_1673 (O_1673,N_19840,N_19995);
nand UO_1674 (O_1674,N_19990,N_19878);
or UO_1675 (O_1675,N_19932,N_19879);
and UO_1676 (O_1676,N_19841,N_19966);
nor UO_1677 (O_1677,N_19984,N_19936);
or UO_1678 (O_1678,N_19949,N_19927);
and UO_1679 (O_1679,N_19942,N_19927);
nand UO_1680 (O_1680,N_19912,N_19993);
or UO_1681 (O_1681,N_19958,N_19863);
nand UO_1682 (O_1682,N_19848,N_19840);
and UO_1683 (O_1683,N_19910,N_19964);
nor UO_1684 (O_1684,N_19943,N_19858);
nor UO_1685 (O_1685,N_19946,N_19847);
nor UO_1686 (O_1686,N_19936,N_19939);
nand UO_1687 (O_1687,N_19946,N_19859);
nor UO_1688 (O_1688,N_19963,N_19905);
or UO_1689 (O_1689,N_19922,N_19840);
or UO_1690 (O_1690,N_19855,N_19881);
nand UO_1691 (O_1691,N_19991,N_19958);
or UO_1692 (O_1692,N_19873,N_19858);
nor UO_1693 (O_1693,N_19940,N_19969);
nand UO_1694 (O_1694,N_19885,N_19987);
or UO_1695 (O_1695,N_19847,N_19898);
nand UO_1696 (O_1696,N_19955,N_19937);
nand UO_1697 (O_1697,N_19866,N_19901);
nand UO_1698 (O_1698,N_19879,N_19916);
nor UO_1699 (O_1699,N_19966,N_19884);
nor UO_1700 (O_1700,N_19949,N_19938);
nand UO_1701 (O_1701,N_19909,N_19953);
or UO_1702 (O_1702,N_19984,N_19904);
or UO_1703 (O_1703,N_19876,N_19981);
or UO_1704 (O_1704,N_19882,N_19869);
and UO_1705 (O_1705,N_19890,N_19841);
nand UO_1706 (O_1706,N_19966,N_19859);
and UO_1707 (O_1707,N_19988,N_19931);
nor UO_1708 (O_1708,N_19949,N_19939);
nor UO_1709 (O_1709,N_19880,N_19886);
and UO_1710 (O_1710,N_19871,N_19846);
and UO_1711 (O_1711,N_19914,N_19969);
or UO_1712 (O_1712,N_19863,N_19855);
or UO_1713 (O_1713,N_19969,N_19908);
nor UO_1714 (O_1714,N_19960,N_19954);
and UO_1715 (O_1715,N_19930,N_19947);
and UO_1716 (O_1716,N_19988,N_19979);
or UO_1717 (O_1717,N_19856,N_19907);
and UO_1718 (O_1718,N_19969,N_19954);
nand UO_1719 (O_1719,N_19985,N_19864);
or UO_1720 (O_1720,N_19904,N_19850);
or UO_1721 (O_1721,N_19966,N_19952);
nand UO_1722 (O_1722,N_19864,N_19974);
nand UO_1723 (O_1723,N_19917,N_19879);
xnor UO_1724 (O_1724,N_19993,N_19981);
nor UO_1725 (O_1725,N_19997,N_19859);
xor UO_1726 (O_1726,N_19957,N_19865);
nand UO_1727 (O_1727,N_19849,N_19923);
and UO_1728 (O_1728,N_19950,N_19901);
and UO_1729 (O_1729,N_19949,N_19917);
nor UO_1730 (O_1730,N_19973,N_19852);
and UO_1731 (O_1731,N_19909,N_19920);
and UO_1732 (O_1732,N_19912,N_19986);
nor UO_1733 (O_1733,N_19873,N_19978);
xnor UO_1734 (O_1734,N_19841,N_19924);
nor UO_1735 (O_1735,N_19891,N_19856);
nor UO_1736 (O_1736,N_19922,N_19861);
nor UO_1737 (O_1737,N_19939,N_19866);
nand UO_1738 (O_1738,N_19871,N_19954);
and UO_1739 (O_1739,N_19875,N_19976);
and UO_1740 (O_1740,N_19929,N_19900);
xnor UO_1741 (O_1741,N_19843,N_19948);
and UO_1742 (O_1742,N_19983,N_19966);
or UO_1743 (O_1743,N_19942,N_19960);
or UO_1744 (O_1744,N_19975,N_19942);
or UO_1745 (O_1745,N_19950,N_19966);
nand UO_1746 (O_1746,N_19931,N_19909);
nand UO_1747 (O_1747,N_19985,N_19973);
and UO_1748 (O_1748,N_19951,N_19992);
nor UO_1749 (O_1749,N_19983,N_19863);
or UO_1750 (O_1750,N_19859,N_19921);
nand UO_1751 (O_1751,N_19847,N_19959);
nor UO_1752 (O_1752,N_19942,N_19872);
nor UO_1753 (O_1753,N_19922,N_19850);
and UO_1754 (O_1754,N_19879,N_19980);
nand UO_1755 (O_1755,N_19940,N_19884);
nand UO_1756 (O_1756,N_19846,N_19993);
nand UO_1757 (O_1757,N_19848,N_19935);
xnor UO_1758 (O_1758,N_19902,N_19876);
nand UO_1759 (O_1759,N_19971,N_19941);
nand UO_1760 (O_1760,N_19926,N_19920);
xor UO_1761 (O_1761,N_19928,N_19936);
nand UO_1762 (O_1762,N_19896,N_19883);
nor UO_1763 (O_1763,N_19877,N_19940);
or UO_1764 (O_1764,N_19932,N_19891);
or UO_1765 (O_1765,N_19977,N_19962);
and UO_1766 (O_1766,N_19855,N_19932);
nor UO_1767 (O_1767,N_19965,N_19944);
and UO_1768 (O_1768,N_19980,N_19969);
nor UO_1769 (O_1769,N_19894,N_19988);
or UO_1770 (O_1770,N_19848,N_19887);
nand UO_1771 (O_1771,N_19950,N_19944);
nand UO_1772 (O_1772,N_19908,N_19999);
nand UO_1773 (O_1773,N_19867,N_19937);
xor UO_1774 (O_1774,N_19910,N_19978);
or UO_1775 (O_1775,N_19862,N_19872);
and UO_1776 (O_1776,N_19973,N_19957);
and UO_1777 (O_1777,N_19894,N_19964);
nor UO_1778 (O_1778,N_19927,N_19850);
xnor UO_1779 (O_1779,N_19873,N_19914);
nand UO_1780 (O_1780,N_19946,N_19863);
nor UO_1781 (O_1781,N_19859,N_19870);
nand UO_1782 (O_1782,N_19871,N_19884);
nand UO_1783 (O_1783,N_19953,N_19920);
and UO_1784 (O_1784,N_19975,N_19935);
and UO_1785 (O_1785,N_19965,N_19998);
or UO_1786 (O_1786,N_19886,N_19965);
and UO_1787 (O_1787,N_19997,N_19918);
nor UO_1788 (O_1788,N_19929,N_19844);
nand UO_1789 (O_1789,N_19954,N_19867);
and UO_1790 (O_1790,N_19854,N_19861);
and UO_1791 (O_1791,N_19876,N_19987);
nor UO_1792 (O_1792,N_19962,N_19995);
or UO_1793 (O_1793,N_19948,N_19853);
nor UO_1794 (O_1794,N_19940,N_19960);
or UO_1795 (O_1795,N_19894,N_19879);
or UO_1796 (O_1796,N_19935,N_19860);
nand UO_1797 (O_1797,N_19932,N_19972);
or UO_1798 (O_1798,N_19959,N_19941);
nor UO_1799 (O_1799,N_19904,N_19973);
or UO_1800 (O_1800,N_19904,N_19841);
nand UO_1801 (O_1801,N_19950,N_19958);
nor UO_1802 (O_1802,N_19962,N_19930);
nand UO_1803 (O_1803,N_19961,N_19977);
or UO_1804 (O_1804,N_19841,N_19972);
or UO_1805 (O_1805,N_19842,N_19874);
and UO_1806 (O_1806,N_19845,N_19974);
nand UO_1807 (O_1807,N_19927,N_19875);
and UO_1808 (O_1808,N_19986,N_19864);
and UO_1809 (O_1809,N_19944,N_19884);
xnor UO_1810 (O_1810,N_19877,N_19848);
or UO_1811 (O_1811,N_19987,N_19955);
nor UO_1812 (O_1812,N_19947,N_19906);
and UO_1813 (O_1813,N_19887,N_19955);
or UO_1814 (O_1814,N_19971,N_19999);
or UO_1815 (O_1815,N_19871,N_19895);
nand UO_1816 (O_1816,N_19914,N_19964);
xnor UO_1817 (O_1817,N_19880,N_19978);
nand UO_1818 (O_1818,N_19955,N_19876);
and UO_1819 (O_1819,N_19847,N_19900);
nor UO_1820 (O_1820,N_19944,N_19932);
nor UO_1821 (O_1821,N_19913,N_19923);
or UO_1822 (O_1822,N_19904,N_19979);
or UO_1823 (O_1823,N_19985,N_19920);
nor UO_1824 (O_1824,N_19973,N_19999);
nand UO_1825 (O_1825,N_19953,N_19869);
nor UO_1826 (O_1826,N_19900,N_19846);
nand UO_1827 (O_1827,N_19867,N_19878);
and UO_1828 (O_1828,N_19971,N_19997);
or UO_1829 (O_1829,N_19886,N_19919);
or UO_1830 (O_1830,N_19943,N_19932);
or UO_1831 (O_1831,N_19988,N_19872);
xnor UO_1832 (O_1832,N_19872,N_19951);
nand UO_1833 (O_1833,N_19928,N_19899);
nor UO_1834 (O_1834,N_19952,N_19985);
nand UO_1835 (O_1835,N_19921,N_19957);
nand UO_1836 (O_1836,N_19905,N_19869);
nor UO_1837 (O_1837,N_19911,N_19976);
or UO_1838 (O_1838,N_19853,N_19919);
nor UO_1839 (O_1839,N_19984,N_19880);
nor UO_1840 (O_1840,N_19908,N_19938);
xor UO_1841 (O_1841,N_19864,N_19841);
nand UO_1842 (O_1842,N_19848,N_19867);
nor UO_1843 (O_1843,N_19961,N_19913);
nand UO_1844 (O_1844,N_19979,N_19915);
nor UO_1845 (O_1845,N_19930,N_19885);
nor UO_1846 (O_1846,N_19856,N_19917);
and UO_1847 (O_1847,N_19946,N_19919);
and UO_1848 (O_1848,N_19985,N_19896);
nand UO_1849 (O_1849,N_19990,N_19867);
nor UO_1850 (O_1850,N_19898,N_19906);
nor UO_1851 (O_1851,N_19906,N_19923);
nand UO_1852 (O_1852,N_19972,N_19934);
nor UO_1853 (O_1853,N_19884,N_19989);
nor UO_1854 (O_1854,N_19954,N_19955);
or UO_1855 (O_1855,N_19952,N_19923);
and UO_1856 (O_1856,N_19919,N_19971);
or UO_1857 (O_1857,N_19928,N_19921);
and UO_1858 (O_1858,N_19883,N_19840);
or UO_1859 (O_1859,N_19858,N_19848);
nor UO_1860 (O_1860,N_19915,N_19896);
nand UO_1861 (O_1861,N_19891,N_19914);
or UO_1862 (O_1862,N_19890,N_19983);
xnor UO_1863 (O_1863,N_19862,N_19998);
nor UO_1864 (O_1864,N_19940,N_19930);
nor UO_1865 (O_1865,N_19975,N_19973);
or UO_1866 (O_1866,N_19848,N_19903);
nor UO_1867 (O_1867,N_19947,N_19938);
or UO_1868 (O_1868,N_19879,N_19982);
and UO_1869 (O_1869,N_19886,N_19949);
xor UO_1870 (O_1870,N_19844,N_19909);
nor UO_1871 (O_1871,N_19851,N_19993);
or UO_1872 (O_1872,N_19958,N_19881);
nand UO_1873 (O_1873,N_19926,N_19969);
xor UO_1874 (O_1874,N_19877,N_19876);
and UO_1875 (O_1875,N_19889,N_19850);
or UO_1876 (O_1876,N_19932,N_19905);
or UO_1877 (O_1877,N_19876,N_19863);
or UO_1878 (O_1878,N_19849,N_19840);
nor UO_1879 (O_1879,N_19896,N_19968);
nor UO_1880 (O_1880,N_19865,N_19986);
nand UO_1881 (O_1881,N_19861,N_19935);
nand UO_1882 (O_1882,N_19911,N_19885);
and UO_1883 (O_1883,N_19885,N_19847);
nand UO_1884 (O_1884,N_19951,N_19973);
nand UO_1885 (O_1885,N_19971,N_19847);
and UO_1886 (O_1886,N_19969,N_19855);
and UO_1887 (O_1887,N_19855,N_19922);
nor UO_1888 (O_1888,N_19977,N_19981);
and UO_1889 (O_1889,N_19940,N_19904);
or UO_1890 (O_1890,N_19859,N_19911);
and UO_1891 (O_1891,N_19864,N_19931);
nand UO_1892 (O_1892,N_19925,N_19947);
or UO_1893 (O_1893,N_19955,N_19856);
nor UO_1894 (O_1894,N_19886,N_19874);
and UO_1895 (O_1895,N_19910,N_19913);
nor UO_1896 (O_1896,N_19965,N_19894);
xor UO_1897 (O_1897,N_19977,N_19911);
and UO_1898 (O_1898,N_19932,N_19895);
and UO_1899 (O_1899,N_19841,N_19846);
and UO_1900 (O_1900,N_19848,N_19913);
nand UO_1901 (O_1901,N_19992,N_19943);
xnor UO_1902 (O_1902,N_19887,N_19891);
nor UO_1903 (O_1903,N_19999,N_19864);
nand UO_1904 (O_1904,N_19863,N_19881);
or UO_1905 (O_1905,N_19958,N_19924);
and UO_1906 (O_1906,N_19849,N_19954);
xor UO_1907 (O_1907,N_19889,N_19956);
or UO_1908 (O_1908,N_19902,N_19996);
nand UO_1909 (O_1909,N_19964,N_19959);
or UO_1910 (O_1910,N_19882,N_19881);
or UO_1911 (O_1911,N_19930,N_19963);
nand UO_1912 (O_1912,N_19865,N_19984);
and UO_1913 (O_1913,N_19970,N_19863);
and UO_1914 (O_1914,N_19967,N_19943);
nor UO_1915 (O_1915,N_19874,N_19911);
nor UO_1916 (O_1916,N_19931,N_19895);
nand UO_1917 (O_1917,N_19906,N_19957);
and UO_1918 (O_1918,N_19936,N_19913);
nand UO_1919 (O_1919,N_19992,N_19904);
and UO_1920 (O_1920,N_19909,N_19971);
or UO_1921 (O_1921,N_19959,N_19912);
or UO_1922 (O_1922,N_19909,N_19875);
nand UO_1923 (O_1923,N_19865,N_19922);
or UO_1924 (O_1924,N_19916,N_19962);
nor UO_1925 (O_1925,N_19985,N_19852);
nor UO_1926 (O_1926,N_19910,N_19912);
xor UO_1927 (O_1927,N_19967,N_19973);
nand UO_1928 (O_1928,N_19843,N_19848);
and UO_1929 (O_1929,N_19879,N_19859);
nand UO_1930 (O_1930,N_19993,N_19964);
nor UO_1931 (O_1931,N_19992,N_19978);
or UO_1932 (O_1932,N_19920,N_19889);
xor UO_1933 (O_1933,N_19840,N_19935);
nand UO_1934 (O_1934,N_19856,N_19909);
or UO_1935 (O_1935,N_19870,N_19953);
nand UO_1936 (O_1936,N_19854,N_19867);
nor UO_1937 (O_1937,N_19996,N_19944);
nand UO_1938 (O_1938,N_19987,N_19947);
nand UO_1939 (O_1939,N_19927,N_19884);
and UO_1940 (O_1940,N_19853,N_19869);
xnor UO_1941 (O_1941,N_19882,N_19904);
or UO_1942 (O_1942,N_19969,N_19970);
or UO_1943 (O_1943,N_19952,N_19890);
and UO_1944 (O_1944,N_19913,N_19997);
nand UO_1945 (O_1945,N_19891,N_19993);
and UO_1946 (O_1946,N_19999,N_19983);
nor UO_1947 (O_1947,N_19874,N_19978);
nand UO_1948 (O_1948,N_19855,N_19848);
or UO_1949 (O_1949,N_19864,N_19991);
nand UO_1950 (O_1950,N_19875,N_19914);
or UO_1951 (O_1951,N_19868,N_19855);
and UO_1952 (O_1952,N_19994,N_19988);
nand UO_1953 (O_1953,N_19982,N_19893);
or UO_1954 (O_1954,N_19845,N_19908);
and UO_1955 (O_1955,N_19882,N_19991);
nand UO_1956 (O_1956,N_19861,N_19999);
and UO_1957 (O_1957,N_19867,N_19915);
or UO_1958 (O_1958,N_19869,N_19844);
nand UO_1959 (O_1959,N_19941,N_19990);
nor UO_1960 (O_1960,N_19890,N_19991);
nand UO_1961 (O_1961,N_19975,N_19903);
nand UO_1962 (O_1962,N_19919,N_19875);
nand UO_1963 (O_1963,N_19870,N_19904);
or UO_1964 (O_1964,N_19993,N_19866);
or UO_1965 (O_1965,N_19972,N_19859);
and UO_1966 (O_1966,N_19963,N_19953);
nand UO_1967 (O_1967,N_19992,N_19956);
nand UO_1968 (O_1968,N_19876,N_19998);
nand UO_1969 (O_1969,N_19889,N_19909);
nand UO_1970 (O_1970,N_19883,N_19884);
and UO_1971 (O_1971,N_19878,N_19905);
nor UO_1972 (O_1972,N_19990,N_19902);
nor UO_1973 (O_1973,N_19853,N_19976);
xor UO_1974 (O_1974,N_19980,N_19974);
nand UO_1975 (O_1975,N_19946,N_19907);
nand UO_1976 (O_1976,N_19856,N_19885);
or UO_1977 (O_1977,N_19870,N_19858);
nor UO_1978 (O_1978,N_19844,N_19934);
or UO_1979 (O_1979,N_19902,N_19913);
nand UO_1980 (O_1980,N_19892,N_19951);
xor UO_1981 (O_1981,N_19934,N_19909);
xor UO_1982 (O_1982,N_19959,N_19885);
nor UO_1983 (O_1983,N_19903,N_19907);
and UO_1984 (O_1984,N_19999,N_19975);
or UO_1985 (O_1985,N_19891,N_19933);
nand UO_1986 (O_1986,N_19911,N_19974);
or UO_1987 (O_1987,N_19844,N_19930);
and UO_1988 (O_1988,N_19940,N_19914);
or UO_1989 (O_1989,N_19864,N_19971);
or UO_1990 (O_1990,N_19941,N_19992);
nand UO_1991 (O_1991,N_19986,N_19982);
xor UO_1992 (O_1992,N_19958,N_19989);
nor UO_1993 (O_1993,N_19872,N_19963);
xnor UO_1994 (O_1994,N_19890,N_19971);
nand UO_1995 (O_1995,N_19911,N_19846);
and UO_1996 (O_1996,N_19904,N_19925);
and UO_1997 (O_1997,N_19927,N_19995);
nor UO_1998 (O_1998,N_19997,N_19910);
or UO_1999 (O_1999,N_19888,N_19997);
nand UO_2000 (O_2000,N_19879,N_19935);
xnor UO_2001 (O_2001,N_19938,N_19995);
nor UO_2002 (O_2002,N_19929,N_19982);
and UO_2003 (O_2003,N_19885,N_19918);
or UO_2004 (O_2004,N_19923,N_19986);
or UO_2005 (O_2005,N_19991,N_19954);
nand UO_2006 (O_2006,N_19840,N_19903);
and UO_2007 (O_2007,N_19921,N_19910);
and UO_2008 (O_2008,N_19897,N_19909);
nor UO_2009 (O_2009,N_19919,N_19928);
nor UO_2010 (O_2010,N_19993,N_19965);
xnor UO_2011 (O_2011,N_19867,N_19932);
and UO_2012 (O_2012,N_19862,N_19883);
or UO_2013 (O_2013,N_19880,N_19986);
xor UO_2014 (O_2014,N_19983,N_19843);
nor UO_2015 (O_2015,N_19894,N_19959);
and UO_2016 (O_2016,N_19935,N_19850);
or UO_2017 (O_2017,N_19864,N_19883);
and UO_2018 (O_2018,N_19932,N_19954);
and UO_2019 (O_2019,N_19947,N_19885);
nand UO_2020 (O_2020,N_19975,N_19848);
or UO_2021 (O_2021,N_19956,N_19842);
or UO_2022 (O_2022,N_19845,N_19907);
and UO_2023 (O_2023,N_19972,N_19885);
nand UO_2024 (O_2024,N_19998,N_19941);
and UO_2025 (O_2025,N_19844,N_19970);
nor UO_2026 (O_2026,N_19852,N_19960);
nand UO_2027 (O_2027,N_19910,N_19897);
and UO_2028 (O_2028,N_19943,N_19934);
nor UO_2029 (O_2029,N_19911,N_19991);
xnor UO_2030 (O_2030,N_19991,N_19852);
and UO_2031 (O_2031,N_19896,N_19866);
nor UO_2032 (O_2032,N_19856,N_19923);
nor UO_2033 (O_2033,N_19928,N_19855);
or UO_2034 (O_2034,N_19850,N_19895);
and UO_2035 (O_2035,N_19907,N_19928);
nor UO_2036 (O_2036,N_19978,N_19995);
and UO_2037 (O_2037,N_19871,N_19992);
nor UO_2038 (O_2038,N_19906,N_19862);
nor UO_2039 (O_2039,N_19946,N_19930);
and UO_2040 (O_2040,N_19983,N_19895);
nor UO_2041 (O_2041,N_19875,N_19992);
or UO_2042 (O_2042,N_19982,N_19895);
or UO_2043 (O_2043,N_19935,N_19926);
nand UO_2044 (O_2044,N_19861,N_19888);
and UO_2045 (O_2045,N_19953,N_19866);
nand UO_2046 (O_2046,N_19876,N_19847);
or UO_2047 (O_2047,N_19902,N_19972);
and UO_2048 (O_2048,N_19860,N_19964);
nor UO_2049 (O_2049,N_19954,N_19887);
or UO_2050 (O_2050,N_19983,N_19887);
xnor UO_2051 (O_2051,N_19921,N_19875);
and UO_2052 (O_2052,N_19871,N_19995);
or UO_2053 (O_2053,N_19933,N_19869);
nand UO_2054 (O_2054,N_19916,N_19866);
nand UO_2055 (O_2055,N_19931,N_19932);
and UO_2056 (O_2056,N_19974,N_19950);
or UO_2057 (O_2057,N_19910,N_19879);
or UO_2058 (O_2058,N_19915,N_19868);
or UO_2059 (O_2059,N_19912,N_19963);
and UO_2060 (O_2060,N_19900,N_19995);
nand UO_2061 (O_2061,N_19876,N_19922);
nor UO_2062 (O_2062,N_19983,N_19936);
or UO_2063 (O_2063,N_19921,N_19977);
nor UO_2064 (O_2064,N_19970,N_19901);
and UO_2065 (O_2065,N_19937,N_19863);
nor UO_2066 (O_2066,N_19874,N_19937);
nor UO_2067 (O_2067,N_19895,N_19958);
xnor UO_2068 (O_2068,N_19998,N_19967);
nand UO_2069 (O_2069,N_19868,N_19957);
xnor UO_2070 (O_2070,N_19856,N_19865);
and UO_2071 (O_2071,N_19865,N_19962);
and UO_2072 (O_2072,N_19877,N_19935);
nand UO_2073 (O_2073,N_19977,N_19966);
or UO_2074 (O_2074,N_19918,N_19967);
nand UO_2075 (O_2075,N_19892,N_19862);
xor UO_2076 (O_2076,N_19950,N_19849);
nand UO_2077 (O_2077,N_19948,N_19876);
nand UO_2078 (O_2078,N_19848,N_19869);
xnor UO_2079 (O_2079,N_19968,N_19900);
xor UO_2080 (O_2080,N_19958,N_19956);
and UO_2081 (O_2081,N_19942,N_19903);
or UO_2082 (O_2082,N_19989,N_19866);
nor UO_2083 (O_2083,N_19933,N_19978);
nand UO_2084 (O_2084,N_19902,N_19958);
nor UO_2085 (O_2085,N_19841,N_19947);
nor UO_2086 (O_2086,N_19922,N_19882);
nand UO_2087 (O_2087,N_19893,N_19846);
and UO_2088 (O_2088,N_19999,N_19865);
nor UO_2089 (O_2089,N_19990,N_19949);
xor UO_2090 (O_2090,N_19917,N_19960);
nand UO_2091 (O_2091,N_19854,N_19967);
and UO_2092 (O_2092,N_19845,N_19941);
and UO_2093 (O_2093,N_19883,N_19870);
nor UO_2094 (O_2094,N_19945,N_19926);
nand UO_2095 (O_2095,N_19949,N_19992);
nor UO_2096 (O_2096,N_19991,N_19862);
and UO_2097 (O_2097,N_19852,N_19986);
or UO_2098 (O_2098,N_19931,N_19970);
and UO_2099 (O_2099,N_19871,N_19965);
nand UO_2100 (O_2100,N_19984,N_19902);
nand UO_2101 (O_2101,N_19997,N_19977);
nor UO_2102 (O_2102,N_19874,N_19883);
xnor UO_2103 (O_2103,N_19967,N_19913);
nor UO_2104 (O_2104,N_19894,N_19847);
nor UO_2105 (O_2105,N_19981,N_19983);
nor UO_2106 (O_2106,N_19863,N_19852);
nor UO_2107 (O_2107,N_19943,N_19926);
nor UO_2108 (O_2108,N_19945,N_19869);
or UO_2109 (O_2109,N_19846,N_19986);
nand UO_2110 (O_2110,N_19981,N_19961);
or UO_2111 (O_2111,N_19910,N_19983);
nand UO_2112 (O_2112,N_19978,N_19856);
or UO_2113 (O_2113,N_19916,N_19983);
nand UO_2114 (O_2114,N_19979,N_19953);
or UO_2115 (O_2115,N_19994,N_19949);
or UO_2116 (O_2116,N_19845,N_19885);
and UO_2117 (O_2117,N_19939,N_19965);
and UO_2118 (O_2118,N_19846,N_19844);
and UO_2119 (O_2119,N_19901,N_19952);
nor UO_2120 (O_2120,N_19912,N_19841);
or UO_2121 (O_2121,N_19952,N_19845);
nand UO_2122 (O_2122,N_19895,N_19888);
nor UO_2123 (O_2123,N_19923,N_19893);
and UO_2124 (O_2124,N_19867,N_19965);
nand UO_2125 (O_2125,N_19923,N_19890);
and UO_2126 (O_2126,N_19904,N_19970);
xnor UO_2127 (O_2127,N_19902,N_19854);
nor UO_2128 (O_2128,N_19924,N_19916);
or UO_2129 (O_2129,N_19845,N_19997);
nor UO_2130 (O_2130,N_19954,N_19891);
or UO_2131 (O_2131,N_19874,N_19876);
and UO_2132 (O_2132,N_19966,N_19939);
nor UO_2133 (O_2133,N_19955,N_19924);
and UO_2134 (O_2134,N_19878,N_19953);
nor UO_2135 (O_2135,N_19917,N_19913);
and UO_2136 (O_2136,N_19849,N_19935);
nand UO_2137 (O_2137,N_19969,N_19942);
and UO_2138 (O_2138,N_19999,N_19845);
nor UO_2139 (O_2139,N_19875,N_19874);
nor UO_2140 (O_2140,N_19912,N_19978);
or UO_2141 (O_2141,N_19874,N_19897);
and UO_2142 (O_2142,N_19841,N_19879);
nand UO_2143 (O_2143,N_19999,N_19986);
nand UO_2144 (O_2144,N_19915,N_19961);
or UO_2145 (O_2145,N_19983,N_19996);
and UO_2146 (O_2146,N_19874,N_19924);
or UO_2147 (O_2147,N_19868,N_19862);
or UO_2148 (O_2148,N_19941,N_19866);
xor UO_2149 (O_2149,N_19891,N_19877);
nor UO_2150 (O_2150,N_19970,N_19952);
nand UO_2151 (O_2151,N_19946,N_19999);
nand UO_2152 (O_2152,N_19874,N_19864);
nor UO_2153 (O_2153,N_19925,N_19958);
and UO_2154 (O_2154,N_19893,N_19875);
nor UO_2155 (O_2155,N_19959,N_19899);
and UO_2156 (O_2156,N_19983,N_19912);
xnor UO_2157 (O_2157,N_19958,N_19922);
or UO_2158 (O_2158,N_19850,N_19947);
nor UO_2159 (O_2159,N_19845,N_19996);
or UO_2160 (O_2160,N_19994,N_19942);
and UO_2161 (O_2161,N_19941,N_19977);
and UO_2162 (O_2162,N_19949,N_19852);
nor UO_2163 (O_2163,N_19842,N_19938);
xnor UO_2164 (O_2164,N_19853,N_19974);
nor UO_2165 (O_2165,N_19888,N_19890);
nand UO_2166 (O_2166,N_19890,N_19929);
xnor UO_2167 (O_2167,N_19842,N_19969);
nor UO_2168 (O_2168,N_19862,N_19894);
or UO_2169 (O_2169,N_19918,N_19905);
nand UO_2170 (O_2170,N_19918,N_19874);
nor UO_2171 (O_2171,N_19845,N_19947);
and UO_2172 (O_2172,N_19893,N_19983);
nand UO_2173 (O_2173,N_19969,N_19906);
xor UO_2174 (O_2174,N_19971,N_19929);
nor UO_2175 (O_2175,N_19840,N_19864);
or UO_2176 (O_2176,N_19846,N_19952);
nand UO_2177 (O_2177,N_19927,N_19984);
xnor UO_2178 (O_2178,N_19978,N_19849);
or UO_2179 (O_2179,N_19989,N_19957);
nor UO_2180 (O_2180,N_19850,N_19950);
and UO_2181 (O_2181,N_19888,N_19948);
or UO_2182 (O_2182,N_19864,N_19887);
nand UO_2183 (O_2183,N_19935,N_19973);
and UO_2184 (O_2184,N_19970,N_19936);
xor UO_2185 (O_2185,N_19994,N_19850);
or UO_2186 (O_2186,N_19850,N_19906);
nand UO_2187 (O_2187,N_19884,N_19933);
nor UO_2188 (O_2188,N_19956,N_19908);
and UO_2189 (O_2189,N_19961,N_19968);
nor UO_2190 (O_2190,N_19940,N_19915);
nand UO_2191 (O_2191,N_19985,N_19901);
or UO_2192 (O_2192,N_19996,N_19981);
or UO_2193 (O_2193,N_19926,N_19919);
or UO_2194 (O_2194,N_19877,N_19916);
nand UO_2195 (O_2195,N_19964,N_19991);
nand UO_2196 (O_2196,N_19957,N_19849);
nor UO_2197 (O_2197,N_19923,N_19891);
nand UO_2198 (O_2198,N_19998,N_19957);
xnor UO_2199 (O_2199,N_19844,N_19894);
or UO_2200 (O_2200,N_19976,N_19922);
and UO_2201 (O_2201,N_19863,N_19845);
nand UO_2202 (O_2202,N_19871,N_19861);
nor UO_2203 (O_2203,N_19925,N_19914);
xnor UO_2204 (O_2204,N_19923,N_19980);
nand UO_2205 (O_2205,N_19881,N_19947);
and UO_2206 (O_2206,N_19927,N_19991);
and UO_2207 (O_2207,N_19943,N_19851);
and UO_2208 (O_2208,N_19925,N_19977);
and UO_2209 (O_2209,N_19959,N_19952);
nand UO_2210 (O_2210,N_19981,N_19962);
nand UO_2211 (O_2211,N_19848,N_19997);
xnor UO_2212 (O_2212,N_19948,N_19897);
or UO_2213 (O_2213,N_19983,N_19950);
nor UO_2214 (O_2214,N_19974,N_19878);
nand UO_2215 (O_2215,N_19863,N_19878);
and UO_2216 (O_2216,N_19904,N_19990);
nand UO_2217 (O_2217,N_19845,N_19851);
and UO_2218 (O_2218,N_19880,N_19923);
nor UO_2219 (O_2219,N_19931,N_19992);
nor UO_2220 (O_2220,N_19917,N_19948);
nor UO_2221 (O_2221,N_19956,N_19855);
nand UO_2222 (O_2222,N_19960,N_19912);
nor UO_2223 (O_2223,N_19934,N_19942);
and UO_2224 (O_2224,N_19973,N_19906);
and UO_2225 (O_2225,N_19883,N_19944);
xor UO_2226 (O_2226,N_19889,N_19989);
nand UO_2227 (O_2227,N_19958,N_19933);
nor UO_2228 (O_2228,N_19859,N_19896);
nand UO_2229 (O_2229,N_19879,N_19928);
nor UO_2230 (O_2230,N_19968,N_19898);
nand UO_2231 (O_2231,N_19953,N_19874);
xnor UO_2232 (O_2232,N_19860,N_19933);
nand UO_2233 (O_2233,N_19932,N_19924);
and UO_2234 (O_2234,N_19913,N_19875);
or UO_2235 (O_2235,N_19960,N_19935);
and UO_2236 (O_2236,N_19851,N_19865);
or UO_2237 (O_2237,N_19917,N_19965);
nor UO_2238 (O_2238,N_19982,N_19952);
xnor UO_2239 (O_2239,N_19906,N_19907);
xnor UO_2240 (O_2240,N_19991,N_19878);
and UO_2241 (O_2241,N_19923,N_19854);
nand UO_2242 (O_2242,N_19908,N_19920);
nand UO_2243 (O_2243,N_19935,N_19936);
nand UO_2244 (O_2244,N_19986,N_19921);
nand UO_2245 (O_2245,N_19885,N_19948);
nor UO_2246 (O_2246,N_19957,N_19872);
and UO_2247 (O_2247,N_19863,N_19841);
and UO_2248 (O_2248,N_19996,N_19843);
or UO_2249 (O_2249,N_19845,N_19975);
xnor UO_2250 (O_2250,N_19987,N_19911);
or UO_2251 (O_2251,N_19986,N_19877);
nor UO_2252 (O_2252,N_19958,N_19966);
xnor UO_2253 (O_2253,N_19990,N_19866);
nand UO_2254 (O_2254,N_19938,N_19849);
and UO_2255 (O_2255,N_19881,N_19880);
or UO_2256 (O_2256,N_19898,N_19914);
and UO_2257 (O_2257,N_19960,N_19903);
nand UO_2258 (O_2258,N_19932,N_19923);
nand UO_2259 (O_2259,N_19886,N_19957);
and UO_2260 (O_2260,N_19969,N_19935);
nor UO_2261 (O_2261,N_19981,N_19854);
nor UO_2262 (O_2262,N_19875,N_19933);
nand UO_2263 (O_2263,N_19853,N_19999);
nor UO_2264 (O_2264,N_19850,N_19841);
xnor UO_2265 (O_2265,N_19840,N_19942);
or UO_2266 (O_2266,N_19983,N_19858);
and UO_2267 (O_2267,N_19974,N_19959);
or UO_2268 (O_2268,N_19866,N_19954);
xor UO_2269 (O_2269,N_19926,N_19930);
or UO_2270 (O_2270,N_19968,N_19915);
or UO_2271 (O_2271,N_19990,N_19991);
nor UO_2272 (O_2272,N_19930,N_19998);
or UO_2273 (O_2273,N_19849,N_19952);
or UO_2274 (O_2274,N_19978,N_19955);
or UO_2275 (O_2275,N_19957,N_19857);
or UO_2276 (O_2276,N_19948,N_19964);
nor UO_2277 (O_2277,N_19846,N_19958);
nor UO_2278 (O_2278,N_19968,N_19935);
xnor UO_2279 (O_2279,N_19850,N_19902);
nor UO_2280 (O_2280,N_19859,N_19866);
xnor UO_2281 (O_2281,N_19994,N_19877);
or UO_2282 (O_2282,N_19976,N_19960);
nor UO_2283 (O_2283,N_19888,N_19848);
xnor UO_2284 (O_2284,N_19908,N_19968);
xor UO_2285 (O_2285,N_19881,N_19892);
nor UO_2286 (O_2286,N_19915,N_19935);
nor UO_2287 (O_2287,N_19889,N_19975);
nand UO_2288 (O_2288,N_19847,N_19990);
nand UO_2289 (O_2289,N_19969,N_19884);
xnor UO_2290 (O_2290,N_19980,N_19913);
xor UO_2291 (O_2291,N_19897,N_19855);
xor UO_2292 (O_2292,N_19898,N_19955);
nor UO_2293 (O_2293,N_19898,N_19843);
or UO_2294 (O_2294,N_19925,N_19871);
nor UO_2295 (O_2295,N_19861,N_19962);
xnor UO_2296 (O_2296,N_19981,N_19954);
xor UO_2297 (O_2297,N_19897,N_19883);
and UO_2298 (O_2298,N_19852,N_19847);
or UO_2299 (O_2299,N_19990,N_19974);
nor UO_2300 (O_2300,N_19873,N_19881);
and UO_2301 (O_2301,N_19843,N_19868);
xor UO_2302 (O_2302,N_19973,N_19940);
or UO_2303 (O_2303,N_19910,N_19985);
or UO_2304 (O_2304,N_19955,N_19922);
or UO_2305 (O_2305,N_19901,N_19967);
nand UO_2306 (O_2306,N_19951,N_19871);
and UO_2307 (O_2307,N_19996,N_19957);
or UO_2308 (O_2308,N_19930,N_19877);
or UO_2309 (O_2309,N_19894,N_19852);
nor UO_2310 (O_2310,N_19841,N_19910);
xor UO_2311 (O_2311,N_19957,N_19972);
or UO_2312 (O_2312,N_19995,N_19895);
xor UO_2313 (O_2313,N_19995,N_19872);
xor UO_2314 (O_2314,N_19965,N_19952);
nand UO_2315 (O_2315,N_19906,N_19937);
or UO_2316 (O_2316,N_19930,N_19928);
nor UO_2317 (O_2317,N_19859,N_19914);
or UO_2318 (O_2318,N_19878,N_19915);
and UO_2319 (O_2319,N_19998,N_19927);
xnor UO_2320 (O_2320,N_19903,N_19869);
and UO_2321 (O_2321,N_19928,N_19914);
nand UO_2322 (O_2322,N_19887,N_19938);
xnor UO_2323 (O_2323,N_19969,N_19957);
nand UO_2324 (O_2324,N_19970,N_19967);
and UO_2325 (O_2325,N_19972,N_19938);
nand UO_2326 (O_2326,N_19894,N_19936);
or UO_2327 (O_2327,N_19843,N_19867);
nand UO_2328 (O_2328,N_19878,N_19977);
nand UO_2329 (O_2329,N_19873,N_19967);
nor UO_2330 (O_2330,N_19915,N_19856);
nand UO_2331 (O_2331,N_19977,N_19891);
or UO_2332 (O_2332,N_19907,N_19847);
xnor UO_2333 (O_2333,N_19964,N_19983);
or UO_2334 (O_2334,N_19842,N_19994);
nand UO_2335 (O_2335,N_19902,N_19967);
and UO_2336 (O_2336,N_19897,N_19995);
or UO_2337 (O_2337,N_19941,N_19873);
nand UO_2338 (O_2338,N_19959,N_19953);
and UO_2339 (O_2339,N_19899,N_19991);
and UO_2340 (O_2340,N_19921,N_19907);
nand UO_2341 (O_2341,N_19985,N_19965);
and UO_2342 (O_2342,N_19919,N_19975);
and UO_2343 (O_2343,N_19921,N_19949);
xor UO_2344 (O_2344,N_19894,N_19892);
nand UO_2345 (O_2345,N_19945,N_19859);
xor UO_2346 (O_2346,N_19907,N_19881);
nor UO_2347 (O_2347,N_19928,N_19849);
nor UO_2348 (O_2348,N_19850,N_19991);
or UO_2349 (O_2349,N_19904,N_19903);
nand UO_2350 (O_2350,N_19919,N_19964);
nand UO_2351 (O_2351,N_19911,N_19916);
or UO_2352 (O_2352,N_19866,N_19961);
nor UO_2353 (O_2353,N_19893,N_19874);
and UO_2354 (O_2354,N_19912,N_19973);
nand UO_2355 (O_2355,N_19904,N_19894);
nand UO_2356 (O_2356,N_19958,N_19911);
nand UO_2357 (O_2357,N_19848,N_19950);
xor UO_2358 (O_2358,N_19970,N_19956);
and UO_2359 (O_2359,N_19921,N_19940);
nor UO_2360 (O_2360,N_19993,N_19998);
and UO_2361 (O_2361,N_19871,N_19851);
and UO_2362 (O_2362,N_19877,N_19945);
nor UO_2363 (O_2363,N_19914,N_19998);
nor UO_2364 (O_2364,N_19941,N_19901);
nand UO_2365 (O_2365,N_19993,N_19845);
and UO_2366 (O_2366,N_19888,N_19914);
nor UO_2367 (O_2367,N_19906,N_19846);
nand UO_2368 (O_2368,N_19841,N_19886);
and UO_2369 (O_2369,N_19900,N_19982);
nand UO_2370 (O_2370,N_19949,N_19959);
and UO_2371 (O_2371,N_19911,N_19999);
nand UO_2372 (O_2372,N_19960,N_19879);
or UO_2373 (O_2373,N_19860,N_19958);
or UO_2374 (O_2374,N_19851,N_19923);
nand UO_2375 (O_2375,N_19977,N_19910);
or UO_2376 (O_2376,N_19977,N_19959);
nand UO_2377 (O_2377,N_19959,N_19926);
and UO_2378 (O_2378,N_19858,N_19902);
and UO_2379 (O_2379,N_19842,N_19922);
and UO_2380 (O_2380,N_19887,N_19921);
and UO_2381 (O_2381,N_19971,N_19978);
nand UO_2382 (O_2382,N_19856,N_19972);
nand UO_2383 (O_2383,N_19851,N_19902);
or UO_2384 (O_2384,N_19932,N_19853);
or UO_2385 (O_2385,N_19847,N_19972);
nand UO_2386 (O_2386,N_19933,N_19932);
and UO_2387 (O_2387,N_19898,N_19897);
nor UO_2388 (O_2388,N_19955,N_19930);
and UO_2389 (O_2389,N_19947,N_19897);
or UO_2390 (O_2390,N_19943,N_19960);
nand UO_2391 (O_2391,N_19854,N_19908);
nand UO_2392 (O_2392,N_19966,N_19954);
and UO_2393 (O_2393,N_19841,N_19915);
and UO_2394 (O_2394,N_19977,N_19976);
nor UO_2395 (O_2395,N_19944,N_19864);
nand UO_2396 (O_2396,N_19965,N_19947);
nand UO_2397 (O_2397,N_19919,N_19999);
and UO_2398 (O_2398,N_19987,N_19900);
xor UO_2399 (O_2399,N_19923,N_19929);
and UO_2400 (O_2400,N_19899,N_19844);
nand UO_2401 (O_2401,N_19890,N_19990);
nand UO_2402 (O_2402,N_19952,N_19928);
and UO_2403 (O_2403,N_19965,N_19987);
nand UO_2404 (O_2404,N_19895,N_19922);
and UO_2405 (O_2405,N_19922,N_19925);
and UO_2406 (O_2406,N_19965,N_19881);
or UO_2407 (O_2407,N_19976,N_19970);
or UO_2408 (O_2408,N_19938,N_19926);
or UO_2409 (O_2409,N_19859,N_19897);
nor UO_2410 (O_2410,N_19932,N_19998);
nor UO_2411 (O_2411,N_19939,N_19885);
and UO_2412 (O_2412,N_19867,N_19888);
or UO_2413 (O_2413,N_19936,N_19853);
nor UO_2414 (O_2414,N_19887,N_19967);
and UO_2415 (O_2415,N_19921,N_19931);
nand UO_2416 (O_2416,N_19907,N_19938);
and UO_2417 (O_2417,N_19924,N_19976);
or UO_2418 (O_2418,N_19881,N_19851);
xor UO_2419 (O_2419,N_19989,N_19843);
nand UO_2420 (O_2420,N_19885,N_19862);
nor UO_2421 (O_2421,N_19903,N_19882);
nand UO_2422 (O_2422,N_19927,N_19900);
xor UO_2423 (O_2423,N_19978,N_19894);
nor UO_2424 (O_2424,N_19896,N_19862);
and UO_2425 (O_2425,N_19870,N_19993);
or UO_2426 (O_2426,N_19950,N_19891);
and UO_2427 (O_2427,N_19868,N_19886);
or UO_2428 (O_2428,N_19980,N_19845);
or UO_2429 (O_2429,N_19847,N_19911);
nor UO_2430 (O_2430,N_19883,N_19968);
nor UO_2431 (O_2431,N_19867,N_19889);
or UO_2432 (O_2432,N_19885,N_19891);
nand UO_2433 (O_2433,N_19896,N_19996);
nor UO_2434 (O_2434,N_19854,N_19946);
nand UO_2435 (O_2435,N_19945,N_19974);
xnor UO_2436 (O_2436,N_19951,N_19935);
and UO_2437 (O_2437,N_19971,N_19952);
nor UO_2438 (O_2438,N_19923,N_19905);
xor UO_2439 (O_2439,N_19973,N_19861);
nand UO_2440 (O_2440,N_19989,N_19891);
nor UO_2441 (O_2441,N_19875,N_19888);
nor UO_2442 (O_2442,N_19979,N_19916);
nor UO_2443 (O_2443,N_19907,N_19895);
nand UO_2444 (O_2444,N_19921,N_19961);
nor UO_2445 (O_2445,N_19961,N_19947);
and UO_2446 (O_2446,N_19969,N_19899);
and UO_2447 (O_2447,N_19927,N_19937);
nand UO_2448 (O_2448,N_19889,N_19861);
nor UO_2449 (O_2449,N_19951,N_19867);
or UO_2450 (O_2450,N_19872,N_19939);
and UO_2451 (O_2451,N_19949,N_19925);
and UO_2452 (O_2452,N_19867,N_19858);
or UO_2453 (O_2453,N_19876,N_19859);
or UO_2454 (O_2454,N_19984,N_19848);
or UO_2455 (O_2455,N_19976,N_19931);
or UO_2456 (O_2456,N_19936,N_19991);
nor UO_2457 (O_2457,N_19914,N_19977);
nor UO_2458 (O_2458,N_19995,N_19986);
or UO_2459 (O_2459,N_19931,N_19929);
and UO_2460 (O_2460,N_19865,N_19928);
or UO_2461 (O_2461,N_19946,N_19910);
nor UO_2462 (O_2462,N_19946,N_19862);
nand UO_2463 (O_2463,N_19915,N_19969);
xor UO_2464 (O_2464,N_19904,N_19867);
nand UO_2465 (O_2465,N_19925,N_19903);
xnor UO_2466 (O_2466,N_19925,N_19917);
and UO_2467 (O_2467,N_19927,N_19986);
nand UO_2468 (O_2468,N_19975,N_19972);
nand UO_2469 (O_2469,N_19859,N_19913);
or UO_2470 (O_2470,N_19896,N_19857);
nand UO_2471 (O_2471,N_19868,N_19999);
and UO_2472 (O_2472,N_19840,N_19992);
xnor UO_2473 (O_2473,N_19997,N_19958);
xor UO_2474 (O_2474,N_19962,N_19858);
xnor UO_2475 (O_2475,N_19842,N_19863);
nor UO_2476 (O_2476,N_19940,N_19938);
nand UO_2477 (O_2477,N_19905,N_19938);
nand UO_2478 (O_2478,N_19844,N_19954);
nor UO_2479 (O_2479,N_19993,N_19884);
and UO_2480 (O_2480,N_19985,N_19868);
and UO_2481 (O_2481,N_19989,N_19908);
and UO_2482 (O_2482,N_19905,N_19995);
or UO_2483 (O_2483,N_19887,N_19949);
nor UO_2484 (O_2484,N_19922,N_19867);
and UO_2485 (O_2485,N_19962,N_19872);
nor UO_2486 (O_2486,N_19939,N_19988);
xor UO_2487 (O_2487,N_19990,N_19870);
or UO_2488 (O_2488,N_19864,N_19938);
nor UO_2489 (O_2489,N_19910,N_19887);
nor UO_2490 (O_2490,N_19945,N_19920);
nand UO_2491 (O_2491,N_19899,N_19933);
or UO_2492 (O_2492,N_19878,N_19927);
nor UO_2493 (O_2493,N_19953,N_19978);
and UO_2494 (O_2494,N_19996,N_19960);
nand UO_2495 (O_2495,N_19911,N_19988);
nand UO_2496 (O_2496,N_19996,N_19977);
and UO_2497 (O_2497,N_19893,N_19901);
and UO_2498 (O_2498,N_19970,N_19984);
nor UO_2499 (O_2499,N_19943,N_19977);
endmodule