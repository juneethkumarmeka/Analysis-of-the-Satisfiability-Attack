module basic_1000_10000_1500_20_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_396,In_728);
and U1 (N_1,In_761,In_104);
and U2 (N_2,In_779,In_3);
nor U3 (N_3,In_833,In_380);
and U4 (N_4,In_116,In_307);
xnor U5 (N_5,In_40,In_2);
nor U6 (N_6,In_676,In_288);
xor U7 (N_7,In_648,In_846);
and U8 (N_8,In_128,In_285);
nor U9 (N_9,In_952,In_91);
nor U10 (N_10,In_967,In_826);
or U11 (N_11,In_989,In_312);
nand U12 (N_12,In_339,In_503);
nor U13 (N_13,In_680,In_295);
or U14 (N_14,In_379,In_386);
nand U15 (N_15,In_519,In_161);
and U16 (N_16,In_12,In_460);
nand U17 (N_17,In_287,In_303);
or U18 (N_18,In_257,In_335);
nand U19 (N_19,In_462,In_271);
and U20 (N_20,In_583,In_100);
nand U21 (N_21,In_572,In_406);
or U22 (N_22,In_475,In_507);
nand U23 (N_23,In_914,In_997);
or U24 (N_24,In_927,In_515);
or U25 (N_25,In_336,In_796);
and U26 (N_26,In_535,In_357);
nand U27 (N_27,In_117,In_421);
nor U28 (N_28,In_979,In_227);
nand U29 (N_29,In_463,In_646);
and U30 (N_30,In_478,In_407);
or U31 (N_31,In_970,In_539);
nand U32 (N_32,In_935,In_780);
nand U33 (N_33,In_494,In_882);
xnor U34 (N_34,In_769,In_650);
nand U35 (N_35,In_317,In_436);
xnor U36 (N_36,In_690,In_345);
or U37 (N_37,In_936,In_305);
xnor U38 (N_38,In_652,In_181);
and U39 (N_39,In_66,In_713);
nor U40 (N_40,In_84,In_381);
nand U41 (N_41,In_455,In_415);
nor U42 (N_42,In_487,In_541);
or U43 (N_43,In_189,In_258);
nor U44 (N_44,In_965,In_332);
nor U45 (N_45,In_738,In_166);
or U46 (N_46,In_47,In_289);
nor U47 (N_47,In_701,In_638);
nor U48 (N_48,In_996,In_919);
or U49 (N_49,In_270,In_810);
nor U50 (N_50,In_746,In_759);
nand U51 (N_51,In_851,In_981);
and U52 (N_52,In_279,In_51);
and U53 (N_53,In_887,In_580);
xnor U54 (N_54,In_20,In_502);
and U55 (N_55,In_448,In_586);
xnor U56 (N_56,In_318,In_777);
nor U57 (N_57,In_784,In_624);
or U58 (N_58,In_226,In_392);
and U59 (N_59,In_955,In_957);
or U60 (N_60,In_71,In_528);
and U61 (N_61,In_958,In_825);
or U62 (N_62,In_221,In_251);
or U63 (N_63,In_488,In_642);
nand U64 (N_64,In_69,In_15);
and U65 (N_65,In_217,In_457);
nand U66 (N_66,In_53,In_361);
and U67 (N_67,In_671,In_425);
and U68 (N_68,In_194,In_19);
nand U69 (N_69,In_554,In_588);
or U70 (N_70,In_772,In_504);
nor U71 (N_71,In_155,In_950);
xor U72 (N_72,In_182,In_630);
or U73 (N_73,In_862,In_120);
nor U74 (N_74,In_685,In_450);
nor U75 (N_75,In_605,In_860);
or U76 (N_76,In_716,In_677);
and U77 (N_77,In_449,In_75);
xor U78 (N_78,In_103,In_290);
nor U79 (N_79,In_923,In_467);
nor U80 (N_80,In_234,In_571);
nand U81 (N_81,In_172,In_253);
nor U82 (N_82,In_980,In_340);
nor U83 (N_83,In_831,In_248);
or U84 (N_84,In_698,In_484);
nand U85 (N_85,In_758,In_64);
nor U86 (N_86,In_751,In_578);
or U87 (N_87,In_865,In_138);
and U88 (N_88,In_293,In_562);
nand U89 (N_89,In_900,In_830);
nor U90 (N_90,In_394,In_978);
or U91 (N_91,In_669,In_343);
nor U92 (N_92,In_323,In_230);
nand U93 (N_93,In_885,In_39);
nor U94 (N_94,In_992,In_156);
nor U95 (N_95,In_988,In_843);
xor U96 (N_96,In_24,In_247);
or U97 (N_97,In_619,In_41);
nor U98 (N_98,In_417,In_430);
or U99 (N_99,In_294,In_135);
and U100 (N_100,In_274,In_960);
or U101 (N_101,In_577,In_543);
or U102 (N_102,In_917,In_351);
and U103 (N_103,In_414,In_260);
or U104 (N_104,In_801,In_125);
and U105 (N_105,In_940,In_358);
nand U106 (N_106,In_880,In_835);
or U107 (N_107,In_232,In_949);
xor U108 (N_108,In_842,In_441);
nor U109 (N_109,In_276,In_327);
nor U110 (N_110,In_495,In_68);
nor U111 (N_111,In_492,In_781);
nor U112 (N_112,In_569,In_454);
nand U113 (N_113,In_590,In_889);
and U114 (N_114,In_344,In_410);
or U115 (N_115,In_333,In_96);
nor U116 (N_116,In_942,In_284);
nand U117 (N_117,In_299,In_141);
or U118 (N_118,In_579,In_309);
or U119 (N_119,In_458,In_218);
or U120 (N_120,In_982,In_177);
or U121 (N_121,In_124,In_849);
nand U122 (N_122,In_99,In_250);
and U123 (N_123,In_614,In_371);
or U124 (N_124,In_239,In_57);
nand U125 (N_125,In_385,In_121);
or U126 (N_126,In_898,In_192);
nor U127 (N_127,In_438,In_593);
nor U128 (N_128,In_640,In_850);
and U129 (N_129,In_62,In_520);
nor U130 (N_130,In_498,In_757);
nor U131 (N_131,In_211,In_373);
xor U132 (N_132,In_665,In_983);
nor U133 (N_133,In_760,In_473);
nor U134 (N_134,In_87,In_545);
and U135 (N_135,In_552,In_891);
or U136 (N_136,In_721,In_868);
nand U137 (N_137,In_237,In_749);
and U138 (N_138,In_635,In_718);
and U139 (N_139,In_97,In_773);
or U140 (N_140,In_328,In_229);
nand U141 (N_141,In_643,In_301);
or U142 (N_142,In_555,In_703);
and U143 (N_143,In_506,In_240);
nor U144 (N_144,In_338,In_266);
and U145 (N_145,In_612,In_395);
nand U146 (N_146,In_311,In_252);
or U147 (N_147,In_966,In_876);
or U148 (N_148,In_601,In_819);
nand U149 (N_149,In_574,In_521);
or U150 (N_150,In_7,In_163);
nand U151 (N_151,In_342,In_522);
nor U152 (N_152,In_402,In_34);
nor U153 (N_153,In_179,In_264);
or U154 (N_154,In_742,In_720);
xor U155 (N_155,In_167,In_514);
nand U156 (N_156,In_687,In_783);
nor U157 (N_157,In_752,In_736);
nand U158 (N_158,In_468,In_233);
or U159 (N_159,In_602,In_59);
nand U160 (N_160,In_178,In_176);
nand U161 (N_161,In_13,In_532);
nand U162 (N_162,In_998,In_723);
nor U163 (N_163,In_472,In_527);
nand U164 (N_164,In_304,In_364);
or U165 (N_165,In_81,In_717);
and U166 (N_166,In_821,In_112);
nand U167 (N_167,In_744,In_409);
and U168 (N_168,In_60,In_429);
nor U169 (N_169,In_215,In_461);
or U170 (N_170,In_667,In_146);
nand U171 (N_171,In_213,In_707);
nor U172 (N_172,In_452,In_416);
or U173 (N_173,In_873,In_205);
nand U174 (N_174,In_105,In_5);
xnor U175 (N_175,In_610,In_670);
and U176 (N_176,In_209,In_65);
nand U177 (N_177,In_929,In_72);
nor U178 (N_178,In_423,In_765);
or U179 (N_179,In_735,In_383);
nor U180 (N_180,In_754,In_613);
nand U181 (N_181,In_444,In_730);
xor U182 (N_182,In_54,In_788);
nor U183 (N_183,In_489,In_168);
xor U184 (N_184,In_975,In_208);
xnor U185 (N_185,In_422,In_994);
and U186 (N_186,In_679,In_536);
nor U187 (N_187,In_948,In_434);
or U188 (N_188,In_298,In_805);
or U189 (N_189,In_786,In_193);
xor U190 (N_190,In_734,In_594);
or U191 (N_191,In_426,In_322);
xor U192 (N_192,In_755,In_627);
and U193 (N_193,In_611,In_661);
and U194 (N_194,In_896,In_911);
nand U195 (N_195,In_326,In_915);
nor U196 (N_196,In_88,In_265);
or U197 (N_197,In_497,In_49);
nand U198 (N_198,In_102,In_477);
nand U199 (N_199,In_775,In_171);
or U200 (N_200,In_798,In_726);
nor U201 (N_201,In_145,In_664);
and U202 (N_202,In_523,In_715);
nor U203 (N_203,In_482,In_341);
nand U204 (N_204,In_870,In_795);
or U205 (N_205,In_771,In_848);
and U206 (N_206,In_618,In_890);
nor U207 (N_207,In_280,In_656);
or U208 (N_208,In_154,In_678);
xnor U209 (N_209,In_45,In_708);
nor U210 (N_210,In_297,In_724);
nor U211 (N_211,In_872,In_725);
nand U212 (N_212,In_479,In_518);
nor U213 (N_213,In_604,In_587);
or U214 (N_214,In_273,In_115);
and U215 (N_215,In_313,In_499);
or U216 (N_216,In_241,In_645);
nand U217 (N_217,In_249,In_706);
nand U218 (N_218,In_954,In_691);
nor U219 (N_219,In_324,In_354);
nand U220 (N_220,In_681,In_733);
and U221 (N_221,In_400,In_52);
and U222 (N_222,In_334,In_557);
or U223 (N_223,In_42,In_470);
nor U224 (N_224,In_930,In_858);
or U225 (N_225,In_30,In_537);
nand U226 (N_226,In_660,In_516);
nor U227 (N_227,In_634,In_568);
or U228 (N_228,In_712,In_158);
xor U229 (N_229,In_35,In_946);
and U230 (N_230,In_440,In_187);
nand U231 (N_231,In_362,In_620);
nor U232 (N_232,In_17,In_933);
or U233 (N_233,In_534,In_617);
nand U234 (N_234,In_413,In_107);
xnor U235 (N_235,In_861,In_790);
and U236 (N_236,In_762,In_325);
nor U237 (N_237,In_808,In_216);
xnor U238 (N_238,In_391,In_902);
nor U239 (N_239,In_609,In_531);
and U240 (N_240,In_228,In_697);
nor U241 (N_241,In_883,In_699);
and U242 (N_242,In_93,In_491);
and U243 (N_243,In_644,In_722);
or U244 (N_244,In_390,In_812);
nand U245 (N_245,In_855,In_196);
or U246 (N_246,In_33,In_576);
xnor U247 (N_247,In_442,In_944);
xnor U248 (N_248,In_231,In_180);
nand U249 (N_249,In_615,In_985);
nand U250 (N_250,In_23,In_223);
nor U251 (N_251,In_129,In_126);
nand U252 (N_252,In_791,In_131);
and U253 (N_253,In_346,In_575);
nor U254 (N_254,In_530,In_82);
or U255 (N_255,In_26,In_505);
and U256 (N_256,In_797,In_419);
nor U257 (N_257,In_672,In_269);
nand U258 (N_258,In_511,In_431);
nand U259 (N_259,In_37,In_320);
or U260 (N_260,In_76,In_608);
and U261 (N_261,In_149,In_824);
or U262 (N_262,In_695,In_401);
nor U263 (N_263,In_106,In_355);
nand U264 (N_264,In_943,In_404);
nor U265 (N_265,In_893,In_939);
nor U266 (N_266,In_398,In_673);
and U267 (N_267,In_551,In_43);
and U268 (N_268,In_356,In_418);
and U269 (N_269,In_631,In_89);
nor U270 (N_270,In_600,In_389);
or U271 (N_271,In_86,In_793);
nor U272 (N_272,In_971,In_603);
and U273 (N_273,In_828,In_159);
and U274 (N_274,In_741,In_922);
or U275 (N_275,In_913,In_711);
nor U276 (N_276,In_877,In_483);
and U277 (N_277,In_403,In_259);
nor U278 (N_278,In_369,In_83);
and U279 (N_279,In_525,In_973);
nand U280 (N_280,In_903,In_529);
and U281 (N_281,In_210,In_969);
or U282 (N_282,In_838,In_689);
xnor U283 (N_283,In_567,In_654);
nand U284 (N_284,In_839,In_219);
nor U285 (N_285,In_606,In_315);
or U286 (N_286,In_55,In_827);
or U287 (N_287,In_991,In_80);
nor U288 (N_288,In_85,In_548);
nand U289 (N_289,In_675,In_925);
and U290 (N_290,In_501,In_98);
nand U291 (N_291,In_151,In_435);
or U292 (N_292,In_823,In_330);
and U293 (N_293,In_888,In_466);
xnor U294 (N_294,In_702,In_683);
or U295 (N_295,In_292,In_244);
nor U296 (N_296,In_77,In_961);
nand U297 (N_297,In_186,In_682);
or U298 (N_298,In_195,In_73);
xnor U299 (N_299,In_490,In_832);
nand U300 (N_300,In_127,In_261);
nand U301 (N_301,In_553,In_353);
xnor U302 (N_302,In_533,In_766);
nor U303 (N_303,In_433,In_909);
nor U304 (N_304,In_142,In_352);
nor U305 (N_305,In_542,In_739);
nor U306 (N_306,In_109,In_753);
or U307 (N_307,In_393,In_694);
nand U308 (N_308,In_316,In_427);
nand U309 (N_309,In_509,In_254);
nor U310 (N_310,In_864,In_837);
xor U311 (N_311,In_496,In_686);
xor U312 (N_312,In_987,In_941);
or U313 (N_313,In_918,In_8);
nor U314 (N_314,In_485,In_243);
or U315 (N_315,In_756,In_693);
nor U316 (N_316,In_133,In_731);
nor U317 (N_317,In_729,In_546);
nor U318 (N_318,In_140,In_79);
or U319 (N_319,In_692,In_714);
nor U320 (N_320,In_118,In_225);
and U321 (N_321,In_770,In_986);
nand U322 (N_322,In_908,In_46);
nand U323 (N_323,In_147,In_659);
nor U324 (N_324,In_246,In_916);
nand U325 (N_325,In_275,In_148);
or U326 (N_326,In_28,In_905);
nor U327 (N_327,In_370,In_36);
nor U328 (N_328,In_170,In_150);
and U329 (N_329,In_408,In_513);
nand U330 (N_330,In_817,In_108);
or U331 (N_331,In_710,In_840);
and U332 (N_332,In_558,In_337);
and U333 (N_333,In_561,In_464);
xnor U334 (N_334,In_856,In_945);
nand U335 (N_335,In_844,In_727);
or U336 (N_336,In_447,In_74);
and U337 (N_337,In_964,In_700);
or U338 (N_338,In_607,In_405);
or U339 (N_339,In_816,In_32);
nand U340 (N_340,In_412,In_397);
xor U341 (N_341,In_589,In_633);
nand U342 (N_342,In_214,In_663);
or U343 (N_343,In_550,In_592);
nor U344 (N_344,In_122,In_382);
nand U345 (N_345,In_931,In_547);
or U346 (N_346,In_300,In_188);
nor U347 (N_347,In_480,In_570);
and U348 (N_348,In_465,In_165);
nand U349 (N_349,In_655,In_157);
nand U350 (N_350,In_367,In_329);
nor U351 (N_351,In_348,In_822);
and U352 (N_352,In_999,In_424);
and U353 (N_353,In_212,In_10);
nor U354 (N_354,In_684,In_508);
nand U355 (N_355,In_29,In_926);
nor U356 (N_356,In_474,In_278);
or U357 (N_357,In_110,In_794);
or U358 (N_358,In_559,In_556);
or U359 (N_359,In_61,In_1);
xor U360 (N_360,In_375,In_544);
nor U361 (N_361,In_591,In_625);
xor U362 (N_362,In_596,In_44);
nand U363 (N_363,In_818,In_932);
and U364 (N_364,In_920,In_928);
nand U365 (N_365,In_820,In_892);
or U366 (N_366,In_696,In_976);
nand U367 (N_367,In_310,In_829);
or U368 (N_368,In_884,In_21);
nor U369 (N_369,In_14,In_549);
or U370 (N_370,In_160,In_481);
xor U371 (N_371,In_173,In_709);
nor U372 (N_372,In_349,In_688);
or U373 (N_373,In_743,In_581);
nand U374 (N_374,In_119,In_114);
xor U375 (N_375,In_296,In_901);
or U376 (N_376,In_500,In_984);
and U377 (N_377,In_63,In_811);
xor U378 (N_378,In_183,In_560);
and U379 (N_379,In_869,In_847);
nand U380 (N_380,In_621,In_804);
nor U381 (N_381,In_657,In_169);
and U382 (N_382,In_732,In_953);
or U383 (N_383,In_658,In_439);
nor U384 (N_384,In_368,In_245);
and U385 (N_385,In_962,In_787);
nor U386 (N_386,In_564,In_207);
nor U387 (N_387,In_622,In_347);
and U388 (N_388,In_653,In_137);
nor U389 (N_389,In_747,In_968);
xnor U390 (N_390,In_912,In_972);
nor U391 (N_391,In_649,In_242);
and U392 (N_392,In_859,In_123);
nand U393 (N_393,In_277,In_774);
or U394 (N_394,In_778,In_934);
and U395 (N_395,In_456,In_651);
or U396 (N_396,In_866,In_420);
and U397 (N_397,In_493,In_977);
nor U398 (N_398,In_512,In_374);
nor U399 (N_399,In_906,In_308);
and U400 (N_400,In_446,In_803);
nor U401 (N_401,In_863,In_582);
nor U402 (N_402,In_789,In_800);
xor U403 (N_403,In_291,In_360);
and U404 (N_404,In_302,In_428);
nor U405 (N_405,In_50,In_867);
or U406 (N_406,In_378,In_25);
and U407 (N_407,In_938,In_262);
nor U408 (N_408,In_70,In_90);
nor U409 (N_409,In_597,In_281);
nor U410 (N_410,In_267,In_584);
nand U411 (N_411,In_22,In_399);
nor U412 (N_412,In_206,In_459);
and U413 (N_413,In_854,In_897);
or U414 (N_414,In_197,In_802);
nand U415 (N_415,In_152,In_875);
and U416 (N_416,In_134,In_282);
nand U417 (N_417,In_517,In_0);
and U418 (N_418,In_616,In_599);
or U419 (N_419,In_937,In_814);
nor U420 (N_420,In_144,In_471);
and U421 (N_421,In_359,In_185);
nor U422 (N_422,In_190,In_95);
xor U423 (N_423,In_283,In_737);
nor U424 (N_424,In_768,In_895);
nand U425 (N_425,In_628,In_268);
and U426 (N_426,In_874,In_815);
or U427 (N_427,In_573,In_639);
and U428 (N_428,In_745,In_437);
or U429 (N_429,In_164,In_16);
and U430 (N_430,In_878,In_384);
nor U431 (N_431,In_56,In_524);
nand U432 (N_432,In_910,In_974);
nand U433 (N_433,In_4,In_799);
and U434 (N_434,In_879,In_963);
and U435 (N_435,In_852,In_222);
xor U436 (N_436,In_411,In_764);
nor U437 (N_437,In_132,In_841);
and U438 (N_438,In_566,In_11);
xnor U439 (N_439,In_674,In_139);
or U440 (N_440,In_363,In_748);
and U441 (N_441,In_377,In_255);
nor U442 (N_442,In_306,In_924);
and U443 (N_443,In_387,In_871);
nand U444 (N_444,In_94,In_785);
nand U445 (N_445,In_198,In_956);
or U446 (N_446,In_813,In_263);
nand U447 (N_447,In_204,In_238);
or U448 (N_448,In_27,In_947);
and U449 (N_449,In_623,In_486);
xor U450 (N_450,In_993,In_443);
nand U451 (N_451,In_331,In_598);
nand U452 (N_452,In_767,In_153);
nor U453 (N_453,In_907,In_538);
xnor U454 (N_454,In_563,In_113);
nand U455 (N_455,In_236,In_809);
nor U456 (N_456,In_432,In_224);
or U457 (N_457,In_641,In_6);
nor U458 (N_458,In_705,In_632);
or U459 (N_459,In_202,In_565);
xnor U460 (N_460,In_130,In_162);
nand U461 (N_461,In_101,In_782);
and U462 (N_462,In_58,In_662);
and U463 (N_463,In_200,In_199);
or U464 (N_464,In_807,In_453);
xor U465 (N_465,In_886,In_629);
nand U466 (N_466,In_388,In_78);
or U467 (N_467,In_48,In_365);
or U468 (N_468,In_595,In_951);
nor U469 (N_469,In_451,In_366);
nor U470 (N_470,In_857,In_92);
nand U471 (N_471,In_31,In_668);
and U472 (N_472,In_445,In_143);
or U473 (N_473,In_9,In_881);
nand U474 (N_474,In_853,In_995);
and U475 (N_475,In_836,In_256);
nor U476 (N_476,In_372,In_272);
xor U477 (N_477,In_845,In_203);
or U478 (N_478,In_184,In_191);
or U479 (N_479,In_314,In_469);
or U480 (N_480,In_626,In_319);
nor U481 (N_481,In_637,In_526);
and U482 (N_482,In_636,In_174);
or U483 (N_483,In_220,In_286);
nand U484 (N_484,In_235,In_776);
and U485 (N_485,In_899,In_921);
or U486 (N_486,In_18,In_763);
and U487 (N_487,In_201,In_476);
or U488 (N_488,In_894,In_834);
nand U489 (N_489,In_990,In_540);
nor U490 (N_490,In_750,In_704);
nand U491 (N_491,In_792,In_38);
nor U492 (N_492,In_376,In_175);
xor U493 (N_493,In_647,In_350);
nor U494 (N_494,In_321,In_510);
and U495 (N_495,In_666,In_806);
or U496 (N_496,In_740,In_585);
and U497 (N_497,In_111,In_719);
nand U498 (N_498,In_904,In_136);
nor U499 (N_499,In_67,In_959);
or U500 (N_500,N_458,N_395);
nand U501 (N_501,N_238,N_472);
and U502 (N_502,N_175,N_144);
or U503 (N_503,N_283,N_66);
and U504 (N_504,N_61,N_162);
xnor U505 (N_505,N_236,N_269);
or U506 (N_506,N_439,N_332);
nor U507 (N_507,N_156,N_229);
xor U508 (N_508,N_306,N_99);
or U509 (N_509,N_113,N_145);
nor U510 (N_510,N_482,N_307);
nand U511 (N_511,N_267,N_53);
and U512 (N_512,N_25,N_250);
or U513 (N_513,N_52,N_379);
nor U514 (N_514,N_481,N_302);
or U515 (N_515,N_87,N_410);
xor U516 (N_516,N_319,N_153);
or U517 (N_517,N_290,N_494);
and U518 (N_518,N_178,N_261);
and U519 (N_519,N_445,N_488);
nand U520 (N_520,N_108,N_173);
xnor U521 (N_521,N_293,N_308);
nor U522 (N_522,N_164,N_100);
or U523 (N_523,N_352,N_259);
nand U524 (N_524,N_461,N_230);
and U525 (N_525,N_205,N_22);
nand U526 (N_526,N_30,N_318);
and U527 (N_527,N_96,N_313);
nand U528 (N_528,N_465,N_184);
xor U529 (N_529,N_412,N_105);
nor U530 (N_530,N_43,N_430);
nand U531 (N_531,N_92,N_137);
and U532 (N_532,N_69,N_389);
nand U533 (N_533,N_6,N_323);
nand U534 (N_534,N_322,N_51);
nor U535 (N_535,N_299,N_365);
nor U536 (N_536,N_377,N_115);
or U537 (N_537,N_274,N_271);
nor U538 (N_538,N_235,N_8);
or U539 (N_539,N_157,N_484);
nor U540 (N_540,N_139,N_218);
nor U541 (N_541,N_45,N_462);
xor U542 (N_542,N_194,N_232);
and U543 (N_543,N_106,N_351);
nand U544 (N_544,N_109,N_372);
xnor U545 (N_545,N_129,N_317);
and U546 (N_546,N_95,N_163);
or U547 (N_547,N_493,N_166);
or U548 (N_548,N_496,N_403);
nor U549 (N_549,N_33,N_368);
or U550 (N_550,N_260,N_247);
nand U551 (N_551,N_233,N_471);
nor U552 (N_552,N_442,N_191);
and U553 (N_553,N_470,N_91);
or U554 (N_554,N_441,N_126);
nand U555 (N_555,N_32,N_466);
or U556 (N_556,N_492,N_304);
or U557 (N_557,N_35,N_281);
nor U558 (N_558,N_160,N_56);
nor U559 (N_559,N_231,N_480);
nand U560 (N_560,N_397,N_330);
nor U561 (N_561,N_84,N_57);
or U562 (N_562,N_150,N_219);
or U563 (N_563,N_415,N_331);
and U564 (N_564,N_263,N_252);
and U565 (N_565,N_190,N_158);
and U566 (N_566,N_15,N_82);
and U567 (N_567,N_434,N_420);
nor U568 (N_568,N_272,N_49);
nand U569 (N_569,N_414,N_54);
xnor U570 (N_570,N_183,N_343);
nor U571 (N_571,N_483,N_294);
and U572 (N_572,N_94,N_3);
or U573 (N_573,N_459,N_79);
nor U574 (N_574,N_417,N_380);
nand U575 (N_575,N_86,N_453);
nand U576 (N_576,N_476,N_170);
nand U577 (N_577,N_149,N_19);
nor U578 (N_578,N_348,N_279);
nand U579 (N_579,N_103,N_98);
nand U580 (N_580,N_288,N_136);
nand U581 (N_581,N_432,N_207);
and U582 (N_582,N_310,N_320);
nor U583 (N_583,N_206,N_76);
nor U584 (N_584,N_489,N_63);
or U585 (N_585,N_311,N_371);
nand U586 (N_586,N_112,N_258);
nor U587 (N_587,N_449,N_309);
and U588 (N_588,N_133,N_303);
and U589 (N_589,N_182,N_291);
or U590 (N_590,N_196,N_242);
nand U591 (N_591,N_44,N_192);
xnor U592 (N_592,N_188,N_64);
and U593 (N_593,N_295,N_48);
xor U594 (N_594,N_354,N_347);
nor U595 (N_595,N_77,N_336);
nor U596 (N_596,N_431,N_401);
or U597 (N_597,N_287,N_324);
and U598 (N_598,N_436,N_181);
or U599 (N_599,N_81,N_240);
xnor U600 (N_600,N_71,N_18);
or U601 (N_601,N_333,N_68);
xnor U602 (N_602,N_358,N_60);
or U603 (N_603,N_378,N_262);
and U604 (N_604,N_425,N_382);
nand U605 (N_605,N_142,N_475);
nand U606 (N_606,N_407,N_346);
xor U607 (N_607,N_135,N_411);
or U608 (N_608,N_152,N_400);
nor U609 (N_609,N_366,N_315);
nor U610 (N_610,N_121,N_67);
nand U611 (N_611,N_120,N_486);
and U612 (N_612,N_58,N_289);
nand U613 (N_613,N_131,N_355);
and U614 (N_614,N_189,N_419);
or U615 (N_615,N_344,N_93);
nand U616 (N_616,N_208,N_424);
or U617 (N_617,N_360,N_85);
and U618 (N_618,N_443,N_187);
and U619 (N_619,N_448,N_423);
and U620 (N_620,N_186,N_416);
nor U621 (N_621,N_123,N_7);
nor U622 (N_622,N_463,N_88);
or U623 (N_623,N_59,N_50);
and U624 (N_624,N_89,N_171);
or U625 (N_625,N_199,N_14);
nor U626 (N_626,N_101,N_128);
or U627 (N_627,N_327,N_270);
and U628 (N_628,N_177,N_473);
or U629 (N_629,N_364,N_405);
xnor U630 (N_630,N_334,N_427);
xor U631 (N_631,N_214,N_321);
nor U632 (N_632,N_143,N_107);
and U633 (N_633,N_110,N_337);
or U634 (N_634,N_141,N_256);
nand U635 (N_635,N_363,N_174);
nand U636 (N_636,N_339,N_396);
or U637 (N_637,N_350,N_159);
nor U638 (N_638,N_345,N_385);
and U639 (N_639,N_83,N_198);
and U640 (N_640,N_392,N_176);
or U641 (N_641,N_210,N_435);
and U642 (N_642,N_454,N_217);
xor U643 (N_643,N_329,N_42);
or U644 (N_644,N_125,N_316);
nor U645 (N_645,N_387,N_241);
nor U646 (N_646,N_147,N_296);
nor U647 (N_647,N_362,N_179);
nor U648 (N_648,N_478,N_468);
nand U649 (N_649,N_220,N_114);
or U650 (N_650,N_65,N_234);
nand U651 (N_651,N_124,N_104);
nand U652 (N_652,N_276,N_464);
and U653 (N_653,N_383,N_16);
nand U654 (N_654,N_97,N_278);
xor U655 (N_655,N_226,N_237);
or U656 (N_656,N_469,N_495);
xor U657 (N_657,N_390,N_228);
and U658 (N_658,N_292,N_402);
nor U659 (N_659,N_499,N_282);
nand U660 (N_660,N_404,N_211);
and U661 (N_661,N_4,N_491);
and U662 (N_662,N_391,N_168);
and U663 (N_663,N_13,N_127);
xor U664 (N_664,N_409,N_254);
nand U665 (N_665,N_202,N_398);
nor U666 (N_666,N_451,N_2);
nand U667 (N_667,N_455,N_422);
nor U668 (N_668,N_349,N_312);
or U669 (N_669,N_46,N_41);
nand U670 (N_670,N_340,N_298);
nand U671 (N_671,N_119,N_10);
and U672 (N_672,N_386,N_172);
xnor U673 (N_673,N_452,N_399);
and U674 (N_674,N_75,N_193);
nor U675 (N_675,N_264,N_356);
nand U676 (N_676,N_457,N_221);
nand U677 (N_677,N_155,N_17);
and U678 (N_678,N_72,N_34);
and U679 (N_679,N_116,N_255);
nor U680 (N_680,N_151,N_134);
xnor U681 (N_681,N_169,N_253);
or U682 (N_682,N_243,N_456);
nand U683 (N_683,N_90,N_200);
and U684 (N_684,N_239,N_227);
or U685 (N_685,N_165,N_146);
and U686 (N_686,N_111,N_338);
nor U687 (N_687,N_209,N_428);
and U688 (N_688,N_273,N_224);
or U689 (N_689,N_195,N_213);
nor U690 (N_690,N_370,N_359);
and U691 (N_691,N_197,N_353);
nand U692 (N_692,N_29,N_225);
or U693 (N_693,N_118,N_0);
nand U694 (N_694,N_490,N_249);
and U695 (N_695,N_180,N_265);
and U696 (N_696,N_479,N_438);
nand U697 (N_697,N_117,N_440);
nor U698 (N_698,N_450,N_437);
or U699 (N_699,N_5,N_216);
xor U700 (N_700,N_497,N_55);
xor U701 (N_701,N_381,N_23);
nor U702 (N_702,N_426,N_122);
or U703 (N_703,N_148,N_314);
nor U704 (N_704,N_342,N_284);
nor U705 (N_705,N_375,N_393);
nor U706 (N_706,N_203,N_361);
nand U707 (N_707,N_498,N_305);
nand U708 (N_708,N_80,N_12);
and U709 (N_709,N_413,N_40);
and U710 (N_710,N_467,N_27);
or U711 (N_711,N_37,N_376);
xnor U712 (N_712,N_28,N_300);
and U713 (N_713,N_477,N_408);
and U714 (N_714,N_102,N_47);
or U715 (N_715,N_1,N_132);
or U716 (N_716,N_447,N_21);
or U717 (N_717,N_373,N_31);
nor U718 (N_718,N_268,N_36);
nand U719 (N_719,N_301,N_277);
nor U720 (N_720,N_245,N_11);
nand U721 (N_721,N_9,N_201);
or U722 (N_722,N_154,N_248);
nand U723 (N_723,N_62,N_39);
nor U724 (N_724,N_328,N_266);
nor U725 (N_725,N_223,N_326);
nor U726 (N_726,N_429,N_275);
and U727 (N_727,N_130,N_257);
or U728 (N_728,N_444,N_487);
nor U729 (N_729,N_369,N_285);
or U730 (N_730,N_138,N_244);
or U731 (N_731,N_161,N_140);
nand U732 (N_732,N_185,N_251);
or U733 (N_733,N_24,N_78);
nand U734 (N_734,N_418,N_70);
and U735 (N_735,N_394,N_286);
or U736 (N_736,N_222,N_204);
or U737 (N_737,N_384,N_421);
or U738 (N_738,N_446,N_406);
nor U739 (N_739,N_212,N_167);
xor U740 (N_740,N_341,N_246);
and U741 (N_741,N_73,N_474);
nor U742 (N_742,N_20,N_38);
or U743 (N_743,N_485,N_460);
or U744 (N_744,N_433,N_357);
or U745 (N_745,N_297,N_388);
and U746 (N_746,N_74,N_325);
or U747 (N_747,N_374,N_215);
or U748 (N_748,N_367,N_26);
and U749 (N_749,N_280,N_335);
and U750 (N_750,N_416,N_470);
nor U751 (N_751,N_472,N_411);
nor U752 (N_752,N_105,N_423);
nand U753 (N_753,N_137,N_367);
and U754 (N_754,N_4,N_100);
or U755 (N_755,N_17,N_29);
nor U756 (N_756,N_34,N_168);
and U757 (N_757,N_358,N_209);
or U758 (N_758,N_196,N_319);
nor U759 (N_759,N_306,N_182);
or U760 (N_760,N_296,N_417);
or U761 (N_761,N_91,N_408);
or U762 (N_762,N_371,N_174);
or U763 (N_763,N_207,N_451);
or U764 (N_764,N_300,N_382);
or U765 (N_765,N_336,N_126);
nand U766 (N_766,N_446,N_261);
nor U767 (N_767,N_491,N_197);
or U768 (N_768,N_139,N_350);
nand U769 (N_769,N_155,N_300);
nor U770 (N_770,N_357,N_160);
and U771 (N_771,N_459,N_51);
and U772 (N_772,N_337,N_328);
and U773 (N_773,N_228,N_423);
nor U774 (N_774,N_308,N_244);
xnor U775 (N_775,N_204,N_376);
or U776 (N_776,N_129,N_38);
xnor U777 (N_777,N_67,N_311);
nand U778 (N_778,N_252,N_385);
or U779 (N_779,N_496,N_463);
nand U780 (N_780,N_484,N_126);
or U781 (N_781,N_117,N_244);
and U782 (N_782,N_223,N_152);
xor U783 (N_783,N_357,N_241);
and U784 (N_784,N_339,N_63);
or U785 (N_785,N_292,N_35);
or U786 (N_786,N_399,N_320);
and U787 (N_787,N_488,N_3);
nor U788 (N_788,N_234,N_103);
nand U789 (N_789,N_394,N_111);
nor U790 (N_790,N_45,N_458);
and U791 (N_791,N_446,N_214);
or U792 (N_792,N_48,N_65);
nand U793 (N_793,N_13,N_67);
nand U794 (N_794,N_22,N_377);
nand U795 (N_795,N_298,N_176);
or U796 (N_796,N_144,N_304);
nor U797 (N_797,N_295,N_122);
and U798 (N_798,N_173,N_10);
or U799 (N_799,N_207,N_365);
nor U800 (N_800,N_448,N_466);
nor U801 (N_801,N_226,N_366);
nand U802 (N_802,N_104,N_105);
xnor U803 (N_803,N_69,N_482);
xor U804 (N_804,N_310,N_330);
or U805 (N_805,N_427,N_142);
or U806 (N_806,N_80,N_174);
and U807 (N_807,N_379,N_383);
or U808 (N_808,N_412,N_407);
nor U809 (N_809,N_131,N_73);
and U810 (N_810,N_4,N_25);
nand U811 (N_811,N_489,N_189);
or U812 (N_812,N_476,N_30);
or U813 (N_813,N_362,N_148);
and U814 (N_814,N_455,N_4);
nand U815 (N_815,N_222,N_156);
or U816 (N_816,N_199,N_370);
nor U817 (N_817,N_484,N_491);
and U818 (N_818,N_156,N_430);
nor U819 (N_819,N_353,N_266);
or U820 (N_820,N_247,N_431);
nand U821 (N_821,N_316,N_379);
nor U822 (N_822,N_270,N_467);
nand U823 (N_823,N_11,N_411);
nor U824 (N_824,N_183,N_421);
and U825 (N_825,N_5,N_49);
nor U826 (N_826,N_305,N_495);
and U827 (N_827,N_276,N_126);
or U828 (N_828,N_496,N_392);
nand U829 (N_829,N_105,N_444);
xor U830 (N_830,N_168,N_259);
and U831 (N_831,N_445,N_267);
nand U832 (N_832,N_21,N_177);
nand U833 (N_833,N_136,N_15);
or U834 (N_834,N_491,N_201);
nor U835 (N_835,N_0,N_203);
or U836 (N_836,N_266,N_84);
xor U837 (N_837,N_160,N_364);
and U838 (N_838,N_281,N_148);
xor U839 (N_839,N_175,N_277);
nand U840 (N_840,N_295,N_455);
or U841 (N_841,N_147,N_384);
and U842 (N_842,N_95,N_19);
nor U843 (N_843,N_419,N_227);
nor U844 (N_844,N_27,N_346);
and U845 (N_845,N_60,N_442);
xnor U846 (N_846,N_370,N_124);
or U847 (N_847,N_6,N_15);
xnor U848 (N_848,N_318,N_445);
nor U849 (N_849,N_344,N_112);
xor U850 (N_850,N_332,N_33);
and U851 (N_851,N_221,N_97);
nor U852 (N_852,N_280,N_162);
nand U853 (N_853,N_407,N_67);
nand U854 (N_854,N_250,N_479);
nand U855 (N_855,N_263,N_333);
nor U856 (N_856,N_345,N_21);
xor U857 (N_857,N_475,N_137);
nand U858 (N_858,N_374,N_267);
nand U859 (N_859,N_290,N_492);
or U860 (N_860,N_347,N_108);
and U861 (N_861,N_282,N_378);
nand U862 (N_862,N_72,N_158);
xnor U863 (N_863,N_25,N_5);
nand U864 (N_864,N_386,N_459);
nor U865 (N_865,N_457,N_107);
nand U866 (N_866,N_259,N_30);
nand U867 (N_867,N_177,N_402);
nand U868 (N_868,N_63,N_62);
nand U869 (N_869,N_366,N_456);
nor U870 (N_870,N_293,N_228);
and U871 (N_871,N_155,N_414);
nor U872 (N_872,N_181,N_162);
or U873 (N_873,N_220,N_128);
nor U874 (N_874,N_312,N_124);
nor U875 (N_875,N_195,N_435);
nor U876 (N_876,N_372,N_406);
or U877 (N_877,N_114,N_102);
or U878 (N_878,N_295,N_21);
or U879 (N_879,N_331,N_216);
nand U880 (N_880,N_199,N_245);
xnor U881 (N_881,N_380,N_424);
nor U882 (N_882,N_65,N_290);
or U883 (N_883,N_142,N_74);
or U884 (N_884,N_375,N_105);
and U885 (N_885,N_430,N_399);
nand U886 (N_886,N_96,N_397);
nor U887 (N_887,N_431,N_112);
or U888 (N_888,N_257,N_412);
or U889 (N_889,N_446,N_76);
nor U890 (N_890,N_63,N_497);
nand U891 (N_891,N_97,N_198);
and U892 (N_892,N_470,N_148);
and U893 (N_893,N_97,N_414);
and U894 (N_894,N_226,N_236);
or U895 (N_895,N_222,N_445);
nor U896 (N_896,N_48,N_381);
nor U897 (N_897,N_418,N_365);
nor U898 (N_898,N_298,N_170);
nor U899 (N_899,N_312,N_114);
or U900 (N_900,N_240,N_42);
xor U901 (N_901,N_493,N_193);
or U902 (N_902,N_449,N_96);
xor U903 (N_903,N_490,N_269);
or U904 (N_904,N_297,N_280);
nand U905 (N_905,N_489,N_303);
xor U906 (N_906,N_29,N_129);
xor U907 (N_907,N_108,N_367);
and U908 (N_908,N_301,N_457);
or U909 (N_909,N_155,N_338);
xor U910 (N_910,N_493,N_96);
nand U911 (N_911,N_116,N_382);
nor U912 (N_912,N_352,N_331);
nand U913 (N_913,N_249,N_94);
nor U914 (N_914,N_369,N_243);
nor U915 (N_915,N_259,N_214);
and U916 (N_916,N_146,N_293);
or U917 (N_917,N_263,N_183);
xor U918 (N_918,N_94,N_369);
nor U919 (N_919,N_31,N_338);
nand U920 (N_920,N_417,N_161);
or U921 (N_921,N_235,N_170);
xor U922 (N_922,N_62,N_470);
xor U923 (N_923,N_141,N_251);
or U924 (N_924,N_413,N_220);
nor U925 (N_925,N_335,N_454);
nand U926 (N_926,N_38,N_246);
nand U927 (N_927,N_382,N_478);
and U928 (N_928,N_372,N_260);
and U929 (N_929,N_428,N_404);
and U930 (N_930,N_376,N_197);
and U931 (N_931,N_39,N_408);
and U932 (N_932,N_17,N_408);
nor U933 (N_933,N_284,N_53);
and U934 (N_934,N_8,N_269);
nand U935 (N_935,N_425,N_328);
nor U936 (N_936,N_329,N_49);
and U937 (N_937,N_134,N_43);
nor U938 (N_938,N_163,N_108);
and U939 (N_939,N_477,N_364);
nand U940 (N_940,N_285,N_310);
nand U941 (N_941,N_388,N_237);
xnor U942 (N_942,N_12,N_265);
and U943 (N_943,N_166,N_473);
nand U944 (N_944,N_432,N_190);
nand U945 (N_945,N_134,N_89);
or U946 (N_946,N_417,N_60);
xor U947 (N_947,N_191,N_163);
nand U948 (N_948,N_91,N_64);
and U949 (N_949,N_8,N_478);
and U950 (N_950,N_407,N_267);
nor U951 (N_951,N_87,N_324);
and U952 (N_952,N_452,N_24);
or U953 (N_953,N_319,N_358);
nor U954 (N_954,N_365,N_192);
xnor U955 (N_955,N_408,N_396);
and U956 (N_956,N_206,N_323);
nand U957 (N_957,N_68,N_310);
nand U958 (N_958,N_339,N_105);
xor U959 (N_959,N_358,N_85);
xnor U960 (N_960,N_470,N_249);
or U961 (N_961,N_192,N_382);
and U962 (N_962,N_73,N_6);
nand U963 (N_963,N_447,N_342);
nor U964 (N_964,N_438,N_204);
nor U965 (N_965,N_92,N_143);
or U966 (N_966,N_390,N_80);
and U967 (N_967,N_416,N_426);
xor U968 (N_968,N_249,N_428);
or U969 (N_969,N_179,N_496);
or U970 (N_970,N_271,N_395);
and U971 (N_971,N_188,N_330);
xor U972 (N_972,N_236,N_461);
nand U973 (N_973,N_47,N_457);
or U974 (N_974,N_348,N_445);
xnor U975 (N_975,N_365,N_476);
and U976 (N_976,N_402,N_469);
nand U977 (N_977,N_192,N_255);
or U978 (N_978,N_467,N_247);
and U979 (N_979,N_471,N_77);
nand U980 (N_980,N_228,N_458);
nand U981 (N_981,N_17,N_136);
or U982 (N_982,N_489,N_262);
nor U983 (N_983,N_27,N_119);
xnor U984 (N_984,N_231,N_331);
nor U985 (N_985,N_170,N_276);
xor U986 (N_986,N_264,N_253);
and U987 (N_987,N_352,N_306);
nor U988 (N_988,N_156,N_490);
and U989 (N_989,N_441,N_250);
nor U990 (N_990,N_14,N_455);
or U991 (N_991,N_290,N_120);
or U992 (N_992,N_197,N_388);
or U993 (N_993,N_25,N_305);
nand U994 (N_994,N_348,N_24);
nor U995 (N_995,N_275,N_124);
nand U996 (N_996,N_208,N_255);
nand U997 (N_997,N_37,N_271);
nor U998 (N_998,N_11,N_428);
nor U999 (N_999,N_343,N_275);
nor U1000 (N_1000,N_698,N_717);
and U1001 (N_1001,N_814,N_898);
or U1002 (N_1002,N_637,N_792);
nand U1003 (N_1003,N_530,N_825);
and U1004 (N_1004,N_708,N_782);
nand U1005 (N_1005,N_917,N_905);
nor U1006 (N_1006,N_998,N_646);
nand U1007 (N_1007,N_872,N_846);
and U1008 (N_1008,N_980,N_714);
nor U1009 (N_1009,N_855,N_536);
nor U1010 (N_1010,N_906,N_934);
and U1011 (N_1011,N_654,N_693);
or U1012 (N_1012,N_716,N_658);
and U1013 (N_1013,N_868,N_900);
xor U1014 (N_1014,N_890,N_884);
nand U1015 (N_1015,N_971,N_920);
nor U1016 (N_1016,N_700,N_542);
and U1017 (N_1017,N_728,N_889);
nand U1018 (N_1018,N_957,N_937);
nand U1019 (N_1019,N_922,N_573);
and U1020 (N_1020,N_778,N_696);
nor U1021 (N_1021,N_932,N_781);
and U1022 (N_1022,N_999,N_552);
nor U1023 (N_1023,N_647,N_771);
or U1024 (N_1024,N_861,N_968);
or U1025 (N_1025,N_801,N_925);
xnor U1026 (N_1026,N_657,N_697);
and U1027 (N_1027,N_732,N_711);
or U1028 (N_1028,N_503,N_736);
or U1029 (N_1029,N_683,N_733);
or U1030 (N_1030,N_887,N_507);
nor U1031 (N_1031,N_961,N_543);
nand U1032 (N_1032,N_946,N_881);
nor U1033 (N_1033,N_726,N_505);
nor U1034 (N_1034,N_833,N_895);
and U1035 (N_1035,N_611,N_854);
or U1036 (N_1036,N_523,N_525);
and U1037 (N_1037,N_877,N_715);
or U1038 (N_1038,N_620,N_858);
or U1039 (N_1039,N_982,N_883);
nor U1040 (N_1040,N_915,N_516);
and U1041 (N_1041,N_882,N_607);
or U1042 (N_1042,N_967,N_737);
or U1043 (N_1043,N_864,N_991);
and U1044 (N_1044,N_772,N_554);
nand U1045 (N_1045,N_688,N_706);
nand U1046 (N_1046,N_558,N_763);
nand U1047 (N_1047,N_633,N_798);
nand U1048 (N_1048,N_911,N_591);
and U1049 (N_1049,N_839,N_666);
nor U1050 (N_1050,N_867,N_750);
nor U1051 (N_1051,N_533,N_759);
xor U1052 (N_1052,N_643,N_694);
nand U1053 (N_1053,N_945,N_606);
and U1054 (N_1054,N_602,N_913);
and U1055 (N_1055,N_594,N_539);
nor U1056 (N_1056,N_595,N_585);
nor U1057 (N_1057,N_838,N_894);
and U1058 (N_1058,N_546,N_995);
or U1059 (N_1059,N_599,N_757);
or U1060 (N_1060,N_849,N_756);
nand U1061 (N_1061,N_878,N_586);
or U1062 (N_1062,N_691,N_788);
nor U1063 (N_1063,N_689,N_972);
xnor U1064 (N_1064,N_789,N_670);
nand U1065 (N_1065,N_580,N_935);
and U1066 (N_1066,N_876,N_812);
or U1067 (N_1067,N_804,N_893);
nand U1068 (N_1068,N_619,N_818);
and U1069 (N_1069,N_744,N_648);
or U1070 (N_1070,N_928,N_745);
nand U1071 (N_1071,N_988,N_909);
nand U1072 (N_1072,N_635,N_755);
xor U1073 (N_1073,N_966,N_835);
or U1074 (N_1074,N_952,N_681);
nand U1075 (N_1075,N_764,N_799);
nand U1076 (N_1076,N_582,N_743);
and U1077 (N_1077,N_983,N_532);
nor U1078 (N_1078,N_871,N_767);
and U1079 (N_1079,N_807,N_931);
nand U1080 (N_1080,N_664,N_929);
xor U1081 (N_1081,N_748,N_687);
and U1082 (N_1082,N_830,N_981);
xor U1083 (N_1083,N_653,N_685);
or U1084 (N_1084,N_762,N_615);
xnor U1085 (N_1085,N_550,N_941);
nor U1086 (N_1086,N_553,N_556);
and U1087 (N_1087,N_891,N_568);
or U1088 (N_1088,N_590,N_600);
nand U1089 (N_1089,N_531,N_985);
nand U1090 (N_1090,N_528,N_730);
nand U1091 (N_1091,N_690,N_583);
or U1092 (N_1092,N_522,N_650);
and U1093 (N_1093,N_823,N_832);
nor U1094 (N_1094,N_754,N_672);
nor U1095 (N_1095,N_951,N_848);
xnor U1096 (N_1096,N_721,N_742);
nor U1097 (N_1097,N_963,N_626);
and U1098 (N_1098,N_660,N_910);
nor U1099 (N_1099,N_773,N_571);
nand U1100 (N_1100,N_955,N_628);
and U1101 (N_1101,N_785,N_609);
and U1102 (N_1102,N_776,N_962);
nor U1103 (N_1103,N_822,N_912);
nand U1104 (N_1104,N_797,N_500);
nor U1105 (N_1105,N_819,N_720);
and U1106 (N_1106,N_779,N_636);
and U1107 (N_1107,N_766,N_671);
nand U1108 (N_1108,N_598,N_749);
nor U1109 (N_1109,N_984,N_914);
xor U1110 (N_1110,N_897,N_551);
nor U1111 (N_1111,N_559,N_975);
nand U1112 (N_1112,N_712,N_622);
or U1113 (N_1113,N_735,N_701);
or U1114 (N_1114,N_753,N_526);
nand U1115 (N_1115,N_751,N_997);
nand U1116 (N_1116,N_682,N_747);
or U1117 (N_1117,N_645,N_659);
and U1118 (N_1118,N_509,N_677);
xor U1119 (N_1119,N_589,N_875);
and U1120 (N_1120,N_727,N_758);
or U1121 (N_1121,N_515,N_723);
or U1122 (N_1122,N_692,N_888);
nand U1123 (N_1123,N_641,N_565);
nor U1124 (N_1124,N_857,N_806);
nor U1125 (N_1125,N_899,N_713);
xor U1126 (N_1126,N_593,N_977);
or U1127 (N_1127,N_567,N_936);
xor U1128 (N_1128,N_793,N_725);
and U1129 (N_1129,N_517,N_502);
and U1130 (N_1130,N_555,N_731);
xor U1131 (N_1131,N_684,N_673);
and U1132 (N_1132,N_902,N_805);
xor U1133 (N_1133,N_661,N_824);
nand U1134 (N_1134,N_640,N_790);
nand U1135 (N_1135,N_649,N_579);
nand U1136 (N_1136,N_993,N_739);
nand U1137 (N_1137,N_561,N_613);
or U1138 (N_1138,N_724,N_841);
nor U1139 (N_1139,N_614,N_852);
and U1140 (N_1140,N_588,N_575);
or U1141 (N_1141,N_919,N_821);
and U1142 (N_1142,N_879,N_809);
and U1143 (N_1143,N_632,N_547);
nand U1144 (N_1144,N_978,N_520);
or U1145 (N_1145,N_534,N_663);
xor U1146 (N_1146,N_752,N_581);
or U1147 (N_1147,N_501,N_512);
nand U1148 (N_1148,N_513,N_540);
nand U1149 (N_1149,N_638,N_662);
or U1150 (N_1150,N_942,N_803);
and U1151 (N_1151,N_959,N_786);
nand U1152 (N_1152,N_836,N_976);
nand U1153 (N_1153,N_578,N_992);
or U1154 (N_1154,N_885,N_856);
nand U1155 (N_1155,N_570,N_777);
or U1156 (N_1156,N_973,N_722);
nand U1157 (N_1157,N_535,N_618);
and U1158 (N_1158,N_979,N_873);
nor U1159 (N_1159,N_802,N_826);
and U1160 (N_1160,N_970,N_617);
nand U1161 (N_1161,N_947,N_990);
and U1162 (N_1162,N_655,N_907);
or U1163 (N_1163,N_859,N_544);
nand U1164 (N_1164,N_880,N_705);
and U1165 (N_1165,N_511,N_770);
or U1166 (N_1166,N_800,N_903);
or U1167 (N_1167,N_939,N_860);
nand U1168 (N_1168,N_704,N_923);
xor U1169 (N_1169,N_538,N_796);
nor U1170 (N_1170,N_908,N_729);
and U1171 (N_1171,N_949,N_597);
nor U1172 (N_1172,N_557,N_549);
nand U1173 (N_1173,N_791,N_930);
xor U1174 (N_1174,N_631,N_676);
nor U1175 (N_1175,N_510,N_639);
nand U1176 (N_1176,N_996,N_624);
nor U1177 (N_1177,N_869,N_740);
and U1178 (N_1178,N_844,N_831);
and U1179 (N_1179,N_629,N_506);
and U1180 (N_1180,N_940,N_545);
xor U1181 (N_1181,N_760,N_668);
and U1182 (N_1182,N_675,N_795);
or U1183 (N_1183,N_933,N_562);
nor U1184 (N_1184,N_518,N_870);
and U1185 (N_1185,N_850,N_783);
and U1186 (N_1186,N_974,N_563);
or U1187 (N_1187,N_572,N_954);
and U1188 (N_1188,N_642,N_828);
and U1189 (N_1189,N_519,N_808);
nor U1190 (N_1190,N_769,N_987);
xor U1191 (N_1191,N_938,N_667);
and U1192 (N_1192,N_634,N_956);
and U1193 (N_1193,N_574,N_950);
nor U1194 (N_1194,N_699,N_719);
or U1195 (N_1195,N_810,N_576);
nand U1196 (N_1196,N_953,N_521);
and U1197 (N_1197,N_840,N_741);
nor U1198 (N_1198,N_596,N_508);
or U1199 (N_1199,N_612,N_794);
and U1200 (N_1200,N_948,N_710);
and U1201 (N_1201,N_811,N_765);
xor U1202 (N_1202,N_866,N_843);
or U1203 (N_1203,N_603,N_817);
or U1204 (N_1204,N_829,N_665);
nor U1205 (N_1205,N_592,N_761);
nor U1206 (N_1206,N_921,N_842);
nor U1207 (N_1207,N_605,N_504);
nor U1208 (N_1208,N_738,N_560);
nor U1209 (N_1209,N_827,N_678);
nor U1210 (N_1210,N_916,N_627);
or U1211 (N_1211,N_703,N_610);
and U1212 (N_1212,N_564,N_541);
nand U1213 (N_1213,N_865,N_718);
and U1214 (N_1214,N_958,N_679);
nand U1215 (N_1215,N_680,N_768);
and U1216 (N_1216,N_625,N_892);
nor U1217 (N_1217,N_815,N_816);
and U1218 (N_1218,N_537,N_604);
and U1219 (N_1219,N_548,N_695);
or U1220 (N_1220,N_652,N_847);
or U1221 (N_1221,N_514,N_960);
xnor U1222 (N_1222,N_845,N_964);
nor U1223 (N_1223,N_837,N_621);
nor U1224 (N_1224,N_709,N_584);
nor U1225 (N_1225,N_608,N_623);
nand U1226 (N_1226,N_834,N_896);
nand U1227 (N_1227,N_886,N_820);
xor U1228 (N_1228,N_702,N_986);
nor U1229 (N_1229,N_863,N_904);
nor U1230 (N_1230,N_569,N_924);
or U1231 (N_1231,N_577,N_813);
or U1232 (N_1232,N_529,N_601);
and U1233 (N_1233,N_874,N_616);
nand U1234 (N_1234,N_965,N_784);
nor U1235 (N_1235,N_994,N_674);
nor U1236 (N_1236,N_587,N_524);
or U1237 (N_1237,N_775,N_644);
xor U1238 (N_1238,N_774,N_918);
or U1239 (N_1239,N_734,N_707);
nor U1240 (N_1240,N_656,N_901);
nand U1241 (N_1241,N_787,N_780);
xor U1242 (N_1242,N_989,N_969);
and U1243 (N_1243,N_862,N_851);
nand U1244 (N_1244,N_566,N_527);
nand U1245 (N_1245,N_944,N_746);
xor U1246 (N_1246,N_686,N_927);
nor U1247 (N_1247,N_853,N_943);
nand U1248 (N_1248,N_630,N_926);
nor U1249 (N_1249,N_669,N_651);
nand U1250 (N_1250,N_694,N_989);
xor U1251 (N_1251,N_860,N_780);
or U1252 (N_1252,N_718,N_879);
or U1253 (N_1253,N_841,N_877);
nor U1254 (N_1254,N_763,N_835);
nand U1255 (N_1255,N_569,N_540);
and U1256 (N_1256,N_727,N_941);
nor U1257 (N_1257,N_572,N_859);
and U1258 (N_1258,N_612,N_881);
or U1259 (N_1259,N_976,N_818);
and U1260 (N_1260,N_899,N_522);
or U1261 (N_1261,N_612,N_622);
and U1262 (N_1262,N_549,N_530);
or U1263 (N_1263,N_582,N_919);
and U1264 (N_1264,N_504,N_925);
and U1265 (N_1265,N_535,N_842);
nor U1266 (N_1266,N_838,N_833);
nor U1267 (N_1267,N_734,N_885);
nor U1268 (N_1268,N_883,N_544);
xnor U1269 (N_1269,N_530,N_771);
or U1270 (N_1270,N_833,N_535);
or U1271 (N_1271,N_812,N_946);
and U1272 (N_1272,N_537,N_588);
nor U1273 (N_1273,N_598,N_704);
xor U1274 (N_1274,N_623,N_812);
nand U1275 (N_1275,N_717,N_761);
or U1276 (N_1276,N_865,N_713);
nand U1277 (N_1277,N_591,N_954);
or U1278 (N_1278,N_608,N_956);
nor U1279 (N_1279,N_846,N_674);
nand U1280 (N_1280,N_686,N_595);
or U1281 (N_1281,N_719,N_985);
and U1282 (N_1282,N_513,N_877);
nand U1283 (N_1283,N_781,N_616);
nor U1284 (N_1284,N_671,N_721);
nor U1285 (N_1285,N_687,N_549);
or U1286 (N_1286,N_762,N_581);
xnor U1287 (N_1287,N_799,N_756);
nand U1288 (N_1288,N_658,N_757);
and U1289 (N_1289,N_548,N_812);
nor U1290 (N_1290,N_760,N_501);
or U1291 (N_1291,N_618,N_722);
or U1292 (N_1292,N_979,N_770);
and U1293 (N_1293,N_728,N_670);
nor U1294 (N_1294,N_963,N_960);
nor U1295 (N_1295,N_520,N_885);
or U1296 (N_1296,N_710,N_680);
nor U1297 (N_1297,N_691,N_693);
nand U1298 (N_1298,N_846,N_615);
nor U1299 (N_1299,N_600,N_649);
or U1300 (N_1300,N_608,N_803);
nand U1301 (N_1301,N_546,N_704);
xnor U1302 (N_1302,N_835,N_944);
or U1303 (N_1303,N_717,N_720);
xnor U1304 (N_1304,N_695,N_704);
and U1305 (N_1305,N_629,N_790);
and U1306 (N_1306,N_905,N_649);
and U1307 (N_1307,N_686,N_987);
nand U1308 (N_1308,N_524,N_744);
or U1309 (N_1309,N_917,N_733);
nand U1310 (N_1310,N_840,N_813);
xor U1311 (N_1311,N_625,N_739);
nand U1312 (N_1312,N_852,N_577);
nor U1313 (N_1313,N_565,N_804);
and U1314 (N_1314,N_530,N_653);
xor U1315 (N_1315,N_938,N_597);
or U1316 (N_1316,N_878,N_635);
or U1317 (N_1317,N_772,N_719);
nand U1318 (N_1318,N_591,N_518);
or U1319 (N_1319,N_971,N_600);
nor U1320 (N_1320,N_792,N_737);
and U1321 (N_1321,N_804,N_903);
or U1322 (N_1322,N_932,N_764);
xnor U1323 (N_1323,N_850,N_834);
or U1324 (N_1324,N_975,N_596);
nand U1325 (N_1325,N_519,N_993);
and U1326 (N_1326,N_913,N_740);
or U1327 (N_1327,N_925,N_776);
or U1328 (N_1328,N_616,N_676);
or U1329 (N_1329,N_798,N_782);
nor U1330 (N_1330,N_575,N_580);
nand U1331 (N_1331,N_756,N_603);
or U1332 (N_1332,N_553,N_712);
nand U1333 (N_1333,N_861,N_504);
and U1334 (N_1334,N_560,N_732);
nor U1335 (N_1335,N_646,N_521);
or U1336 (N_1336,N_989,N_635);
or U1337 (N_1337,N_579,N_813);
or U1338 (N_1338,N_660,N_964);
and U1339 (N_1339,N_760,N_997);
or U1340 (N_1340,N_917,N_919);
nor U1341 (N_1341,N_624,N_768);
nor U1342 (N_1342,N_790,N_523);
and U1343 (N_1343,N_902,N_543);
nand U1344 (N_1344,N_749,N_886);
and U1345 (N_1345,N_834,N_855);
or U1346 (N_1346,N_888,N_618);
nor U1347 (N_1347,N_752,N_650);
xor U1348 (N_1348,N_807,N_912);
nand U1349 (N_1349,N_550,N_925);
or U1350 (N_1350,N_713,N_837);
nand U1351 (N_1351,N_983,N_912);
or U1352 (N_1352,N_695,N_888);
and U1353 (N_1353,N_972,N_737);
and U1354 (N_1354,N_681,N_753);
and U1355 (N_1355,N_868,N_740);
nor U1356 (N_1356,N_736,N_918);
or U1357 (N_1357,N_972,N_531);
nand U1358 (N_1358,N_820,N_828);
and U1359 (N_1359,N_952,N_582);
or U1360 (N_1360,N_700,N_994);
xnor U1361 (N_1361,N_713,N_554);
or U1362 (N_1362,N_780,N_570);
xnor U1363 (N_1363,N_777,N_896);
and U1364 (N_1364,N_718,N_826);
and U1365 (N_1365,N_517,N_684);
and U1366 (N_1366,N_684,N_759);
or U1367 (N_1367,N_763,N_707);
or U1368 (N_1368,N_616,N_895);
nor U1369 (N_1369,N_972,N_574);
and U1370 (N_1370,N_951,N_814);
or U1371 (N_1371,N_688,N_979);
nand U1372 (N_1372,N_605,N_610);
nor U1373 (N_1373,N_529,N_786);
or U1374 (N_1374,N_883,N_502);
or U1375 (N_1375,N_761,N_892);
nand U1376 (N_1376,N_641,N_789);
xor U1377 (N_1377,N_916,N_667);
or U1378 (N_1378,N_878,N_611);
nand U1379 (N_1379,N_812,N_651);
or U1380 (N_1380,N_856,N_970);
or U1381 (N_1381,N_526,N_808);
or U1382 (N_1382,N_584,N_624);
and U1383 (N_1383,N_980,N_589);
or U1384 (N_1384,N_598,N_893);
nand U1385 (N_1385,N_771,N_775);
nand U1386 (N_1386,N_954,N_772);
or U1387 (N_1387,N_984,N_513);
nand U1388 (N_1388,N_750,N_799);
nor U1389 (N_1389,N_785,N_577);
or U1390 (N_1390,N_630,N_936);
and U1391 (N_1391,N_935,N_661);
xor U1392 (N_1392,N_828,N_548);
nand U1393 (N_1393,N_534,N_685);
nor U1394 (N_1394,N_881,N_992);
xnor U1395 (N_1395,N_870,N_871);
or U1396 (N_1396,N_706,N_596);
and U1397 (N_1397,N_841,N_538);
nand U1398 (N_1398,N_562,N_815);
or U1399 (N_1399,N_691,N_734);
nand U1400 (N_1400,N_697,N_569);
or U1401 (N_1401,N_828,N_791);
nor U1402 (N_1402,N_735,N_560);
nor U1403 (N_1403,N_840,N_652);
or U1404 (N_1404,N_959,N_997);
nand U1405 (N_1405,N_907,N_791);
nand U1406 (N_1406,N_986,N_902);
or U1407 (N_1407,N_686,N_904);
or U1408 (N_1408,N_953,N_924);
nor U1409 (N_1409,N_960,N_909);
nor U1410 (N_1410,N_637,N_784);
and U1411 (N_1411,N_932,N_704);
or U1412 (N_1412,N_593,N_683);
nand U1413 (N_1413,N_504,N_973);
or U1414 (N_1414,N_907,N_723);
or U1415 (N_1415,N_551,N_937);
xor U1416 (N_1416,N_553,N_962);
nor U1417 (N_1417,N_916,N_986);
nor U1418 (N_1418,N_724,N_997);
nor U1419 (N_1419,N_559,N_552);
and U1420 (N_1420,N_611,N_559);
or U1421 (N_1421,N_950,N_964);
and U1422 (N_1422,N_848,N_930);
nand U1423 (N_1423,N_524,N_618);
and U1424 (N_1424,N_620,N_752);
and U1425 (N_1425,N_541,N_925);
or U1426 (N_1426,N_903,N_588);
xnor U1427 (N_1427,N_725,N_704);
or U1428 (N_1428,N_820,N_644);
and U1429 (N_1429,N_787,N_822);
and U1430 (N_1430,N_653,N_918);
and U1431 (N_1431,N_899,N_763);
or U1432 (N_1432,N_612,N_522);
nor U1433 (N_1433,N_841,N_525);
or U1434 (N_1434,N_515,N_867);
and U1435 (N_1435,N_531,N_869);
nand U1436 (N_1436,N_828,N_605);
and U1437 (N_1437,N_967,N_616);
nand U1438 (N_1438,N_784,N_785);
nor U1439 (N_1439,N_888,N_705);
nor U1440 (N_1440,N_601,N_866);
or U1441 (N_1441,N_715,N_950);
and U1442 (N_1442,N_755,N_972);
nand U1443 (N_1443,N_964,N_898);
xor U1444 (N_1444,N_733,N_713);
xnor U1445 (N_1445,N_566,N_962);
nor U1446 (N_1446,N_818,N_558);
nand U1447 (N_1447,N_614,N_720);
or U1448 (N_1448,N_933,N_545);
and U1449 (N_1449,N_659,N_720);
nand U1450 (N_1450,N_683,N_688);
xnor U1451 (N_1451,N_678,N_602);
and U1452 (N_1452,N_565,N_892);
nor U1453 (N_1453,N_555,N_613);
nor U1454 (N_1454,N_697,N_524);
or U1455 (N_1455,N_573,N_602);
or U1456 (N_1456,N_882,N_902);
nor U1457 (N_1457,N_685,N_573);
nor U1458 (N_1458,N_836,N_604);
nand U1459 (N_1459,N_864,N_729);
and U1460 (N_1460,N_509,N_985);
nor U1461 (N_1461,N_563,N_665);
nor U1462 (N_1462,N_550,N_921);
or U1463 (N_1463,N_728,N_571);
nand U1464 (N_1464,N_732,N_642);
or U1465 (N_1465,N_600,N_880);
or U1466 (N_1466,N_722,N_514);
nor U1467 (N_1467,N_897,N_553);
nand U1468 (N_1468,N_552,N_645);
and U1469 (N_1469,N_557,N_776);
or U1470 (N_1470,N_548,N_921);
nor U1471 (N_1471,N_579,N_917);
nor U1472 (N_1472,N_954,N_976);
and U1473 (N_1473,N_565,N_580);
nand U1474 (N_1474,N_888,N_521);
and U1475 (N_1475,N_951,N_695);
xnor U1476 (N_1476,N_932,N_858);
or U1477 (N_1477,N_847,N_895);
and U1478 (N_1478,N_978,N_803);
or U1479 (N_1479,N_665,N_571);
nor U1480 (N_1480,N_550,N_907);
or U1481 (N_1481,N_610,N_545);
nor U1482 (N_1482,N_886,N_939);
and U1483 (N_1483,N_514,N_803);
or U1484 (N_1484,N_867,N_538);
or U1485 (N_1485,N_859,N_699);
and U1486 (N_1486,N_710,N_575);
or U1487 (N_1487,N_520,N_939);
or U1488 (N_1488,N_723,N_713);
nor U1489 (N_1489,N_704,N_577);
or U1490 (N_1490,N_591,N_525);
or U1491 (N_1491,N_526,N_604);
and U1492 (N_1492,N_605,N_764);
or U1493 (N_1493,N_623,N_930);
nand U1494 (N_1494,N_678,N_522);
nor U1495 (N_1495,N_611,N_826);
or U1496 (N_1496,N_906,N_772);
and U1497 (N_1497,N_998,N_791);
nor U1498 (N_1498,N_522,N_681);
nor U1499 (N_1499,N_917,N_740);
nor U1500 (N_1500,N_1479,N_1221);
and U1501 (N_1501,N_1443,N_1145);
nor U1502 (N_1502,N_1257,N_1112);
and U1503 (N_1503,N_1031,N_1357);
and U1504 (N_1504,N_1407,N_1067);
nor U1505 (N_1505,N_1464,N_1450);
nand U1506 (N_1506,N_1051,N_1455);
nor U1507 (N_1507,N_1389,N_1060);
nor U1508 (N_1508,N_1436,N_1243);
and U1509 (N_1509,N_1196,N_1131);
nor U1510 (N_1510,N_1096,N_1488);
and U1511 (N_1511,N_1003,N_1093);
nor U1512 (N_1512,N_1302,N_1033);
xor U1513 (N_1513,N_1429,N_1063);
xnor U1514 (N_1514,N_1348,N_1168);
nand U1515 (N_1515,N_1207,N_1198);
or U1516 (N_1516,N_1122,N_1329);
nand U1517 (N_1517,N_1249,N_1078);
xor U1518 (N_1518,N_1177,N_1269);
nand U1519 (N_1519,N_1283,N_1366);
and U1520 (N_1520,N_1396,N_1181);
nand U1521 (N_1521,N_1182,N_1330);
and U1522 (N_1522,N_1360,N_1367);
or U1523 (N_1523,N_1020,N_1244);
and U1524 (N_1524,N_1337,N_1164);
nor U1525 (N_1525,N_1327,N_1304);
and U1526 (N_1526,N_1212,N_1085);
xor U1527 (N_1527,N_1483,N_1072);
and U1528 (N_1528,N_1150,N_1363);
and U1529 (N_1529,N_1176,N_1158);
nand U1530 (N_1530,N_1490,N_1333);
and U1531 (N_1531,N_1377,N_1321);
and U1532 (N_1532,N_1376,N_1385);
or U1533 (N_1533,N_1365,N_1448);
or U1534 (N_1534,N_1265,N_1192);
nand U1535 (N_1535,N_1125,N_1190);
and U1536 (N_1536,N_1328,N_1166);
nand U1537 (N_1537,N_1447,N_1395);
nor U1538 (N_1538,N_1191,N_1154);
nand U1539 (N_1539,N_1011,N_1410);
nand U1540 (N_1540,N_1276,N_1120);
or U1541 (N_1541,N_1287,N_1040);
nor U1542 (N_1542,N_1292,N_1345);
or U1543 (N_1543,N_1170,N_1424);
nand U1544 (N_1544,N_1398,N_1107);
nor U1545 (N_1545,N_1126,N_1194);
nand U1546 (N_1546,N_1038,N_1057);
nand U1547 (N_1547,N_1384,N_1435);
nand U1548 (N_1548,N_1458,N_1134);
xnor U1549 (N_1549,N_1471,N_1338);
nand U1550 (N_1550,N_1076,N_1108);
nor U1551 (N_1551,N_1390,N_1266);
nor U1552 (N_1552,N_1024,N_1316);
nor U1553 (N_1553,N_1061,N_1252);
nor U1554 (N_1554,N_1449,N_1086);
nand U1555 (N_1555,N_1326,N_1437);
and U1556 (N_1556,N_1016,N_1215);
and U1557 (N_1557,N_1273,N_1318);
and U1558 (N_1558,N_1115,N_1233);
nor U1559 (N_1559,N_1383,N_1049);
nand U1560 (N_1560,N_1001,N_1209);
nor U1561 (N_1561,N_1402,N_1079);
nand U1562 (N_1562,N_1046,N_1497);
or U1563 (N_1563,N_1225,N_1082);
nand U1564 (N_1564,N_1347,N_1098);
or U1565 (N_1565,N_1071,N_1184);
or U1566 (N_1566,N_1434,N_1064);
or U1567 (N_1567,N_1091,N_1080);
and U1568 (N_1568,N_1454,N_1341);
nor U1569 (N_1569,N_1281,N_1132);
nor U1570 (N_1570,N_1226,N_1043);
or U1571 (N_1571,N_1439,N_1431);
or U1572 (N_1572,N_1259,N_1297);
or U1573 (N_1573,N_1013,N_1161);
and U1574 (N_1574,N_1419,N_1314);
or U1575 (N_1575,N_1460,N_1427);
nor U1576 (N_1576,N_1416,N_1110);
nor U1577 (N_1577,N_1124,N_1202);
and U1578 (N_1578,N_1359,N_1343);
nor U1579 (N_1579,N_1401,N_1068);
nor U1580 (N_1580,N_1008,N_1000);
nand U1581 (N_1581,N_1148,N_1271);
nand U1582 (N_1582,N_1295,N_1426);
nor U1583 (N_1583,N_1279,N_1296);
nand U1584 (N_1584,N_1310,N_1152);
xor U1585 (N_1585,N_1409,N_1397);
nor U1586 (N_1586,N_1356,N_1178);
nand U1587 (N_1587,N_1066,N_1255);
and U1588 (N_1588,N_1189,N_1139);
nand U1589 (N_1589,N_1432,N_1237);
nor U1590 (N_1590,N_1494,N_1324);
and U1591 (N_1591,N_1334,N_1408);
and U1592 (N_1592,N_1232,N_1351);
nor U1593 (N_1593,N_1111,N_1291);
and U1594 (N_1594,N_1456,N_1213);
nand U1595 (N_1595,N_1235,N_1090);
or U1596 (N_1596,N_1224,N_1307);
and U1597 (N_1597,N_1261,N_1153);
nand U1598 (N_1598,N_1228,N_1127);
xor U1599 (N_1599,N_1238,N_1151);
or U1600 (N_1600,N_1109,N_1054);
nor U1601 (N_1601,N_1452,N_1070);
nand U1602 (N_1602,N_1476,N_1149);
and U1603 (N_1603,N_1496,N_1414);
and U1604 (N_1604,N_1270,N_1441);
xnor U1605 (N_1605,N_1413,N_1399);
nor U1606 (N_1606,N_1275,N_1009);
or U1607 (N_1607,N_1286,N_1335);
nor U1608 (N_1608,N_1015,N_1473);
nor U1609 (N_1609,N_1322,N_1141);
and U1610 (N_1610,N_1203,N_1394);
or U1611 (N_1611,N_1218,N_1159);
or U1612 (N_1612,N_1380,N_1251);
and U1613 (N_1613,N_1073,N_1034);
nor U1614 (N_1614,N_1116,N_1463);
nor U1615 (N_1615,N_1174,N_1484);
or U1616 (N_1616,N_1325,N_1133);
nor U1617 (N_1617,N_1263,N_1087);
and U1618 (N_1618,N_1173,N_1155);
and U1619 (N_1619,N_1475,N_1121);
xnor U1620 (N_1620,N_1143,N_1421);
and U1621 (N_1621,N_1032,N_1355);
xor U1622 (N_1622,N_1042,N_1451);
and U1623 (N_1623,N_1467,N_1147);
nand U1624 (N_1624,N_1364,N_1018);
or U1625 (N_1625,N_1320,N_1425);
nand U1626 (N_1626,N_1313,N_1498);
and U1627 (N_1627,N_1388,N_1368);
or U1628 (N_1628,N_1284,N_1470);
and U1629 (N_1629,N_1094,N_1262);
or U1630 (N_1630,N_1246,N_1241);
nand U1631 (N_1631,N_1440,N_1406);
nand U1632 (N_1632,N_1227,N_1478);
nor U1633 (N_1633,N_1250,N_1446);
and U1634 (N_1634,N_1129,N_1391);
xor U1635 (N_1635,N_1231,N_1340);
xnor U1636 (N_1636,N_1010,N_1428);
or U1637 (N_1637,N_1438,N_1422);
nor U1638 (N_1638,N_1106,N_1208);
nor U1639 (N_1639,N_1415,N_1373);
or U1640 (N_1640,N_1021,N_1113);
and U1641 (N_1641,N_1028,N_1358);
nand U1642 (N_1642,N_1216,N_1405);
nand U1643 (N_1643,N_1350,N_1123);
nor U1644 (N_1644,N_1017,N_1240);
nand U1645 (N_1645,N_1387,N_1486);
or U1646 (N_1646,N_1492,N_1099);
or U1647 (N_1647,N_1012,N_1059);
or U1648 (N_1648,N_1005,N_1466);
and U1649 (N_1649,N_1171,N_1206);
or U1650 (N_1650,N_1372,N_1204);
or U1651 (N_1651,N_1056,N_1342);
and U1652 (N_1652,N_1047,N_1362);
nand U1653 (N_1653,N_1323,N_1487);
nor U1654 (N_1654,N_1234,N_1029);
nor U1655 (N_1655,N_1062,N_1392);
or U1656 (N_1656,N_1444,N_1058);
nand U1657 (N_1657,N_1069,N_1393);
nor U1658 (N_1658,N_1433,N_1180);
nor U1659 (N_1659,N_1382,N_1193);
nand U1660 (N_1660,N_1004,N_1400);
and U1661 (N_1661,N_1315,N_1169);
nor U1662 (N_1662,N_1253,N_1274);
nand U1663 (N_1663,N_1239,N_1371);
xnor U1664 (N_1664,N_1481,N_1294);
nor U1665 (N_1665,N_1298,N_1044);
nand U1666 (N_1666,N_1041,N_1205);
xor U1667 (N_1667,N_1077,N_1258);
nor U1668 (N_1668,N_1118,N_1092);
or U1669 (N_1669,N_1370,N_1007);
and U1670 (N_1670,N_1489,N_1197);
nor U1671 (N_1671,N_1344,N_1293);
nand U1672 (N_1672,N_1499,N_1102);
xnor U1673 (N_1673,N_1378,N_1223);
or U1674 (N_1674,N_1285,N_1346);
nand U1675 (N_1675,N_1101,N_1308);
nor U1676 (N_1676,N_1312,N_1306);
or U1677 (N_1677,N_1354,N_1477);
nand U1678 (N_1678,N_1493,N_1201);
or U1679 (N_1679,N_1256,N_1465);
and U1680 (N_1680,N_1163,N_1188);
nand U1681 (N_1681,N_1105,N_1420);
and U1682 (N_1682,N_1290,N_1442);
and U1683 (N_1683,N_1352,N_1055);
nand U1684 (N_1684,N_1211,N_1157);
or U1685 (N_1685,N_1299,N_1319);
nor U1686 (N_1686,N_1461,N_1095);
and U1687 (N_1687,N_1179,N_1187);
nand U1688 (N_1688,N_1305,N_1268);
xnor U1689 (N_1689,N_1272,N_1081);
or U1690 (N_1690,N_1375,N_1374);
or U1691 (N_1691,N_1468,N_1128);
and U1692 (N_1692,N_1183,N_1278);
or U1693 (N_1693,N_1140,N_1472);
and U1694 (N_1694,N_1036,N_1267);
and U1695 (N_1695,N_1411,N_1459);
xnor U1696 (N_1696,N_1156,N_1412);
nand U1697 (N_1697,N_1301,N_1165);
nor U1698 (N_1698,N_1045,N_1303);
nor U1699 (N_1699,N_1023,N_1053);
and U1700 (N_1700,N_1130,N_1491);
and U1701 (N_1701,N_1418,N_1117);
and U1702 (N_1702,N_1014,N_1457);
and U1703 (N_1703,N_1136,N_1264);
nor U1704 (N_1704,N_1311,N_1002);
nand U1705 (N_1705,N_1135,N_1332);
and U1706 (N_1706,N_1138,N_1006);
or U1707 (N_1707,N_1146,N_1100);
or U1708 (N_1708,N_1242,N_1300);
xor U1709 (N_1709,N_1119,N_1217);
nand U1710 (N_1710,N_1289,N_1361);
nand U1711 (N_1711,N_1288,N_1167);
nor U1712 (N_1712,N_1339,N_1025);
and U1713 (N_1713,N_1162,N_1210);
xnor U1714 (N_1714,N_1035,N_1277);
or U1715 (N_1715,N_1219,N_1186);
or U1716 (N_1716,N_1495,N_1030);
nand U1717 (N_1717,N_1474,N_1089);
nand U1718 (N_1718,N_1254,N_1379);
xnor U1719 (N_1719,N_1097,N_1026);
or U1720 (N_1720,N_1220,N_1331);
nand U1721 (N_1721,N_1199,N_1403);
nor U1722 (N_1722,N_1248,N_1386);
and U1723 (N_1723,N_1185,N_1052);
nand U1724 (N_1724,N_1137,N_1480);
nand U1725 (N_1725,N_1430,N_1103);
nand U1726 (N_1726,N_1353,N_1280);
and U1727 (N_1727,N_1230,N_1083);
and U1728 (N_1728,N_1417,N_1027);
and U1729 (N_1729,N_1469,N_1022);
and U1730 (N_1730,N_1445,N_1084);
nor U1731 (N_1731,N_1485,N_1019);
nand U1732 (N_1732,N_1048,N_1037);
or U1733 (N_1733,N_1175,N_1195);
and U1734 (N_1734,N_1065,N_1282);
or U1735 (N_1735,N_1309,N_1039);
nand U1736 (N_1736,N_1245,N_1453);
and U1737 (N_1737,N_1482,N_1349);
nand U1738 (N_1738,N_1088,N_1247);
and U1739 (N_1739,N_1229,N_1214);
nor U1740 (N_1740,N_1222,N_1144);
or U1741 (N_1741,N_1462,N_1336);
xnor U1742 (N_1742,N_1404,N_1114);
or U1743 (N_1743,N_1142,N_1075);
nand U1744 (N_1744,N_1423,N_1172);
nor U1745 (N_1745,N_1381,N_1369);
or U1746 (N_1746,N_1050,N_1074);
or U1747 (N_1747,N_1160,N_1317);
nand U1748 (N_1748,N_1200,N_1104);
nand U1749 (N_1749,N_1236,N_1260);
and U1750 (N_1750,N_1133,N_1387);
nor U1751 (N_1751,N_1057,N_1101);
nor U1752 (N_1752,N_1290,N_1308);
and U1753 (N_1753,N_1253,N_1064);
nor U1754 (N_1754,N_1256,N_1444);
nor U1755 (N_1755,N_1115,N_1496);
nand U1756 (N_1756,N_1451,N_1445);
nand U1757 (N_1757,N_1312,N_1302);
nor U1758 (N_1758,N_1001,N_1188);
nor U1759 (N_1759,N_1004,N_1072);
nand U1760 (N_1760,N_1062,N_1115);
nor U1761 (N_1761,N_1188,N_1404);
or U1762 (N_1762,N_1284,N_1157);
xnor U1763 (N_1763,N_1470,N_1389);
nand U1764 (N_1764,N_1244,N_1348);
nor U1765 (N_1765,N_1076,N_1390);
nor U1766 (N_1766,N_1212,N_1290);
or U1767 (N_1767,N_1275,N_1410);
nor U1768 (N_1768,N_1142,N_1037);
or U1769 (N_1769,N_1498,N_1363);
nor U1770 (N_1770,N_1405,N_1352);
and U1771 (N_1771,N_1017,N_1117);
and U1772 (N_1772,N_1305,N_1424);
xnor U1773 (N_1773,N_1294,N_1174);
or U1774 (N_1774,N_1165,N_1319);
nand U1775 (N_1775,N_1484,N_1298);
or U1776 (N_1776,N_1212,N_1238);
and U1777 (N_1777,N_1289,N_1385);
nand U1778 (N_1778,N_1146,N_1315);
nand U1779 (N_1779,N_1338,N_1257);
or U1780 (N_1780,N_1134,N_1486);
nand U1781 (N_1781,N_1426,N_1318);
and U1782 (N_1782,N_1473,N_1265);
or U1783 (N_1783,N_1027,N_1015);
and U1784 (N_1784,N_1116,N_1342);
nand U1785 (N_1785,N_1498,N_1135);
nor U1786 (N_1786,N_1189,N_1278);
nand U1787 (N_1787,N_1381,N_1111);
or U1788 (N_1788,N_1222,N_1461);
and U1789 (N_1789,N_1063,N_1145);
nor U1790 (N_1790,N_1006,N_1456);
or U1791 (N_1791,N_1043,N_1025);
or U1792 (N_1792,N_1079,N_1204);
or U1793 (N_1793,N_1375,N_1159);
xnor U1794 (N_1794,N_1371,N_1093);
nor U1795 (N_1795,N_1087,N_1190);
or U1796 (N_1796,N_1161,N_1445);
or U1797 (N_1797,N_1414,N_1409);
and U1798 (N_1798,N_1397,N_1022);
and U1799 (N_1799,N_1187,N_1341);
and U1800 (N_1800,N_1131,N_1490);
nor U1801 (N_1801,N_1288,N_1305);
xnor U1802 (N_1802,N_1482,N_1270);
and U1803 (N_1803,N_1249,N_1387);
nand U1804 (N_1804,N_1082,N_1123);
xnor U1805 (N_1805,N_1174,N_1454);
nor U1806 (N_1806,N_1409,N_1327);
xnor U1807 (N_1807,N_1106,N_1402);
and U1808 (N_1808,N_1266,N_1203);
nor U1809 (N_1809,N_1174,N_1168);
or U1810 (N_1810,N_1474,N_1000);
xor U1811 (N_1811,N_1425,N_1499);
and U1812 (N_1812,N_1303,N_1006);
or U1813 (N_1813,N_1138,N_1373);
xor U1814 (N_1814,N_1090,N_1468);
or U1815 (N_1815,N_1003,N_1235);
nand U1816 (N_1816,N_1263,N_1253);
nor U1817 (N_1817,N_1452,N_1107);
xor U1818 (N_1818,N_1470,N_1311);
nand U1819 (N_1819,N_1299,N_1127);
and U1820 (N_1820,N_1137,N_1436);
or U1821 (N_1821,N_1135,N_1005);
nand U1822 (N_1822,N_1000,N_1099);
nor U1823 (N_1823,N_1063,N_1372);
and U1824 (N_1824,N_1049,N_1101);
or U1825 (N_1825,N_1299,N_1070);
nand U1826 (N_1826,N_1202,N_1471);
or U1827 (N_1827,N_1185,N_1158);
xnor U1828 (N_1828,N_1068,N_1359);
nand U1829 (N_1829,N_1172,N_1061);
nor U1830 (N_1830,N_1115,N_1301);
or U1831 (N_1831,N_1117,N_1019);
or U1832 (N_1832,N_1374,N_1390);
nand U1833 (N_1833,N_1276,N_1096);
or U1834 (N_1834,N_1430,N_1019);
nand U1835 (N_1835,N_1446,N_1170);
or U1836 (N_1836,N_1105,N_1223);
nand U1837 (N_1837,N_1273,N_1209);
and U1838 (N_1838,N_1469,N_1411);
nor U1839 (N_1839,N_1167,N_1374);
nor U1840 (N_1840,N_1095,N_1045);
nor U1841 (N_1841,N_1208,N_1259);
nor U1842 (N_1842,N_1212,N_1442);
nand U1843 (N_1843,N_1354,N_1010);
nand U1844 (N_1844,N_1352,N_1367);
and U1845 (N_1845,N_1119,N_1310);
xor U1846 (N_1846,N_1313,N_1142);
or U1847 (N_1847,N_1014,N_1086);
and U1848 (N_1848,N_1029,N_1015);
nand U1849 (N_1849,N_1060,N_1452);
xnor U1850 (N_1850,N_1210,N_1188);
and U1851 (N_1851,N_1172,N_1132);
xnor U1852 (N_1852,N_1177,N_1030);
nor U1853 (N_1853,N_1468,N_1234);
nor U1854 (N_1854,N_1126,N_1417);
and U1855 (N_1855,N_1346,N_1320);
nor U1856 (N_1856,N_1013,N_1066);
or U1857 (N_1857,N_1029,N_1239);
nor U1858 (N_1858,N_1208,N_1471);
nand U1859 (N_1859,N_1471,N_1248);
nor U1860 (N_1860,N_1217,N_1076);
nand U1861 (N_1861,N_1298,N_1412);
nand U1862 (N_1862,N_1091,N_1426);
or U1863 (N_1863,N_1075,N_1369);
and U1864 (N_1864,N_1066,N_1398);
nor U1865 (N_1865,N_1265,N_1176);
nand U1866 (N_1866,N_1000,N_1133);
and U1867 (N_1867,N_1422,N_1004);
and U1868 (N_1868,N_1390,N_1063);
or U1869 (N_1869,N_1177,N_1139);
nand U1870 (N_1870,N_1439,N_1419);
and U1871 (N_1871,N_1064,N_1082);
nand U1872 (N_1872,N_1254,N_1173);
or U1873 (N_1873,N_1065,N_1325);
and U1874 (N_1874,N_1014,N_1178);
nor U1875 (N_1875,N_1204,N_1060);
nor U1876 (N_1876,N_1247,N_1009);
nand U1877 (N_1877,N_1431,N_1228);
xor U1878 (N_1878,N_1235,N_1118);
and U1879 (N_1879,N_1436,N_1312);
xor U1880 (N_1880,N_1218,N_1075);
nor U1881 (N_1881,N_1276,N_1475);
nor U1882 (N_1882,N_1132,N_1004);
xor U1883 (N_1883,N_1171,N_1306);
nand U1884 (N_1884,N_1423,N_1249);
or U1885 (N_1885,N_1225,N_1400);
xor U1886 (N_1886,N_1257,N_1115);
and U1887 (N_1887,N_1244,N_1357);
or U1888 (N_1888,N_1053,N_1205);
and U1889 (N_1889,N_1097,N_1155);
or U1890 (N_1890,N_1139,N_1469);
xor U1891 (N_1891,N_1385,N_1261);
and U1892 (N_1892,N_1147,N_1170);
nand U1893 (N_1893,N_1061,N_1147);
nand U1894 (N_1894,N_1105,N_1264);
xor U1895 (N_1895,N_1214,N_1285);
and U1896 (N_1896,N_1068,N_1013);
or U1897 (N_1897,N_1370,N_1160);
nand U1898 (N_1898,N_1420,N_1071);
nand U1899 (N_1899,N_1065,N_1053);
nand U1900 (N_1900,N_1126,N_1446);
nand U1901 (N_1901,N_1423,N_1436);
nand U1902 (N_1902,N_1266,N_1015);
xnor U1903 (N_1903,N_1443,N_1353);
nor U1904 (N_1904,N_1232,N_1090);
nand U1905 (N_1905,N_1440,N_1263);
and U1906 (N_1906,N_1258,N_1129);
nand U1907 (N_1907,N_1210,N_1271);
or U1908 (N_1908,N_1492,N_1480);
nand U1909 (N_1909,N_1133,N_1347);
and U1910 (N_1910,N_1106,N_1155);
nor U1911 (N_1911,N_1203,N_1140);
nand U1912 (N_1912,N_1237,N_1228);
and U1913 (N_1913,N_1244,N_1238);
and U1914 (N_1914,N_1209,N_1028);
or U1915 (N_1915,N_1372,N_1452);
nand U1916 (N_1916,N_1468,N_1242);
nor U1917 (N_1917,N_1368,N_1375);
nand U1918 (N_1918,N_1181,N_1182);
nor U1919 (N_1919,N_1286,N_1456);
nor U1920 (N_1920,N_1446,N_1318);
or U1921 (N_1921,N_1489,N_1417);
or U1922 (N_1922,N_1388,N_1022);
and U1923 (N_1923,N_1440,N_1386);
nor U1924 (N_1924,N_1004,N_1138);
and U1925 (N_1925,N_1088,N_1394);
nand U1926 (N_1926,N_1298,N_1244);
and U1927 (N_1927,N_1287,N_1499);
nand U1928 (N_1928,N_1217,N_1253);
xnor U1929 (N_1929,N_1390,N_1119);
nor U1930 (N_1930,N_1348,N_1102);
and U1931 (N_1931,N_1017,N_1131);
nor U1932 (N_1932,N_1361,N_1427);
xnor U1933 (N_1933,N_1116,N_1403);
xnor U1934 (N_1934,N_1418,N_1437);
nor U1935 (N_1935,N_1163,N_1303);
and U1936 (N_1936,N_1360,N_1354);
xnor U1937 (N_1937,N_1293,N_1479);
nor U1938 (N_1938,N_1221,N_1428);
or U1939 (N_1939,N_1022,N_1361);
and U1940 (N_1940,N_1363,N_1220);
and U1941 (N_1941,N_1496,N_1244);
nor U1942 (N_1942,N_1189,N_1028);
and U1943 (N_1943,N_1135,N_1008);
nand U1944 (N_1944,N_1106,N_1471);
and U1945 (N_1945,N_1291,N_1192);
nor U1946 (N_1946,N_1020,N_1187);
and U1947 (N_1947,N_1118,N_1096);
nand U1948 (N_1948,N_1278,N_1363);
nand U1949 (N_1949,N_1158,N_1041);
or U1950 (N_1950,N_1063,N_1488);
nand U1951 (N_1951,N_1471,N_1182);
nor U1952 (N_1952,N_1214,N_1073);
and U1953 (N_1953,N_1026,N_1153);
nor U1954 (N_1954,N_1476,N_1245);
or U1955 (N_1955,N_1424,N_1240);
nand U1956 (N_1956,N_1180,N_1320);
nand U1957 (N_1957,N_1417,N_1451);
and U1958 (N_1958,N_1323,N_1267);
or U1959 (N_1959,N_1466,N_1045);
nand U1960 (N_1960,N_1495,N_1496);
or U1961 (N_1961,N_1306,N_1294);
nand U1962 (N_1962,N_1213,N_1401);
and U1963 (N_1963,N_1280,N_1249);
nor U1964 (N_1964,N_1021,N_1038);
or U1965 (N_1965,N_1498,N_1176);
or U1966 (N_1966,N_1125,N_1242);
and U1967 (N_1967,N_1226,N_1217);
and U1968 (N_1968,N_1025,N_1277);
nand U1969 (N_1969,N_1422,N_1183);
nand U1970 (N_1970,N_1151,N_1406);
and U1971 (N_1971,N_1199,N_1061);
or U1972 (N_1972,N_1190,N_1338);
or U1973 (N_1973,N_1230,N_1133);
and U1974 (N_1974,N_1217,N_1445);
nand U1975 (N_1975,N_1294,N_1448);
or U1976 (N_1976,N_1401,N_1182);
or U1977 (N_1977,N_1269,N_1109);
nand U1978 (N_1978,N_1441,N_1089);
nand U1979 (N_1979,N_1205,N_1427);
nor U1980 (N_1980,N_1346,N_1449);
or U1981 (N_1981,N_1406,N_1340);
or U1982 (N_1982,N_1132,N_1043);
nor U1983 (N_1983,N_1496,N_1090);
or U1984 (N_1984,N_1467,N_1152);
nor U1985 (N_1985,N_1079,N_1362);
nor U1986 (N_1986,N_1328,N_1386);
xnor U1987 (N_1987,N_1145,N_1006);
nor U1988 (N_1988,N_1041,N_1369);
and U1989 (N_1989,N_1011,N_1089);
nand U1990 (N_1990,N_1193,N_1105);
or U1991 (N_1991,N_1331,N_1299);
or U1992 (N_1992,N_1079,N_1299);
nor U1993 (N_1993,N_1223,N_1355);
xor U1994 (N_1994,N_1433,N_1297);
nand U1995 (N_1995,N_1447,N_1143);
or U1996 (N_1996,N_1256,N_1178);
or U1997 (N_1997,N_1495,N_1052);
nand U1998 (N_1998,N_1001,N_1170);
nand U1999 (N_1999,N_1195,N_1458);
or U2000 (N_2000,N_1711,N_1837);
and U2001 (N_2001,N_1696,N_1967);
or U2002 (N_2002,N_1574,N_1861);
xor U2003 (N_2003,N_1719,N_1513);
and U2004 (N_2004,N_1564,N_1732);
nor U2005 (N_2005,N_1651,N_1607);
or U2006 (N_2006,N_1899,N_1684);
nor U2007 (N_2007,N_1787,N_1571);
and U2008 (N_2008,N_1643,N_1878);
and U2009 (N_2009,N_1982,N_1912);
and U2010 (N_2010,N_1504,N_1692);
and U2011 (N_2011,N_1802,N_1936);
nor U2012 (N_2012,N_1977,N_1911);
and U2013 (N_2013,N_1636,N_1520);
nand U2014 (N_2014,N_1944,N_1815);
or U2015 (N_2015,N_1949,N_1757);
nor U2016 (N_2016,N_1552,N_1993);
nand U2017 (N_2017,N_1700,N_1540);
and U2018 (N_2018,N_1909,N_1854);
or U2019 (N_2019,N_1502,N_1793);
xnor U2020 (N_2020,N_1928,N_1821);
xor U2021 (N_2021,N_1503,N_1637);
nand U2022 (N_2022,N_1863,N_1976);
nand U2023 (N_2023,N_1649,N_1901);
nand U2024 (N_2024,N_1597,N_1544);
nand U2025 (N_2025,N_1688,N_1683);
and U2026 (N_2026,N_1934,N_1619);
nor U2027 (N_2027,N_1783,N_1691);
and U2028 (N_2028,N_1754,N_1834);
and U2029 (N_2029,N_1748,N_1890);
xor U2030 (N_2030,N_1988,N_1960);
nand U2031 (N_2031,N_1839,N_1717);
nor U2032 (N_2032,N_1616,N_1773);
and U2033 (N_2033,N_1853,N_1781);
nor U2034 (N_2034,N_1566,N_1873);
nand U2035 (N_2035,N_1575,N_1900);
and U2036 (N_2036,N_1841,N_1823);
nand U2037 (N_2037,N_1752,N_1930);
or U2038 (N_2038,N_1868,N_1755);
and U2039 (N_2039,N_1563,N_1908);
xnor U2040 (N_2040,N_1737,N_1756);
nand U2041 (N_2041,N_1595,N_1985);
xor U2042 (N_2042,N_1678,N_1623);
nor U2043 (N_2043,N_1604,N_1672);
nor U2044 (N_2044,N_1689,N_1610);
nor U2045 (N_2045,N_1654,N_1971);
nor U2046 (N_2046,N_1827,N_1903);
or U2047 (N_2047,N_1990,N_1892);
and U2048 (N_2048,N_1989,N_1555);
nand U2049 (N_2049,N_1613,N_1542);
nor U2050 (N_2050,N_1699,N_1921);
or U2051 (N_2051,N_1995,N_1587);
nand U2052 (N_2052,N_1550,N_1582);
xnor U2053 (N_2053,N_1956,N_1716);
or U2054 (N_2054,N_1975,N_1818);
or U2055 (N_2055,N_1655,N_1507);
and U2056 (N_2056,N_1560,N_1685);
nand U2057 (N_2057,N_1686,N_1953);
nand U2058 (N_2058,N_1628,N_1606);
nand U2059 (N_2059,N_1952,N_1541);
or U2060 (N_2060,N_1762,N_1938);
nor U2061 (N_2061,N_1617,N_1573);
xnor U2062 (N_2062,N_1517,N_1519);
nand U2063 (N_2063,N_1926,N_1723);
or U2064 (N_2064,N_1782,N_1799);
nor U2065 (N_2065,N_1728,N_1669);
or U2066 (N_2066,N_1585,N_1648);
nor U2067 (N_2067,N_1736,N_1620);
nor U2068 (N_2068,N_1994,N_1796);
and U2069 (N_2069,N_1786,N_1816);
nand U2070 (N_2070,N_1798,N_1531);
and U2071 (N_2071,N_1652,N_1720);
nor U2072 (N_2072,N_1634,N_1906);
nor U2073 (N_2073,N_1904,N_1920);
nand U2074 (N_2074,N_1891,N_1941);
nand U2075 (N_2075,N_1917,N_1933);
nor U2076 (N_2076,N_1761,N_1803);
nand U2077 (N_2077,N_1614,N_1664);
nand U2078 (N_2078,N_1876,N_1704);
or U2079 (N_2079,N_1851,N_1833);
nand U2080 (N_2080,N_1894,N_1725);
xnor U2081 (N_2081,N_1794,N_1661);
or U2082 (N_2082,N_1624,N_1806);
nor U2083 (N_2083,N_1509,N_1528);
nor U2084 (N_2084,N_1972,N_1826);
and U2085 (N_2085,N_1663,N_1553);
and U2086 (N_2086,N_1644,N_1819);
nand U2087 (N_2087,N_1500,N_1730);
nor U2088 (N_2088,N_1939,N_1998);
nor U2089 (N_2089,N_1775,N_1910);
nor U2090 (N_2090,N_1974,N_1514);
or U2091 (N_2091,N_1742,N_1556);
nand U2092 (N_2092,N_1545,N_1687);
nor U2093 (N_2093,N_1638,N_1847);
nor U2094 (N_2094,N_1522,N_1931);
nor U2095 (N_2095,N_1532,N_1549);
nor U2096 (N_2096,N_1769,N_1872);
and U2097 (N_2097,N_1877,N_1992);
nor U2098 (N_2098,N_1508,N_1800);
and U2099 (N_2099,N_1785,N_1779);
or U2100 (N_2100,N_1832,N_1935);
nor U2101 (N_2101,N_1603,N_1741);
and U2102 (N_2102,N_1801,N_1590);
or U2103 (N_2103,N_1784,N_1647);
and U2104 (N_2104,N_1862,N_1860);
nor U2105 (N_2105,N_1896,N_1665);
nor U2106 (N_2106,N_1721,N_1615);
nor U2107 (N_2107,N_1562,N_1812);
or U2108 (N_2108,N_1797,N_1724);
nand U2109 (N_2109,N_1588,N_1836);
and U2110 (N_2110,N_1602,N_1961);
or U2111 (N_2111,N_1653,N_1970);
and U2112 (N_2112,N_1568,N_1694);
nor U2113 (N_2113,N_1712,N_1771);
nand U2114 (N_2114,N_1848,N_1889);
or U2115 (N_2115,N_1764,N_1829);
and U2116 (N_2116,N_1999,N_1776);
and U2117 (N_2117,N_1518,N_1963);
and U2118 (N_2118,N_1625,N_1580);
nand U2119 (N_2119,N_1957,N_1830);
or U2120 (N_2120,N_1635,N_1902);
nand U2121 (N_2121,N_1825,N_1709);
nand U2122 (N_2122,N_1656,N_1981);
nor U2123 (N_2123,N_1918,N_1991);
nor U2124 (N_2124,N_1701,N_1674);
nor U2125 (N_2125,N_1506,N_1551);
xnor U2126 (N_2126,N_1739,N_1706);
nor U2127 (N_2127,N_1633,N_1630);
nand U2128 (N_2128,N_1817,N_1547);
nor U2129 (N_2129,N_1855,N_1789);
or U2130 (N_2130,N_1707,N_1594);
or U2131 (N_2131,N_1774,N_1584);
xor U2132 (N_2132,N_1919,N_1767);
nand U2133 (N_2133,N_1640,N_1927);
nor U2134 (N_2134,N_1599,N_1576);
nand U2135 (N_2135,N_1768,N_1641);
nand U2136 (N_2136,N_1526,N_1539);
nand U2137 (N_2137,N_1632,N_1697);
nand U2138 (N_2138,N_1505,N_1969);
and U2139 (N_2139,N_1626,N_1954);
xnor U2140 (N_2140,N_1530,N_1759);
or U2141 (N_2141,N_1516,N_1515);
nor U2142 (N_2142,N_1622,N_1790);
and U2143 (N_2143,N_1907,N_1923);
xnor U2144 (N_2144,N_1535,N_1929);
or U2145 (N_2145,N_1766,N_1842);
nand U2146 (N_2146,N_1533,N_1780);
nand U2147 (N_2147,N_1950,N_1888);
nand U2148 (N_2148,N_1852,N_1858);
nor U2149 (N_2149,N_1627,N_1645);
and U2150 (N_2150,N_1940,N_1810);
nor U2151 (N_2151,N_1955,N_1924);
or U2152 (N_2152,N_1824,N_1554);
nor U2153 (N_2153,N_1579,N_1679);
or U2154 (N_2154,N_1512,N_1611);
nor U2155 (N_2155,N_1673,N_1893);
nand U2156 (N_2156,N_1592,N_1844);
or U2157 (N_2157,N_1601,N_1598);
nand U2158 (N_2158,N_1659,N_1753);
nor U2159 (N_2159,N_1879,N_1875);
nor U2160 (N_2160,N_1867,N_1925);
nand U2161 (N_2161,N_1869,N_1979);
nor U2162 (N_2162,N_1968,N_1548);
nand U2163 (N_2163,N_1589,N_1746);
nor U2164 (N_2164,N_1523,N_1572);
and U2165 (N_2165,N_1543,N_1557);
and U2166 (N_2166,N_1942,N_1702);
nor U2167 (N_2167,N_1639,N_1880);
nand U2168 (N_2168,N_1642,N_1561);
and U2169 (N_2169,N_1546,N_1932);
or U2170 (N_2170,N_1612,N_1738);
xnor U2171 (N_2171,N_1629,N_1510);
and U2172 (N_2172,N_1666,N_1814);
and U2173 (N_2173,N_1733,N_1807);
or U2174 (N_2174,N_1850,N_1822);
or U2175 (N_2175,N_1915,N_1859);
nand U2176 (N_2176,N_1914,N_1559);
and U2177 (N_2177,N_1886,N_1600);
nor U2178 (N_2178,N_1865,N_1698);
nand U2179 (N_2179,N_1671,N_1681);
and U2180 (N_2180,N_1758,N_1745);
nor U2181 (N_2181,N_1772,N_1811);
nor U2182 (N_2182,N_1788,N_1727);
nand U2183 (N_2183,N_1805,N_1675);
nor U2184 (N_2184,N_1987,N_1751);
nor U2185 (N_2185,N_1570,N_1715);
and U2186 (N_2186,N_1866,N_1760);
or U2187 (N_2187,N_1650,N_1948);
and U2188 (N_2188,N_1897,N_1770);
and U2189 (N_2189,N_1558,N_1795);
or U2190 (N_2190,N_1578,N_1567);
nand U2191 (N_2191,N_1997,N_1682);
nand U2192 (N_2192,N_1871,N_1605);
or U2193 (N_2193,N_1947,N_1884);
or U2194 (N_2194,N_1905,N_1529);
nand U2195 (N_2195,N_1750,N_1916);
and U2196 (N_2196,N_1621,N_1708);
and U2197 (N_2197,N_1937,N_1521);
or U2198 (N_2198,N_1680,N_1534);
xnor U2199 (N_2199,N_1951,N_1856);
nand U2200 (N_2200,N_1662,N_1966);
nand U2201 (N_2201,N_1962,N_1831);
nor U2202 (N_2202,N_1980,N_1731);
nor U2203 (N_2203,N_1804,N_1735);
and U2204 (N_2204,N_1658,N_1973);
nand U2205 (N_2205,N_1820,N_1922);
or U2206 (N_2206,N_1729,N_1986);
or U2207 (N_2207,N_1596,N_1667);
or U2208 (N_2208,N_1581,N_1808);
nor U2209 (N_2209,N_1591,N_1945);
nor U2210 (N_2210,N_1608,N_1657);
xor U2211 (N_2211,N_1747,N_1857);
xnor U2212 (N_2212,N_1586,N_1714);
nor U2213 (N_2213,N_1718,N_1996);
nor U2214 (N_2214,N_1791,N_1882);
and U2215 (N_2215,N_1946,N_1726);
or U2216 (N_2216,N_1959,N_1722);
or U2217 (N_2217,N_1870,N_1765);
and U2218 (N_2218,N_1843,N_1537);
or U2219 (N_2219,N_1943,N_1792);
and U2220 (N_2220,N_1743,N_1887);
and U2221 (N_2221,N_1569,N_1984);
xnor U2222 (N_2222,N_1744,N_1538);
or U2223 (N_2223,N_1813,N_1846);
nor U2224 (N_2224,N_1670,N_1690);
or U2225 (N_2225,N_1895,N_1646);
nor U2226 (N_2226,N_1828,N_1835);
nor U2227 (N_2227,N_1898,N_1695);
and U2228 (N_2228,N_1618,N_1749);
and U2229 (N_2229,N_1881,N_1978);
and U2230 (N_2230,N_1525,N_1740);
or U2231 (N_2231,N_1913,N_1840);
and U2232 (N_2232,N_1577,N_1677);
nor U2233 (N_2233,N_1536,N_1838);
nor U2234 (N_2234,N_1501,N_1524);
xor U2235 (N_2235,N_1885,N_1864);
nor U2236 (N_2236,N_1809,N_1609);
xnor U2237 (N_2237,N_1660,N_1777);
or U2238 (N_2238,N_1713,N_1583);
and U2239 (N_2239,N_1845,N_1527);
or U2240 (N_2240,N_1705,N_1565);
nor U2241 (N_2241,N_1734,N_1849);
nor U2242 (N_2242,N_1511,N_1693);
or U2243 (N_2243,N_1874,N_1676);
nand U2244 (N_2244,N_1631,N_1983);
nand U2245 (N_2245,N_1965,N_1593);
and U2246 (N_2246,N_1883,N_1964);
and U2247 (N_2247,N_1668,N_1710);
nor U2248 (N_2248,N_1778,N_1703);
or U2249 (N_2249,N_1958,N_1763);
nor U2250 (N_2250,N_1956,N_1838);
and U2251 (N_2251,N_1731,N_1843);
or U2252 (N_2252,N_1732,N_1742);
nand U2253 (N_2253,N_1638,N_1593);
or U2254 (N_2254,N_1710,N_1794);
or U2255 (N_2255,N_1649,N_1583);
or U2256 (N_2256,N_1543,N_1701);
nand U2257 (N_2257,N_1953,N_1806);
and U2258 (N_2258,N_1724,N_1592);
and U2259 (N_2259,N_1625,N_1619);
nand U2260 (N_2260,N_1741,N_1812);
nor U2261 (N_2261,N_1775,N_1806);
xor U2262 (N_2262,N_1802,N_1778);
and U2263 (N_2263,N_1753,N_1859);
and U2264 (N_2264,N_1704,N_1620);
nor U2265 (N_2265,N_1576,N_1521);
nand U2266 (N_2266,N_1787,N_1829);
nor U2267 (N_2267,N_1668,N_1604);
and U2268 (N_2268,N_1643,N_1564);
and U2269 (N_2269,N_1502,N_1840);
and U2270 (N_2270,N_1675,N_1649);
and U2271 (N_2271,N_1525,N_1625);
or U2272 (N_2272,N_1688,N_1501);
and U2273 (N_2273,N_1858,N_1641);
and U2274 (N_2274,N_1538,N_1527);
and U2275 (N_2275,N_1781,N_1922);
nand U2276 (N_2276,N_1685,N_1740);
or U2277 (N_2277,N_1898,N_1931);
or U2278 (N_2278,N_1961,N_1611);
nand U2279 (N_2279,N_1888,N_1809);
nand U2280 (N_2280,N_1976,N_1692);
and U2281 (N_2281,N_1773,N_1969);
xnor U2282 (N_2282,N_1854,N_1877);
nand U2283 (N_2283,N_1578,N_1805);
nand U2284 (N_2284,N_1548,N_1809);
nor U2285 (N_2285,N_1790,N_1911);
and U2286 (N_2286,N_1835,N_1899);
or U2287 (N_2287,N_1734,N_1577);
nor U2288 (N_2288,N_1959,N_1545);
nor U2289 (N_2289,N_1548,N_1504);
and U2290 (N_2290,N_1910,N_1762);
nand U2291 (N_2291,N_1960,N_1968);
or U2292 (N_2292,N_1946,N_1902);
nand U2293 (N_2293,N_1521,N_1987);
nand U2294 (N_2294,N_1539,N_1645);
and U2295 (N_2295,N_1647,N_1569);
or U2296 (N_2296,N_1791,N_1789);
or U2297 (N_2297,N_1963,N_1740);
and U2298 (N_2298,N_1580,N_1936);
xnor U2299 (N_2299,N_1928,N_1892);
or U2300 (N_2300,N_1909,N_1921);
or U2301 (N_2301,N_1711,N_1802);
nor U2302 (N_2302,N_1864,N_1762);
or U2303 (N_2303,N_1880,N_1886);
and U2304 (N_2304,N_1796,N_1941);
nand U2305 (N_2305,N_1621,N_1677);
xor U2306 (N_2306,N_1679,N_1917);
nand U2307 (N_2307,N_1784,N_1880);
and U2308 (N_2308,N_1792,N_1882);
and U2309 (N_2309,N_1959,N_1856);
or U2310 (N_2310,N_1799,N_1706);
or U2311 (N_2311,N_1582,N_1923);
nand U2312 (N_2312,N_1514,N_1691);
and U2313 (N_2313,N_1801,N_1556);
nor U2314 (N_2314,N_1748,N_1558);
and U2315 (N_2315,N_1638,N_1774);
xor U2316 (N_2316,N_1593,N_1589);
nand U2317 (N_2317,N_1819,N_1501);
or U2318 (N_2318,N_1511,N_1913);
nand U2319 (N_2319,N_1944,N_1560);
and U2320 (N_2320,N_1651,N_1869);
nor U2321 (N_2321,N_1666,N_1505);
and U2322 (N_2322,N_1802,N_1570);
and U2323 (N_2323,N_1868,N_1875);
or U2324 (N_2324,N_1605,N_1554);
nand U2325 (N_2325,N_1605,N_1557);
nand U2326 (N_2326,N_1503,N_1727);
xnor U2327 (N_2327,N_1938,N_1765);
and U2328 (N_2328,N_1864,N_1580);
nand U2329 (N_2329,N_1846,N_1606);
or U2330 (N_2330,N_1525,N_1855);
and U2331 (N_2331,N_1549,N_1752);
nand U2332 (N_2332,N_1938,N_1557);
and U2333 (N_2333,N_1836,N_1677);
and U2334 (N_2334,N_1673,N_1571);
nand U2335 (N_2335,N_1887,N_1566);
nand U2336 (N_2336,N_1632,N_1958);
and U2337 (N_2337,N_1500,N_1666);
and U2338 (N_2338,N_1921,N_1702);
and U2339 (N_2339,N_1982,N_1849);
and U2340 (N_2340,N_1558,N_1931);
nand U2341 (N_2341,N_1746,N_1541);
nand U2342 (N_2342,N_1645,N_1849);
xnor U2343 (N_2343,N_1785,N_1626);
nor U2344 (N_2344,N_1544,N_1658);
nor U2345 (N_2345,N_1747,N_1515);
nor U2346 (N_2346,N_1967,N_1626);
or U2347 (N_2347,N_1936,N_1727);
or U2348 (N_2348,N_1932,N_1949);
and U2349 (N_2349,N_1689,N_1551);
xor U2350 (N_2350,N_1567,N_1806);
and U2351 (N_2351,N_1976,N_1804);
nor U2352 (N_2352,N_1870,N_1613);
nand U2353 (N_2353,N_1594,N_1675);
nand U2354 (N_2354,N_1750,N_1628);
xor U2355 (N_2355,N_1545,N_1893);
or U2356 (N_2356,N_1805,N_1510);
and U2357 (N_2357,N_1960,N_1619);
nand U2358 (N_2358,N_1834,N_1555);
nor U2359 (N_2359,N_1888,N_1696);
xor U2360 (N_2360,N_1722,N_1507);
and U2361 (N_2361,N_1931,N_1850);
and U2362 (N_2362,N_1584,N_1566);
or U2363 (N_2363,N_1886,N_1642);
nor U2364 (N_2364,N_1911,N_1902);
or U2365 (N_2365,N_1795,N_1781);
xor U2366 (N_2366,N_1901,N_1664);
nor U2367 (N_2367,N_1982,N_1829);
or U2368 (N_2368,N_1575,N_1869);
or U2369 (N_2369,N_1657,N_1796);
and U2370 (N_2370,N_1736,N_1721);
or U2371 (N_2371,N_1833,N_1744);
and U2372 (N_2372,N_1954,N_1515);
nor U2373 (N_2373,N_1753,N_1758);
and U2374 (N_2374,N_1966,N_1658);
nor U2375 (N_2375,N_1759,N_1778);
or U2376 (N_2376,N_1982,N_1790);
and U2377 (N_2377,N_1861,N_1942);
and U2378 (N_2378,N_1601,N_1804);
nand U2379 (N_2379,N_1663,N_1786);
or U2380 (N_2380,N_1896,N_1989);
or U2381 (N_2381,N_1997,N_1543);
or U2382 (N_2382,N_1554,N_1980);
and U2383 (N_2383,N_1640,N_1834);
or U2384 (N_2384,N_1813,N_1619);
and U2385 (N_2385,N_1834,N_1577);
and U2386 (N_2386,N_1629,N_1807);
and U2387 (N_2387,N_1928,N_1834);
or U2388 (N_2388,N_1756,N_1579);
or U2389 (N_2389,N_1967,N_1992);
and U2390 (N_2390,N_1525,N_1698);
nor U2391 (N_2391,N_1582,N_1660);
nor U2392 (N_2392,N_1816,N_1565);
nand U2393 (N_2393,N_1557,N_1554);
and U2394 (N_2394,N_1585,N_1864);
nor U2395 (N_2395,N_1946,N_1606);
or U2396 (N_2396,N_1623,N_1669);
or U2397 (N_2397,N_1517,N_1958);
nor U2398 (N_2398,N_1746,N_1915);
nor U2399 (N_2399,N_1821,N_1896);
and U2400 (N_2400,N_1864,N_1886);
xnor U2401 (N_2401,N_1988,N_1600);
and U2402 (N_2402,N_1600,N_1648);
nand U2403 (N_2403,N_1889,N_1833);
nand U2404 (N_2404,N_1589,N_1982);
nand U2405 (N_2405,N_1877,N_1905);
or U2406 (N_2406,N_1890,N_1927);
or U2407 (N_2407,N_1724,N_1792);
and U2408 (N_2408,N_1899,N_1647);
nor U2409 (N_2409,N_1833,N_1807);
and U2410 (N_2410,N_1558,N_1900);
or U2411 (N_2411,N_1993,N_1841);
or U2412 (N_2412,N_1897,N_1718);
and U2413 (N_2413,N_1594,N_1507);
or U2414 (N_2414,N_1979,N_1528);
or U2415 (N_2415,N_1596,N_1654);
nor U2416 (N_2416,N_1770,N_1755);
nand U2417 (N_2417,N_1863,N_1883);
and U2418 (N_2418,N_1804,N_1798);
nor U2419 (N_2419,N_1552,N_1568);
nand U2420 (N_2420,N_1999,N_1755);
or U2421 (N_2421,N_1776,N_1781);
or U2422 (N_2422,N_1971,N_1655);
or U2423 (N_2423,N_1959,N_1539);
nand U2424 (N_2424,N_1666,N_1516);
xor U2425 (N_2425,N_1786,N_1911);
xnor U2426 (N_2426,N_1654,N_1681);
and U2427 (N_2427,N_1693,N_1726);
nor U2428 (N_2428,N_1635,N_1880);
nand U2429 (N_2429,N_1973,N_1906);
or U2430 (N_2430,N_1952,N_1865);
nand U2431 (N_2431,N_1766,N_1917);
nand U2432 (N_2432,N_1726,N_1985);
nor U2433 (N_2433,N_1833,N_1862);
nand U2434 (N_2434,N_1649,N_1737);
nor U2435 (N_2435,N_1768,N_1881);
nand U2436 (N_2436,N_1572,N_1864);
nor U2437 (N_2437,N_1801,N_1992);
and U2438 (N_2438,N_1887,N_1983);
nor U2439 (N_2439,N_1537,N_1809);
nand U2440 (N_2440,N_1782,N_1777);
and U2441 (N_2441,N_1923,N_1854);
xnor U2442 (N_2442,N_1841,N_1671);
and U2443 (N_2443,N_1949,N_1593);
or U2444 (N_2444,N_1948,N_1992);
xor U2445 (N_2445,N_1855,N_1858);
or U2446 (N_2446,N_1819,N_1638);
nand U2447 (N_2447,N_1915,N_1814);
or U2448 (N_2448,N_1684,N_1718);
nand U2449 (N_2449,N_1923,N_1876);
and U2450 (N_2450,N_1668,N_1528);
nand U2451 (N_2451,N_1648,N_1748);
nand U2452 (N_2452,N_1728,N_1892);
xnor U2453 (N_2453,N_1826,N_1867);
or U2454 (N_2454,N_1546,N_1841);
xor U2455 (N_2455,N_1652,N_1711);
nand U2456 (N_2456,N_1614,N_1909);
and U2457 (N_2457,N_1990,N_1547);
nand U2458 (N_2458,N_1971,N_1890);
and U2459 (N_2459,N_1897,N_1726);
nor U2460 (N_2460,N_1676,N_1844);
and U2461 (N_2461,N_1701,N_1734);
nand U2462 (N_2462,N_1959,N_1521);
nor U2463 (N_2463,N_1960,N_1865);
nand U2464 (N_2464,N_1930,N_1958);
nor U2465 (N_2465,N_1981,N_1610);
nor U2466 (N_2466,N_1678,N_1608);
and U2467 (N_2467,N_1957,N_1540);
nor U2468 (N_2468,N_1577,N_1930);
nand U2469 (N_2469,N_1842,N_1859);
nor U2470 (N_2470,N_1904,N_1687);
xor U2471 (N_2471,N_1883,N_1843);
nor U2472 (N_2472,N_1725,N_1520);
xor U2473 (N_2473,N_1941,N_1508);
or U2474 (N_2474,N_1514,N_1698);
or U2475 (N_2475,N_1870,N_1519);
or U2476 (N_2476,N_1730,N_1803);
nor U2477 (N_2477,N_1814,N_1508);
or U2478 (N_2478,N_1681,N_1949);
or U2479 (N_2479,N_1969,N_1696);
xnor U2480 (N_2480,N_1797,N_1895);
or U2481 (N_2481,N_1588,N_1515);
nand U2482 (N_2482,N_1881,N_1610);
and U2483 (N_2483,N_1577,N_1658);
nand U2484 (N_2484,N_1823,N_1548);
nand U2485 (N_2485,N_1807,N_1949);
or U2486 (N_2486,N_1908,N_1714);
xnor U2487 (N_2487,N_1818,N_1509);
nor U2488 (N_2488,N_1763,N_1595);
or U2489 (N_2489,N_1932,N_1958);
nor U2490 (N_2490,N_1653,N_1642);
nand U2491 (N_2491,N_1520,N_1828);
nor U2492 (N_2492,N_1844,N_1926);
and U2493 (N_2493,N_1926,N_1579);
nor U2494 (N_2494,N_1505,N_1771);
xnor U2495 (N_2495,N_1920,N_1948);
xor U2496 (N_2496,N_1563,N_1887);
nor U2497 (N_2497,N_1687,N_1588);
nor U2498 (N_2498,N_1935,N_1561);
nand U2499 (N_2499,N_1728,N_1845);
or U2500 (N_2500,N_2109,N_2350);
nand U2501 (N_2501,N_2481,N_2455);
and U2502 (N_2502,N_2184,N_2442);
or U2503 (N_2503,N_2336,N_2141);
and U2504 (N_2504,N_2163,N_2240);
or U2505 (N_2505,N_2100,N_2359);
nor U2506 (N_2506,N_2028,N_2010);
and U2507 (N_2507,N_2454,N_2219);
nand U2508 (N_2508,N_2170,N_2417);
nor U2509 (N_2509,N_2158,N_2257);
xnor U2510 (N_2510,N_2361,N_2200);
nor U2511 (N_2511,N_2444,N_2472);
nor U2512 (N_2512,N_2462,N_2117);
xnor U2513 (N_2513,N_2319,N_2042);
nand U2514 (N_2514,N_2258,N_2285);
xor U2515 (N_2515,N_2494,N_2263);
nor U2516 (N_2516,N_2202,N_2015);
nand U2517 (N_2517,N_2367,N_2495);
nand U2518 (N_2518,N_2372,N_2103);
nand U2519 (N_2519,N_2093,N_2185);
or U2520 (N_2520,N_2133,N_2448);
nand U2521 (N_2521,N_2484,N_2296);
and U2522 (N_2522,N_2204,N_2412);
nor U2523 (N_2523,N_2314,N_2058);
and U2524 (N_2524,N_2247,N_2199);
nand U2525 (N_2525,N_2322,N_2121);
or U2526 (N_2526,N_2421,N_2483);
nor U2527 (N_2527,N_2377,N_2370);
nor U2528 (N_2528,N_2174,N_2497);
nor U2529 (N_2529,N_2392,N_2321);
nor U2530 (N_2530,N_2159,N_2434);
nor U2531 (N_2531,N_2046,N_2292);
nand U2532 (N_2532,N_2362,N_2168);
nand U2533 (N_2533,N_2080,N_2179);
nor U2534 (N_2534,N_2255,N_2413);
and U2535 (N_2535,N_2051,N_2308);
nand U2536 (N_2536,N_2471,N_2301);
or U2537 (N_2537,N_2169,N_2156);
or U2538 (N_2538,N_2279,N_2261);
and U2539 (N_2539,N_2461,N_2001);
nor U2540 (N_2540,N_2379,N_2487);
and U2541 (N_2541,N_2406,N_2091);
nor U2542 (N_2542,N_2333,N_2101);
and U2543 (N_2543,N_2265,N_2467);
nand U2544 (N_2544,N_2127,N_2380);
nor U2545 (N_2545,N_2162,N_2102);
nand U2546 (N_2546,N_2008,N_2346);
or U2547 (N_2547,N_2374,N_2271);
and U2548 (N_2548,N_2254,N_2086);
or U2549 (N_2549,N_2234,N_2335);
and U2550 (N_2550,N_2252,N_2173);
xor U2551 (N_2551,N_2074,N_2171);
nand U2552 (N_2552,N_2192,N_2228);
and U2553 (N_2553,N_2233,N_2390);
and U2554 (N_2554,N_2036,N_2343);
and U2555 (N_2555,N_2437,N_2428);
nor U2556 (N_2556,N_2139,N_2224);
or U2557 (N_2557,N_2191,N_2394);
xor U2558 (N_2558,N_2193,N_2073);
nand U2559 (N_2559,N_2023,N_2099);
nand U2560 (N_2560,N_2026,N_2157);
nor U2561 (N_2561,N_2276,N_2241);
nor U2562 (N_2562,N_2189,N_2423);
nand U2563 (N_2563,N_2107,N_2003);
nor U2564 (N_2564,N_2355,N_2118);
or U2565 (N_2565,N_2386,N_2112);
or U2566 (N_2566,N_2289,N_2356);
nand U2567 (N_2567,N_2070,N_2050);
or U2568 (N_2568,N_2248,N_2340);
nor U2569 (N_2569,N_2106,N_2368);
and U2570 (N_2570,N_2266,N_2024);
nand U2571 (N_2571,N_2014,N_2272);
and U2572 (N_2572,N_2007,N_2396);
nor U2573 (N_2573,N_2165,N_2230);
nand U2574 (N_2574,N_2426,N_2299);
or U2575 (N_2575,N_2161,N_2237);
nor U2576 (N_2576,N_2131,N_2398);
xor U2577 (N_2577,N_2145,N_2357);
or U2578 (N_2578,N_2443,N_2077);
and U2579 (N_2579,N_2498,N_2302);
or U2580 (N_2580,N_2485,N_2383);
and U2581 (N_2581,N_2315,N_2470);
nor U2582 (N_2582,N_2128,N_2281);
nor U2583 (N_2583,N_2060,N_2190);
and U2584 (N_2584,N_2229,N_2166);
nand U2585 (N_2585,N_2277,N_2337);
nand U2586 (N_2586,N_2120,N_2045);
nand U2587 (N_2587,N_2420,N_2135);
nor U2588 (N_2588,N_2071,N_2013);
nand U2589 (N_2589,N_2293,N_2205);
or U2590 (N_2590,N_2125,N_2317);
nand U2591 (N_2591,N_2476,N_2344);
or U2592 (N_2592,N_2463,N_2327);
and U2593 (N_2593,N_2123,N_2197);
nor U2594 (N_2594,N_2178,N_2339);
or U2595 (N_2595,N_2212,N_2399);
nand U2596 (N_2596,N_2387,N_2220);
xor U2597 (N_2597,N_2430,N_2410);
nand U2598 (N_2598,N_2009,N_2020);
and U2599 (N_2599,N_2324,N_2040);
or U2600 (N_2600,N_2114,N_2273);
nor U2601 (N_2601,N_2290,N_2287);
or U2602 (N_2602,N_2280,N_2391);
and U2603 (N_2603,N_2116,N_2130);
nand U2604 (N_2604,N_2416,N_2016);
nand U2605 (N_2605,N_2326,N_2221);
and U2606 (N_2606,N_2492,N_2458);
nor U2607 (N_2607,N_2075,N_2198);
nor U2608 (N_2608,N_2351,N_2404);
nand U2609 (N_2609,N_2218,N_2429);
or U2610 (N_2610,N_2460,N_2294);
nor U2611 (N_2611,N_2039,N_2066);
nand U2612 (N_2612,N_2011,N_2303);
and U2613 (N_2613,N_2088,N_2445);
nor U2614 (N_2614,N_2181,N_2186);
and U2615 (N_2615,N_2160,N_2140);
and U2616 (N_2616,N_2278,N_2262);
nor U2617 (N_2617,N_2243,N_2083);
or U2618 (N_2618,N_2384,N_2411);
and U2619 (N_2619,N_2425,N_2076);
nand U2620 (N_2620,N_2295,N_2403);
or U2621 (N_2621,N_2284,N_2288);
nand U2622 (N_2622,N_2110,N_2473);
or U2623 (N_2623,N_2264,N_2283);
or U2624 (N_2624,N_2490,N_2175);
and U2625 (N_2625,N_2239,N_2354);
or U2626 (N_2626,N_2352,N_2019);
and U2627 (N_2627,N_2424,N_2347);
nand U2628 (N_2628,N_2316,N_2402);
and U2629 (N_2629,N_2095,N_2208);
nor U2630 (N_2630,N_2477,N_2167);
or U2631 (N_2631,N_2201,N_2064);
and U2632 (N_2632,N_2090,N_2496);
and U2633 (N_2633,N_2489,N_2318);
nand U2634 (N_2634,N_2069,N_2297);
and U2635 (N_2635,N_2401,N_2486);
nand U2636 (N_2636,N_2466,N_2005);
and U2637 (N_2637,N_2081,N_2134);
and U2638 (N_2638,N_2018,N_2056);
nor U2639 (N_2639,N_2065,N_2433);
and U2640 (N_2640,N_2482,N_2054);
and U2641 (N_2641,N_2030,N_2222);
and U2642 (N_2642,N_2092,N_2253);
nor U2643 (N_2643,N_2479,N_2098);
nand U2644 (N_2644,N_2311,N_2176);
nor U2645 (N_2645,N_2447,N_2381);
or U2646 (N_2646,N_2022,N_2155);
and U2647 (N_2647,N_2378,N_2478);
nand U2648 (N_2648,N_2027,N_2035);
nor U2649 (N_2649,N_2148,N_2052);
or U2650 (N_2650,N_2451,N_2365);
nand U2651 (N_2651,N_2049,N_2260);
xnor U2652 (N_2652,N_2310,N_2457);
nand U2653 (N_2653,N_2061,N_2236);
or U2654 (N_2654,N_2085,N_2151);
and U2655 (N_2655,N_2067,N_2342);
nand U2656 (N_2656,N_2195,N_2043);
nand U2657 (N_2657,N_2246,N_2366);
nor U2658 (N_2658,N_2154,N_2111);
nor U2659 (N_2659,N_2021,N_2488);
nand U2660 (N_2660,N_2465,N_2360);
nand U2661 (N_2661,N_2491,N_2033);
nor U2662 (N_2662,N_2180,N_2094);
and U2663 (N_2663,N_2144,N_2446);
or U2664 (N_2664,N_2249,N_2017);
xnor U2665 (N_2665,N_2172,N_2480);
or U2666 (N_2666,N_2275,N_2147);
xor U2667 (N_2667,N_2259,N_2215);
and U2668 (N_2668,N_2242,N_2376);
nand U2669 (N_2669,N_2129,N_2382);
or U2670 (N_2670,N_2441,N_2493);
nor U2671 (N_2671,N_2087,N_2320);
nand U2672 (N_2672,N_2137,N_2312);
nand U2673 (N_2673,N_2329,N_2223);
nor U2674 (N_2674,N_2267,N_2300);
nand U2675 (N_2675,N_2364,N_2432);
and U2676 (N_2676,N_2216,N_2375);
and U2677 (N_2677,N_2115,N_2097);
or U2678 (N_2678,N_2213,N_2323);
or U2679 (N_2679,N_2206,N_2025);
nand U2680 (N_2680,N_2328,N_2146);
or U2681 (N_2681,N_2187,N_2459);
and U2682 (N_2682,N_2474,N_2464);
or U2683 (N_2683,N_2126,N_2150);
or U2684 (N_2684,N_2306,N_2291);
or U2685 (N_2685,N_2400,N_2440);
nor U2686 (N_2686,N_2245,N_2389);
nor U2687 (N_2687,N_2143,N_2334);
and U2688 (N_2688,N_2132,N_2227);
nor U2689 (N_2689,N_2068,N_2452);
or U2690 (N_2690,N_2006,N_2079);
nor U2691 (N_2691,N_2053,N_2153);
nand U2692 (N_2692,N_2072,N_2034);
nand U2693 (N_2693,N_2456,N_2244);
xnor U2694 (N_2694,N_2325,N_2251);
and U2695 (N_2695,N_2078,N_2207);
nand U2696 (N_2696,N_2012,N_2371);
or U2697 (N_2697,N_2231,N_2305);
nand U2698 (N_2698,N_2196,N_2286);
or U2699 (N_2699,N_2388,N_2124);
nand U2700 (N_2700,N_2307,N_2149);
nor U2701 (N_2701,N_2453,N_2211);
and U2702 (N_2702,N_2435,N_2209);
nor U2703 (N_2703,N_2108,N_2385);
nand U2704 (N_2704,N_2274,N_2004);
and U2705 (N_2705,N_2415,N_2238);
nor U2706 (N_2706,N_2353,N_2063);
nand U2707 (N_2707,N_2341,N_2450);
and U2708 (N_2708,N_2203,N_2408);
nand U2709 (N_2709,N_2373,N_2183);
nand U2710 (N_2710,N_2304,N_2037);
nand U2711 (N_2711,N_2089,N_2000);
nand U2712 (N_2712,N_2225,N_2029);
and U2713 (N_2713,N_2418,N_2499);
xnor U2714 (N_2714,N_2405,N_2397);
and U2715 (N_2715,N_2041,N_2422);
and U2716 (N_2716,N_2313,N_2439);
or U2717 (N_2717,N_2331,N_2177);
and U2718 (N_2718,N_2369,N_2330);
nand U2719 (N_2719,N_2214,N_2084);
nand U2720 (N_2720,N_2136,N_2194);
and U2721 (N_2721,N_2393,N_2469);
or U2722 (N_2722,N_2407,N_2055);
nand U2723 (N_2723,N_2358,N_2138);
and U2724 (N_2724,N_2096,N_2152);
nor U2725 (N_2725,N_2217,N_2282);
xor U2726 (N_2726,N_2431,N_2250);
nor U2727 (N_2727,N_2235,N_2031);
nor U2728 (N_2728,N_2119,N_2438);
xnor U2729 (N_2729,N_2038,N_2348);
nand U2730 (N_2730,N_2082,N_2338);
or U2731 (N_2731,N_2419,N_2349);
nand U2732 (N_2732,N_2104,N_2182);
and U2733 (N_2733,N_2057,N_2164);
nor U2734 (N_2734,N_2059,N_2298);
nand U2735 (N_2735,N_2047,N_2113);
and U2736 (N_2736,N_2268,N_2436);
or U2737 (N_2737,N_2363,N_2332);
or U2738 (N_2738,N_2468,N_2142);
nand U2739 (N_2739,N_2395,N_2475);
nor U2740 (N_2740,N_2062,N_2414);
and U2741 (N_2741,N_2105,N_2427);
and U2742 (N_2742,N_2188,N_2269);
or U2743 (N_2743,N_2345,N_2048);
or U2744 (N_2744,N_2002,N_2044);
xnor U2745 (N_2745,N_2449,N_2409);
or U2746 (N_2746,N_2032,N_2226);
xnor U2747 (N_2747,N_2122,N_2232);
and U2748 (N_2748,N_2256,N_2270);
and U2749 (N_2749,N_2210,N_2309);
and U2750 (N_2750,N_2441,N_2370);
and U2751 (N_2751,N_2165,N_2178);
and U2752 (N_2752,N_2042,N_2119);
nand U2753 (N_2753,N_2172,N_2228);
xnor U2754 (N_2754,N_2222,N_2027);
and U2755 (N_2755,N_2332,N_2301);
nand U2756 (N_2756,N_2011,N_2085);
and U2757 (N_2757,N_2442,N_2069);
or U2758 (N_2758,N_2261,N_2157);
nand U2759 (N_2759,N_2014,N_2057);
or U2760 (N_2760,N_2223,N_2220);
nor U2761 (N_2761,N_2150,N_2309);
and U2762 (N_2762,N_2266,N_2147);
or U2763 (N_2763,N_2273,N_2340);
nand U2764 (N_2764,N_2155,N_2027);
and U2765 (N_2765,N_2265,N_2089);
and U2766 (N_2766,N_2081,N_2302);
or U2767 (N_2767,N_2312,N_2434);
and U2768 (N_2768,N_2161,N_2223);
nand U2769 (N_2769,N_2063,N_2399);
and U2770 (N_2770,N_2100,N_2142);
or U2771 (N_2771,N_2407,N_2151);
or U2772 (N_2772,N_2128,N_2226);
xor U2773 (N_2773,N_2204,N_2175);
nor U2774 (N_2774,N_2058,N_2085);
or U2775 (N_2775,N_2405,N_2137);
or U2776 (N_2776,N_2188,N_2327);
and U2777 (N_2777,N_2197,N_2271);
nor U2778 (N_2778,N_2104,N_2376);
nor U2779 (N_2779,N_2392,N_2446);
and U2780 (N_2780,N_2132,N_2200);
or U2781 (N_2781,N_2092,N_2285);
or U2782 (N_2782,N_2006,N_2380);
or U2783 (N_2783,N_2360,N_2199);
or U2784 (N_2784,N_2063,N_2275);
nor U2785 (N_2785,N_2417,N_2452);
nor U2786 (N_2786,N_2246,N_2286);
or U2787 (N_2787,N_2486,N_2022);
nand U2788 (N_2788,N_2042,N_2382);
or U2789 (N_2789,N_2449,N_2193);
and U2790 (N_2790,N_2018,N_2262);
and U2791 (N_2791,N_2210,N_2202);
and U2792 (N_2792,N_2296,N_2378);
and U2793 (N_2793,N_2090,N_2479);
nand U2794 (N_2794,N_2127,N_2439);
nand U2795 (N_2795,N_2444,N_2267);
nand U2796 (N_2796,N_2192,N_2417);
and U2797 (N_2797,N_2371,N_2370);
or U2798 (N_2798,N_2070,N_2174);
nand U2799 (N_2799,N_2095,N_2181);
nor U2800 (N_2800,N_2446,N_2286);
and U2801 (N_2801,N_2077,N_2421);
nor U2802 (N_2802,N_2490,N_2007);
or U2803 (N_2803,N_2492,N_2372);
nor U2804 (N_2804,N_2092,N_2045);
nor U2805 (N_2805,N_2007,N_2487);
xor U2806 (N_2806,N_2362,N_2486);
xor U2807 (N_2807,N_2134,N_2303);
nor U2808 (N_2808,N_2480,N_2344);
nor U2809 (N_2809,N_2015,N_2153);
and U2810 (N_2810,N_2476,N_2309);
nand U2811 (N_2811,N_2333,N_2424);
xnor U2812 (N_2812,N_2339,N_2447);
and U2813 (N_2813,N_2181,N_2212);
nand U2814 (N_2814,N_2097,N_2427);
or U2815 (N_2815,N_2335,N_2361);
and U2816 (N_2816,N_2242,N_2258);
nor U2817 (N_2817,N_2147,N_2008);
nand U2818 (N_2818,N_2209,N_2401);
nor U2819 (N_2819,N_2099,N_2304);
xor U2820 (N_2820,N_2190,N_2265);
or U2821 (N_2821,N_2417,N_2197);
nand U2822 (N_2822,N_2248,N_2226);
and U2823 (N_2823,N_2427,N_2268);
or U2824 (N_2824,N_2261,N_2021);
xnor U2825 (N_2825,N_2351,N_2355);
nand U2826 (N_2826,N_2285,N_2389);
nor U2827 (N_2827,N_2419,N_2015);
nor U2828 (N_2828,N_2415,N_2078);
and U2829 (N_2829,N_2380,N_2131);
and U2830 (N_2830,N_2167,N_2217);
nand U2831 (N_2831,N_2390,N_2082);
and U2832 (N_2832,N_2375,N_2285);
or U2833 (N_2833,N_2036,N_2140);
nand U2834 (N_2834,N_2111,N_2046);
nand U2835 (N_2835,N_2268,N_2448);
nand U2836 (N_2836,N_2092,N_2095);
and U2837 (N_2837,N_2201,N_2190);
nor U2838 (N_2838,N_2463,N_2000);
and U2839 (N_2839,N_2183,N_2015);
nand U2840 (N_2840,N_2471,N_2191);
nor U2841 (N_2841,N_2451,N_2494);
nor U2842 (N_2842,N_2041,N_2204);
or U2843 (N_2843,N_2202,N_2266);
nand U2844 (N_2844,N_2356,N_2132);
nand U2845 (N_2845,N_2021,N_2419);
or U2846 (N_2846,N_2329,N_2266);
or U2847 (N_2847,N_2145,N_2232);
or U2848 (N_2848,N_2105,N_2443);
nand U2849 (N_2849,N_2391,N_2003);
nand U2850 (N_2850,N_2293,N_2331);
and U2851 (N_2851,N_2394,N_2083);
nand U2852 (N_2852,N_2388,N_2226);
nor U2853 (N_2853,N_2142,N_2151);
xnor U2854 (N_2854,N_2438,N_2444);
xnor U2855 (N_2855,N_2043,N_2182);
or U2856 (N_2856,N_2360,N_2293);
or U2857 (N_2857,N_2120,N_2168);
nand U2858 (N_2858,N_2435,N_2251);
nor U2859 (N_2859,N_2194,N_2425);
and U2860 (N_2860,N_2232,N_2466);
xnor U2861 (N_2861,N_2059,N_2035);
nor U2862 (N_2862,N_2056,N_2124);
and U2863 (N_2863,N_2455,N_2340);
nor U2864 (N_2864,N_2105,N_2322);
and U2865 (N_2865,N_2318,N_2186);
nand U2866 (N_2866,N_2031,N_2446);
xnor U2867 (N_2867,N_2068,N_2144);
nand U2868 (N_2868,N_2421,N_2389);
nor U2869 (N_2869,N_2438,N_2033);
and U2870 (N_2870,N_2474,N_2413);
or U2871 (N_2871,N_2005,N_2484);
and U2872 (N_2872,N_2070,N_2309);
nor U2873 (N_2873,N_2482,N_2484);
and U2874 (N_2874,N_2110,N_2233);
and U2875 (N_2875,N_2000,N_2328);
and U2876 (N_2876,N_2033,N_2322);
or U2877 (N_2877,N_2373,N_2193);
xor U2878 (N_2878,N_2162,N_2257);
nor U2879 (N_2879,N_2387,N_2350);
or U2880 (N_2880,N_2384,N_2400);
or U2881 (N_2881,N_2078,N_2425);
xnor U2882 (N_2882,N_2392,N_2257);
and U2883 (N_2883,N_2374,N_2428);
and U2884 (N_2884,N_2109,N_2087);
nor U2885 (N_2885,N_2093,N_2286);
xnor U2886 (N_2886,N_2377,N_2091);
nor U2887 (N_2887,N_2264,N_2315);
nor U2888 (N_2888,N_2467,N_2197);
nand U2889 (N_2889,N_2300,N_2205);
nand U2890 (N_2890,N_2139,N_2482);
or U2891 (N_2891,N_2013,N_2080);
or U2892 (N_2892,N_2190,N_2432);
nand U2893 (N_2893,N_2387,N_2008);
nand U2894 (N_2894,N_2272,N_2024);
nor U2895 (N_2895,N_2057,N_2238);
nand U2896 (N_2896,N_2219,N_2440);
and U2897 (N_2897,N_2301,N_2409);
nor U2898 (N_2898,N_2262,N_2384);
nor U2899 (N_2899,N_2301,N_2122);
or U2900 (N_2900,N_2253,N_2076);
or U2901 (N_2901,N_2436,N_2472);
and U2902 (N_2902,N_2221,N_2083);
and U2903 (N_2903,N_2264,N_2334);
or U2904 (N_2904,N_2419,N_2033);
nor U2905 (N_2905,N_2105,N_2206);
and U2906 (N_2906,N_2290,N_2260);
or U2907 (N_2907,N_2482,N_2224);
nor U2908 (N_2908,N_2375,N_2303);
nand U2909 (N_2909,N_2441,N_2276);
nand U2910 (N_2910,N_2055,N_2361);
nor U2911 (N_2911,N_2355,N_2316);
nand U2912 (N_2912,N_2226,N_2067);
or U2913 (N_2913,N_2129,N_2480);
nand U2914 (N_2914,N_2432,N_2407);
nor U2915 (N_2915,N_2451,N_2370);
nand U2916 (N_2916,N_2084,N_2131);
nand U2917 (N_2917,N_2243,N_2200);
xnor U2918 (N_2918,N_2175,N_2328);
and U2919 (N_2919,N_2031,N_2484);
or U2920 (N_2920,N_2151,N_2408);
nor U2921 (N_2921,N_2269,N_2068);
and U2922 (N_2922,N_2419,N_2129);
and U2923 (N_2923,N_2104,N_2450);
nor U2924 (N_2924,N_2264,N_2361);
nand U2925 (N_2925,N_2211,N_2313);
and U2926 (N_2926,N_2331,N_2458);
and U2927 (N_2927,N_2343,N_2023);
xnor U2928 (N_2928,N_2248,N_2299);
nand U2929 (N_2929,N_2002,N_2166);
or U2930 (N_2930,N_2420,N_2488);
nor U2931 (N_2931,N_2192,N_2071);
or U2932 (N_2932,N_2059,N_2003);
and U2933 (N_2933,N_2447,N_2225);
nand U2934 (N_2934,N_2298,N_2125);
and U2935 (N_2935,N_2421,N_2060);
or U2936 (N_2936,N_2137,N_2096);
and U2937 (N_2937,N_2249,N_2332);
nor U2938 (N_2938,N_2401,N_2459);
nand U2939 (N_2939,N_2334,N_2249);
xor U2940 (N_2940,N_2495,N_2368);
and U2941 (N_2941,N_2037,N_2068);
nand U2942 (N_2942,N_2430,N_2415);
and U2943 (N_2943,N_2070,N_2270);
and U2944 (N_2944,N_2293,N_2240);
or U2945 (N_2945,N_2026,N_2001);
and U2946 (N_2946,N_2084,N_2238);
nor U2947 (N_2947,N_2249,N_2006);
or U2948 (N_2948,N_2144,N_2067);
xnor U2949 (N_2949,N_2362,N_2249);
and U2950 (N_2950,N_2000,N_2274);
nor U2951 (N_2951,N_2265,N_2483);
and U2952 (N_2952,N_2214,N_2038);
or U2953 (N_2953,N_2169,N_2015);
and U2954 (N_2954,N_2258,N_2494);
nand U2955 (N_2955,N_2239,N_2148);
nand U2956 (N_2956,N_2427,N_2180);
nor U2957 (N_2957,N_2179,N_2233);
and U2958 (N_2958,N_2215,N_2382);
nand U2959 (N_2959,N_2230,N_2038);
or U2960 (N_2960,N_2431,N_2043);
or U2961 (N_2961,N_2082,N_2466);
or U2962 (N_2962,N_2126,N_2377);
nor U2963 (N_2963,N_2459,N_2188);
or U2964 (N_2964,N_2014,N_2045);
nand U2965 (N_2965,N_2440,N_2420);
nor U2966 (N_2966,N_2464,N_2132);
nand U2967 (N_2967,N_2173,N_2022);
nand U2968 (N_2968,N_2378,N_2394);
xnor U2969 (N_2969,N_2327,N_2113);
nand U2970 (N_2970,N_2488,N_2155);
or U2971 (N_2971,N_2261,N_2353);
and U2972 (N_2972,N_2122,N_2049);
nor U2973 (N_2973,N_2219,N_2107);
nor U2974 (N_2974,N_2128,N_2184);
nand U2975 (N_2975,N_2172,N_2132);
xor U2976 (N_2976,N_2078,N_2472);
and U2977 (N_2977,N_2321,N_2041);
and U2978 (N_2978,N_2377,N_2425);
nor U2979 (N_2979,N_2417,N_2060);
and U2980 (N_2980,N_2131,N_2491);
and U2981 (N_2981,N_2261,N_2491);
or U2982 (N_2982,N_2234,N_2333);
nor U2983 (N_2983,N_2274,N_2153);
nor U2984 (N_2984,N_2388,N_2271);
nor U2985 (N_2985,N_2275,N_2293);
or U2986 (N_2986,N_2331,N_2380);
nand U2987 (N_2987,N_2171,N_2068);
nand U2988 (N_2988,N_2106,N_2097);
and U2989 (N_2989,N_2239,N_2218);
nor U2990 (N_2990,N_2325,N_2150);
and U2991 (N_2991,N_2457,N_2413);
xor U2992 (N_2992,N_2230,N_2264);
nor U2993 (N_2993,N_2438,N_2494);
nor U2994 (N_2994,N_2246,N_2298);
nor U2995 (N_2995,N_2072,N_2452);
xor U2996 (N_2996,N_2110,N_2439);
nand U2997 (N_2997,N_2303,N_2092);
and U2998 (N_2998,N_2348,N_2002);
xor U2999 (N_2999,N_2482,N_2269);
nand U3000 (N_3000,N_2957,N_2796);
or U3001 (N_3001,N_2792,N_2810);
nor U3002 (N_3002,N_2506,N_2913);
and U3003 (N_3003,N_2633,N_2733);
nand U3004 (N_3004,N_2959,N_2614);
nor U3005 (N_3005,N_2599,N_2604);
xnor U3006 (N_3006,N_2942,N_2669);
nor U3007 (N_3007,N_2778,N_2892);
and U3008 (N_3008,N_2522,N_2896);
nand U3009 (N_3009,N_2543,N_2908);
or U3010 (N_3010,N_2759,N_2576);
nor U3011 (N_3011,N_2713,N_2779);
nand U3012 (N_3012,N_2820,N_2680);
or U3013 (N_3013,N_2515,N_2945);
and U3014 (N_3014,N_2620,N_2535);
and U3015 (N_3015,N_2685,N_2590);
or U3016 (N_3016,N_2802,N_2763);
or U3017 (N_3017,N_2617,N_2518);
and U3018 (N_3018,N_2541,N_2902);
xor U3019 (N_3019,N_2901,N_2904);
nand U3020 (N_3020,N_2533,N_2530);
xnor U3021 (N_3021,N_2843,N_2992);
and U3022 (N_3022,N_2740,N_2975);
and U3023 (N_3023,N_2983,N_2721);
and U3024 (N_3024,N_2677,N_2678);
nor U3025 (N_3025,N_2508,N_2972);
xnor U3026 (N_3026,N_2825,N_2690);
nand U3027 (N_3027,N_2723,N_2621);
or U3028 (N_3028,N_2640,N_2840);
or U3029 (N_3029,N_2752,N_2513);
nor U3030 (N_3030,N_2742,N_2847);
or U3031 (N_3031,N_2786,N_2747);
or U3032 (N_3032,N_2775,N_2780);
nand U3033 (N_3033,N_2563,N_2641);
nand U3034 (N_3034,N_2939,N_2603);
nand U3035 (N_3035,N_2666,N_2963);
nor U3036 (N_3036,N_2812,N_2824);
and U3037 (N_3037,N_2708,N_2981);
xor U3038 (N_3038,N_2635,N_2647);
nand U3039 (N_3039,N_2798,N_2863);
nand U3040 (N_3040,N_2996,N_2536);
and U3041 (N_3041,N_2745,N_2800);
or U3042 (N_3042,N_2643,N_2547);
nand U3043 (N_3043,N_2605,N_2671);
nor U3044 (N_3044,N_2804,N_2969);
or U3045 (N_3045,N_2750,N_2806);
and U3046 (N_3046,N_2987,N_2593);
or U3047 (N_3047,N_2550,N_2553);
nand U3048 (N_3048,N_2586,N_2727);
nor U3049 (N_3049,N_2566,N_2882);
xnor U3050 (N_3050,N_2676,N_2537);
and U3051 (N_3051,N_2795,N_2601);
and U3052 (N_3052,N_2661,N_2912);
xnor U3053 (N_3053,N_2670,N_2558);
nor U3054 (N_3054,N_2848,N_2642);
or U3055 (N_3055,N_2735,N_2846);
xor U3056 (N_3056,N_2809,N_2933);
or U3057 (N_3057,N_2832,N_2575);
or U3058 (N_3058,N_2524,N_2934);
xor U3059 (N_3059,N_2585,N_2895);
nand U3060 (N_3060,N_2729,N_2574);
nand U3061 (N_3061,N_2507,N_2916);
xor U3062 (N_3062,N_2597,N_2703);
and U3063 (N_3063,N_2577,N_2738);
and U3064 (N_3064,N_2833,N_2766);
and U3065 (N_3065,N_2954,N_2822);
nor U3066 (N_3066,N_2656,N_2611);
nand U3067 (N_3067,N_2839,N_2819);
nand U3068 (N_3068,N_2551,N_2728);
or U3069 (N_3069,N_2956,N_2925);
nand U3070 (N_3070,N_2868,N_2598);
or U3071 (N_3071,N_2736,N_2869);
and U3072 (N_3072,N_2877,N_2700);
nand U3073 (N_3073,N_2570,N_2788);
nor U3074 (N_3074,N_2865,N_2704);
and U3075 (N_3075,N_2568,N_2973);
nand U3076 (N_3076,N_2658,N_2785);
and U3077 (N_3077,N_2974,N_2517);
and U3078 (N_3078,N_2560,N_2887);
or U3079 (N_3079,N_2582,N_2940);
nor U3080 (N_3080,N_2527,N_2807);
or U3081 (N_3081,N_2862,N_2756);
nand U3082 (N_3082,N_2675,N_2514);
nor U3083 (N_3083,N_2679,N_2503);
nand U3084 (N_3084,N_2993,N_2610);
nand U3085 (N_3085,N_2655,N_2907);
nand U3086 (N_3086,N_2534,N_2794);
nand U3087 (N_3087,N_2707,N_2697);
nand U3088 (N_3088,N_2924,N_2519);
and U3089 (N_3089,N_2761,N_2982);
and U3090 (N_3090,N_2999,N_2571);
nand U3091 (N_3091,N_2732,N_2684);
nor U3092 (N_3092,N_2753,N_2755);
or U3093 (N_3093,N_2837,N_2588);
nand U3094 (N_3094,N_2851,N_2844);
or U3095 (N_3095,N_2965,N_2556);
nor U3096 (N_3096,N_2826,N_2835);
nand U3097 (N_3097,N_2927,N_2538);
nor U3098 (N_3098,N_2627,N_2979);
or U3099 (N_3099,N_2946,N_2579);
nand U3100 (N_3100,N_2856,N_2501);
and U3101 (N_3101,N_2878,N_2572);
and U3102 (N_3102,N_2608,N_2918);
or U3103 (N_3103,N_2711,N_2867);
nand U3104 (N_3104,N_2789,N_2554);
and U3105 (N_3105,N_2782,N_2616);
xor U3106 (N_3106,N_2926,N_2905);
nand U3107 (N_3107,N_2516,N_2718);
or U3108 (N_3108,N_2947,N_2829);
xor U3109 (N_3109,N_2814,N_2891);
nand U3110 (N_3110,N_2623,N_2562);
nand U3111 (N_3111,N_2803,N_2589);
nand U3112 (N_3112,N_2564,N_2739);
nand U3113 (N_3113,N_2984,N_2873);
nand U3114 (N_3114,N_2692,N_2696);
or U3115 (N_3115,N_2950,N_2978);
and U3116 (N_3116,N_2830,N_2784);
xor U3117 (N_3117,N_2706,N_2719);
and U3118 (N_3118,N_2932,N_2660);
or U3119 (N_3119,N_2852,N_2906);
nor U3120 (N_3120,N_2662,N_2646);
nand U3121 (N_3121,N_2966,N_2885);
xnor U3122 (N_3122,N_2857,N_2529);
xnor U3123 (N_3123,N_2970,N_2699);
and U3124 (N_3124,N_2609,N_2651);
nand U3125 (N_3125,N_2871,N_2583);
nand U3126 (N_3126,N_2526,N_2768);
nor U3127 (N_3127,N_2855,N_2613);
or U3128 (N_3128,N_2625,N_2520);
nand U3129 (N_3129,N_2532,N_2607);
xnor U3130 (N_3130,N_2645,N_2580);
xnor U3131 (N_3131,N_2861,N_2751);
nand U3132 (N_3132,N_2995,N_2818);
and U3133 (N_3133,N_2565,N_2767);
nor U3134 (N_3134,N_2790,N_2920);
nor U3135 (N_3135,N_2624,N_2967);
nor U3136 (N_3136,N_2898,N_2687);
and U3137 (N_3137,N_2668,N_2724);
and U3138 (N_3138,N_2900,N_2883);
or U3139 (N_3139,N_2549,N_2673);
xnor U3140 (N_3140,N_2698,N_2841);
nor U3141 (N_3141,N_2716,N_2888);
or U3142 (N_3142,N_2663,N_2858);
and U3143 (N_3143,N_2632,N_2799);
and U3144 (N_3144,N_2705,N_2774);
xor U3145 (N_3145,N_2859,N_2509);
or U3146 (N_3146,N_2941,N_2720);
or U3147 (N_3147,N_2821,N_2815);
or U3148 (N_3148,N_2866,N_2875);
nand U3149 (N_3149,N_2921,N_2702);
xor U3150 (N_3150,N_2985,N_2717);
or U3151 (N_3151,N_2612,N_2665);
or U3152 (N_3152,N_2689,N_2731);
nand U3153 (N_3153,N_2930,N_2636);
nor U3154 (N_3154,N_2893,N_2827);
xor U3155 (N_3155,N_2649,N_2793);
and U3156 (N_3156,N_2850,N_2994);
nor U3157 (N_3157,N_2505,N_2701);
nand U3158 (N_3158,N_2630,N_2960);
or U3159 (N_3159,N_2886,N_2828);
or U3160 (N_3160,N_2584,N_2654);
and U3161 (N_3161,N_2688,N_2917);
nor U3162 (N_3162,N_2652,N_2838);
nor U3163 (N_3163,N_2816,N_2659);
or U3164 (N_3164,N_2639,N_2773);
nand U3165 (N_3165,N_2644,N_2544);
or U3166 (N_3166,N_2769,N_2834);
or U3167 (N_3167,N_2650,N_2929);
nand U3168 (N_3168,N_2854,N_2915);
or U3169 (N_3169,N_2606,N_2914);
nor U3170 (N_3170,N_2626,N_2777);
nand U3171 (N_3171,N_2986,N_2754);
or U3172 (N_3172,N_2964,N_2657);
xnor U3173 (N_3173,N_2845,N_2569);
nand U3174 (N_3174,N_2686,N_2762);
nand U3175 (N_3175,N_2682,N_2743);
nand U3176 (N_3176,N_2504,N_2758);
and U3177 (N_3177,N_2876,N_2931);
and U3178 (N_3178,N_2502,N_2971);
xor U3179 (N_3179,N_2776,N_2765);
nand U3180 (N_3180,N_2722,N_2555);
or U3181 (N_3181,N_2592,N_2938);
and U3182 (N_3182,N_2811,N_2801);
nor U3183 (N_3183,N_2787,N_2922);
and U3184 (N_3184,N_2667,N_2781);
nor U3185 (N_3185,N_2808,N_2889);
and U3186 (N_3186,N_2545,N_2653);
nor U3187 (N_3187,N_2935,N_2602);
nand U3188 (N_3188,N_2622,N_2770);
nand U3189 (N_3189,N_2619,N_2542);
and U3190 (N_3190,N_2923,N_2958);
nor U3191 (N_3191,N_2976,N_2694);
or U3192 (N_3192,N_2990,N_2997);
and U3193 (N_3193,N_2911,N_2587);
and U3194 (N_3194,N_2573,N_2881);
nand U3195 (N_3195,N_2615,N_2962);
xor U3196 (N_3196,N_2521,N_2725);
nand U3197 (N_3197,N_2903,N_2672);
nand U3198 (N_3198,N_2890,N_2581);
nor U3199 (N_3199,N_2548,N_2559);
nor U3200 (N_3200,N_2737,N_2952);
or U3201 (N_3201,N_2634,N_2618);
xor U3202 (N_3202,N_2631,N_2791);
xnor U3203 (N_3203,N_2771,N_2884);
nand U3204 (N_3204,N_2949,N_2961);
nand U3205 (N_3205,N_2951,N_2836);
and U3206 (N_3206,N_2714,N_2757);
nand U3207 (N_3207,N_2936,N_2948);
and U3208 (N_3208,N_2726,N_2748);
nor U3209 (N_3209,N_2648,N_2764);
or U3210 (N_3210,N_2695,N_2709);
nor U3211 (N_3211,N_2674,N_2909);
nand U3212 (N_3212,N_2937,N_2944);
nor U3213 (N_3213,N_2578,N_2989);
xnor U3214 (N_3214,N_2595,N_2817);
and U3215 (N_3215,N_2512,N_2831);
or U3216 (N_3216,N_2943,N_2510);
nand U3217 (N_3217,N_2749,N_2955);
nor U3218 (N_3218,N_2910,N_2741);
and U3219 (N_3219,N_2523,N_2953);
and U3220 (N_3220,N_2664,N_2540);
nand U3221 (N_3221,N_2531,N_2744);
nand U3222 (N_3222,N_2772,N_2879);
nor U3223 (N_3223,N_2710,N_2797);
nand U3224 (N_3224,N_2864,N_2894);
and U3225 (N_3225,N_2628,N_2805);
or U3226 (N_3226,N_2874,N_2683);
or U3227 (N_3227,N_2899,N_2860);
nand U3228 (N_3228,N_2988,N_2968);
or U3229 (N_3229,N_2760,N_2500);
xor U3230 (N_3230,N_2715,N_2880);
or U3231 (N_3231,N_2853,N_2511);
nor U3232 (N_3232,N_2552,N_2557);
and U3233 (N_3233,N_2998,N_2980);
and U3234 (N_3234,N_2977,N_2637);
nor U3235 (N_3235,N_2546,N_2561);
xnor U3236 (N_3236,N_2842,N_2567);
nand U3237 (N_3237,N_2734,N_2928);
or U3238 (N_3238,N_2528,N_2870);
and U3239 (N_3239,N_2746,N_2591);
nor U3240 (N_3240,N_2849,N_2596);
and U3241 (N_3241,N_2600,N_2897);
xnor U3242 (N_3242,N_2872,N_2681);
and U3243 (N_3243,N_2629,N_2730);
nand U3244 (N_3244,N_2638,N_2539);
and U3245 (N_3245,N_2823,N_2712);
nand U3246 (N_3246,N_2594,N_2813);
nor U3247 (N_3247,N_2693,N_2919);
and U3248 (N_3248,N_2691,N_2525);
or U3249 (N_3249,N_2783,N_2991);
nor U3250 (N_3250,N_2549,N_2760);
or U3251 (N_3251,N_2638,N_2780);
and U3252 (N_3252,N_2949,N_2909);
nor U3253 (N_3253,N_2514,N_2686);
nand U3254 (N_3254,N_2954,N_2921);
nor U3255 (N_3255,N_2800,N_2696);
nand U3256 (N_3256,N_2721,N_2645);
nand U3257 (N_3257,N_2533,N_2635);
nor U3258 (N_3258,N_2981,N_2523);
nand U3259 (N_3259,N_2551,N_2506);
nand U3260 (N_3260,N_2750,N_2771);
or U3261 (N_3261,N_2690,N_2937);
and U3262 (N_3262,N_2908,N_2633);
nor U3263 (N_3263,N_2623,N_2531);
or U3264 (N_3264,N_2972,N_2590);
and U3265 (N_3265,N_2831,N_2763);
nor U3266 (N_3266,N_2625,N_2661);
or U3267 (N_3267,N_2605,N_2953);
nand U3268 (N_3268,N_2547,N_2756);
nor U3269 (N_3269,N_2799,N_2831);
nand U3270 (N_3270,N_2821,N_2712);
nand U3271 (N_3271,N_2843,N_2709);
nor U3272 (N_3272,N_2507,N_2579);
nor U3273 (N_3273,N_2555,N_2741);
nor U3274 (N_3274,N_2789,N_2975);
nor U3275 (N_3275,N_2556,N_2670);
nand U3276 (N_3276,N_2921,N_2942);
and U3277 (N_3277,N_2964,N_2820);
nor U3278 (N_3278,N_2873,N_2979);
and U3279 (N_3279,N_2553,N_2883);
or U3280 (N_3280,N_2806,N_2840);
nor U3281 (N_3281,N_2505,N_2923);
or U3282 (N_3282,N_2805,N_2521);
or U3283 (N_3283,N_2546,N_2506);
nor U3284 (N_3284,N_2946,N_2878);
and U3285 (N_3285,N_2877,N_2996);
and U3286 (N_3286,N_2703,N_2866);
xor U3287 (N_3287,N_2800,N_2804);
and U3288 (N_3288,N_2789,N_2548);
and U3289 (N_3289,N_2580,N_2632);
or U3290 (N_3290,N_2911,N_2846);
and U3291 (N_3291,N_2592,N_2613);
xnor U3292 (N_3292,N_2542,N_2857);
nand U3293 (N_3293,N_2698,N_2939);
or U3294 (N_3294,N_2654,N_2515);
or U3295 (N_3295,N_2987,N_2514);
or U3296 (N_3296,N_2659,N_2955);
or U3297 (N_3297,N_2573,N_2765);
or U3298 (N_3298,N_2594,N_2635);
and U3299 (N_3299,N_2558,N_2973);
nand U3300 (N_3300,N_2960,N_2728);
nor U3301 (N_3301,N_2788,N_2524);
nand U3302 (N_3302,N_2719,N_2644);
and U3303 (N_3303,N_2760,N_2755);
or U3304 (N_3304,N_2745,N_2873);
or U3305 (N_3305,N_2985,N_2981);
nor U3306 (N_3306,N_2984,N_2610);
nand U3307 (N_3307,N_2903,N_2951);
xor U3308 (N_3308,N_2934,N_2612);
and U3309 (N_3309,N_2902,N_2783);
nor U3310 (N_3310,N_2820,N_2693);
nor U3311 (N_3311,N_2762,N_2821);
nand U3312 (N_3312,N_2563,N_2965);
and U3313 (N_3313,N_2967,N_2905);
nor U3314 (N_3314,N_2967,N_2769);
and U3315 (N_3315,N_2610,N_2709);
xor U3316 (N_3316,N_2990,N_2871);
nand U3317 (N_3317,N_2937,N_2521);
nand U3318 (N_3318,N_2702,N_2884);
nor U3319 (N_3319,N_2856,N_2899);
nor U3320 (N_3320,N_2921,N_2537);
nand U3321 (N_3321,N_2540,N_2824);
nor U3322 (N_3322,N_2575,N_2672);
nand U3323 (N_3323,N_2701,N_2766);
or U3324 (N_3324,N_2966,N_2733);
or U3325 (N_3325,N_2781,N_2991);
xor U3326 (N_3326,N_2990,N_2730);
and U3327 (N_3327,N_2933,N_2781);
nand U3328 (N_3328,N_2566,N_2551);
and U3329 (N_3329,N_2855,N_2950);
or U3330 (N_3330,N_2853,N_2616);
or U3331 (N_3331,N_2618,N_2932);
or U3332 (N_3332,N_2963,N_2678);
xor U3333 (N_3333,N_2845,N_2811);
or U3334 (N_3334,N_2672,N_2840);
nor U3335 (N_3335,N_2875,N_2547);
and U3336 (N_3336,N_2531,N_2839);
and U3337 (N_3337,N_2995,N_2996);
or U3338 (N_3338,N_2548,N_2621);
nor U3339 (N_3339,N_2556,N_2976);
nor U3340 (N_3340,N_2819,N_2537);
nand U3341 (N_3341,N_2760,N_2509);
and U3342 (N_3342,N_2879,N_2831);
nor U3343 (N_3343,N_2889,N_2679);
or U3344 (N_3344,N_2535,N_2869);
and U3345 (N_3345,N_2763,N_2866);
or U3346 (N_3346,N_2924,N_2704);
or U3347 (N_3347,N_2687,N_2764);
and U3348 (N_3348,N_2526,N_2812);
and U3349 (N_3349,N_2861,N_2919);
nand U3350 (N_3350,N_2831,N_2736);
nor U3351 (N_3351,N_2765,N_2504);
nor U3352 (N_3352,N_2512,N_2716);
nand U3353 (N_3353,N_2525,N_2997);
and U3354 (N_3354,N_2846,N_2816);
nand U3355 (N_3355,N_2968,N_2928);
nor U3356 (N_3356,N_2713,N_2517);
and U3357 (N_3357,N_2920,N_2800);
nand U3358 (N_3358,N_2958,N_2557);
nand U3359 (N_3359,N_2851,N_2657);
or U3360 (N_3360,N_2833,N_2755);
and U3361 (N_3361,N_2978,N_2666);
or U3362 (N_3362,N_2830,N_2941);
nand U3363 (N_3363,N_2858,N_2701);
or U3364 (N_3364,N_2712,N_2737);
or U3365 (N_3365,N_2537,N_2742);
and U3366 (N_3366,N_2788,N_2964);
and U3367 (N_3367,N_2893,N_2906);
xnor U3368 (N_3368,N_2688,N_2928);
or U3369 (N_3369,N_2517,N_2545);
nor U3370 (N_3370,N_2873,N_2803);
or U3371 (N_3371,N_2542,N_2972);
or U3372 (N_3372,N_2589,N_2839);
and U3373 (N_3373,N_2787,N_2902);
nand U3374 (N_3374,N_2535,N_2992);
and U3375 (N_3375,N_2646,N_2508);
or U3376 (N_3376,N_2567,N_2604);
and U3377 (N_3377,N_2627,N_2621);
nand U3378 (N_3378,N_2714,N_2755);
nand U3379 (N_3379,N_2707,N_2742);
nand U3380 (N_3380,N_2902,N_2574);
nand U3381 (N_3381,N_2512,N_2933);
nor U3382 (N_3382,N_2983,N_2994);
nand U3383 (N_3383,N_2697,N_2770);
and U3384 (N_3384,N_2650,N_2958);
or U3385 (N_3385,N_2617,N_2757);
nand U3386 (N_3386,N_2920,N_2601);
nor U3387 (N_3387,N_2765,N_2741);
and U3388 (N_3388,N_2780,N_2618);
nand U3389 (N_3389,N_2867,N_2717);
or U3390 (N_3390,N_2503,N_2934);
and U3391 (N_3391,N_2852,N_2929);
and U3392 (N_3392,N_2587,N_2703);
or U3393 (N_3393,N_2625,N_2802);
or U3394 (N_3394,N_2953,N_2902);
nor U3395 (N_3395,N_2994,N_2737);
or U3396 (N_3396,N_2835,N_2704);
nor U3397 (N_3397,N_2573,N_2850);
nand U3398 (N_3398,N_2579,N_2656);
or U3399 (N_3399,N_2979,N_2765);
nand U3400 (N_3400,N_2904,N_2985);
and U3401 (N_3401,N_2608,N_2692);
or U3402 (N_3402,N_2796,N_2886);
nor U3403 (N_3403,N_2709,N_2639);
and U3404 (N_3404,N_2797,N_2753);
and U3405 (N_3405,N_2552,N_2988);
and U3406 (N_3406,N_2873,N_2587);
nand U3407 (N_3407,N_2984,N_2722);
xnor U3408 (N_3408,N_2834,N_2845);
and U3409 (N_3409,N_2541,N_2531);
or U3410 (N_3410,N_2618,N_2803);
nor U3411 (N_3411,N_2767,N_2852);
or U3412 (N_3412,N_2820,N_2661);
and U3413 (N_3413,N_2946,N_2629);
and U3414 (N_3414,N_2672,N_2555);
nand U3415 (N_3415,N_2537,N_2572);
nand U3416 (N_3416,N_2814,N_2816);
and U3417 (N_3417,N_2983,N_2731);
and U3418 (N_3418,N_2828,N_2747);
nand U3419 (N_3419,N_2944,N_2504);
nor U3420 (N_3420,N_2532,N_2667);
and U3421 (N_3421,N_2640,N_2943);
nor U3422 (N_3422,N_2602,N_2688);
and U3423 (N_3423,N_2750,N_2704);
and U3424 (N_3424,N_2509,N_2715);
or U3425 (N_3425,N_2662,N_2621);
and U3426 (N_3426,N_2590,N_2955);
and U3427 (N_3427,N_2500,N_2576);
xor U3428 (N_3428,N_2918,N_2803);
and U3429 (N_3429,N_2969,N_2926);
nand U3430 (N_3430,N_2941,N_2852);
or U3431 (N_3431,N_2565,N_2546);
and U3432 (N_3432,N_2674,N_2747);
nand U3433 (N_3433,N_2805,N_2825);
xnor U3434 (N_3434,N_2719,N_2825);
or U3435 (N_3435,N_2760,N_2646);
and U3436 (N_3436,N_2721,N_2915);
xor U3437 (N_3437,N_2872,N_2965);
and U3438 (N_3438,N_2750,N_2970);
xnor U3439 (N_3439,N_2735,N_2864);
or U3440 (N_3440,N_2915,N_2929);
or U3441 (N_3441,N_2530,N_2740);
nor U3442 (N_3442,N_2818,N_2898);
nor U3443 (N_3443,N_2943,N_2674);
nand U3444 (N_3444,N_2623,N_2815);
nand U3445 (N_3445,N_2685,N_2894);
and U3446 (N_3446,N_2821,N_2811);
nor U3447 (N_3447,N_2872,N_2570);
nand U3448 (N_3448,N_2829,N_2695);
and U3449 (N_3449,N_2985,N_2744);
nor U3450 (N_3450,N_2538,N_2554);
nand U3451 (N_3451,N_2996,N_2884);
and U3452 (N_3452,N_2767,N_2636);
or U3453 (N_3453,N_2804,N_2585);
nor U3454 (N_3454,N_2526,N_2530);
xnor U3455 (N_3455,N_2646,N_2572);
or U3456 (N_3456,N_2642,N_2742);
and U3457 (N_3457,N_2674,N_2502);
nand U3458 (N_3458,N_2626,N_2746);
xnor U3459 (N_3459,N_2525,N_2752);
and U3460 (N_3460,N_2997,N_2797);
and U3461 (N_3461,N_2896,N_2567);
xnor U3462 (N_3462,N_2635,N_2994);
nand U3463 (N_3463,N_2623,N_2841);
and U3464 (N_3464,N_2689,N_2545);
nor U3465 (N_3465,N_2530,N_2644);
nand U3466 (N_3466,N_2529,N_2786);
nor U3467 (N_3467,N_2948,N_2924);
nor U3468 (N_3468,N_2899,N_2871);
xnor U3469 (N_3469,N_2584,N_2649);
nand U3470 (N_3470,N_2828,N_2603);
xor U3471 (N_3471,N_2561,N_2689);
or U3472 (N_3472,N_2848,N_2831);
xor U3473 (N_3473,N_2934,N_2796);
nand U3474 (N_3474,N_2636,N_2799);
and U3475 (N_3475,N_2856,N_2757);
nor U3476 (N_3476,N_2945,N_2880);
nand U3477 (N_3477,N_2789,N_2541);
nand U3478 (N_3478,N_2645,N_2902);
or U3479 (N_3479,N_2561,N_2647);
or U3480 (N_3480,N_2653,N_2667);
or U3481 (N_3481,N_2982,N_2560);
or U3482 (N_3482,N_2587,N_2846);
and U3483 (N_3483,N_2586,N_2700);
and U3484 (N_3484,N_2759,N_2830);
nand U3485 (N_3485,N_2742,N_2872);
nor U3486 (N_3486,N_2928,N_2831);
nor U3487 (N_3487,N_2554,N_2994);
nor U3488 (N_3488,N_2636,N_2775);
or U3489 (N_3489,N_2722,N_2686);
nand U3490 (N_3490,N_2872,N_2637);
nand U3491 (N_3491,N_2986,N_2971);
nor U3492 (N_3492,N_2866,N_2594);
and U3493 (N_3493,N_2898,N_2993);
nor U3494 (N_3494,N_2966,N_2621);
nor U3495 (N_3495,N_2899,N_2925);
nand U3496 (N_3496,N_2536,N_2795);
nor U3497 (N_3497,N_2719,N_2586);
or U3498 (N_3498,N_2793,N_2885);
nand U3499 (N_3499,N_2807,N_2994);
nor U3500 (N_3500,N_3110,N_3058);
nand U3501 (N_3501,N_3098,N_3106);
and U3502 (N_3502,N_3228,N_3488);
and U3503 (N_3503,N_3116,N_3401);
or U3504 (N_3504,N_3236,N_3458);
or U3505 (N_3505,N_3171,N_3479);
or U3506 (N_3506,N_3427,N_3043);
or U3507 (N_3507,N_3444,N_3338);
nor U3508 (N_3508,N_3426,N_3237);
xor U3509 (N_3509,N_3068,N_3341);
nor U3510 (N_3510,N_3349,N_3142);
or U3511 (N_3511,N_3096,N_3254);
or U3512 (N_3512,N_3198,N_3261);
or U3513 (N_3513,N_3232,N_3084);
and U3514 (N_3514,N_3468,N_3118);
nor U3515 (N_3515,N_3003,N_3137);
nand U3516 (N_3516,N_3248,N_3157);
and U3517 (N_3517,N_3387,N_3329);
and U3518 (N_3518,N_3327,N_3051);
or U3519 (N_3519,N_3060,N_3105);
xnor U3520 (N_3520,N_3224,N_3460);
nor U3521 (N_3521,N_3423,N_3080);
nand U3522 (N_3522,N_3326,N_3112);
and U3523 (N_3523,N_3487,N_3364);
and U3524 (N_3524,N_3025,N_3324);
nor U3525 (N_3525,N_3282,N_3223);
nand U3526 (N_3526,N_3378,N_3314);
or U3527 (N_3527,N_3195,N_3109);
xor U3528 (N_3528,N_3410,N_3264);
nor U3529 (N_3529,N_3303,N_3465);
nor U3530 (N_3530,N_3477,N_3081);
nand U3531 (N_3531,N_3049,N_3186);
and U3532 (N_3532,N_3192,N_3312);
nand U3533 (N_3533,N_3161,N_3104);
nor U3534 (N_3534,N_3339,N_3055);
or U3535 (N_3535,N_3015,N_3222);
xnor U3536 (N_3536,N_3094,N_3021);
nor U3537 (N_3537,N_3149,N_3200);
and U3538 (N_3538,N_3193,N_3010);
or U3539 (N_3539,N_3474,N_3197);
and U3540 (N_3540,N_3485,N_3188);
nand U3541 (N_3541,N_3076,N_3047);
nor U3542 (N_3542,N_3139,N_3185);
nor U3543 (N_3543,N_3159,N_3181);
nand U3544 (N_3544,N_3221,N_3226);
nor U3545 (N_3545,N_3062,N_3398);
and U3546 (N_3546,N_3136,N_3033);
nor U3547 (N_3547,N_3455,N_3376);
nand U3548 (N_3548,N_3438,N_3344);
nand U3549 (N_3549,N_3187,N_3108);
and U3550 (N_3550,N_3151,N_3361);
or U3551 (N_3551,N_3160,N_3127);
or U3552 (N_3552,N_3234,N_3220);
nor U3553 (N_3553,N_3309,N_3391);
nand U3554 (N_3554,N_3004,N_3417);
or U3555 (N_3555,N_3050,N_3090);
or U3556 (N_3556,N_3267,N_3173);
nand U3557 (N_3557,N_3399,N_3331);
nor U3558 (N_3558,N_3300,N_3172);
nor U3559 (N_3559,N_3238,N_3183);
and U3560 (N_3560,N_3233,N_3208);
or U3561 (N_3561,N_3184,N_3352);
nand U3562 (N_3562,N_3253,N_3362);
nand U3563 (N_3563,N_3143,N_3163);
nand U3564 (N_3564,N_3001,N_3346);
or U3565 (N_3565,N_3075,N_3394);
xor U3566 (N_3566,N_3245,N_3316);
nor U3567 (N_3567,N_3054,N_3340);
nand U3568 (N_3568,N_3283,N_3380);
nor U3569 (N_3569,N_3088,N_3069);
and U3570 (N_3570,N_3202,N_3227);
and U3571 (N_3571,N_3445,N_3356);
or U3572 (N_3572,N_3421,N_3247);
and U3573 (N_3573,N_3345,N_3476);
nor U3574 (N_3574,N_3271,N_3342);
nand U3575 (N_3575,N_3408,N_3250);
nor U3576 (N_3576,N_3099,N_3373);
or U3577 (N_3577,N_3306,N_3384);
nor U3578 (N_3578,N_3379,N_3463);
or U3579 (N_3579,N_3168,N_3420);
nor U3580 (N_3580,N_3443,N_3319);
or U3581 (N_3581,N_3404,N_3041);
nor U3582 (N_3582,N_3432,N_3070);
or U3583 (N_3583,N_3255,N_3424);
nand U3584 (N_3584,N_3360,N_3291);
or U3585 (N_3585,N_3037,N_3419);
nand U3586 (N_3586,N_3257,N_3241);
nand U3587 (N_3587,N_3495,N_3467);
nand U3588 (N_3588,N_3019,N_3353);
nor U3589 (N_3589,N_3056,N_3484);
nand U3590 (N_3590,N_3201,N_3311);
and U3591 (N_3591,N_3175,N_3144);
nor U3592 (N_3592,N_3447,N_3170);
nor U3593 (N_3593,N_3497,N_3411);
nand U3594 (N_3594,N_3194,N_3006);
and U3595 (N_3595,N_3454,N_3252);
nor U3596 (N_3596,N_3385,N_3020);
xor U3597 (N_3597,N_3461,N_3328);
or U3598 (N_3598,N_3397,N_3335);
or U3599 (N_3599,N_3087,N_3013);
or U3600 (N_3600,N_3138,N_3350);
and U3601 (N_3601,N_3211,N_3292);
or U3602 (N_3602,N_3403,N_3017);
or U3603 (N_3603,N_3150,N_3266);
nor U3604 (N_3604,N_3035,N_3322);
or U3605 (N_3605,N_3048,N_3207);
and U3606 (N_3606,N_3190,N_3370);
or U3607 (N_3607,N_3204,N_3383);
nand U3608 (N_3608,N_3024,N_3162);
or U3609 (N_3609,N_3212,N_3442);
nor U3610 (N_3610,N_3066,N_3196);
or U3611 (N_3611,N_3005,N_3493);
and U3612 (N_3612,N_3242,N_3141);
or U3613 (N_3613,N_3028,N_3158);
nor U3614 (N_3614,N_3434,N_3274);
nor U3615 (N_3615,N_3128,N_3030);
or U3616 (N_3616,N_3293,N_3124);
nor U3617 (N_3617,N_3453,N_3176);
and U3618 (N_3618,N_3012,N_3011);
xnor U3619 (N_3619,N_3085,N_3435);
and U3620 (N_3620,N_3036,N_3456);
nor U3621 (N_3621,N_3365,N_3336);
nand U3622 (N_3622,N_3032,N_3416);
xor U3623 (N_3623,N_3466,N_3273);
nor U3624 (N_3624,N_3103,N_3215);
and U3625 (N_3625,N_3262,N_3289);
or U3626 (N_3626,N_3126,N_3179);
nand U3627 (N_3627,N_3483,N_3014);
or U3628 (N_3628,N_3489,N_3371);
nor U3629 (N_3629,N_3083,N_3079);
or U3630 (N_3630,N_3229,N_3459);
xnor U3631 (N_3631,N_3061,N_3074);
nand U3632 (N_3632,N_3486,N_3270);
nor U3633 (N_3633,N_3042,N_3122);
or U3634 (N_3634,N_3205,N_3097);
or U3635 (N_3635,N_3225,N_3167);
and U3636 (N_3636,N_3462,N_3480);
or U3637 (N_3637,N_3147,N_3357);
nand U3638 (N_3638,N_3372,N_3431);
and U3639 (N_3639,N_3114,N_3191);
nand U3640 (N_3640,N_3287,N_3498);
xnor U3641 (N_3641,N_3057,N_3433);
xnor U3642 (N_3642,N_3165,N_3089);
nand U3643 (N_3643,N_3016,N_3246);
nor U3644 (N_3644,N_3240,N_3132);
nor U3645 (N_3645,N_3217,N_3490);
xor U3646 (N_3646,N_3276,N_3153);
nand U3647 (N_3647,N_3308,N_3077);
xor U3648 (N_3648,N_3405,N_3382);
or U3649 (N_3649,N_3140,N_3148);
xnor U3650 (N_3650,N_3354,N_3482);
or U3651 (N_3651,N_3156,N_3359);
and U3652 (N_3652,N_3235,N_3279);
or U3653 (N_3653,N_3491,N_3072);
xnor U3654 (N_3654,N_3164,N_3386);
and U3655 (N_3655,N_3304,N_3064);
or U3656 (N_3656,N_3392,N_3121);
or U3657 (N_3657,N_3358,N_3218);
nor U3658 (N_3658,N_3281,N_3259);
and U3659 (N_3659,N_3374,N_3430);
nand U3660 (N_3660,N_3120,N_3101);
and U3661 (N_3661,N_3294,N_3154);
nor U3662 (N_3662,N_3332,N_3366);
nand U3663 (N_3663,N_3038,N_3189);
nor U3664 (N_3664,N_3313,N_3395);
xnor U3665 (N_3665,N_3134,N_3451);
and U3666 (N_3666,N_3214,N_3368);
nand U3667 (N_3667,N_3039,N_3310);
nor U3668 (N_3668,N_3166,N_3067);
or U3669 (N_3669,N_3330,N_3268);
or U3670 (N_3670,N_3470,N_3182);
nand U3671 (N_3671,N_3251,N_3305);
nand U3672 (N_3672,N_3412,N_3146);
or U3673 (N_3673,N_3478,N_3422);
nand U3674 (N_3674,N_3078,N_3402);
and U3675 (N_3675,N_3249,N_3135);
and U3676 (N_3676,N_3206,N_3073);
nand U3677 (N_3677,N_3496,N_3317);
and U3678 (N_3678,N_3063,N_3230);
nor U3679 (N_3679,N_3469,N_3355);
nor U3680 (N_3680,N_3007,N_3428);
or U3681 (N_3681,N_3439,N_3113);
and U3682 (N_3682,N_3026,N_3290);
and U3683 (N_3683,N_3034,N_3213);
or U3684 (N_3684,N_3130,N_3333);
nor U3685 (N_3685,N_3231,N_3278);
nor U3686 (N_3686,N_3334,N_3133);
or U3687 (N_3687,N_3337,N_3446);
or U3688 (N_3688,N_3301,N_3390);
and U3689 (N_3689,N_3095,N_3022);
xnor U3690 (N_3690,N_3369,N_3053);
nand U3691 (N_3691,N_3436,N_3396);
or U3692 (N_3692,N_3473,N_3448);
nor U3693 (N_3693,N_3044,N_3320);
nor U3694 (N_3694,N_3351,N_3244);
nor U3695 (N_3695,N_3272,N_3377);
and U3696 (N_3696,N_3343,N_3307);
nor U3697 (N_3697,N_3256,N_3288);
xor U3698 (N_3698,N_3027,N_3023);
nand U3699 (N_3699,N_3131,N_3449);
xor U3700 (N_3700,N_3409,N_3177);
and U3701 (N_3701,N_3029,N_3180);
or U3702 (N_3702,N_3002,N_3123);
nand U3703 (N_3703,N_3243,N_3111);
nor U3704 (N_3704,N_3275,N_3031);
nand U3705 (N_3705,N_3302,N_3009);
xnor U3706 (N_3706,N_3318,N_3429);
and U3707 (N_3707,N_3492,N_3375);
or U3708 (N_3708,N_3415,N_3046);
or U3709 (N_3709,N_3125,N_3152);
xnor U3710 (N_3710,N_3155,N_3315);
nand U3711 (N_3711,N_3363,N_3296);
xnor U3712 (N_3712,N_3381,N_3457);
nor U3713 (N_3713,N_3102,N_3100);
and U3714 (N_3714,N_3092,N_3440);
and U3715 (N_3715,N_3000,N_3239);
and U3716 (N_3716,N_3117,N_3414);
nor U3717 (N_3717,N_3284,N_3219);
or U3718 (N_3718,N_3472,N_3286);
nand U3719 (N_3719,N_3425,N_3107);
or U3720 (N_3720,N_3052,N_3299);
and U3721 (N_3721,N_3119,N_3367);
and U3722 (N_3722,N_3325,N_3040);
and U3723 (N_3723,N_3169,N_3086);
and U3724 (N_3724,N_3263,N_3413);
nor U3725 (N_3725,N_3091,N_3494);
xnor U3726 (N_3726,N_3285,N_3203);
xnor U3727 (N_3727,N_3209,N_3348);
xor U3728 (N_3728,N_3059,N_3323);
and U3729 (N_3729,N_3045,N_3297);
and U3730 (N_3730,N_3216,N_3321);
nor U3731 (N_3731,N_3178,N_3277);
nor U3732 (N_3732,N_3093,N_3008);
nor U3733 (N_3733,N_3407,N_3260);
or U3734 (N_3734,N_3452,N_3471);
or U3735 (N_3735,N_3441,N_3258);
nor U3736 (N_3736,N_3210,N_3418);
nand U3737 (N_3737,N_3071,N_3145);
or U3738 (N_3738,N_3388,N_3199);
xor U3739 (N_3739,N_3464,N_3389);
or U3740 (N_3740,N_3082,N_3018);
nand U3741 (N_3741,N_3265,N_3347);
and U3742 (N_3742,N_3393,N_3298);
and U3743 (N_3743,N_3295,N_3450);
or U3744 (N_3744,N_3475,N_3269);
nor U3745 (N_3745,N_3280,N_3129);
and U3746 (N_3746,N_3115,N_3174);
xor U3747 (N_3747,N_3065,N_3437);
nor U3748 (N_3748,N_3406,N_3481);
nand U3749 (N_3749,N_3400,N_3499);
and U3750 (N_3750,N_3050,N_3081);
and U3751 (N_3751,N_3157,N_3163);
nand U3752 (N_3752,N_3304,N_3441);
nand U3753 (N_3753,N_3438,N_3425);
or U3754 (N_3754,N_3424,N_3174);
nor U3755 (N_3755,N_3151,N_3001);
nor U3756 (N_3756,N_3060,N_3126);
nand U3757 (N_3757,N_3313,N_3373);
nor U3758 (N_3758,N_3199,N_3414);
and U3759 (N_3759,N_3449,N_3239);
and U3760 (N_3760,N_3084,N_3370);
xnor U3761 (N_3761,N_3437,N_3391);
and U3762 (N_3762,N_3474,N_3216);
and U3763 (N_3763,N_3428,N_3236);
or U3764 (N_3764,N_3479,N_3038);
nor U3765 (N_3765,N_3118,N_3307);
or U3766 (N_3766,N_3487,N_3194);
nor U3767 (N_3767,N_3391,N_3319);
and U3768 (N_3768,N_3018,N_3414);
and U3769 (N_3769,N_3125,N_3046);
or U3770 (N_3770,N_3064,N_3300);
nor U3771 (N_3771,N_3132,N_3176);
nand U3772 (N_3772,N_3276,N_3198);
nor U3773 (N_3773,N_3093,N_3319);
or U3774 (N_3774,N_3364,N_3174);
and U3775 (N_3775,N_3463,N_3421);
or U3776 (N_3776,N_3089,N_3484);
and U3777 (N_3777,N_3047,N_3475);
and U3778 (N_3778,N_3481,N_3055);
or U3779 (N_3779,N_3263,N_3127);
or U3780 (N_3780,N_3320,N_3110);
nand U3781 (N_3781,N_3224,N_3336);
or U3782 (N_3782,N_3232,N_3049);
nand U3783 (N_3783,N_3276,N_3190);
nor U3784 (N_3784,N_3312,N_3329);
nand U3785 (N_3785,N_3397,N_3261);
nand U3786 (N_3786,N_3030,N_3255);
nand U3787 (N_3787,N_3000,N_3245);
nor U3788 (N_3788,N_3334,N_3181);
nor U3789 (N_3789,N_3087,N_3214);
nor U3790 (N_3790,N_3454,N_3103);
and U3791 (N_3791,N_3115,N_3041);
or U3792 (N_3792,N_3033,N_3059);
nand U3793 (N_3793,N_3254,N_3196);
and U3794 (N_3794,N_3405,N_3067);
nand U3795 (N_3795,N_3429,N_3116);
or U3796 (N_3796,N_3441,N_3048);
xnor U3797 (N_3797,N_3425,N_3137);
nand U3798 (N_3798,N_3064,N_3109);
xor U3799 (N_3799,N_3078,N_3186);
nor U3800 (N_3800,N_3103,N_3330);
xnor U3801 (N_3801,N_3330,N_3328);
and U3802 (N_3802,N_3135,N_3459);
or U3803 (N_3803,N_3437,N_3097);
nor U3804 (N_3804,N_3397,N_3040);
or U3805 (N_3805,N_3312,N_3241);
nand U3806 (N_3806,N_3036,N_3134);
nand U3807 (N_3807,N_3228,N_3030);
nor U3808 (N_3808,N_3026,N_3279);
or U3809 (N_3809,N_3252,N_3070);
and U3810 (N_3810,N_3337,N_3251);
or U3811 (N_3811,N_3404,N_3075);
xnor U3812 (N_3812,N_3442,N_3431);
or U3813 (N_3813,N_3127,N_3444);
nor U3814 (N_3814,N_3403,N_3299);
and U3815 (N_3815,N_3105,N_3309);
nand U3816 (N_3816,N_3080,N_3445);
nand U3817 (N_3817,N_3477,N_3383);
nand U3818 (N_3818,N_3168,N_3441);
and U3819 (N_3819,N_3079,N_3009);
or U3820 (N_3820,N_3083,N_3008);
or U3821 (N_3821,N_3273,N_3437);
nor U3822 (N_3822,N_3357,N_3292);
nand U3823 (N_3823,N_3362,N_3421);
and U3824 (N_3824,N_3073,N_3261);
or U3825 (N_3825,N_3187,N_3235);
and U3826 (N_3826,N_3405,N_3132);
nor U3827 (N_3827,N_3302,N_3353);
nor U3828 (N_3828,N_3101,N_3303);
nand U3829 (N_3829,N_3014,N_3120);
nand U3830 (N_3830,N_3109,N_3181);
nor U3831 (N_3831,N_3421,N_3470);
nand U3832 (N_3832,N_3156,N_3390);
nor U3833 (N_3833,N_3098,N_3462);
nor U3834 (N_3834,N_3218,N_3259);
nor U3835 (N_3835,N_3345,N_3313);
and U3836 (N_3836,N_3436,N_3223);
or U3837 (N_3837,N_3496,N_3144);
or U3838 (N_3838,N_3447,N_3129);
or U3839 (N_3839,N_3210,N_3388);
xor U3840 (N_3840,N_3230,N_3259);
nor U3841 (N_3841,N_3384,N_3187);
xnor U3842 (N_3842,N_3067,N_3424);
nand U3843 (N_3843,N_3452,N_3164);
and U3844 (N_3844,N_3430,N_3283);
nor U3845 (N_3845,N_3094,N_3210);
or U3846 (N_3846,N_3071,N_3383);
nor U3847 (N_3847,N_3099,N_3228);
nor U3848 (N_3848,N_3136,N_3005);
and U3849 (N_3849,N_3339,N_3278);
or U3850 (N_3850,N_3487,N_3241);
or U3851 (N_3851,N_3309,N_3015);
or U3852 (N_3852,N_3375,N_3441);
and U3853 (N_3853,N_3422,N_3434);
nand U3854 (N_3854,N_3338,N_3252);
or U3855 (N_3855,N_3142,N_3210);
xor U3856 (N_3856,N_3199,N_3280);
or U3857 (N_3857,N_3077,N_3339);
nor U3858 (N_3858,N_3181,N_3483);
nor U3859 (N_3859,N_3014,N_3400);
nand U3860 (N_3860,N_3385,N_3003);
and U3861 (N_3861,N_3214,N_3104);
nand U3862 (N_3862,N_3451,N_3194);
nor U3863 (N_3863,N_3172,N_3180);
nand U3864 (N_3864,N_3059,N_3418);
and U3865 (N_3865,N_3408,N_3285);
and U3866 (N_3866,N_3493,N_3026);
nor U3867 (N_3867,N_3337,N_3381);
xnor U3868 (N_3868,N_3209,N_3428);
and U3869 (N_3869,N_3246,N_3125);
xnor U3870 (N_3870,N_3153,N_3306);
nor U3871 (N_3871,N_3438,N_3108);
or U3872 (N_3872,N_3071,N_3093);
nand U3873 (N_3873,N_3040,N_3305);
and U3874 (N_3874,N_3396,N_3292);
xnor U3875 (N_3875,N_3273,N_3255);
and U3876 (N_3876,N_3351,N_3319);
nor U3877 (N_3877,N_3490,N_3316);
or U3878 (N_3878,N_3355,N_3295);
nor U3879 (N_3879,N_3234,N_3160);
nand U3880 (N_3880,N_3094,N_3405);
and U3881 (N_3881,N_3449,N_3011);
or U3882 (N_3882,N_3050,N_3123);
and U3883 (N_3883,N_3309,N_3041);
xnor U3884 (N_3884,N_3200,N_3333);
or U3885 (N_3885,N_3180,N_3155);
nor U3886 (N_3886,N_3477,N_3220);
nand U3887 (N_3887,N_3319,N_3348);
nor U3888 (N_3888,N_3157,N_3097);
or U3889 (N_3889,N_3244,N_3197);
or U3890 (N_3890,N_3012,N_3495);
or U3891 (N_3891,N_3170,N_3463);
nor U3892 (N_3892,N_3498,N_3199);
nand U3893 (N_3893,N_3318,N_3146);
nor U3894 (N_3894,N_3350,N_3422);
nor U3895 (N_3895,N_3013,N_3335);
and U3896 (N_3896,N_3406,N_3444);
or U3897 (N_3897,N_3468,N_3398);
and U3898 (N_3898,N_3485,N_3313);
or U3899 (N_3899,N_3240,N_3146);
nand U3900 (N_3900,N_3186,N_3220);
nor U3901 (N_3901,N_3238,N_3258);
and U3902 (N_3902,N_3224,N_3498);
and U3903 (N_3903,N_3426,N_3069);
nand U3904 (N_3904,N_3037,N_3241);
and U3905 (N_3905,N_3148,N_3423);
or U3906 (N_3906,N_3364,N_3269);
and U3907 (N_3907,N_3195,N_3104);
or U3908 (N_3908,N_3366,N_3164);
and U3909 (N_3909,N_3321,N_3030);
and U3910 (N_3910,N_3190,N_3430);
and U3911 (N_3911,N_3475,N_3318);
or U3912 (N_3912,N_3082,N_3478);
and U3913 (N_3913,N_3116,N_3373);
nor U3914 (N_3914,N_3077,N_3447);
xor U3915 (N_3915,N_3188,N_3169);
nor U3916 (N_3916,N_3086,N_3084);
nor U3917 (N_3917,N_3172,N_3163);
or U3918 (N_3918,N_3184,N_3442);
or U3919 (N_3919,N_3042,N_3471);
nand U3920 (N_3920,N_3306,N_3430);
nor U3921 (N_3921,N_3275,N_3014);
or U3922 (N_3922,N_3084,N_3153);
or U3923 (N_3923,N_3466,N_3033);
xnor U3924 (N_3924,N_3157,N_3394);
nand U3925 (N_3925,N_3411,N_3223);
nor U3926 (N_3926,N_3253,N_3461);
and U3927 (N_3927,N_3230,N_3228);
xor U3928 (N_3928,N_3245,N_3093);
nand U3929 (N_3929,N_3339,N_3380);
xnor U3930 (N_3930,N_3051,N_3388);
and U3931 (N_3931,N_3047,N_3234);
and U3932 (N_3932,N_3116,N_3363);
or U3933 (N_3933,N_3071,N_3207);
nor U3934 (N_3934,N_3394,N_3242);
nor U3935 (N_3935,N_3413,N_3091);
and U3936 (N_3936,N_3004,N_3007);
and U3937 (N_3937,N_3452,N_3255);
or U3938 (N_3938,N_3496,N_3018);
and U3939 (N_3939,N_3140,N_3164);
or U3940 (N_3940,N_3433,N_3379);
or U3941 (N_3941,N_3243,N_3317);
nand U3942 (N_3942,N_3471,N_3362);
nand U3943 (N_3943,N_3091,N_3353);
xnor U3944 (N_3944,N_3188,N_3033);
nor U3945 (N_3945,N_3318,N_3440);
nor U3946 (N_3946,N_3127,N_3065);
and U3947 (N_3947,N_3179,N_3272);
nand U3948 (N_3948,N_3387,N_3124);
and U3949 (N_3949,N_3414,N_3119);
nand U3950 (N_3950,N_3212,N_3263);
or U3951 (N_3951,N_3196,N_3139);
xor U3952 (N_3952,N_3226,N_3281);
nor U3953 (N_3953,N_3211,N_3296);
nand U3954 (N_3954,N_3215,N_3180);
xor U3955 (N_3955,N_3178,N_3067);
nand U3956 (N_3956,N_3451,N_3322);
xor U3957 (N_3957,N_3434,N_3398);
nor U3958 (N_3958,N_3172,N_3446);
nand U3959 (N_3959,N_3073,N_3083);
nor U3960 (N_3960,N_3090,N_3457);
nor U3961 (N_3961,N_3121,N_3185);
or U3962 (N_3962,N_3419,N_3408);
nor U3963 (N_3963,N_3011,N_3094);
nand U3964 (N_3964,N_3323,N_3245);
nor U3965 (N_3965,N_3312,N_3327);
and U3966 (N_3966,N_3284,N_3475);
and U3967 (N_3967,N_3206,N_3373);
nor U3968 (N_3968,N_3248,N_3043);
nand U3969 (N_3969,N_3000,N_3218);
and U3970 (N_3970,N_3075,N_3430);
and U3971 (N_3971,N_3443,N_3000);
nor U3972 (N_3972,N_3040,N_3144);
xor U3973 (N_3973,N_3310,N_3041);
nand U3974 (N_3974,N_3435,N_3076);
and U3975 (N_3975,N_3031,N_3038);
nand U3976 (N_3976,N_3071,N_3485);
xnor U3977 (N_3977,N_3466,N_3282);
or U3978 (N_3978,N_3236,N_3476);
nand U3979 (N_3979,N_3297,N_3494);
nor U3980 (N_3980,N_3136,N_3472);
or U3981 (N_3981,N_3172,N_3273);
nor U3982 (N_3982,N_3315,N_3415);
and U3983 (N_3983,N_3293,N_3276);
or U3984 (N_3984,N_3388,N_3128);
or U3985 (N_3985,N_3400,N_3311);
nand U3986 (N_3986,N_3116,N_3016);
nand U3987 (N_3987,N_3055,N_3382);
and U3988 (N_3988,N_3369,N_3233);
nand U3989 (N_3989,N_3203,N_3272);
and U3990 (N_3990,N_3098,N_3435);
xnor U3991 (N_3991,N_3157,N_3219);
nor U3992 (N_3992,N_3220,N_3226);
nor U3993 (N_3993,N_3288,N_3230);
nand U3994 (N_3994,N_3190,N_3477);
nor U3995 (N_3995,N_3150,N_3112);
and U3996 (N_3996,N_3434,N_3008);
or U3997 (N_3997,N_3494,N_3431);
and U3998 (N_3998,N_3206,N_3062);
nand U3999 (N_3999,N_3485,N_3207);
and U4000 (N_4000,N_3532,N_3523);
nand U4001 (N_4001,N_3706,N_3726);
and U4002 (N_4002,N_3646,N_3853);
or U4003 (N_4003,N_3510,N_3651);
nor U4004 (N_4004,N_3633,N_3722);
xnor U4005 (N_4005,N_3834,N_3689);
nor U4006 (N_4006,N_3643,N_3863);
nand U4007 (N_4007,N_3754,N_3644);
nand U4008 (N_4008,N_3824,N_3731);
and U4009 (N_4009,N_3681,N_3894);
nand U4010 (N_4010,N_3612,N_3957);
xnor U4011 (N_4011,N_3514,N_3635);
and U4012 (N_4012,N_3971,N_3539);
and U4013 (N_4013,N_3768,N_3799);
nor U4014 (N_4014,N_3691,N_3941);
and U4015 (N_4015,N_3989,N_3950);
nand U4016 (N_4016,N_3877,N_3794);
or U4017 (N_4017,N_3571,N_3773);
and U4018 (N_4018,N_3800,N_3584);
nor U4019 (N_4019,N_3869,N_3710);
nand U4020 (N_4020,N_3966,N_3636);
nor U4021 (N_4021,N_3870,N_3900);
or U4022 (N_4022,N_3958,N_3830);
nand U4023 (N_4023,N_3991,N_3601);
nor U4024 (N_4024,N_3923,N_3888);
nor U4025 (N_4025,N_3924,N_3516);
nand U4026 (N_4026,N_3956,N_3945);
nand U4027 (N_4027,N_3567,N_3547);
and U4028 (N_4028,N_3952,N_3666);
xnor U4029 (N_4029,N_3831,N_3909);
nor U4030 (N_4030,N_3778,N_3916);
nand U4031 (N_4031,N_3901,N_3718);
nor U4032 (N_4032,N_3746,N_3749);
nor U4033 (N_4033,N_3913,N_3594);
and U4034 (N_4034,N_3565,N_3714);
nand U4035 (N_4035,N_3673,N_3719);
or U4036 (N_4036,N_3994,N_3763);
nand U4037 (N_4037,N_3562,N_3784);
or U4038 (N_4038,N_3979,N_3887);
or U4039 (N_4039,N_3798,N_3968);
nand U4040 (N_4040,N_3850,N_3802);
nor U4041 (N_4041,N_3732,N_3744);
xor U4042 (N_4042,N_3934,N_3915);
or U4043 (N_4043,N_3609,N_3815);
or U4044 (N_4044,N_3506,N_3883);
or U4045 (N_4045,N_3629,N_3791);
nand U4046 (N_4046,N_3825,N_3587);
nand U4047 (N_4047,N_3965,N_3751);
nand U4048 (N_4048,N_3769,N_3588);
nand U4049 (N_4049,N_3875,N_3623);
or U4050 (N_4050,N_3728,N_3683);
xnor U4051 (N_4051,N_3876,N_3697);
xnor U4052 (N_4052,N_3835,N_3858);
and U4053 (N_4053,N_3550,N_3503);
or U4054 (N_4054,N_3812,N_3625);
nand U4055 (N_4055,N_3943,N_3692);
or U4056 (N_4056,N_3804,N_3723);
and U4057 (N_4057,N_3712,N_3809);
and U4058 (N_4058,N_3650,N_3843);
nand U4059 (N_4059,N_3573,N_3603);
nand U4060 (N_4060,N_3828,N_3688);
and U4061 (N_4061,N_3929,N_3578);
and U4062 (N_4062,N_3551,N_3590);
and U4063 (N_4063,N_3600,N_3679);
nand U4064 (N_4064,N_3884,N_3842);
nand U4065 (N_4065,N_3713,N_3517);
and U4066 (N_4066,N_3944,N_3806);
nand U4067 (N_4067,N_3608,N_3509);
nand U4068 (N_4068,N_3793,N_3949);
nand U4069 (N_4069,N_3583,N_3621);
and U4070 (N_4070,N_3709,N_3559);
nor U4071 (N_4071,N_3935,N_3841);
and U4072 (N_4072,N_3823,N_3797);
nand U4073 (N_4073,N_3922,N_3693);
and U4074 (N_4074,N_3617,N_3885);
nor U4075 (N_4075,N_3739,N_3839);
and U4076 (N_4076,N_3519,N_3589);
or U4077 (N_4077,N_3611,N_3661);
or U4078 (N_4078,N_3969,N_3792);
and U4079 (N_4079,N_3618,N_3535);
or U4080 (N_4080,N_3524,N_3970);
nor U4081 (N_4081,N_3964,N_3647);
nand U4082 (N_4082,N_3730,N_3844);
or U4083 (N_4083,N_3538,N_3640);
nand U4084 (N_4084,N_3564,N_3978);
nor U4085 (N_4085,N_3715,N_3988);
and U4086 (N_4086,N_3753,N_3639);
nand U4087 (N_4087,N_3933,N_3557);
or U4088 (N_4088,N_3817,N_3743);
nor U4089 (N_4089,N_3748,N_3593);
nand U4090 (N_4090,N_3585,N_3946);
and U4091 (N_4091,N_3654,N_3504);
or U4092 (N_4092,N_3724,N_3615);
or U4093 (N_4093,N_3826,N_3833);
nand U4094 (N_4094,N_3528,N_3680);
and U4095 (N_4095,N_3677,N_3602);
xor U4096 (N_4096,N_3694,N_3541);
nor U4097 (N_4097,N_3796,N_3747);
nand U4098 (N_4098,N_3790,N_3906);
nand U4099 (N_4099,N_3955,N_3967);
nand U4100 (N_4100,N_3983,N_3904);
and U4101 (N_4101,N_3700,N_3903);
and U4102 (N_4102,N_3605,N_3663);
and U4103 (N_4103,N_3648,N_3820);
xnor U4104 (N_4104,N_3776,N_3918);
nand U4105 (N_4105,N_3921,N_3622);
nor U4106 (N_4106,N_3781,N_3813);
nand U4107 (N_4107,N_3656,N_3727);
and U4108 (N_4108,N_3576,N_3995);
nand U4109 (N_4109,N_3865,N_3675);
nor U4110 (N_4110,N_3986,N_3740);
xor U4111 (N_4111,N_3686,N_3897);
nand U4112 (N_4112,N_3822,N_3772);
or U4113 (N_4113,N_3599,N_3597);
nand U4114 (N_4114,N_3866,N_3999);
and U4115 (N_4115,N_3627,N_3992);
nand U4116 (N_4116,N_3515,N_3533);
and U4117 (N_4117,N_3761,N_3981);
nor U4118 (N_4118,N_3849,N_3771);
nor U4119 (N_4119,N_3948,N_3872);
nand U4120 (N_4120,N_3513,N_3954);
nor U4121 (N_4121,N_3745,N_3716);
and U4122 (N_4122,N_3898,N_3641);
and U4123 (N_4123,N_3705,N_3674);
nand U4124 (N_4124,N_3810,N_3568);
or U4125 (N_4125,N_3630,N_3840);
or U4126 (N_4126,N_3676,N_3982);
or U4127 (N_4127,N_3520,N_3667);
nor U4128 (N_4128,N_3546,N_3811);
nor U4129 (N_4129,N_3878,N_3805);
nand U4130 (N_4130,N_3638,N_3501);
and U4131 (N_4131,N_3801,N_3757);
nor U4132 (N_4132,N_3848,N_3660);
nand U4133 (N_4133,N_3917,N_3882);
or U4134 (N_4134,N_3814,N_3736);
or U4135 (N_4135,N_3649,N_3920);
nor U4136 (N_4136,N_3684,N_3711);
and U4137 (N_4137,N_3614,N_3556);
or U4138 (N_4138,N_3536,N_3755);
nand U4139 (N_4139,N_3540,N_3655);
nor U4140 (N_4140,N_3819,N_3760);
and U4141 (N_4141,N_3975,N_3505);
nor U4142 (N_4142,N_3893,N_3807);
nand U4143 (N_4143,N_3832,N_3996);
nor U4144 (N_4144,N_3560,N_3642);
nand U4145 (N_4145,N_3972,N_3671);
xor U4146 (N_4146,N_3664,N_3857);
and U4147 (N_4147,N_3765,N_3668);
or U4148 (N_4148,N_3997,N_3717);
or U4149 (N_4149,N_3976,N_3953);
nor U4150 (N_4150,N_3572,N_3659);
nand U4151 (N_4151,N_3852,N_3931);
nand U4152 (N_4152,N_3657,N_3725);
or U4153 (N_4153,N_3879,N_3598);
or U4154 (N_4154,N_3553,N_3637);
or U4155 (N_4155,N_3595,N_3847);
nor U4156 (N_4156,N_3534,N_3702);
nor U4157 (N_4157,N_3742,N_3787);
xor U4158 (N_4158,N_3558,N_3905);
nor U4159 (N_4159,N_3912,N_3961);
nor U4160 (N_4160,N_3604,N_3549);
nand U4161 (N_4161,N_3616,N_3669);
and U4162 (N_4162,N_3586,N_3704);
nor U4163 (N_4163,N_3938,N_3708);
xnor U4164 (N_4164,N_3764,N_3838);
or U4165 (N_4165,N_3891,N_3774);
and U4166 (N_4166,N_3930,N_3543);
nor U4167 (N_4167,N_3856,N_3579);
nor U4168 (N_4168,N_3974,N_3864);
and U4169 (N_4169,N_3699,N_3570);
nand U4170 (N_4170,N_3619,N_3735);
and U4171 (N_4171,N_3738,N_3846);
nand U4172 (N_4172,N_3977,N_3741);
or U4173 (N_4173,N_3932,N_3620);
nor U4174 (N_4174,N_3963,N_3581);
or U4175 (N_4175,N_3770,N_3928);
nand U4176 (N_4176,N_3626,N_3707);
xnor U4177 (N_4177,N_3569,N_3818);
and U4178 (N_4178,N_3628,N_3613);
nor U4179 (N_4179,N_3854,N_3881);
nand U4180 (N_4180,N_3574,N_3591);
xor U4181 (N_4181,N_3703,N_3960);
or U4182 (N_4182,N_3526,N_3874);
or U4183 (N_4183,N_3662,N_3829);
xnor U4184 (N_4184,N_3859,N_3511);
nand U4185 (N_4185,N_3733,N_3939);
and U4186 (N_4186,N_3721,N_3632);
xor U4187 (N_4187,N_3789,N_3527);
nor U4188 (N_4188,N_3993,N_3782);
or U4189 (N_4189,N_3767,N_3634);
or U4190 (N_4190,N_3554,N_3984);
xnor U4191 (N_4191,N_3803,N_3752);
xnor U4192 (N_4192,N_3895,N_3959);
xor U4193 (N_4193,N_3867,N_3665);
nor U4194 (N_4194,N_3592,N_3899);
nor U4195 (N_4195,N_3507,N_3690);
nand U4196 (N_4196,N_3582,N_3563);
nor U4197 (N_4197,N_3672,N_3777);
xor U4198 (N_4198,N_3508,N_3947);
or U4199 (N_4199,N_3980,N_3737);
and U4200 (N_4200,N_3762,N_3892);
and U4201 (N_4201,N_3911,N_3908);
nor U4202 (N_4202,N_3645,N_3512);
and U4203 (N_4203,N_3502,N_3610);
and U4204 (N_4204,N_3500,N_3889);
and U4205 (N_4205,N_3973,N_3886);
nor U4206 (N_4206,N_3862,N_3577);
or U4207 (N_4207,N_3682,N_3548);
xor U4208 (N_4208,N_3606,N_3775);
and U4209 (N_4209,N_3537,N_3871);
nand U4210 (N_4210,N_3529,N_3836);
nand U4211 (N_4211,N_3990,N_3518);
nor U4212 (N_4212,N_3919,N_3914);
nand U4213 (N_4213,N_3545,N_3542);
and U4214 (N_4214,N_3937,N_3696);
nand U4215 (N_4215,N_3851,N_3998);
and U4216 (N_4216,N_3780,N_3631);
xor U4217 (N_4217,N_3766,N_3873);
or U4218 (N_4218,N_3907,N_3624);
xor U4219 (N_4219,N_3607,N_3795);
xor U4220 (N_4220,N_3720,N_3868);
and U4221 (N_4221,N_3522,N_3530);
nand U4222 (N_4222,N_3652,N_3962);
or U4223 (N_4223,N_3951,N_3936);
and U4224 (N_4224,N_3927,N_3925);
or U4225 (N_4225,N_3544,N_3940);
nor U4226 (N_4226,N_3756,N_3926);
and U4227 (N_4227,N_3580,N_3758);
nor U4228 (N_4228,N_3896,N_3816);
nand U4229 (N_4229,N_3678,N_3561);
xnor U4230 (N_4230,N_3687,N_3890);
nand U4231 (N_4231,N_3785,N_3942);
nand U4232 (N_4232,N_3521,N_3575);
nand U4233 (N_4233,N_3552,N_3786);
xor U4234 (N_4234,N_3779,N_3658);
or U4235 (N_4235,N_3734,N_3987);
nand U4236 (N_4236,N_3985,N_3729);
nand U4237 (N_4237,N_3525,N_3788);
and U4238 (N_4238,N_3860,N_3759);
nand U4239 (N_4239,N_3880,N_3861);
or U4240 (N_4240,N_3902,N_3855);
xnor U4241 (N_4241,N_3685,N_3783);
and U4242 (N_4242,N_3596,N_3837);
and U4243 (N_4243,N_3845,N_3821);
nand U4244 (N_4244,N_3653,N_3827);
and U4245 (N_4245,N_3555,N_3750);
nor U4246 (N_4246,N_3531,N_3910);
nor U4247 (N_4247,N_3566,N_3698);
and U4248 (N_4248,N_3695,N_3808);
nor U4249 (N_4249,N_3701,N_3670);
nand U4250 (N_4250,N_3700,N_3866);
or U4251 (N_4251,N_3954,N_3681);
nand U4252 (N_4252,N_3509,N_3697);
or U4253 (N_4253,N_3934,N_3583);
nor U4254 (N_4254,N_3749,N_3775);
nand U4255 (N_4255,N_3931,N_3884);
nand U4256 (N_4256,N_3960,N_3542);
nand U4257 (N_4257,N_3767,N_3700);
nor U4258 (N_4258,N_3942,N_3643);
nand U4259 (N_4259,N_3979,N_3748);
nand U4260 (N_4260,N_3831,N_3983);
nand U4261 (N_4261,N_3930,N_3616);
nand U4262 (N_4262,N_3969,N_3757);
nor U4263 (N_4263,N_3850,N_3522);
or U4264 (N_4264,N_3563,N_3790);
and U4265 (N_4265,N_3938,N_3593);
xnor U4266 (N_4266,N_3682,N_3837);
or U4267 (N_4267,N_3870,N_3889);
xnor U4268 (N_4268,N_3641,N_3866);
and U4269 (N_4269,N_3817,N_3537);
or U4270 (N_4270,N_3569,N_3612);
nand U4271 (N_4271,N_3522,N_3764);
or U4272 (N_4272,N_3919,N_3823);
and U4273 (N_4273,N_3960,N_3799);
xnor U4274 (N_4274,N_3852,N_3705);
and U4275 (N_4275,N_3730,N_3725);
xnor U4276 (N_4276,N_3967,N_3987);
and U4277 (N_4277,N_3562,N_3761);
nor U4278 (N_4278,N_3717,N_3870);
nand U4279 (N_4279,N_3581,N_3645);
xor U4280 (N_4280,N_3566,N_3666);
nand U4281 (N_4281,N_3696,N_3760);
and U4282 (N_4282,N_3719,N_3988);
or U4283 (N_4283,N_3792,N_3532);
and U4284 (N_4284,N_3622,N_3607);
nor U4285 (N_4285,N_3888,N_3660);
and U4286 (N_4286,N_3733,N_3816);
and U4287 (N_4287,N_3901,N_3765);
and U4288 (N_4288,N_3821,N_3565);
nor U4289 (N_4289,N_3808,N_3782);
or U4290 (N_4290,N_3983,N_3594);
xnor U4291 (N_4291,N_3871,N_3990);
nand U4292 (N_4292,N_3666,N_3914);
nand U4293 (N_4293,N_3876,N_3863);
xnor U4294 (N_4294,N_3762,N_3852);
or U4295 (N_4295,N_3959,N_3986);
nand U4296 (N_4296,N_3623,N_3645);
xor U4297 (N_4297,N_3514,N_3565);
or U4298 (N_4298,N_3939,N_3938);
and U4299 (N_4299,N_3859,N_3825);
and U4300 (N_4300,N_3813,N_3751);
or U4301 (N_4301,N_3933,N_3958);
or U4302 (N_4302,N_3775,N_3905);
and U4303 (N_4303,N_3739,N_3727);
or U4304 (N_4304,N_3856,N_3857);
xnor U4305 (N_4305,N_3730,N_3519);
or U4306 (N_4306,N_3739,N_3687);
or U4307 (N_4307,N_3876,N_3891);
nor U4308 (N_4308,N_3843,N_3562);
or U4309 (N_4309,N_3948,N_3549);
nand U4310 (N_4310,N_3876,N_3931);
xnor U4311 (N_4311,N_3557,N_3960);
nor U4312 (N_4312,N_3703,N_3808);
xnor U4313 (N_4313,N_3875,N_3622);
xor U4314 (N_4314,N_3693,N_3588);
nor U4315 (N_4315,N_3770,N_3946);
nor U4316 (N_4316,N_3879,N_3594);
nand U4317 (N_4317,N_3698,N_3935);
nand U4318 (N_4318,N_3808,N_3754);
nand U4319 (N_4319,N_3822,N_3937);
and U4320 (N_4320,N_3990,N_3815);
nor U4321 (N_4321,N_3696,N_3981);
nand U4322 (N_4322,N_3910,N_3687);
and U4323 (N_4323,N_3982,N_3971);
or U4324 (N_4324,N_3610,N_3688);
xor U4325 (N_4325,N_3682,N_3981);
nor U4326 (N_4326,N_3573,N_3506);
or U4327 (N_4327,N_3641,N_3806);
nand U4328 (N_4328,N_3806,N_3771);
or U4329 (N_4329,N_3607,N_3534);
xnor U4330 (N_4330,N_3674,N_3597);
nand U4331 (N_4331,N_3511,N_3923);
or U4332 (N_4332,N_3855,N_3823);
or U4333 (N_4333,N_3739,N_3924);
nand U4334 (N_4334,N_3861,N_3502);
and U4335 (N_4335,N_3787,N_3517);
or U4336 (N_4336,N_3509,N_3589);
and U4337 (N_4337,N_3525,N_3803);
or U4338 (N_4338,N_3615,N_3854);
nor U4339 (N_4339,N_3793,N_3731);
nor U4340 (N_4340,N_3917,N_3894);
nor U4341 (N_4341,N_3574,N_3706);
nor U4342 (N_4342,N_3735,N_3826);
nor U4343 (N_4343,N_3738,N_3732);
and U4344 (N_4344,N_3960,N_3517);
xnor U4345 (N_4345,N_3706,N_3740);
nand U4346 (N_4346,N_3604,N_3949);
or U4347 (N_4347,N_3842,N_3598);
nand U4348 (N_4348,N_3644,N_3566);
and U4349 (N_4349,N_3865,N_3887);
nand U4350 (N_4350,N_3522,N_3932);
and U4351 (N_4351,N_3563,N_3760);
xnor U4352 (N_4352,N_3819,N_3698);
nor U4353 (N_4353,N_3534,N_3596);
and U4354 (N_4354,N_3946,N_3544);
nor U4355 (N_4355,N_3802,N_3513);
nand U4356 (N_4356,N_3775,N_3760);
and U4357 (N_4357,N_3798,N_3759);
or U4358 (N_4358,N_3575,N_3975);
nor U4359 (N_4359,N_3720,N_3922);
nor U4360 (N_4360,N_3966,N_3517);
or U4361 (N_4361,N_3841,N_3733);
and U4362 (N_4362,N_3534,N_3524);
and U4363 (N_4363,N_3721,N_3891);
and U4364 (N_4364,N_3563,N_3943);
nor U4365 (N_4365,N_3957,N_3919);
or U4366 (N_4366,N_3506,N_3570);
nand U4367 (N_4367,N_3775,N_3591);
nor U4368 (N_4368,N_3990,N_3534);
or U4369 (N_4369,N_3972,N_3527);
or U4370 (N_4370,N_3638,N_3995);
or U4371 (N_4371,N_3932,N_3899);
and U4372 (N_4372,N_3647,N_3801);
nand U4373 (N_4373,N_3542,N_3513);
and U4374 (N_4374,N_3885,N_3753);
and U4375 (N_4375,N_3715,N_3623);
or U4376 (N_4376,N_3882,N_3892);
nor U4377 (N_4377,N_3879,N_3543);
nand U4378 (N_4378,N_3939,N_3695);
nor U4379 (N_4379,N_3948,N_3862);
and U4380 (N_4380,N_3946,N_3959);
nand U4381 (N_4381,N_3670,N_3642);
nor U4382 (N_4382,N_3862,N_3958);
nor U4383 (N_4383,N_3557,N_3978);
or U4384 (N_4384,N_3802,N_3601);
nor U4385 (N_4385,N_3986,N_3742);
nand U4386 (N_4386,N_3799,N_3547);
xnor U4387 (N_4387,N_3588,N_3976);
xor U4388 (N_4388,N_3631,N_3623);
nand U4389 (N_4389,N_3518,N_3598);
xor U4390 (N_4390,N_3814,N_3964);
nor U4391 (N_4391,N_3991,N_3715);
and U4392 (N_4392,N_3704,N_3745);
nor U4393 (N_4393,N_3744,N_3598);
nor U4394 (N_4394,N_3751,N_3653);
nor U4395 (N_4395,N_3633,N_3773);
or U4396 (N_4396,N_3674,N_3738);
and U4397 (N_4397,N_3801,N_3897);
nor U4398 (N_4398,N_3818,N_3513);
and U4399 (N_4399,N_3853,N_3692);
nand U4400 (N_4400,N_3570,N_3851);
nor U4401 (N_4401,N_3992,N_3822);
nand U4402 (N_4402,N_3771,N_3571);
and U4403 (N_4403,N_3647,N_3822);
nand U4404 (N_4404,N_3574,N_3951);
nand U4405 (N_4405,N_3528,N_3768);
and U4406 (N_4406,N_3637,N_3577);
and U4407 (N_4407,N_3787,N_3922);
and U4408 (N_4408,N_3527,N_3841);
or U4409 (N_4409,N_3609,N_3769);
and U4410 (N_4410,N_3815,N_3742);
nor U4411 (N_4411,N_3592,N_3943);
and U4412 (N_4412,N_3731,N_3625);
nand U4413 (N_4413,N_3662,N_3768);
or U4414 (N_4414,N_3570,N_3777);
nand U4415 (N_4415,N_3731,N_3902);
or U4416 (N_4416,N_3522,N_3508);
or U4417 (N_4417,N_3924,N_3750);
or U4418 (N_4418,N_3666,N_3546);
nor U4419 (N_4419,N_3803,N_3630);
nor U4420 (N_4420,N_3730,N_3828);
xnor U4421 (N_4421,N_3730,N_3830);
nor U4422 (N_4422,N_3668,N_3770);
xnor U4423 (N_4423,N_3611,N_3688);
xnor U4424 (N_4424,N_3804,N_3775);
and U4425 (N_4425,N_3971,N_3915);
and U4426 (N_4426,N_3563,N_3735);
nand U4427 (N_4427,N_3811,N_3762);
and U4428 (N_4428,N_3926,N_3798);
xor U4429 (N_4429,N_3729,N_3989);
or U4430 (N_4430,N_3534,N_3921);
nand U4431 (N_4431,N_3879,N_3768);
nand U4432 (N_4432,N_3685,N_3660);
nand U4433 (N_4433,N_3575,N_3589);
and U4434 (N_4434,N_3763,N_3560);
nor U4435 (N_4435,N_3584,N_3501);
nand U4436 (N_4436,N_3525,N_3889);
xor U4437 (N_4437,N_3953,N_3736);
nand U4438 (N_4438,N_3934,N_3754);
or U4439 (N_4439,N_3553,N_3774);
nor U4440 (N_4440,N_3583,N_3615);
and U4441 (N_4441,N_3623,N_3635);
or U4442 (N_4442,N_3620,N_3641);
or U4443 (N_4443,N_3934,N_3987);
nor U4444 (N_4444,N_3838,N_3695);
and U4445 (N_4445,N_3676,N_3991);
and U4446 (N_4446,N_3694,N_3832);
and U4447 (N_4447,N_3976,N_3507);
nand U4448 (N_4448,N_3993,N_3885);
nand U4449 (N_4449,N_3762,N_3726);
nand U4450 (N_4450,N_3930,N_3789);
and U4451 (N_4451,N_3814,N_3989);
or U4452 (N_4452,N_3974,N_3510);
nand U4453 (N_4453,N_3861,N_3713);
nor U4454 (N_4454,N_3950,N_3952);
nor U4455 (N_4455,N_3911,N_3993);
nand U4456 (N_4456,N_3503,N_3796);
nor U4457 (N_4457,N_3643,N_3803);
and U4458 (N_4458,N_3697,N_3569);
or U4459 (N_4459,N_3923,N_3862);
nor U4460 (N_4460,N_3785,N_3943);
and U4461 (N_4461,N_3679,N_3690);
nand U4462 (N_4462,N_3747,N_3961);
and U4463 (N_4463,N_3902,N_3617);
nand U4464 (N_4464,N_3951,N_3810);
or U4465 (N_4465,N_3698,N_3524);
nor U4466 (N_4466,N_3882,N_3726);
nor U4467 (N_4467,N_3663,N_3512);
or U4468 (N_4468,N_3732,N_3769);
or U4469 (N_4469,N_3527,N_3831);
nor U4470 (N_4470,N_3590,N_3895);
or U4471 (N_4471,N_3773,N_3570);
xnor U4472 (N_4472,N_3946,N_3987);
nand U4473 (N_4473,N_3982,N_3554);
xnor U4474 (N_4474,N_3660,N_3779);
and U4475 (N_4475,N_3616,N_3787);
or U4476 (N_4476,N_3599,N_3954);
or U4477 (N_4477,N_3768,N_3666);
or U4478 (N_4478,N_3871,N_3955);
nand U4479 (N_4479,N_3534,N_3923);
nor U4480 (N_4480,N_3531,N_3713);
nand U4481 (N_4481,N_3827,N_3795);
and U4482 (N_4482,N_3825,N_3582);
or U4483 (N_4483,N_3787,N_3508);
and U4484 (N_4484,N_3688,N_3559);
or U4485 (N_4485,N_3736,N_3684);
nand U4486 (N_4486,N_3688,N_3871);
and U4487 (N_4487,N_3795,N_3685);
xnor U4488 (N_4488,N_3797,N_3892);
or U4489 (N_4489,N_3901,N_3925);
nand U4490 (N_4490,N_3906,N_3830);
nor U4491 (N_4491,N_3881,N_3635);
or U4492 (N_4492,N_3916,N_3733);
xor U4493 (N_4493,N_3533,N_3781);
and U4494 (N_4494,N_3891,N_3848);
nand U4495 (N_4495,N_3689,N_3600);
or U4496 (N_4496,N_3728,N_3931);
xnor U4497 (N_4497,N_3576,N_3881);
nor U4498 (N_4498,N_3625,N_3830);
or U4499 (N_4499,N_3881,N_3855);
nor U4500 (N_4500,N_4162,N_4414);
and U4501 (N_4501,N_4298,N_4057);
nor U4502 (N_4502,N_4263,N_4142);
and U4503 (N_4503,N_4035,N_4327);
nor U4504 (N_4504,N_4079,N_4369);
nor U4505 (N_4505,N_4264,N_4288);
xnor U4506 (N_4506,N_4297,N_4405);
nor U4507 (N_4507,N_4480,N_4393);
and U4508 (N_4508,N_4144,N_4166);
or U4509 (N_4509,N_4147,N_4056);
nor U4510 (N_4510,N_4175,N_4285);
nand U4511 (N_4511,N_4330,N_4435);
nand U4512 (N_4512,N_4068,N_4363);
or U4513 (N_4513,N_4458,N_4312);
or U4514 (N_4514,N_4492,N_4477);
or U4515 (N_4515,N_4049,N_4470);
and U4516 (N_4516,N_4321,N_4491);
nand U4517 (N_4517,N_4307,N_4239);
xnor U4518 (N_4518,N_4004,N_4257);
nor U4519 (N_4519,N_4357,N_4100);
or U4520 (N_4520,N_4053,N_4333);
nor U4521 (N_4521,N_4037,N_4343);
or U4522 (N_4522,N_4001,N_4188);
nand U4523 (N_4523,N_4459,N_4489);
nand U4524 (N_4524,N_4226,N_4006);
and U4525 (N_4525,N_4326,N_4398);
nor U4526 (N_4526,N_4216,N_4420);
or U4527 (N_4527,N_4427,N_4411);
nor U4528 (N_4528,N_4048,N_4268);
and U4529 (N_4529,N_4418,N_4483);
nor U4530 (N_4530,N_4221,N_4030);
nor U4531 (N_4531,N_4373,N_4442);
or U4532 (N_4532,N_4388,N_4095);
and U4533 (N_4533,N_4109,N_4067);
xnor U4534 (N_4534,N_4238,N_4089);
nand U4535 (N_4535,N_4410,N_4482);
and U4536 (N_4536,N_4206,N_4218);
or U4537 (N_4537,N_4200,N_4033);
nand U4538 (N_4538,N_4335,N_4361);
nand U4539 (N_4539,N_4495,N_4207);
nor U4540 (N_4540,N_4422,N_4378);
nor U4541 (N_4541,N_4087,N_4242);
and U4542 (N_4542,N_4341,N_4250);
and U4543 (N_4543,N_4261,N_4043);
nor U4544 (N_4544,N_4047,N_4260);
nand U4545 (N_4545,N_4417,N_4404);
or U4546 (N_4546,N_4097,N_4432);
nor U4547 (N_4547,N_4408,N_4292);
and U4548 (N_4548,N_4413,N_4428);
nor U4549 (N_4549,N_4457,N_4134);
or U4550 (N_4550,N_4069,N_4039);
nand U4551 (N_4551,N_4101,N_4277);
nand U4552 (N_4552,N_4340,N_4186);
nor U4553 (N_4553,N_4396,N_4415);
and U4554 (N_4554,N_4274,N_4122);
or U4555 (N_4555,N_4083,N_4024);
nand U4556 (N_4556,N_4368,N_4283);
nor U4557 (N_4557,N_4262,N_4441);
and U4558 (N_4558,N_4365,N_4303);
nor U4559 (N_4559,N_4085,N_4296);
nand U4560 (N_4560,N_4461,N_4042);
and U4561 (N_4561,N_4005,N_4193);
nand U4562 (N_4562,N_4464,N_4252);
and U4563 (N_4563,N_4187,N_4247);
xor U4564 (N_4564,N_4012,N_4301);
xnor U4565 (N_4565,N_4081,N_4355);
nor U4566 (N_4566,N_4382,N_4389);
or U4567 (N_4567,N_4044,N_4350);
nand U4568 (N_4568,N_4176,N_4183);
or U4569 (N_4569,N_4476,N_4407);
and U4570 (N_4570,N_4496,N_4267);
and U4571 (N_4571,N_4342,N_4468);
nand U4572 (N_4572,N_4270,N_4258);
xnor U4573 (N_4573,N_4169,N_4107);
nor U4574 (N_4574,N_4161,N_4402);
nand U4575 (N_4575,N_4205,N_4148);
and U4576 (N_4576,N_4106,N_4019);
nor U4577 (N_4577,N_4153,N_4438);
nor U4578 (N_4578,N_4062,N_4290);
nand U4579 (N_4579,N_4434,N_4214);
or U4580 (N_4580,N_4469,N_4452);
and U4581 (N_4581,N_4278,N_4356);
or U4582 (N_4582,N_4454,N_4123);
xnor U4583 (N_4583,N_4137,N_4338);
nand U4584 (N_4584,N_4008,N_4478);
or U4585 (N_4585,N_4167,N_4103);
and U4586 (N_4586,N_4099,N_4446);
nor U4587 (N_4587,N_4104,N_4170);
or U4588 (N_4588,N_4299,N_4329);
and U4589 (N_4589,N_4244,N_4151);
or U4590 (N_4590,N_4400,N_4286);
and U4591 (N_4591,N_4310,N_4054);
nor U4592 (N_4592,N_4051,N_4248);
nor U4593 (N_4593,N_4111,N_4311);
or U4594 (N_4594,N_4347,N_4178);
or U4595 (N_4595,N_4465,N_4474);
nand U4596 (N_4596,N_4066,N_4451);
nand U4597 (N_4597,N_4021,N_4376);
or U4598 (N_4598,N_4105,N_4015);
xor U4599 (N_4599,N_4390,N_4196);
or U4600 (N_4600,N_4145,N_4318);
and U4601 (N_4601,N_4453,N_4426);
or U4602 (N_4602,N_4171,N_4332);
nor U4603 (N_4603,N_4098,N_4040);
or U4604 (N_4604,N_4395,N_4377);
and U4605 (N_4605,N_4366,N_4433);
and U4606 (N_4606,N_4460,N_4023);
nor U4607 (N_4607,N_4336,N_4279);
or U4608 (N_4608,N_4423,N_4437);
xor U4609 (N_4609,N_4241,N_4273);
and U4610 (N_4610,N_4352,N_4182);
and U4611 (N_4611,N_4466,N_4319);
nand U4612 (N_4612,N_4157,N_4113);
and U4613 (N_4613,N_4281,N_4499);
and U4614 (N_4614,N_4163,N_4050);
nor U4615 (N_4615,N_4275,N_4082);
nor U4616 (N_4616,N_4059,N_4463);
xor U4617 (N_4617,N_4253,N_4197);
and U4618 (N_4618,N_4225,N_4091);
nand U4619 (N_4619,N_4237,N_4013);
nand U4620 (N_4620,N_4036,N_4394);
and U4621 (N_4621,N_4306,N_4320);
or U4622 (N_4622,N_4031,N_4351);
nor U4623 (N_4623,N_4076,N_4429);
and U4624 (N_4624,N_4245,N_4118);
nor U4625 (N_4625,N_4077,N_4117);
nor U4626 (N_4626,N_4086,N_4128);
nor U4627 (N_4627,N_4072,N_4450);
or U4628 (N_4628,N_4265,N_4313);
nand U4629 (N_4629,N_4359,N_4269);
or U4630 (N_4630,N_4022,N_4133);
or U4631 (N_4631,N_4135,N_4322);
and U4632 (N_4632,N_4165,N_4075);
or U4633 (N_4633,N_4029,N_4445);
nor U4634 (N_4634,N_4129,N_4156);
xor U4635 (N_4635,N_4490,N_4488);
xor U4636 (N_4636,N_4412,N_4325);
or U4637 (N_4637,N_4345,N_4360);
and U4638 (N_4638,N_4154,N_4014);
and U4639 (N_4639,N_4358,N_4112);
nor U4640 (N_4640,N_4314,N_4479);
and U4641 (N_4641,N_4094,N_4127);
nor U4642 (N_4642,N_4164,N_4073);
nand U4643 (N_4643,N_4372,N_4026);
or U4644 (N_4644,N_4271,N_4254);
or U4645 (N_4645,N_4449,N_4240);
nand U4646 (N_4646,N_4397,N_4304);
nand U4647 (N_4647,N_4071,N_4189);
nand U4648 (N_4648,N_4431,N_4191);
or U4649 (N_4649,N_4204,N_4143);
or U4650 (N_4650,N_4090,N_4473);
or U4651 (N_4651,N_4231,N_4302);
or U4652 (N_4652,N_4291,N_4421);
and U4653 (N_4653,N_4331,N_4305);
nor U4654 (N_4654,N_4403,N_4084);
or U4655 (N_4655,N_4308,N_4370);
xnor U4656 (N_4656,N_4456,N_4354);
nand U4657 (N_4657,N_4080,N_4472);
and U4658 (N_4658,N_4177,N_4102);
nand U4659 (N_4659,N_4309,N_4436);
or U4660 (N_4660,N_4346,N_4210);
nand U4661 (N_4661,N_4141,N_4293);
or U4662 (N_4662,N_4481,N_4055);
nand U4663 (N_4663,N_4150,N_4401);
nor U4664 (N_4664,N_4045,N_4131);
nand U4665 (N_4665,N_4364,N_4295);
nand U4666 (N_4666,N_4194,N_4018);
or U4667 (N_4667,N_4052,N_4494);
nand U4668 (N_4668,N_4058,N_4259);
or U4669 (N_4669,N_4255,N_4092);
and U4670 (N_4670,N_4236,N_4223);
xor U4671 (N_4671,N_4149,N_4243);
nor U4672 (N_4672,N_4228,N_4116);
xnor U4673 (N_4673,N_4027,N_4201);
xor U4674 (N_4674,N_4110,N_4120);
xnor U4675 (N_4675,N_4185,N_4416);
nor U4676 (N_4676,N_4070,N_4374);
or U4677 (N_4677,N_4246,N_4020);
xnor U4678 (N_4678,N_4168,N_4475);
nor U4679 (N_4679,N_4230,N_4152);
nor U4680 (N_4680,N_4443,N_4190);
nor U4681 (N_4681,N_4034,N_4146);
or U4682 (N_4682,N_4287,N_4344);
nand U4683 (N_4683,N_4000,N_4140);
xor U4684 (N_4684,N_4003,N_4017);
or U4685 (N_4685,N_4184,N_4229);
nand U4686 (N_4686,N_4375,N_4115);
nand U4687 (N_4687,N_4016,N_4493);
nor U4688 (N_4688,N_4339,N_4195);
and U4689 (N_4689,N_4119,N_4316);
or U4690 (N_4690,N_4497,N_4011);
or U4691 (N_4691,N_4455,N_4289);
nand U4692 (N_4692,N_4323,N_4172);
and U4693 (N_4693,N_4007,N_4208);
nor U4694 (N_4694,N_4219,N_4041);
nor U4695 (N_4695,N_4160,N_4462);
nor U4696 (N_4696,N_4284,N_4392);
xor U4697 (N_4697,N_4276,N_4317);
nor U4698 (N_4698,N_4383,N_4233);
nor U4699 (N_4699,N_4385,N_4155);
nor U4700 (N_4700,N_4124,N_4213);
xnor U4701 (N_4701,N_4010,N_4487);
and U4702 (N_4702,N_4439,N_4471);
and U4703 (N_4703,N_4061,N_4215);
nor U4704 (N_4704,N_4063,N_4114);
nor U4705 (N_4705,N_4108,N_4399);
nand U4706 (N_4706,N_4430,N_4379);
xnor U4707 (N_4707,N_4498,N_4159);
or U4708 (N_4708,N_4444,N_4136);
nor U4709 (N_4709,N_4315,N_4209);
and U4710 (N_4710,N_4180,N_4025);
xor U4711 (N_4711,N_4386,N_4222);
xnor U4712 (N_4712,N_4220,N_4234);
nand U4713 (N_4713,N_4002,N_4130);
or U4714 (N_4714,N_4380,N_4485);
or U4715 (N_4715,N_4046,N_4280);
and U4716 (N_4716,N_4235,N_4174);
nand U4717 (N_4717,N_4484,N_4353);
and U4718 (N_4718,N_4424,N_4387);
and U4719 (N_4719,N_4202,N_4266);
and U4720 (N_4720,N_4324,N_4078);
nor U4721 (N_4721,N_4009,N_4032);
nor U4722 (N_4722,N_4065,N_4381);
nor U4723 (N_4723,N_4419,N_4282);
nor U4724 (N_4724,N_4334,N_4028);
or U4725 (N_4725,N_4227,N_4349);
and U4726 (N_4726,N_4447,N_4440);
xnor U4727 (N_4727,N_4181,N_4212);
nand U4728 (N_4728,N_4198,N_4448);
nor U4729 (N_4729,N_4224,N_4272);
and U4730 (N_4730,N_4060,N_4337);
nand U4731 (N_4731,N_4249,N_4074);
or U4732 (N_4732,N_4300,N_4406);
and U4733 (N_4733,N_4348,N_4409);
or U4734 (N_4734,N_4088,N_4138);
nor U4735 (N_4735,N_4179,N_4367);
or U4736 (N_4736,N_4371,N_4126);
or U4737 (N_4737,N_4064,N_4232);
nor U4738 (N_4738,N_4121,N_4486);
nand U4739 (N_4739,N_4192,N_4132);
and U4740 (N_4740,N_4425,N_4256);
and U4741 (N_4741,N_4362,N_4251);
and U4742 (N_4742,N_4038,N_4467);
xnor U4743 (N_4743,N_4211,N_4203);
xor U4744 (N_4744,N_4125,N_4158);
xnor U4745 (N_4745,N_4217,N_4173);
nand U4746 (N_4746,N_4096,N_4384);
or U4747 (N_4747,N_4294,N_4139);
nand U4748 (N_4748,N_4093,N_4391);
nor U4749 (N_4749,N_4328,N_4199);
and U4750 (N_4750,N_4208,N_4456);
or U4751 (N_4751,N_4494,N_4078);
and U4752 (N_4752,N_4468,N_4153);
and U4753 (N_4753,N_4183,N_4390);
nand U4754 (N_4754,N_4450,N_4404);
nand U4755 (N_4755,N_4114,N_4360);
and U4756 (N_4756,N_4408,N_4187);
or U4757 (N_4757,N_4028,N_4279);
nor U4758 (N_4758,N_4054,N_4011);
nand U4759 (N_4759,N_4032,N_4373);
nand U4760 (N_4760,N_4485,N_4135);
or U4761 (N_4761,N_4216,N_4288);
xor U4762 (N_4762,N_4078,N_4346);
nand U4763 (N_4763,N_4021,N_4463);
or U4764 (N_4764,N_4067,N_4359);
xnor U4765 (N_4765,N_4402,N_4392);
or U4766 (N_4766,N_4166,N_4205);
nor U4767 (N_4767,N_4191,N_4172);
or U4768 (N_4768,N_4203,N_4082);
nand U4769 (N_4769,N_4249,N_4490);
nor U4770 (N_4770,N_4129,N_4183);
or U4771 (N_4771,N_4169,N_4477);
nand U4772 (N_4772,N_4411,N_4288);
xnor U4773 (N_4773,N_4474,N_4319);
xnor U4774 (N_4774,N_4301,N_4485);
nand U4775 (N_4775,N_4269,N_4112);
nor U4776 (N_4776,N_4262,N_4045);
and U4777 (N_4777,N_4205,N_4490);
nand U4778 (N_4778,N_4070,N_4223);
or U4779 (N_4779,N_4489,N_4029);
and U4780 (N_4780,N_4022,N_4475);
nand U4781 (N_4781,N_4198,N_4445);
or U4782 (N_4782,N_4093,N_4398);
nor U4783 (N_4783,N_4462,N_4119);
and U4784 (N_4784,N_4455,N_4155);
nand U4785 (N_4785,N_4238,N_4311);
nor U4786 (N_4786,N_4403,N_4247);
or U4787 (N_4787,N_4041,N_4092);
and U4788 (N_4788,N_4147,N_4210);
nor U4789 (N_4789,N_4100,N_4353);
and U4790 (N_4790,N_4090,N_4489);
or U4791 (N_4791,N_4346,N_4131);
nor U4792 (N_4792,N_4177,N_4402);
and U4793 (N_4793,N_4439,N_4006);
and U4794 (N_4794,N_4142,N_4047);
nand U4795 (N_4795,N_4138,N_4176);
and U4796 (N_4796,N_4089,N_4384);
nand U4797 (N_4797,N_4171,N_4211);
nand U4798 (N_4798,N_4231,N_4033);
and U4799 (N_4799,N_4386,N_4003);
nand U4800 (N_4800,N_4315,N_4024);
nor U4801 (N_4801,N_4046,N_4406);
or U4802 (N_4802,N_4203,N_4277);
nand U4803 (N_4803,N_4043,N_4317);
or U4804 (N_4804,N_4105,N_4143);
nand U4805 (N_4805,N_4237,N_4095);
and U4806 (N_4806,N_4462,N_4355);
or U4807 (N_4807,N_4309,N_4472);
or U4808 (N_4808,N_4206,N_4061);
and U4809 (N_4809,N_4281,N_4129);
nor U4810 (N_4810,N_4135,N_4447);
nand U4811 (N_4811,N_4273,N_4049);
nor U4812 (N_4812,N_4462,N_4347);
nand U4813 (N_4813,N_4324,N_4059);
nor U4814 (N_4814,N_4348,N_4229);
nor U4815 (N_4815,N_4171,N_4053);
nor U4816 (N_4816,N_4358,N_4497);
nand U4817 (N_4817,N_4467,N_4457);
or U4818 (N_4818,N_4070,N_4257);
and U4819 (N_4819,N_4172,N_4490);
and U4820 (N_4820,N_4428,N_4129);
nor U4821 (N_4821,N_4321,N_4258);
nor U4822 (N_4822,N_4359,N_4385);
nand U4823 (N_4823,N_4438,N_4052);
nor U4824 (N_4824,N_4160,N_4494);
nor U4825 (N_4825,N_4177,N_4382);
xor U4826 (N_4826,N_4496,N_4233);
nor U4827 (N_4827,N_4111,N_4041);
and U4828 (N_4828,N_4490,N_4295);
or U4829 (N_4829,N_4297,N_4115);
nand U4830 (N_4830,N_4474,N_4295);
nor U4831 (N_4831,N_4149,N_4100);
nand U4832 (N_4832,N_4052,N_4431);
or U4833 (N_4833,N_4179,N_4043);
nand U4834 (N_4834,N_4019,N_4148);
and U4835 (N_4835,N_4010,N_4463);
xnor U4836 (N_4836,N_4372,N_4200);
xnor U4837 (N_4837,N_4077,N_4481);
nand U4838 (N_4838,N_4197,N_4141);
xor U4839 (N_4839,N_4482,N_4098);
and U4840 (N_4840,N_4370,N_4242);
and U4841 (N_4841,N_4076,N_4176);
nand U4842 (N_4842,N_4264,N_4349);
or U4843 (N_4843,N_4327,N_4214);
nor U4844 (N_4844,N_4423,N_4178);
and U4845 (N_4845,N_4323,N_4446);
or U4846 (N_4846,N_4111,N_4173);
and U4847 (N_4847,N_4405,N_4369);
nand U4848 (N_4848,N_4311,N_4141);
nor U4849 (N_4849,N_4337,N_4294);
xor U4850 (N_4850,N_4228,N_4440);
or U4851 (N_4851,N_4467,N_4149);
and U4852 (N_4852,N_4344,N_4372);
nor U4853 (N_4853,N_4136,N_4135);
nor U4854 (N_4854,N_4302,N_4363);
and U4855 (N_4855,N_4334,N_4254);
or U4856 (N_4856,N_4420,N_4199);
nor U4857 (N_4857,N_4206,N_4279);
nand U4858 (N_4858,N_4373,N_4088);
nor U4859 (N_4859,N_4251,N_4422);
or U4860 (N_4860,N_4464,N_4313);
nor U4861 (N_4861,N_4298,N_4259);
nor U4862 (N_4862,N_4429,N_4180);
nand U4863 (N_4863,N_4184,N_4471);
xor U4864 (N_4864,N_4391,N_4483);
or U4865 (N_4865,N_4355,N_4364);
nor U4866 (N_4866,N_4275,N_4187);
nor U4867 (N_4867,N_4387,N_4016);
and U4868 (N_4868,N_4258,N_4032);
nor U4869 (N_4869,N_4167,N_4232);
nor U4870 (N_4870,N_4101,N_4187);
and U4871 (N_4871,N_4333,N_4076);
nor U4872 (N_4872,N_4478,N_4000);
or U4873 (N_4873,N_4126,N_4295);
nor U4874 (N_4874,N_4236,N_4174);
nor U4875 (N_4875,N_4268,N_4097);
xnor U4876 (N_4876,N_4168,N_4176);
nor U4877 (N_4877,N_4287,N_4288);
nand U4878 (N_4878,N_4141,N_4395);
xnor U4879 (N_4879,N_4436,N_4188);
or U4880 (N_4880,N_4089,N_4123);
nor U4881 (N_4881,N_4342,N_4061);
nand U4882 (N_4882,N_4009,N_4112);
nor U4883 (N_4883,N_4440,N_4139);
and U4884 (N_4884,N_4460,N_4172);
nor U4885 (N_4885,N_4164,N_4057);
and U4886 (N_4886,N_4186,N_4030);
or U4887 (N_4887,N_4205,N_4316);
nor U4888 (N_4888,N_4430,N_4292);
nor U4889 (N_4889,N_4267,N_4133);
or U4890 (N_4890,N_4461,N_4372);
nand U4891 (N_4891,N_4074,N_4321);
nor U4892 (N_4892,N_4178,N_4417);
nand U4893 (N_4893,N_4037,N_4242);
nand U4894 (N_4894,N_4427,N_4217);
nor U4895 (N_4895,N_4458,N_4471);
nand U4896 (N_4896,N_4314,N_4429);
nor U4897 (N_4897,N_4418,N_4387);
or U4898 (N_4898,N_4383,N_4428);
or U4899 (N_4899,N_4362,N_4055);
or U4900 (N_4900,N_4004,N_4119);
nand U4901 (N_4901,N_4139,N_4230);
nor U4902 (N_4902,N_4196,N_4163);
and U4903 (N_4903,N_4404,N_4185);
nand U4904 (N_4904,N_4145,N_4105);
nor U4905 (N_4905,N_4121,N_4288);
and U4906 (N_4906,N_4085,N_4221);
and U4907 (N_4907,N_4431,N_4392);
or U4908 (N_4908,N_4464,N_4156);
or U4909 (N_4909,N_4218,N_4474);
nor U4910 (N_4910,N_4291,N_4020);
nor U4911 (N_4911,N_4188,N_4098);
nand U4912 (N_4912,N_4359,N_4307);
and U4913 (N_4913,N_4075,N_4259);
nand U4914 (N_4914,N_4085,N_4332);
xor U4915 (N_4915,N_4354,N_4228);
or U4916 (N_4916,N_4370,N_4095);
and U4917 (N_4917,N_4032,N_4374);
or U4918 (N_4918,N_4012,N_4470);
xnor U4919 (N_4919,N_4033,N_4359);
and U4920 (N_4920,N_4339,N_4238);
and U4921 (N_4921,N_4054,N_4283);
and U4922 (N_4922,N_4013,N_4268);
and U4923 (N_4923,N_4119,N_4275);
and U4924 (N_4924,N_4268,N_4276);
nor U4925 (N_4925,N_4269,N_4331);
nand U4926 (N_4926,N_4162,N_4159);
and U4927 (N_4927,N_4361,N_4411);
nor U4928 (N_4928,N_4124,N_4187);
nand U4929 (N_4929,N_4480,N_4069);
and U4930 (N_4930,N_4491,N_4106);
xor U4931 (N_4931,N_4166,N_4394);
and U4932 (N_4932,N_4483,N_4238);
or U4933 (N_4933,N_4447,N_4325);
nand U4934 (N_4934,N_4461,N_4137);
nand U4935 (N_4935,N_4004,N_4075);
nor U4936 (N_4936,N_4169,N_4414);
nor U4937 (N_4937,N_4246,N_4196);
or U4938 (N_4938,N_4307,N_4381);
and U4939 (N_4939,N_4459,N_4329);
or U4940 (N_4940,N_4462,N_4223);
nor U4941 (N_4941,N_4489,N_4283);
nand U4942 (N_4942,N_4486,N_4433);
nor U4943 (N_4943,N_4406,N_4257);
and U4944 (N_4944,N_4013,N_4214);
nor U4945 (N_4945,N_4192,N_4142);
nor U4946 (N_4946,N_4401,N_4404);
nand U4947 (N_4947,N_4364,N_4265);
nand U4948 (N_4948,N_4097,N_4074);
nand U4949 (N_4949,N_4079,N_4261);
nand U4950 (N_4950,N_4065,N_4443);
nand U4951 (N_4951,N_4259,N_4417);
nor U4952 (N_4952,N_4136,N_4007);
and U4953 (N_4953,N_4275,N_4169);
or U4954 (N_4954,N_4432,N_4083);
or U4955 (N_4955,N_4152,N_4114);
and U4956 (N_4956,N_4000,N_4173);
nand U4957 (N_4957,N_4015,N_4310);
nor U4958 (N_4958,N_4465,N_4319);
and U4959 (N_4959,N_4163,N_4364);
and U4960 (N_4960,N_4004,N_4435);
nor U4961 (N_4961,N_4054,N_4165);
xor U4962 (N_4962,N_4242,N_4273);
nand U4963 (N_4963,N_4295,N_4300);
nand U4964 (N_4964,N_4137,N_4127);
nand U4965 (N_4965,N_4158,N_4445);
or U4966 (N_4966,N_4055,N_4452);
or U4967 (N_4967,N_4122,N_4046);
nand U4968 (N_4968,N_4047,N_4036);
and U4969 (N_4969,N_4362,N_4397);
and U4970 (N_4970,N_4446,N_4205);
or U4971 (N_4971,N_4275,N_4130);
and U4972 (N_4972,N_4011,N_4074);
nor U4973 (N_4973,N_4429,N_4366);
nor U4974 (N_4974,N_4311,N_4083);
or U4975 (N_4975,N_4403,N_4288);
nor U4976 (N_4976,N_4050,N_4328);
or U4977 (N_4977,N_4193,N_4353);
nor U4978 (N_4978,N_4164,N_4189);
or U4979 (N_4979,N_4013,N_4457);
or U4980 (N_4980,N_4424,N_4334);
and U4981 (N_4981,N_4022,N_4412);
nand U4982 (N_4982,N_4428,N_4278);
and U4983 (N_4983,N_4065,N_4157);
nand U4984 (N_4984,N_4278,N_4458);
and U4985 (N_4985,N_4450,N_4025);
or U4986 (N_4986,N_4167,N_4229);
nor U4987 (N_4987,N_4431,N_4071);
or U4988 (N_4988,N_4308,N_4187);
or U4989 (N_4989,N_4019,N_4186);
nor U4990 (N_4990,N_4458,N_4196);
xor U4991 (N_4991,N_4116,N_4435);
xnor U4992 (N_4992,N_4077,N_4400);
nor U4993 (N_4993,N_4172,N_4373);
or U4994 (N_4994,N_4396,N_4171);
or U4995 (N_4995,N_4291,N_4118);
or U4996 (N_4996,N_4123,N_4112);
xor U4997 (N_4997,N_4167,N_4160);
or U4998 (N_4998,N_4053,N_4165);
nor U4999 (N_4999,N_4062,N_4417);
nand U5000 (N_5000,N_4911,N_4829);
or U5001 (N_5001,N_4797,N_4771);
nand U5002 (N_5002,N_4934,N_4683);
nand U5003 (N_5003,N_4700,N_4912);
xor U5004 (N_5004,N_4687,N_4809);
nor U5005 (N_5005,N_4898,N_4983);
or U5006 (N_5006,N_4563,N_4559);
or U5007 (N_5007,N_4997,N_4815);
and U5008 (N_5008,N_4804,N_4745);
or U5009 (N_5009,N_4637,N_4754);
or U5010 (N_5010,N_4602,N_4735);
xor U5011 (N_5011,N_4633,N_4694);
nor U5012 (N_5012,N_4778,N_4676);
nand U5013 (N_5013,N_4550,N_4509);
and U5014 (N_5014,N_4684,N_4674);
or U5015 (N_5015,N_4869,N_4503);
nand U5016 (N_5016,N_4526,N_4714);
or U5017 (N_5017,N_4678,N_4675);
and U5018 (N_5018,N_4650,N_4781);
and U5019 (N_5019,N_4647,N_4662);
or U5020 (N_5020,N_4729,N_4882);
nor U5021 (N_5021,N_4588,N_4517);
nand U5022 (N_5022,N_4669,N_4639);
nand U5023 (N_5023,N_4516,N_4715);
nor U5024 (N_5024,N_4646,N_4685);
xnor U5025 (N_5025,N_4734,N_4884);
or U5026 (N_5026,N_4680,N_4738);
nor U5027 (N_5027,N_4641,N_4594);
xnor U5028 (N_5028,N_4887,N_4741);
nor U5029 (N_5029,N_4962,N_4765);
nand U5030 (N_5030,N_4762,N_4742);
and U5031 (N_5031,N_4699,N_4940);
and U5032 (N_5032,N_4536,N_4944);
xnor U5033 (N_5033,N_4508,N_4877);
or U5034 (N_5034,N_4981,N_4579);
and U5035 (N_5035,N_4892,N_4920);
nand U5036 (N_5036,N_4896,N_4914);
and U5037 (N_5037,N_4853,N_4731);
or U5038 (N_5038,N_4736,N_4987);
nand U5039 (N_5039,N_4514,N_4640);
nand U5040 (N_5040,N_4984,N_4750);
nor U5041 (N_5041,N_4743,N_4522);
nand U5042 (N_5042,N_4897,N_4936);
nand U5043 (N_5043,N_4533,N_4638);
or U5044 (N_5044,N_4881,N_4631);
or U5045 (N_5045,N_4969,N_4998);
and U5046 (N_5046,N_4860,N_4696);
or U5047 (N_5047,N_4621,N_4603);
nand U5048 (N_5048,N_4827,N_4961);
and U5049 (N_5049,N_4649,N_4672);
or U5050 (N_5050,N_4501,N_4928);
nor U5051 (N_5051,N_4906,N_4768);
and U5052 (N_5052,N_4937,N_4993);
nand U5053 (N_5053,N_4706,N_4659);
nand U5054 (N_5054,N_4774,N_4578);
nor U5055 (N_5055,N_4632,N_4851);
or U5056 (N_5056,N_4560,N_4974);
nand U5057 (N_5057,N_4883,N_4849);
nor U5058 (N_5058,N_4544,N_4740);
and U5059 (N_5059,N_4572,N_4567);
or U5060 (N_5060,N_4819,N_4710);
and U5061 (N_5061,N_4994,N_4599);
and U5062 (N_5062,N_4653,N_4553);
xor U5063 (N_5063,N_4719,N_4657);
xnor U5064 (N_5064,N_4842,N_4956);
nor U5065 (N_5065,N_4606,N_4978);
or U5066 (N_5066,N_4798,N_4592);
or U5067 (N_5067,N_4830,N_4823);
and U5068 (N_5068,N_4615,N_4532);
xnor U5069 (N_5069,N_4670,N_4689);
and U5070 (N_5070,N_4652,N_4767);
nor U5071 (N_5071,N_4889,N_4612);
or U5072 (N_5072,N_4856,N_4966);
or U5073 (N_5073,N_4635,N_4586);
and U5074 (N_5074,N_4521,N_4913);
and U5075 (N_5075,N_4510,N_4890);
xnor U5076 (N_5076,N_4569,N_4697);
nor U5077 (N_5077,N_4616,N_4540);
and U5078 (N_5078,N_4548,N_4874);
nor U5079 (N_5079,N_4749,N_4930);
and U5080 (N_5080,N_4722,N_4645);
and U5081 (N_5081,N_4753,N_4891);
nor U5082 (N_5082,N_4529,N_4844);
xnor U5083 (N_5083,N_4904,N_4907);
and U5084 (N_5084,N_4926,N_4681);
and U5085 (N_5085,N_4927,N_4582);
or U5086 (N_5086,N_4573,N_4859);
or U5087 (N_5087,N_4776,N_4607);
nand U5088 (N_5088,N_4620,N_4992);
and U5089 (N_5089,N_4964,N_4996);
and U5090 (N_5090,N_4702,N_4895);
and U5091 (N_5091,N_4583,N_4933);
and U5092 (N_5092,N_4945,N_4538);
nor U5093 (N_5093,N_4793,N_4910);
nor U5094 (N_5094,N_4668,N_4663);
nand U5095 (N_5095,N_4923,N_4542);
nand U5096 (N_5096,N_4739,N_4925);
xnor U5097 (N_5097,N_4772,N_4718);
or U5098 (N_5098,N_4677,N_4766);
and U5099 (N_5099,N_4693,N_4564);
and U5100 (N_5100,N_4888,N_4712);
nand U5101 (N_5101,N_4834,N_4973);
nor U5102 (N_5102,N_4979,N_4975);
and U5103 (N_5103,N_4642,N_4737);
nor U5104 (N_5104,N_4957,N_4561);
nor U5105 (N_5105,N_4502,N_4939);
nor U5106 (N_5106,N_4751,N_4618);
and U5107 (N_5107,N_4917,N_4900);
nor U5108 (N_5108,N_4658,N_4811);
and U5109 (N_5109,N_4716,N_4713);
nand U5110 (N_5110,N_4506,N_4777);
and U5111 (N_5111,N_4980,N_4717);
and U5112 (N_5112,N_4839,N_4574);
nor U5113 (N_5113,N_4836,N_4868);
or U5114 (N_5114,N_4761,N_4899);
or U5115 (N_5115,N_4863,N_4817);
nor U5116 (N_5116,N_4661,N_4565);
or U5117 (N_5117,N_4703,N_4585);
nand U5118 (N_5118,N_4549,N_4660);
nor U5119 (N_5119,N_4947,N_4946);
or U5120 (N_5120,N_4725,N_4673);
nor U5121 (N_5121,N_4518,N_4595);
and U5122 (N_5122,N_4950,N_4908);
and U5123 (N_5123,N_4786,N_4760);
nand U5124 (N_5124,N_4795,N_4698);
or U5125 (N_5125,N_4810,N_4959);
or U5126 (N_5126,N_4577,N_4512);
and U5127 (N_5127,N_4770,N_4831);
and U5128 (N_5128,N_4686,N_4720);
nor U5129 (N_5129,N_4613,N_4779);
nor U5130 (N_5130,N_4858,N_4708);
nand U5131 (N_5131,N_4832,N_4644);
or U5132 (N_5132,N_4611,N_4626);
nor U5133 (N_5133,N_4985,N_4921);
xor U5134 (N_5134,N_4692,N_4733);
nor U5135 (N_5135,N_4801,N_4763);
and U5136 (N_5136,N_4535,N_4791);
nor U5137 (N_5137,N_4551,N_4794);
nand U5138 (N_5138,N_4614,N_4664);
and U5139 (N_5139,N_4955,N_4759);
and U5140 (N_5140,N_4816,N_4593);
nor U5141 (N_5141,N_4843,N_4800);
xnor U5142 (N_5142,N_4705,N_4654);
or U5143 (N_5143,N_4787,N_4557);
nand U5144 (N_5144,N_4723,N_4814);
or U5145 (N_5145,N_4513,N_4524);
nor U5146 (N_5146,N_4840,N_4825);
and U5147 (N_5147,N_4972,N_4805);
or U5148 (N_5148,N_4764,N_4875);
xnor U5149 (N_5149,N_4905,N_4584);
nor U5150 (N_5150,N_4855,N_4628);
and U5151 (N_5151,N_4527,N_4758);
nor U5152 (N_5152,N_4977,N_4732);
nor U5153 (N_5153,N_4789,N_4576);
nand U5154 (N_5154,N_4534,N_4556);
nor U5155 (N_5155,N_4589,N_4775);
or U5156 (N_5156,N_4748,N_4916);
nand U5157 (N_5157,N_4721,N_4546);
nand U5158 (N_5158,N_4873,N_4727);
or U5159 (N_5159,N_4982,N_4746);
xor U5160 (N_5160,N_4545,N_4773);
nor U5161 (N_5161,N_4971,N_4943);
nor U5162 (N_5162,N_4951,N_4901);
nand U5163 (N_5163,N_4651,N_4818);
nand U5164 (N_5164,N_4837,N_4991);
nand U5165 (N_5165,N_4598,N_4531);
or U5166 (N_5166,N_4643,N_4747);
nand U5167 (N_5167,N_4803,N_4679);
or U5168 (N_5168,N_4952,N_4730);
and U5169 (N_5169,N_4528,N_4802);
xor U5170 (N_5170,N_4799,N_4580);
and U5171 (N_5171,N_4871,N_4539);
or U5172 (N_5172,N_4519,N_4854);
xor U5173 (N_5173,N_4924,N_4541);
xor U5174 (N_5174,N_4530,N_4704);
or U5175 (N_5175,N_4948,N_4828);
nor U5176 (N_5176,N_4630,N_4820);
and U5177 (N_5177,N_4846,N_4622);
nor U5178 (N_5178,N_4756,N_4507);
or U5179 (N_5179,N_4782,N_4941);
or U5180 (N_5180,N_4590,N_4596);
nand U5181 (N_5181,N_4505,N_4629);
nand U5182 (N_5182,N_4575,N_4990);
and U5183 (N_5183,N_4624,N_4995);
and U5184 (N_5184,N_4667,N_4872);
nor U5185 (N_5185,N_4909,N_4893);
and U5186 (N_5186,N_4543,N_4806);
or U5187 (N_5187,N_4812,N_4808);
and U5188 (N_5188,N_4835,N_4848);
nand U5189 (N_5189,N_4520,N_4619);
or U5190 (N_5190,N_4857,N_4822);
nand U5191 (N_5191,N_4785,N_4965);
nor U5192 (N_5192,N_4511,N_4870);
nand U5193 (N_5193,N_4688,N_4999);
and U5194 (N_5194,N_4783,N_4655);
or U5195 (N_5195,N_4671,N_4558);
xor U5196 (N_5196,N_4562,N_4932);
and U5197 (N_5197,N_4591,N_4570);
nor U5198 (N_5198,N_4833,N_4942);
and U5199 (N_5199,N_4864,N_4623);
nor U5200 (N_5200,N_4744,N_4821);
or U5201 (N_5201,N_4537,N_4691);
nand U5202 (N_5202,N_4610,N_4571);
nor U5203 (N_5203,N_4515,N_4903);
or U5204 (N_5204,N_4807,N_4666);
and U5205 (N_5205,N_4784,N_4880);
nand U5206 (N_5206,N_4636,N_4931);
xor U5207 (N_5207,N_4879,N_4970);
nor U5208 (N_5208,N_4597,N_4780);
nor U5209 (N_5209,N_4963,N_4876);
and U5210 (N_5210,N_4792,N_4755);
and U5211 (N_5211,N_4886,N_4852);
nand U5212 (N_5212,N_4915,N_4841);
nand U5213 (N_5213,N_4790,N_4690);
or U5214 (N_5214,N_4525,N_4878);
nor U5215 (N_5215,N_4902,N_4701);
nor U5216 (N_5216,N_4867,N_4866);
or U5217 (N_5217,N_4554,N_4935);
or U5218 (N_5218,N_4552,N_4796);
nor U5219 (N_5219,N_4711,N_4949);
nand U5220 (N_5220,N_4605,N_4919);
and U5221 (N_5221,N_4968,N_4601);
nand U5222 (N_5222,N_4728,N_4625);
nor U5223 (N_5223,N_4617,N_4695);
and U5224 (N_5224,N_4707,N_4865);
xnor U5225 (N_5225,N_4523,N_4788);
nand U5226 (N_5226,N_4634,N_4862);
nand U5227 (N_5227,N_4500,N_4954);
nor U5228 (N_5228,N_4838,N_4918);
xnor U5229 (N_5229,N_4845,N_4769);
nand U5230 (N_5230,N_4555,N_4976);
or U5231 (N_5231,N_4608,N_4953);
and U5232 (N_5232,N_4587,N_4988);
and U5233 (N_5233,N_4504,N_4894);
nor U5234 (N_5234,N_4627,N_4568);
nor U5235 (N_5235,N_4960,N_4682);
nand U5236 (N_5236,N_4813,N_4989);
nand U5237 (N_5237,N_4566,N_4958);
or U5238 (N_5238,N_4604,N_4922);
and U5239 (N_5239,N_4724,N_4967);
nand U5240 (N_5240,N_4726,N_4757);
or U5241 (N_5241,N_4656,N_4600);
nor U5242 (N_5242,N_4709,N_4752);
or U5243 (N_5243,N_4847,N_4938);
nor U5244 (N_5244,N_4665,N_4826);
xnor U5245 (N_5245,N_4861,N_4581);
nor U5246 (N_5246,N_4547,N_4648);
nor U5247 (N_5247,N_4929,N_4850);
xnor U5248 (N_5248,N_4986,N_4885);
and U5249 (N_5249,N_4824,N_4609);
nand U5250 (N_5250,N_4821,N_4670);
or U5251 (N_5251,N_4841,N_4560);
and U5252 (N_5252,N_4605,N_4827);
or U5253 (N_5253,N_4530,N_4528);
or U5254 (N_5254,N_4821,N_4901);
or U5255 (N_5255,N_4754,N_4831);
or U5256 (N_5256,N_4844,N_4537);
and U5257 (N_5257,N_4643,N_4991);
and U5258 (N_5258,N_4986,N_4739);
nand U5259 (N_5259,N_4712,N_4846);
nor U5260 (N_5260,N_4899,N_4742);
and U5261 (N_5261,N_4812,N_4565);
nand U5262 (N_5262,N_4653,N_4630);
and U5263 (N_5263,N_4510,N_4962);
and U5264 (N_5264,N_4559,N_4757);
and U5265 (N_5265,N_4613,N_4603);
xnor U5266 (N_5266,N_4598,N_4953);
and U5267 (N_5267,N_4645,N_4616);
nor U5268 (N_5268,N_4815,N_4982);
nor U5269 (N_5269,N_4894,N_4831);
and U5270 (N_5270,N_4827,N_4933);
or U5271 (N_5271,N_4648,N_4595);
nor U5272 (N_5272,N_4867,N_4679);
or U5273 (N_5273,N_4651,N_4606);
or U5274 (N_5274,N_4542,N_4968);
nor U5275 (N_5275,N_4975,N_4841);
nand U5276 (N_5276,N_4562,N_4953);
and U5277 (N_5277,N_4973,N_4613);
or U5278 (N_5278,N_4789,N_4863);
and U5279 (N_5279,N_4794,N_4672);
and U5280 (N_5280,N_4664,N_4801);
or U5281 (N_5281,N_4678,N_4611);
nor U5282 (N_5282,N_4567,N_4807);
nor U5283 (N_5283,N_4669,N_4540);
and U5284 (N_5284,N_4652,N_4832);
xnor U5285 (N_5285,N_4583,N_4724);
and U5286 (N_5286,N_4907,N_4820);
or U5287 (N_5287,N_4952,N_4940);
nor U5288 (N_5288,N_4618,N_4928);
or U5289 (N_5289,N_4699,N_4903);
or U5290 (N_5290,N_4795,N_4998);
xnor U5291 (N_5291,N_4765,N_4949);
nor U5292 (N_5292,N_4837,N_4956);
nor U5293 (N_5293,N_4527,N_4923);
xor U5294 (N_5294,N_4672,N_4858);
nand U5295 (N_5295,N_4651,N_4614);
and U5296 (N_5296,N_4673,N_4574);
or U5297 (N_5297,N_4694,N_4656);
and U5298 (N_5298,N_4862,N_4742);
nand U5299 (N_5299,N_4742,N_4826);
nand U5300 (N_5300,N_4817,N_4540);
and U5301 (N_5301,N_4960,N_4730);
or U5302 (N_5302,N_4728,N_4614);
xor U5303 (N_5303,N_4861,N_4805);
nand U5304 (N_5304,N_4681,N_4921);
nor U5305 (N_5305,N_4933,N_4908);
nand U5306 (N_5306,N_4744,N_4849);
or U5307 (N_5307,N_4904,N_4501);
nand U5308 (N_5308,N_4752,N_4872);
or U5309 (N_5309,N_4710,N_4584);
and U5310 (N_5310,N_4789,N_4903);
or U5311 (N_5311,N_4977,N_4767);
and U5312 (N_5312,N_4790,N_4640);
nand U5313 (N_5313,N_4765,N_4604);
nand U5314 (N_5314,N_4817,N_4826);
nor U5315 (N_5315,N_4894,N_4780);
or U5316 (N_5316,N_4543,N_4689);
nand U5317 (N_5317,N_4703,N_4573);
nor U5318 (N_5318,N_4687,N_4828);
or U5319 (N_5319,N_4584,N_4908);
and U5320 (N_5320,N_4845,N_4698);
nand U5321 (N_5321,N_4677,N_4502);
nor U5322 (N_5322,N_4844,N_4963);
nor U5323 (N_5323,N_4519,N_4980);
nor U5324 (N_5324,N_4788,N_4890);
and U5325 (N_5325,N_4825,N_4846);
and U5326 (N_5326,N_4897,N_4549);
and U5327 (N_5327,N_4566,N_4586);
and U5328 (N_5328,N_4806,N_4680);
xnor U5329 (N_5329,N_4815,N_4956);
or U5330 (N_5330,N_4995,N_4783);
and U5331 (N_5331,N_4527,N_4559);
nor U5332 (N_5332,N_4596,N_4836);
nand U5333 (N_5333,N_4560,N_4697);
or U5334 (N_5334,N_4577,N_4924);
or U5335 (N_5335,N_4642,N_4722);
xor U5336 (N_5336,N_4895,N_4804);
or U5337 (N_5337,N_4710,N_4975);
nor U5338 (N_5338,N_4599,N_4500);
and U5339 (N_5339,N_4854,N_4909);
xor U5340 (N_5340,N_4727,N_4535);
and U5341 (N_5341,N_4567,N_4584);
nor U5342 (N_5342,N_4872,N_4688);
xnor U5343 (N_5343,N_4649,N_4794);
and U5344 (N_5344,N_4609,N_4980);
and U5345 (N_5345,N_4743,N_4545);
nand U5346 (N_5346,N_4822,N_4660);
nor U5347 (N_5347,N_4646,N_4531);
nand U5348 (N_5348,N_4687,N_4615);
nor U5349 (N_5349,N_4802,N_4796);
or U5350 (N_5350,N_4721,N_4967);
nand U5351 (N_5351,N_4793,N_4897);
or U5352 (N_5352,N_4729,N_4563);
or U5353 (N_5353,N_4863,N_4738);
xnor U5354 (N_5354,N_4552,N_4768);
xor U5355 (N_5355,N_4566,N_4806);
nor U5356 (N_5356,N_4661,N_4584);
nor U5357 (N_5357,N_4661,N_4751);
nand U5358 (N_5358,N_4993,N_4888);
or U5359 (N_5359,N_4596,N_4926);
nor U5360 (N_5360,N_4730,N_4687);
nand U5361 (N_5361,N_4611,N_4742);
and U5362 (N_5362,N_4914,N_4929);
xnor U5363 (N_5363,N_4855,N_4643);
nand U5364 (N_5364,N_4596,N_4665);
nand U5365 (N_5365,N_4749,N_4925);
xor U5366 (N_5366,N_4604,N_4545);
xnor U5367 (N_5367,N_4809,N_4876);
nand U5368 (N_5368,N_4807,N_4701);
and U5369 (N_5369,N_4975,N_4509);
nand U5370 (N_5370,N_4720,N_4561);
nor U5371 (N_5371,N_4961,N_4580);
nor U5372 (N_5372,N_4938,N_4810);
xnor U5373 (N_5373,N_4508,N_4685);
nand U5374 (N_5374,N_4724,N_4668);
or U5375 (N_5375,N_4977,N_4548);
nor U5376 (N_5376,N_4841,N_4837);
or U5377 (N_5377,N_4620,N_4909);
nand U5378 (N_5378,N_4646,N_4542);
nand U5379 (N_5379,N_4538,N_4548);
and U5380 (N_5380,N_4670,N_4644);
nand U5381 (N_5381,N_4919,N_4687);
or U5382 (N_5382,N_4947,N_4787);
and U5383 (N_5383,N_4639,N_4672);
nand U5384 (N_5384,N_4682,N_4931);
xnor U5385 (N_5385,N_4518,N_4636);
nand U5386 (N_5386,N_4951,N_4800);
or U5387 (N_5387,N_4671,N_4761);
nand U5388 (N_5388,N_4569,N_4824);
nand U5389 (N_5389,N_4938,N_4944);
nor U5390 (N_5390,N_4587,N_4509);
nand U5391 (N_5391,N_4948,N_4714);
nor U5392 (N_5392,N_4758,N_4890);
and U5393 (N_5393,N_4686,N_4891);
xor U5394 (N_5394,N_4930,N_4507);
nand U5395 (N_5395,N_4859,N_4875);
and U5396 (N_5396,N_4654,N_4902);
nor U5397 (N_5397,N_4926,N_4573);
nand U5398 (N_5398,N_4908,N_4794);
nor U5399 (N_5399,N_4908,N_4678);
and U5400 (N_5400,N_4810,N_4554);
and U5401 (N_5401,N_4501,N_4804);
nand U5402 (N_5402,N_4964,N_4590);
and U5403 (N_5403,N_4933,N_4608);
nand U5404 (N_5404,N_4616,N_4757);
nand U5405 (N_5405,N_4797,N_4977);
nor U5406 (N_5406,N_4518,N_4863);
and U5407 (N_5407,N_4956,N_4660);
nor U5408 (N_5408,N_4990,N_4583);
or U5409 (N_5409,N_4600,N_4834);
nand U5410 (N_5410,N_4809,N_4804);
xnor U5411 (N_5411,N_4890,N_4648);
nor U5412 (N_5412,N_4959,N_4737);
and U5413 (N_5413,N_4605,N_4635);
nand U5414 (N_5414,N_4981,N_4607);
or U5415 (N_5415,N_4793,N_4675);
or U5416 (N_5416,N_4503,N_4863);
nand U5417 (N_5417,N_4745,N_4547);
and U5418 (N_5418,N_4812,N_4743);
or U5419 (N_5419,N_4609,N_4893);
nand U5420 (N_5420,N_4941,N_4730);
nand U5421 (N_5421,N_4927,N_4806);
or U5422 (N_5422,N_4883,N_4965);
nor U5423 (N_5423,N_4816,N_4944);
or U5424 (N_5424,N_4674,N_4580);
and U5425 (N_5425,N_4584,N_4711);
or U5426 (N_5426,N_4695,N_4863);
or U5427 (N_5427,N_4903,N_4952);
xnor U5428 (N_5428,N_4605,N_4843);
nor U5429 (N_5429,N_4526,N_4771);
or U5430 (N_5430,N_4518,N_4613);
nor U5431 (N_5431,N_4708,N_4523);
nand U5432 (N_5432,N_4573,N_4638);
nand U5433 (N_5433,N_4513,N_4742);
nand U5434 (N_5434,N_4839,N_4624);
nand U5435 (N_5435,N_4867,N_4803);
nand U5436 (N_5436,N_4808,N_4532);
nand U5437 (N_5437,N_4906,N_4885);
xnor U5438 (N_5438,N_4733,N_4941);
nand U5439 (N_5439,N_4933,N_4805);
and U5440 (N_5440,N_4710,N_4602);
nand U5441 (N_5441,N_4962,N_4950);
or U5442 (N_5442,N_4956,N_4866);
nand U5443 (N_5443,N_4787,N_4649);
nor U5444 (N_5444,N_4834,N_4539);
nor U5445 (N_5445,N_4505,N_4695);
nand U5446 (N_5446,N_4715,N_4957);
and U5447 (N_5447,N_4751,N_4627);
and U5448 (N_5448,N_4926,N_4788);
nor U5449 (N_5449,N_4689,N_4821);
nand U5450 (N_5450,N_4921,N_4823);
nor U5451 (N_5451,N_4745,N_4587);
nand U5452 (N_5452,N_4872,N_4689);
and U5453 (N_5453,N_4690,N_4570);
nand U5454 (N_5454,N_4889,N_4524);
or U5455 (N_5455,N_4625,N_4962);
or U5456 (N_5456,N_4619,N_4894);
nand U5457 (N_5457,N_4954,N_4737);
nor U5458 (N_5458,N_4858,N_4503);
nor U5459 (N_5459,N_4820,N_4649);
and U5460 (N_5460,N_4973,N_4816);
nor U5461 (N_5461,N_4970,N_4678);
nand U5462 (N_5462,N_4586,N_4501);
nand U5463 (N_5463,N_4671,N_4816);
or U5464 (N_5464,N_4918,N_4709);
and U5465 (N_5465,N_4884,N_4689);
nor U5466 (N_5466,N_4626,N_4613);
nand U5467 (N_5467,N_4614,N_4522);
and U5468 (N_5468,N_4536,N_4896);
nand U5469 (N_5469,N_4691,N_4505);
or U5470 (N_5470,N_4677,N_4534);
and U5471 (N_5471,N_4688,N_4560);
nand U5472 (N_5472,N_4640,N_4761);
nand U5473 (N_5473,N_4899,N_4516);
nand U5474 (N_5474,N_4570,N_4876);
or U5475 (N_5475,N_4863,N_4857);
or U5476 (N_5476,N_4685,N_4581);
or U5477 (N_5477,N_4711,N_4572);
nand U5478 (N_5478,N_4590,N_4553);
nand U5479 (N_5479,N_4623,N_4775);
or U5480 (N_5480,N_4963,N_4979);
xor U5481 (N_5481,N_4812,N_4966);
xor U5482 (N_5482,N_4568,N_4527);
nand U5483 (N_5483,N_4704,N_4896);
and U5484 (N_5484,N_4989,N_4643);
and U5485 (N_5485,N_4597,N_4697);
nor U5486 (N_5486,N_4972,N_4913);
nand U5487 (N_5487,N_4850,N_4912);
nor U5488 (N_5488,N_4689,N_4549);
nand U5489 (N_5489,N_4593,N_4698);
nand U5490 (N_5490,N_4599,N_4935);
nand U5491 (N_5491,N_4781,N_4804);
nand U5492 (N_5492,N_4950,N_4570);
nor U5493 (N_5493,N_4979,N_4992);
nand U5494 (N_5494,N_4728,N_4973);
nor U5495 (N_5495,N_4557,N_4870);
nand U5496 (N_5496,N_4670,N_4665);
nor U5497 (N_5497,N_4553,N_4556);
and U5498 (N_5498,N_4867,N_4706);
nor U5499 (N_5499,N_4757,N_4752);
xor U5500 (N_5500,N_5130,N_5327);
nor U5501 (N_5501,N_5056,N_5418);
and U5502 (N_5502,N_5334,N_5459);
nor U5503 (N_5503,N_5426,N_5373);
nor U5504 (N_5504,N_5076,N_5149);
and U5505 (N_5505,N_5068,N_5018);
nor U5506 (N_5506,N_5410,N_5131);
nand U5507 (N_5507,N_5361,N_5235);
xor U5508 (N_5508,N_5041,N_5246);
nor U5509 (N_5509,N_5178,N_5071);
or U5510 (N_5510,N_5431,N_5318);
and U5511 (N_5511,N_5374,N_5198);
and U5512 (N_5512,N_5357,N_5103);
nand U5513 (N_5513,N_5417,N_5155);
and U5514 (N_5514,N_5030,N_5263);
nand U5515 (N_5515,N_5013,N_5218);
nor U5516 (N_5516,N_5236,N_5256);
xor U5517 (N_5517,N_5341,N_5368);
and U5518 (N_5518,N_5465,N_5183);
and U5519 (N_5519,N_5480,N_5483);
nor U5520 (N_5520,N_5231,N_5194);
and U5521 (N_5521,N_5355,N_5358);
nor U5522 (N_5522,N_5162,N_5296);
nand U5523 (N_5523,N_5190,N_5458);
nor U5524 (N_5524,N_5478,N_5299);
nand U5525 (N_5525,N_5436,N_5451);
and U5526 (N_5526,N_5192,N_5435);
nand U5527 (N_5527,N_5234,N_5464);
and U5528 (N_5528,N_5012,N_5281);
and U5529 (N_5529,N_5081,N_5058);
or U5530 (N_5530,N_5269,N_5353);
nor U5531 (N_5531,N_5019,N_5031);
or U5532 (N_5532,N_5287,N_5101);
and U5533 (N_5533,N_5278,N_5216);
nand U5534 (N_5534,N_5224,N_5188);
or U5535 (N_5535,N_5348,N_5365);
nor U5536 (N_5536,N_5481,N_5331);
nand U5537 (N_5537,N_5199,N_5185);
and U5538 (N_5538,N_5412,N_5051);
xor U5539 (N_5539,N_5083,N_5364);
or U5540 (N_5540,N_5390,N_5320);
and U5541 (N_5541,N_5238,N_5028);
nand U5542 (N_5542,N_5105,N_5266);
nor U5543 (N_5543,N_5273,N_5466);
nor U5544 (N_5544,N_5042,N_5387);
and U5545 (N_5545,N_5469,N_5289);
nand U5546 (N_5546,N_5453,N_5124);
nor U5547 (N_5547,N_5401,N_5180);
nand U5548 (N_5548,N_5247,N_5409);
nand U5549 (N_5549,N_5326,N_5118);
nor U5550 (N_5550,N_5148,N_5021);
nor U5551 (N_5551,N_5027,N_5475);
nor U5552 (N_5552,N_5448,N_5277);
nand U5553 (N_5553,N_5145,N_5422);
nor U5554 (N_5554,N_5170,N_5315);
or U5555 (N_5555,N_5322,N_5164);
or U5556 (N_5556,N_5097,N_5311);
and U5557 (N_5557,N_5074,N_5110);
nor U5558 (N_5558,N_5008,N_5065);
or U5559 (N_5559,N_5457,N_5053);
xor U5560 (N_5560,N_5111,N_5154);
nand U5561 (N_5561,N_5034,N_5203);
and U5562 (N_5562,N_5158,N_5383);
nand U5563 (N_5563,N_5079,N_5182);
xor U5564 (N_5564,N_5086,N_5445);
and U5565 (N_5565,N_5474,N_5352);
nand U5566 (N_5566,N_5085,N_5020);
and U5567 (N_5567,N_5156,N_5078);
nand U5568 (N_5568,N_5191,N_5408);
or U5569 (N_5569,N_5228,N_5347);
and U5570 (N_5570,N_5396,N_5283);
or U5571 (N_5571,N_5036,N_5276);
nand U5572 (N_5572,N_5169,N_5195);
nand U5573 (N_5573,N_5305,N_5395);
and U5574 (N_5574,N_5415,N_5439);
or U5575 (N_5575,N_5039,N_5398);
nor U5576 (N_5576,N_5279,N_5212);
nor U5577 (N_5577,N_5225,N_5485);
xnor U5578 (N_5578,N_5217,N_5179);
and U5579 (N_5579,N_5015,N_5397);
nand U5580 (N_5580,N_5386,N_5423);
nand U5581 (N_5581,N_5389,N_5215);
xnor U5582 (N_5582,N_5437,N_5119);
xnor U5583 (N_5583,N_5023,N_5494);
or U5584 (N_5584,N_5239,N_5159);
or U5585 (N_5585,N_5025,N_5092);
or U5586 (N_5586,N_5425,N_5443);
or U5587 (N_5587,N_5297,N_5440);
nand U5588 (N_5588,N_5282,N_5112);
nor U5589 (N_5589,N_5043,N_5167);
nand U5590 (N_5590,N_5172,N_5360);
and U5591 (N_5591,N_5377,N_5244);
and U5592 (N_5592,N_5161,N_5223);
xor U5593 (N_5593,N_5399,N_5057);
or U5594 (N_5594,N_5454,N_5343);
or U5595 (N_5595,N_5120,N_5226);
and U5596 (N_5596,N_5173,N_5220);
nor U5597 (N_5597,N_5370,N_5432);
nand U5598 (N_5598,N_5006,N_5288);
or U5599 (N_5599,N_5460,N_5496);
or U5600 (N_5600,N_5104,N_5292);
and U5601 (N_5601,N_5487,N_5301);
nor U5602 (N_5602,N_5227,N_5242);
or U5603 (N_5603,N_5241,N_5163);
or U5604 (N_5604,N_5424,N_5325);
and U5605 (N_5605,N_5003,N_5196);
xnor U5606 (N_5606,N_5243,N_5367);
nand U5607 (N_5607,N_5047,N_5268);
nand U5608 (N_5608,N_5264,N_5251);
and U5609 (N_5609,N_5142,N_5147);
nor U5610 (N_5610,N_5267,N_5314);
nand U5611 (N_5611,N_5116,N_5486);
and U5612 (N_5612,N_5088,N_5274);
and U5613 (N_5613,N_5403,N_5202);
and U5614 (N_5614,N_5113,N_5321);
xnor U5615 (N_5615,N_5265,N_5477);
nor U5616 (N_5616,N_5095,N_5333);
or U5617 (N_5617,N_5467,N_5309);
xnor U5618 (N_5618,N_5446,N_5463);
nor U5619 (N_5619,N_5029,N_5392);
nand U5620 (N_5620,N_5050,N_5026);
xor U5621 (N_5621,N_5302,N_5349);
nand U5622 (N_5622,N_5254,N_5004);
and U5623 (N_5623,N_5313,N_5052);
nand U5624 (N_5624,N_5329,N_5328);
or U5625 (N_5625,N_5488,N_5099);
xnor U5626 (N_5626,N_5260,N_5186);
xnor U5627 (N_5627,N_5100,N_5259);
nor U5628 (N_5628,N_5064,N_5298);
and U5629 (N_5629,N_5080,N_5175);
or U5630 (N_5630,N_5232,N_5022);
and U5631 (N_5631,N_5339,N_5428);
or U5632 (N_5632,N_5461,N_5093);
nand U5633 (N_5633,N_5109,N_5338);
or U5634 (N_5634,N_5310,N_5354);
or U5635 (N_5635,N_5084,N_5127);
or U5636 (N_5636,N_5014,N_5449);
xor U5637 (N_5637,N_5070,N_5204);
or U5638 (N_5638,N_5157,N_5306);
or U5639 (N_5639,N_5121,N_5324);
nor U5640 (N_5640,N_5429,N_5344);
and U5641 (N_5641,N_5427,N_5498);
and U5642 (N_5642,N_5146,N_5342);
and U5643 (N_5643,N_5055,N_5197);
or U5644 (N_5644,N_5107,N_5420);
or U5645 (N_5645,N_5416,N_5010);
nor U5646 (N_5646,N_5211,N_5054);
nand U5647 (N_5647,N_5441,N_5316);
nand U5648 (N_5648,N_5049,N_5400);
nor U5649 (N_5649,N_5061,N_5059);
nor U5650 (N_5650,N_5117,N_5002);
and U5651 (N_5651,N_5304,N_5438);
nor U5652 (N_5652,N_5271,N_5140);
and U5653 (N_5653,N_5375,N_5378);
and U5654 (N_5654,N_5497,N_5152);
nand U5655 (N_5655,N_5011,N_5005);
nand U5656 (N_5656,N_5262,N_5484);
and U5657 (N_5657,N_5444,N_5091);
and U5658 (N_5658,N_5363,N_5181);
and U5659 (N_5659,N_5307,N_5456);
and U5660 (N_5660,N_5369,N_5123);
or U5661 (N_5661,N_5108,N_5136);
or U5662 (N_5662,N_5040,N_5362);
nor U5663 (N_5663,N_5490,N_5144);
nor U5664 (N_5664,N_5024,N_5221);
nor U5665 (N_5665,N_5351,N_5413);
nand U5666 (N_5666,N_5174,N_5141);
nor U5667 (N_5667,N_5462,N_5404);
nand U5668 (N_5668,N_5046,N_5405);
nand U5669 (N_5669,N_5308,N_5001);
nor U5670 (N_5670,N_5499,N_5143);
nand U5671 (N_5671,N_5138,N_5200);
or U5672 (N_5672,N_5229,N_5294);
nand U5673 (N_5673,N_5044,N_5115);
or U5674 (N_5674,N_5470,N_5219);
nor U5675 (N_5675,N_5222,N_5132);
and U5676 (N_5676,N_5067,N_5208);
and U5677 (N_5677,N_5082,N_5066);
xor U5678 (N_5678,N_5102,N_5150);
and U5679 (N_5679,N_5411,N_5009);
and U5680 (N_5680,N_5037,N_5258);
nand U5681 (N_5681,N_5089,N_5332);
or U5682 (N_5682,N_5381,N_5252);
or U5683 (N_5683,N_5330,N_5371);
or U5684 (N_5684,N_5380,N_5184);
or U5685 (N_5685,N_5452,N_5048);
nand U5686 (N_5686,N_5151,N_5176);
or U5687 (N_5687,N_5290,N_5393);
nand U5688 (N_5688,N_5319,N_5414);
nor U5689 (N_5689,N_5033,N_5245);
nor U5690 (N_5690,N_5072,N_5153);
and U5691 (N_5691,N_5406,N_5201);
nor U5692 (N_5692,N_5255,N_5275);
or U5693 (N_5693,N_5489,N_5233);
nand U5694 (N_5694,N_5062,N_5468);
nand U5695 (N_5695,N_5295,N_5210);
and U5696 (N_5696,N_5135,N_5394);
and U5697 (N_5697,N_5372,N_5060);
nand U5698 (N_5698,N_5359,N_5090);
and U5699 (N_5699,N_5495,N_5165);
and U5700 (N_5700,N_5126,N_5479);
xor U5701 (N_5701,N_5442,N_5493);
nand U5702 (N_5702,N_5000,N_5379);
and U5703 (N_5703,N_5473,N_5434);
nand U5704 (N_5704,N_5016,N_5482);
nand U5705 (N_5705,N_5450,N_5291);
nor U5706 (N_5706,N_5139,N_5335);
nand U5707 (N_5707,N_5098,N_5069);
nor U5708 (N_5708,N_5077,N_5407);
xor U5709 (N_5709,N_5376,N_5171);
nor U5710 (N_5710,N_5356,N_5384);
nand U5711 (N_5711,N_5166,N_5471);
and U5712 (N_5712,N_5286,N_5207);
xnor U5713 (N_5713,N_5209,N_5382);
and U5714 (N_5714,N_5350,N_5447);
nor U5715 (N_5715,N_5230,N_5094);
and U5716 (N_5716,N_5300,N_5293);
or U5717 (N_5717,N_5492,N_5240);
nor U5718 (N_5718,N_5032,N_5237);
or U5719 (N_5719,N_5187,N_5075);
nor U5720 (N_5720,N_5129,N_5491);
or U5721 (N_5721,N_5137,N_5270);
xnor U5722 (N_5722,N_5336,N_5285);
or U5723 (N_5723,N_5402,N_5337);
nand U5724 (N_5724,N_5193,N_5340);
and U5725 (N_5725,N_5160,N_5280);
nand U5726 (N_5726,N_5063,N_5248);
or U5727 (N_5727,N_5323,N_5205);
or U5728 (N_5728,N_5472,N_5114);
or U5729 (N_5729,N_5038,N_5096);
and U5730 (N_5730,N_5249,N_5168);
and U5731 (N_5731,N_5177,N_5303);
or U5732 (N_5732,N_5433,N_5250);
xnor U5733 (N_5733,N_5128,N_5346);
and U5734 (N_5734,N_5284,N_5133);
and U5735 (N_5735,N_5206,N_5261);
nor U5736 (N_5736,N_5122,N_5045);
nor U5737 (N_5737,N_5189,N_5430);
nand U5738 (N_5738,N_5419,N_5214);
and U5739 (N_5739,N_5125,N_5134);
or U5740 (N_5740,N_5391,N_5345);
xor U5741 (N_5741,N_5455,N_5017);
nor U5742 (N_5742,N_5366,N_5073);
nor U5743 (N_5743,N_5007,N_5253);
and U5744 (N_5744,N_5087,N_5106);
nor U5745 (N_5745,N_5385,N_5035);
nor U5746 (N_5746,N_5476,N_5317);
nand U5747 (N_5747,N_5421,N_5388);
xor U5748 (N_5748,N_5312,N_5257);
and U5749 (N_5749,N_5213,N_5272);
and U5750 (N_5750,N_5224,N_5378);
nand U5751 (N_5751,N_5420,N_5260);
or U5752 (N_5752,N_5058,N_5167);
nand U5753 (N_5753,N_5222,N_5362);
nor U5754 (N_5754,N_5044,N_5298);
or U5755 (N_5755,N_5426,N_5404);
nand U5756 (N_5756,N_5091,N_5217);
nand U5757 (N_5757,N_5144,N_5043);
nor U5758 (N_5758,N_5476,N_5213);
and U5759 (N_5759,N_5262,N_5340);
nor U5760 (N_5760,N_5120,N_5123);
nand U5761 (N_5761,N_5061,N_5405);
nand U5762 (N_5762,N_5136,N_5297);
nand U5763 (N_5763,N_5421,N_5101);
xor U5764 (N_5764,N_5437,N_5474);
or U5765 (N_5765,N_5010,N_5051);
or U5766 (N_5766,N_5414,N_5449);
nand U5767 (N_5767,N_5199,N_5426);
nor U5768 (N_5768,N_5416,N_5447);
nand U5769 (N_5769,N_5344,N_5302);
or U5770 (N_5770,N_5032,N_5246);
and U5771 (N_5771,N_5339,N_5327);
nand U5772 (N_5772,N_5208,N_5007);
and U5773 (N_5773,N_5387,N_5419);
xor U5774 (N_5774,N_5086,N_5489);
or U5775 (N_5775,N_5145,N_5401);
or U5776 (N_5776,N_5150,N_5205);
nand U5777 (N_5777,N_5008,N_5186);
nor U5778 (N_5778,N_5295,N_5427);
xnor U5779 (N_5779,N_5183,N_5217);
and U5780 (N_5780,N_5418,N_5011);
or U5781 (N_5781,N_5472,N_5434);
or U5782 (N_5782,N_5079,N_5434);
nand U5783 (N_5783,N_5191,N_5472);
or U5784 (N_5784,N_5086,N_5363);
nor U5785 (N_5785,N_5229,N_5337);
nor U5786 (N_5786,N_5031,N_5323);
nand U5787 (N_5787,N_5274,N_5422);
nand U5788 (N_5788,N_5026,N_5339);
xnor U5789 (N_5789,N_5193,N_5268);
xnor U5790 (N_5790,N_5132,N_5418);
xnor U5791 (N_5791,N_5370,N_5112);
nand U5792 (N_5792,N_5212,N_5243);
and U5793 (N_5793,N_5332,N_5179);
or U5794 (N_5794,N_5299,N_5003);
nand U5795 (N_5795,N_5138,N_5397);
or U5796 (N_5796,N_5433,N_5295);
or U5797 (N_5797,N_5113,N_5377);
or U5798 (N_5798,N_5070,N_5265);
nand U5799 (N_5799,N_5188,N_5076);
nor U5800 (N_5800,N_5026,N_5412);
nor U5801 (N_5801,N_5272,N_5316);
or U5802 (N_5802,N_5445,N_5390);
or U5803 (N_5803,N_5077,N_5280);
nand U5804 (N_5804,N_5069,N_5007);
xor U5805 (N_5805,N_5021,N_5381);
or U5806 (N_5806,N_5484,N_5300);
xnor U5807 (N_5807,N_5487,N_5230);
and U5808 (N_5808,N_5398,N_5437);
or U5809 (N_5809,N_5443,N_5202);
and U5810 (N_5810,N_5316,N_5148);
and U5811 (N_5811,N_5038,N_5276);
xor U5812 (N_5812,N_5352,N_5200);
xnor U5813 (N_5813,N_5359,N_5495);
xor U5814 (N_5814,N_5157,N_5268);
nor U5815 (N_5815,N_5171,N_5381);
and U5816 (N_5816,N_5243,N_5001);
and U5817 (N_5817,N_5262,N_5372);
nand U5818 (N_5818,N_5155,N_5305);
nand U5819 (N_5819,N_5249,N_5328);
nand U5820 (N_5820,N_5122,N_5249);
nand U5821 (N_5821,N_5391,N_5078);
and U5822 (N_5822,N_5468,N_5251);
and U5823 (N_5823,N_5106,N_5347);
and U5824 (N_5824,N_5210,N_5258);
or U5825 (N_5825,N_5038,N_5089);
nor U5826 (N_5826,N_5372,N_5289);
nand U5827 (N_5827,N_5309,N_5157);
or U5828 (N_5828,N_5227,N_5280);
nor U5829 (N_5829,N_5284,N_5095);
nand U5830 (N_5830,N_5210,N_5352);
nor U5831 (N_5831,N_5403,N_5416);
nor U5832 (N_5832,N_5354,N_5186);
nand U5833 (N_5833,N_5181,N_5067);
xor U5834 (N_5834,N_5447,N_5042);
nor U5835 (N_5835,N_5314,N_5381);
nor U5836 (N_5836,N_5040,N_5391);
nand U5837 (N_5837,N_5005,N_5293);
nand U5838 (N_5838,N_5141,N_5415);
nand U5839 (N_5839,N_5447,N_5221);
xnor U5840 (N_5840,N_5269,N_5446);
nor U5841 (N_5841,N_5113,N_5320);
and U5842 (N_5842,N_5099,N_5429);
nand U5843 (N_5843,N_5346,N_5430);
nand U5844 (N_5844,N_5172,N_5223);
nor U5845 (N_5845,N_5343,N_5336);
nor U5846 (N_5846,N_5212,N_5091);
xor U5847 (N_5847,N_5070,N_5482);
nor U5848 (N_5848,N_5302,N_5283);
and U5849 (N_5849,N_5187,N_5236);
nor U5850 (N_5850,N_5438,N_5293);
and U5851 (N_5851,N_5093,N_5211);
nand U5852 (N_5852,N_5043,N_5444);
xor U5853 (N_5853,N_5351,N_5140);
xor U5854 (N_5854,N_5194,N_5201);
nor U5855 (N_5855,N_5331,N_5223);
nand U5856 (N_5856,N_5438,N_5346);
nor U5857 (N_5857,N_5099,N_5042);
nor U5858 (N_5858,N_5266,N_5097);
and U5859 (N_5859,N_5309,N_5143);
and U5860 (N_5860,N_5148,N_5292);
nand U5861 (N_5861,N_5493,N_5105);
nand U5862 (N_5862,N_5176,N_5431);
and U5863 (N_5863,N_5308,N_5458);
nand U5864 (N_5864,N_5038,N_5218);
and U5865 (N_5865,N_5497,N_5085);
nand U5866 (N_5866,N_5260,N_5067);
xor U5867 (N_5867,N_5419,N_5455);
or U5868 (N_5868,N_5340,N_5327);
nand U5869 (N_5869,N_5170,N_5049);
xor U5870 (N_5870,N_5200,N_5306);
and U5871 (N_5871,N_5374,N_5185);
nand U5872 (N_5872,N_5370,N_5258);
nor U5873 (N_5873,N_5006,N_5493);
or U5874 (N_5874,N_5467,N_5375);
or U5875 (N_5875,N_5408,N_5489);
nand U5876 (N_5876,N_5126,N_5122);
and U5877 (N_5877,N_5389,N_5351);
and U5878 (N_5878,N_5364,N_5112);
nand U5879 (N_5879,N_5250,N_5124);
or U5880 (N_5880,N_5376,N_5137);
and U5881 (N_5881,N_5256,N_5022);
and U5882 (N_5882,N_5114,N_5142);
xor U5883 (N_5883,N_5436,N_5372);
and U5884 (N_5884,N_5265,N_5146);
nand U5885 (N_5885,N_5053,N_5491);
or U5886 (N_5886,N_5200,N_5298);
or U5887 (N_5887,N_5215,N_5237);
xnor U5888 (N_5888,N_5176,N_5244);
and U5889 (N_5889,N_5186,N_5352);
nand U5890 (N_5890,N_5385,N_5205);
xnor U5891 (N_5891,N_5419,N_5452);
nand U5892 (N_5892,N_5373,N_5177);
nor U5893 (N_5893,N_5143,N_5166);
nor U5894 (N_5894,N_5073,N_5355);
nor U5895 (N_5895,N_5190,N_5480);
nand U5896 (N_5896,N_5364,N_5021);
nor U5897 (N_5897,N_5026,N_5356);
xnor U5898 (N_5898,N_5455,N_5408);
nand U5899 (N_5899,N_5266,N_5430);
xnor U5900 (N_5900,N_5160,N_5393);
or U5901 (N_5901,N_5080,N_5126);
nor U5902 (N_5902,N_5146,N_5460);
nor U5903 (N_5903,N_5201,N_5138);
nor U5904 (N_5904,N_5161,N_5469);
nand U5905 (N_5905,N_5474,N_5357);
or U5906 (N_5906,N_5466,N_5371);
nand U5907 (N_5907,N_5190,N_5140);
or U5908 (N_5908,N_5217,N_5340);
nand U5909 (N_5909,N_5169,N_5378);
xor U5910 (N_5910,N_5326,N_5036);
and U5911 (N_5911,N_5285,N_5352);
and U5912 (N_5912,N_5259,N_5287);
xnor U5913 (N_5913,N_5030,N_5321);
and U5914 (N_5914,N_5042,N_5082);
or U5915 (N_5915,N_5465,N_5185);
or U5916 (N_5916,N_5292,N_5095);
nand U5917 (N_5917,N_5048,N_5119);
or U5918 (N_5918,N_5185,N_5314);
and U5919 (N_5919,N_5048,N_5237);
or U5920 (N_5920,N_5008,N_5185);
and U5921 (N_5921,N_5305,N_5312);
or U5922 (N_5922,N_5066,N_5210);
nand U5923 (N_5923,N_5364,N_5105);
xnor U5924 (N_5924,N_5150,N_5066);
and U5925 (N_5925,N_5188,N_5299);
or U5926 (N_5926,N_5021,N_5444);
nor U5927 (N_5927,N_5313,N_5230);
xor U5928 (N_5928,N_5186,N_5170);
or U5929 (N_5929,N_5238,N_5413);
xnor U5930 (N_5930,N_5194,N_5381);
nand U5931 (N_5931,N_5046,N_5114);
nor U5932 (N_5932,N_5477,N_5388);
or U5933 (N_5933,N_5063,N_5411);
or U5934 (N_5934,N_5132,N_5403);
and U5935 (N_5935,N_5158,N_5238);
xnor U5936 (N_5936,N_5378,N_5270);
nor U5937 (N_5937,N_5026,N_5199);
nand U5938 (N_5938,N_5248,N_5430);
nand U5939 (N_5939,N_5238,N_5032);
or U5940 (N_5940,N_5142,N_5173);
nor U5941 (N_5941,N_5216,N_5063);
nor U5942 (N_5942,N_5236,N_5315);
nand U5943 (N_5943,N_5123,N_5433);
or U5944 (N_5944,N_5217,N_5241);
nor U5945 (N_5945,N_5288,N_5017);
or U5946 (N_5946,N_5215,N_5405);
and U5947 (N_5947,N_5440,N_5076);
nand U5948 (N_5948,N_5118,N_5199);
nor U5949 (N_5949,N_5064,N_5367);
nand U5950 (N_5950,N_5173,N_5429);
or U5951 (N_5951,N_5098,N_5381);
xnor U5952 (N_5952,N_5011,N_5134);
nand U5953 (N_5953,N_5095,N_5454);
or U5954 (N_5954,N_5276,N_5103);
and U5955 (N_5955,N_5280,N_5382);
nor U5956 (N_5956,N_5268,N_5411);
nand U5957 (N_5957,N_5120,N_5485);
nand U5958 (N_5958,N_5403,N_5147);
nand U5959 (N_5959,N_5193,N_5044);
nand U5960 (N_5960,N_5217,N_5022);
xor U5961 (N_5961,N_5332,N_5181);
or U5962 (N_5962,N_5462,N_5366);
nand U5963 (N_5963,N_5315,N_5291);
and U5964 (N_5964,N_5061,N_5131);
nor U5965 (N_5965,N_5013,N_5030);
nand U5966 (N_5966,N_5105,N_5122);
nor U5967 (N_5967,N_5234,N_5354);
nor U5968 (N_5968,N_5471,N_5089);
nand U5969 (N_5969,N_5243,N_5029);
or U5970 (N_5970,N_5272,N_5394);
or U5971 (N_5971,N_5294,N_5379);
nand U5972 (N_5972,N_5258,N_5403);
or U5973 (N_5973,N_5482,N_5416);
and U5974 (N_5974,N_5415,N_5485);
or U5975 (N_5975,N_5151,N_5171);
nor U5976 (N_5976,N_5259,N_5044);
nor U5977 (N_5977,N_5465,N_5178);
nor U5978 (N_5978,N_5225,N_5244);
nand U5979 (N_5979,N_5491,N_5158);
xor U5980 (N_5980,N_5208,N_5256);
or U5981 (N_5981,N_5252,N_5287);
and U5982 (N_5982,N_5440,N_5291);
nor U5983 (N_5983,N_5200,N_5165);
nand U5984 (N_5984,N_5389,N_5052);
xnor U5985 (N_5985,N_5043,N_5495);
or U5986 (N_5986,N_5336,N_5018);
or U5987 (N_5987,N_5468,N_5403);
xnor U5988 (N_5988,N_5043,N_5053);
nor U5989 (N_5989,N_5308,N_5447);
or U5990 (N_5990,N_5397,N_5031);
nor U5991 (N_5991,N_5003,N_5070);
and U5992 (N_5992,N_5412,N_5311);
nor U5993 (N_5993,N_5470,N_5006);
or U5994 (N_5994,N_5200,N_5076);
or U5995 (N_5995,N_5064,N_5035);
nand U5996 (N_5996,N_5328,N_5027);
or U5997 (N_5997,N_5083,N_5190);
nand U5998 (N_5998,N_5156,N_5079);
nor U5999 (N_5999,N_5151,N_5403);
nor U6000 (N_6000,N_5718,N_5768);
or U6001 (N_6001,N_5717,N_5748);
nor U6002 (N_6002,N_5599,N_5891);
and U6003 (N_6003,N_5851,N_5726);
nand U6004 (N_6004,N_5847,N_5517);
nor U6005 (N_6005,N_5567,N_5700);
nand U6006 (N_6006,N_5984,N_5765);
and U6007 (N_6007,N_5929,N_5829);
nand U6008 (N_6008,N_5825,N_5990);
nor U6009 (N_6009,N_5772,N_5606);
nand U6010 (N_6010,N_5594,N_5711);
or U6011 (N_6011,N_5786,N_5611);
nor U6012 (N_6012,N_5960,N_5645);
nand U6013 (N_6013,N_5977,N_5673);
nor U6014 (N_6014,N_5539,N_5643);
or U6015 (N_6015,N_5674,N_5936);
nor U6016 (N_6016,N_5879,N_5756);
xor U6017 (N_6017,N_5721,N_5881);
nor U6018 (N_6018,N_5576,N_5918);
xor U6019 (N_6019,N_5789,N_5507);
nor U6020 (N_6020,N_5608,N_5665);
and U6021 (N_6021,N_5569,N_5828);
xor U6022 (N_6022,N_5981,N_5761);
nor U6023 (N_6023,N_5757,N_5512);
or U6024 (N_6024,N_5893,N_5842);
nor U6025 (N_6025,N_5745,N_5776);
nor U6026 (N_6026,N_5978,N_5667);
nor U6027 (N_6027,N_5950,N_5582);
nand U6028 (N_6028,N_5848,N_5875);
nor U6029 (N_6029,N_5737,N_5729);
nand U6030 (N_6030,N_5971,N_5937);
and U6031 (N_6031,N_5953,N_5760);
or U6032 (N_6032,N_5513,N_5672);
or U6033 (N_6033,N_5540,N_5652);
nand U6034 (N_6034,N_5784,N_5750);
nand U6035 (N_6035,N_5863,N_5986);
or U6036 (N_6036,N_5722,N_5574);
nand U6037 (N_6037,N_5558,N_5769);
or U6038 (N_6038,N_5532,N_5708);
nor U6039 (N_6039,N_5754,N_5653);
nor U6040 (N_6040,N_5980,N_5735);
or U6041 (N_6041,N_5728,N_5840);
nand U6042 (N_6042,N_5808,N_5676);
nor U6043 (N_6043,N_5796,N_5697);
nand U6044 (N_6044,N_5633,N_5523);
or U6045 (N_6045,N_5962,N_5689);
and U6046 (N_6046,N_5823,N_5560);
nor U6047 (N_6047,N_5668,N_5682);
and U6048 (N_6048,N_5510,N_5675);
xnor U6049 (N_6049,N_5688,N_5749);
nand U6050 (N_6050,N_5855,N_5989);
nand U6051 (N_6051,N_5519,N_5629);
xor U6052 (N_6052,N_5931,N_5886);
nor U6053 (N_6053,N_5988,N_5764);
nor U6054 (N_6054,N_5501,N_5854);
and U6055 (N_6055,N_5910,N_5927);
xnor U6056 (N_6056,N_5883,N_5954);
xor U6057 (N_6057,N_5834,N_5841);
nand U6058 (N_6058,N_5712,N_5811);
nor U6059 (N_6059,N_5544,N_5755);
or U6060 (N_6060,N_5715,N_5511);
or U6061 (N_6061,N_5999,N_5552);
xor U6062 (N_6062,N_5763,N_5723);
or U6063 (N_6063,N_5659,N_5586);
or U6064 (N_6064,N_5790,N_5565);
and U6065 (N_6065,N_5778,N_5583);
or U6066 (N_6066,N_5982,N_5710);
or U6067 (N_6067,N_5610,N_5615);
or U6068 (N_6068,N_5970,N_5899);
nor U6069 (N_6069,N_5976,N_5955);
xnor U6070 (N_6070,N_5827,N_5740);
and U6071 (N_6071,N_5767,N_5656);
xnor U6072 (N_6072,N_5619,N_5521);
nand U6073 (N_6073,N_5613,N_5838);
nor U6074 (N_6074,N_5742,N_5877);
or U6075 (N_6075,N_5520,N_5914);
or U6076 (N_6076,N_5733,N_5546);
and U6077 (N_6077,N_5900,N_5975);
xnor U6078 (N_6078,N_5527,N_5731);
or U6079 (N_6079,N_5518,N_5683);
xor U6080 (N_6080,N_5911,N_5632);
xnor U6081 (N_6081,N_5807,N_5938);
nor U6082 (N_6082,N_5669,N_5525);
nor U6083 (N_6083,N_5624,N_5584);
nor U6084 (N_6084,N_5866,N_5695);
xor U6085 (N_6085,N_5921,N_5942);
and U6086 (N_6086,N_5535,N_5932);
nand U6087 (N_6087,N_5903,N_5941);
and U6088 (N_6088,N_5744,N_5800);
or U6089 (N_6089,N_5892,N_5782);
nor U6090 (N_6090,N_5826,N_5531);
or U6091 (N_6091,N_5766,N_5538);
xnor U6092 (N_6092,N_5515,N_5861);
nor U6093 (N_6093,N_5878,N_5617);
nand U6094 (N_6094,N_5551,N_5704);
nand U6095 (N_6095,N_5578,N_5743);
nor U6096 (N_6096,N_5905,N_5758);
xnor U6097 (N_6097,N_5654,N_5549);
nand U6098 (N_6098,N_5801,N_5602);
and U6099 (N_6099,N_5880,N_5563);
nand U6100 (N_6100,N_5943,N_5849);
nor U6101 (N_6101,N_5741,N_5588);
nand U6102 (N_6102,N_5966,N_5636);
or U6103 (N_6103,N_5592,N_5865);
xnor U6104 (N_6104,N_5612,N_5607);
and U6105 (N_6105,N_5868,N_5634);
xnor U6106 (N_6106,N_5631,N_5939);
nand U6107 (N_6107,N_5662,N_5997);
nand U6108 (N_6108,N_5664,N_5788);
xnor U6109 (N_6109,N_5920,N_5884);
nor U6110 (N_6110,N_5770,N_5803);
nor U6111 (N_6111,N_5548,N_5876);
nand U6112 (N_6112,N_5922,N_5725);
or U6113 (N_6113,N_5746,N_5820);
and U6114 (N_6114,N_5916,N_5888);
nor U6115 (N_6115,N_5555,N_5590);
nand U6116 (N_6116,N_5844,N_5651);
nor U6117 (N_6117,N_5577,N_5979);
nor U6118 (N_6118,N_5638,N_5974);
nor U6119 (N_6119,N_5951,N_5564);
nand U6120 (N_6120,N_5618,N_5783);
or U6121 (N_6121,N_5542,N_5566);
xnor U6122 (N_6122,N_5500,N_5625);
nand U6123 (N_6123,N_5573,N_5589);
nor U6124 (N_6124,N_5568,N_5570);
nand U6125 (N_6125,N_5736,N_5707);
nand U6126 (N_6126,N_5983,N_5541);
and U6127 (N_6127,N_5909,N_5926);
and U6128 (N_6128,N_5965,N_5593);
nor U6129 (N_6129,N_5830,N_5889);
nand U6130 (N_6130,N_5524,N_5835);
and U6131 (N_6131,N_5747,N_5896);
or U6132 (N_6132,N_5773,N_5732);
nand U6133 (N_6133,N_5814,N_5973);
and U6134 (N_6134,N_5604,N_5522);
nor U6135 (N_6135,N_5639,N_5684);
or U6136 (N_6136,N_5930,N_5821);
nand U6137 (N_6137,N_5692,N_5819);
nand U6138 (N_6138,N_5804,N_5640);
nand U6139 (N_6139,N_5996,N_5813);
or U6140 (N_6140,N_5843,N_5856);
or U6141 (N_6141,N_5598,N_5575);
and U6142 (N_6142,N_5958,N_5809);
and U6143 (N_6143,N_5714,N_5822);
nand U6144 (N_6144,N_5724,N_5759);
nand U6145 (N_6145,N_5526,N_5690);
and U6146 (N_6146,N_5536,N_5648);
xnor U6147 (N_6147,N_5562,N_5882);
xnor U6148 (N_6148,N_5727,N_5857);
nor U6149 (N_6149,N_5952,N_5687);
nor U6150 (N_6150,N_5706,N_5816);
nor U6151 (N_6151,N_5508,N_5793);
or U6152 (N_6152,N_5553,N_5908);
nor U6153 (N_6153,N_5812,N_5533);
or U6154 (N_6154,N_5680,N_5585);
nor U6155 (N_6155,N_5571,N_5719);
xor U6156 (N_6156,N_5663,N_5798);
and U6157 (N_6157,N_5545,N_5795);
xnor U6158 (N_6158,N_5956,N_5913);
nor U6159 (N_6159,N_5806,N_5605);
and U6160 (N_6160,N_5928,N_5963);
xor U6161 (N_6161,N_5556,N_5968);
nand U6162 (N_6162,N_5991,N_5890);
and U6163 (N_6163,N_5959,N_5529);
nor U6164 (N_6164,N_5658,N_5751);
nand U6165 (N_6165,N_5785,N_5677);
and U6166 (N_6166,N_5509,N_5912);
nand U6167 (N_6167,N_5904,N_5693);
and U6168 (N_6168,N_5600,N_5972);
nor U6169 (N_6169,N_5753,N_5915);
nor U6170 (N_6170,N_5699,N_5833);
nor U6171 (N_6171,N_5873,N_5623);
xnor U6172 (N_6172,N_5872,N_5994);
or U6173 (N_6173,N_5992,N_5995);
nand U6174 (N_6174,N_5815,N_5595);
and U6175 (N_6175,N_5702,N_5924);
nor U6176 (N_6176,N_5635,N_5557);
nand U6177 (N_6177,N_5628,N_5777);
nor U6178 (N_6178,N_5637,N_5596);
nor U6179 (N_6179,N_5630,N_5505);
and U6180 (N_6180,N_5858,N_5794);
and U6181 (N_6181,N_5603,N_5679);
and U6182 (N_6182,N_5839,N_5894);
and U6183 (N_6183,N_5661,N_5528);
nand U6184 (N_6184,N_5622,N_5620);
or U6185 (N_6185,N_5944,N_5832);
and U6186 (N_6186,N_5587,N_5871);
xnor U6187 (N_6187,N_5898,N_5897);
and U6188 (N_6188,N_5933,N_5597);
and U6189 (N_6189,N_5534,N_5993);
and U6190 (N_6190,N_5846,N_5670);
and U6191 (N_6191,N_5734,N_5650);
xnor U6192 (N_6192,N_5961,N_5626);
nor U6193 (N_6193,N_5649,N_5967);
and U6194 (N_6194,N_5681,N_5859);
and U6195 (N_6195,N_5616,N_5694);
nor U6196 (N_6196,N_5591,N_5647);
or U6197 (N_6197,N_5837,N_5779);
nand U6198 (N_6198,N_5709,N_5579);
nand U6199 (N_6199,N_5907,N_5957);
nor U6200 (N_6200,N_5543,N_5701);
and U6201 (N_6201,N_5506,N_5642);
or U6202 (N_6202,N_5720,N_5799);
and U6203 (N_6203,N_5781,N_5810);
or U6204 (N_6204,N_5787,N_5655);
or U6205 (N_6205,N_5739,N_5686);
or U6206 (N_6206,N_5831,N_5947);
nand U6207 (N_6207,N_5660,N_5940);
nand U6208 (N_6208,N_5887,N_5581);
and U6209 (N_6209,N_5818,N_5987);
nand U6210 (N_6210,N_5852,N_5762);
nand U6211 (N_6211,N_5964,N_5901);
nor U6212 (N_6212,N_5845,N_5713);
nand U6213 (N_6213,N_5621,N_5514);
nand U6214 (N_6214,N_5752,N_5666);
and U6215 (N_6215,N_5530,N_5774);
nor U6216 (N_6216,N_5644,N_5895);
or U6217 (N_6217,N_5985,N_5730);
xor U6218 (N_6218,N_5862,N_5547);
nand U6219 (N_6219,N_5646,N_5853);
nand U6220 (N_6220,N_5925,N_5923);
nand U6221 (N_6221,N_5738,N_5703);
and U6222 (N_6222,N_5867,N_5797);
xor U6223 (N_6223,N_5572,N_5554);
nand U6224 (N_6224,N_5580,N_5516);
nor U6225 (N_6225,N_5691,N_5869);
nor U6226 (N_6226,N_5864,N_5906);
nor U6227 (N_6227,N_5969,N_5627);
and U6228 (N_6228,N_5885,N_5559);
xor U6229 (N_6229,N_5537,N_5919);
nor U6230 (N_6230,N_5802,N_5775);
and U6231 (N_6231,N_5698,N_5641);
or U6232 (N_6232,N_5998,N_5860);
xnor U6233 (N_6233,N_5792,N_5945);
nand U6234 (N_6234,N_5657,N_5817);
nand U6235 (N_6235,N_5870,N_5902);
or U6236 (N_6236,N_5949,N_5696);
and U6237 (N_6237,N_5503,N_5685);
nor U6238 (N_6238,N_5609,N_5874);
or U6239 (N_6239,N_5502,N_5671);
nor U6240 (N_6240,N_5678,N_5836);
or U6241 (N_6241,N_5771,N_5705);
and U6242 (N_6242,N_5850,N_5504);
nand U6243 (N_6243,N_5824,N_5780);
nand U6244 (N_6244,N_5716,N_5791);
or U6245 (N_6245,N_5934,N_5917);
nor U6246 (N_6246,N_5550,N_5601);
or U6247 (N_6247,N_5561,N_5946);
nor U6248 (N_6248,N_5805,N_5935);
xor U6249 (N_6249,N_5614,N_5948);
nand U6250 (N_6250,N_5511,N_5631);
nand U6251 (N_6251,N_5944,N_5516);
and U6252 (N_6252,N_5558,N_5990);
or U6253 (N_6253,N_5669,N_5999);
or U6254 (N_6254,N_5861,N_5987);
nand U6255 (N_6255,N_5668,N_5600);
or U6256 (N_6256,N_5572,N_5932);
or U6257 (N_6257,N_5967,N_5746);
nor U6258 (N_6258,N_5899,N_5664);
xor U6259 (N_6259,N_5762,N_5701);
nor U6260 (N_6260,N_5592,N_5789);
and U6261 (N_6261,N_5930,N_5854);
xor U6262 (N_6262,N_5724,N_5746);
nand U6263 (N_6263,N_5929,N_5547);
and U6264 (N_6264,N_5784,N_5975);
nand U6265 (N_6265,N_5988,N_5628);
and U6266 (N_6266,N_5690,N_5929);
nor U6267 (N_6267,N_5750,N_5827);
and U6268 (N_6268,N_5627,N_5889);
nand U6269 (N_6269,N_5608,N_5991);
nor U6270 (N_6270,N_5701,N_5615);
nand U6271 (N_6271,N_5542,N_5713);
and U6272 (N_6272,N_5510,N_5645);
and U6273 (N_6273,N_5659,N_5927);
nor U6274 (N_6274,N_5553,N_5769);
nor U6275 (N_6275,N_5848,N_5720);
nand U6276 (N_6276,N_5987,N_5775);
nor U6277 (N_6277,N_5700,N_5927);
and U6278 (N_6278,N_5677,N_5635);
and U6279 (N_6279,N_5838,N_5820);
nor U6280 (N_6280,N_5552,N_5706);
and U6281 (N_6281,N_5915,N_5822);
xor U6282 (N_6282,N_5858,N_5893);
nand U6283 (N_6283,N_5696,N_5579);
or U6284 (N_6284,N_5840,N_5749);
nand U6285 (N_6285,N_5701,N_5717);
and U6286 (N_6286,N_5743,N_5952);
and U6287 (N_6287,N_5625,N_5628);
and U6288 (N_6288,N_5891,N_5992);
nand U6289 (N_6289,N_5603,N_5811);
and U6290 (N_6290,N_5552,N_5584);
nor U6291 (N_6291,N_5572,N_5965);
nand U6292 (N_6292,N_5847,N_5552);
nor U6293 (N_6293,N_5834,N_5867);
nor U6294 (N_6294,N_5726,N_5751);
xor U6295 (N_6295,N_5588,N_5844);
nor U6296 (N_6296,N_5580,N_5537);
and U6297 (N_6297,N_5544,N_5973);
and U6298 (N_6298,N_5929,N_5664);
or U6299 (N_6299,N_5545,N_5909);
or U6300 (N_6300,N_5933,N_5801);
nor U6301 (N_6301,N_5562,N_5958);
nand U6302 (N_6302,N_5793,N_5656);
or U6303 (N_6303,N_5588,N_5698);
or U6304 (N_6304,N_5812,N_5953);
or U6305 (N_6305,N_5547,N_5682);
and U6306 (N_6306,N_5885,N_5562);
nor U6307 (N_6307,N_5681,N_5629);
nor U6308 (N_6308,N_5694,N_5737);
xnor U6309 (N_6309,N_5580,N_5796);
nor U6310 (N_6310,N_5638,N_5663);
or U6311 (N_6311,N_5858,N_5822);
nand U6312 (N_6312,N_5793,N_5569);
and U6313 (N_6313,N_5852,N_5747);
nand U6314 (N_6314,N_5920,N_5927);
nor U6315 (N_6315,N_5991,N_5788);
or U6316 (N_6316,N_5768,N_5744);
or U6317 (N_6317,N_5517,N_5944);
xnor U6318 (N_6318,N_5654,N_5913);
nor U6319 (N_6319,N_5570,N_5519);
nor U6320 (N_6320,N_5922,N_5987);
and U6321 (N_6321,N_5531,N_5996);
or U6322 (N_6322,N_5826,N_5541);
and U6323 (N_6323,N_5794,N_5811);
and U6324 (N_6324,N_5616,N_5925);
nand U6325 (N_6325,N_5554,N_5725);
nor U6326 (N_6326,N_5700,N_5514);
nand U6327 (N_6327,N_5843,N_5948);
nand U6328 (N_6328,N_5737,N_5749);
nand U6329 (N_6329,N_5687,N_5944);
nand U6330 (N_6330,N_5710,N_5721);
xnor U6331 (N_6331,N_5900,N_5669);
nand U6332 (N_6332,N_5531,N_5716);
nand U6333 (N_6333,N_5990,N_5760);
nor U6334 (N_6334,N_5771,N_5821);
and U6335 (N_6335,N_5746,N_5946);
nand U6336 (N_6336,N_5934,N_5751);
and U6337 (N_6337,N_5707,N_5926);
nor U6338 (N_6338,N_5732,N_5915);
nor U6339 (N_6339,N_5628,N_5524);
nor U6340 (N_6340,N_5626,N_5537);
or U6341 (N_6341,N_5760,N_5729);
nand U6342 (N_6342,N_5746,N_5881);
or U6343 (N_6343,N_5877,N_5564);
and U6344 (N_6344,N_5599,N_5744);
nor U6345 (N_6345,N_5896,N_5846);
and U6346 (N_6346,N_5993,N_5585);
or U6347 (N_6347,N_5554,N_5882);
or U6348 (N_6348,N_5679,N_5665);
and U6349 (N_6349,N_5810,N_5584);
and U6350 (N_6350,N_5704,N_5547);
nand U6351 (N_6351,N_5707,N_5647);
nor U6352 (N_6352,N_5702,N_5639);
nor U6353 (N_6353,N_5859,N_5529);
and U6354 (N_6354,N_5839,N_5717);
xor U6355 (N_6355,N_5865,N_5966);
and U6356 (N_6356,N_5820,N_5853);
nand U6357 (N_6357,N_5549,N_5777);
xor U6358 (N_6358,N_5789,N_5969);
and U6359 (N_6359,N_5750,N_5848);
and U6360 (N_6360,N_5780,N_5639);
nand U6361 (N_6361,N_5886,N_5520);
nand U6362 (N_6362,N_5832,N_5713);
and U6363 (N_6363,N_5555,N_5876);
nand U6364 (N_6364,N_5797,N_5511);
nor U6365 (N_6365,N_5805,N_5672);
and U6366 (N_6366,N_5850,N_5907);
nor U6367 (N_6367,N_5811,N_5943);
or U6368 (N_6368,N_5778,N_5980);
nand U6369 (N_6369,N_5891,N_5788);
nand U6370 (N_6370,N_5834,N_5733);
xor U6371 (N_6371,N_5772,N_5504);
xnor U6372 (N_6372,N_5966,N_5985);
nand U6373 (N_6373,N_5773,N_5849);
nand U6374 (N_6374,N_5854,N_5944);
nand U6375 (N_6375,N_5550,N_5589);
nor U6376 (N_6376,N_5727,N_5516);
and U6377 (N_6377,N_5520,N_5824);
or U6378 (N_6378,N_5798,N_5550);
and U6379 (N_6379,N_5686,N_5531);
and U6380 (N_6380,N_5735,N_5885);
and U6381 (N_6381,N_5929,N_5610);
nor U6382 (N_6382,N_5963,N_5723);
or U6383 (N_6383,N_5649,N_5979);
nand U6384 (N_6384,N_5721,N_5764);
nand U6385 (N_6385,N_5666,N_5877);
nor U6386 (N_6386,N_5575,N_5622);
and U6387 (N_6387,N_5573,N_5610);
or U6388 (N_6388,N_5964,N_5987);
xor U6389 (N_6389,N_5831,N_5696);
nand U6390 (N_6390,N_5848,N_5515);
xor U6391 (N_6391,N_5897,N_5610);
nand U6392 (N_6392,N_5709,N_5560);
and U6393 (N_6393,N_5940,N_5897);
nor U6394 (N_6394,N_5928,N_5508);
or U6395 (N_6395,N_5976,N_5756);
xnor U6396 (N_6396,N_5546,N_5633);
nand U6397 (N_6397,N_5787,N_5657);
or U6398 (N_6398,N_5838,N_5739);
nand U6399 (N_6399,N_5861,N_5684);
xor U6400 (N_6400,N_5552,N_5663);
or U6401 (N_6401,N_5816,N_5687);
and U6402 (N_6402,N_5849,N_5730);
and U6403 (N_6403,N_5834,N_5517);
and U6404 (N_6404,N_5652,N_5719);
nor U6405 (N_6405,N_5587,N_5613);
or U6406 (N_6406,N_5631,N_5557);
and U6407 (N_6407,N_5656,N_5899);
nand U6408 (N_6408,N_5919,N_5640);
nand U6409 (N_6409,N_5946,N_5596);
nand U6410 (N_6410,N_5933,N_5836);
nor U6411 (N_6411,N_5531,N_5869);
nand U6412 (N_6412,N_5621,N_5897);
nand U6413 (N_6413,N_5686,N_5599);
nor U6414 (N_6414,N_5544,N_5700);
nor U6415 (N_6415,N_5598,N_5908);
or U6416 (N_6416,N_5822,N_5849);
or U6417 (N_6417,N_5598,N_5527);
xnor U6418 (N_6418,N_5589,N_5872);
xor U6419 (N_6419,N_5535,N_5846);
nor U6420 (N_6420,N_5552,N_5760);
nand U6421 (N_6421,N_5679,N_5567);
nand U6422 (N_6422,N_5684,N_5842);
nand U6423 (N_6423,N_5813,N_5880);
nor U6424 (N_6424,N_5932,N_5993);
and U6425 (N_6425,N_5965,N_5643);
xnor U6426 (N_6426,N_5626,N_5804);
nor U6427 (N_6427,N_5729,N_5694);
nand U6428 (N_6428,N_5807,N_5848);
nand U6429 (N_6429,N_5967,N_5605);
and U6430 (N_6430,N_5544,N_5826);
nand U6431 (N_6431,N_5765,N_5881);
xor U6432 (N_6432,N_5710,N_5560);
or U6433 (N_6433,N_5959,N_5844);
or U6434 (N_6434,N_5652,N_5699);
or U6435 (N_6435,N_5690,N_5702);
nand U6436 (N_6436,N_5966,N_5835);
or U6437 (N_6437,N_5785,N_5671);
nor U6438 (N_6438,N_5540,N_5891);
nor U6439 (N_6439,N_5681,N_5796);
nand U6440 (N_6440,N_5501,N_5537);
nand U6441 (N_6441,N_5915,N_5584);
nor U6442 (N_6442,N_5705,N_5653);
or U6443 (N_6443,N_5551,N_5946);
nand U6444 (N_6444,N_5630,N_5523);
and U6445 (N_6445,N_5971,N_5801);
nor U6446 (N_6446,N_5783,N_5666);
and U6447 (N_6447,N_5534,N_5545);
nor U6448 (N_6448,N_5740,N_5659);
or U6449 (N_6449,N_5567,N_5654);
nand U6450 (N_6450,N_5533,N_5859);
nand U6451 (N_6451,N_5963,N_5833);
xor U6452 (N_6452,N_5550,N_5713);
nand U6453 (N_6453,N_5842,N_5620);
nor U6454 (N_6454,N_5666,N_5818);
nor U6455 (N_6455,N_5679,N_5838);
nand U6456 (N_6456,N_5612,N_5911);
or U6457 (N_6457,N_5962,N_5838);
nand U6458 (N_6458,N_5626,N_5943);
and U6459 (N_6459,N_5619,N_5840);
and U6460 (N_6460,N_5534,N_5666);
and U6461 (N_6461,N_5824,N_5790);
nand U6462 (N_6462,N_5778,N_5997);
xnor U6463 (N_6463,N_5562,N_5544);
xnor U6464 (N_6464,N_5955,N_5635);
and U6465 (N_6465,N_5548,N_5868);
nor U6466 (N_6466,N_5678,N_5698);
xnor U6467 (N_6467,N_5867,N_5774);
xnor U6468 (N_6468,N_5775,N_5743);
or U6469 (N_6469,N_5543,N_5649);
nor U6470 (N_6470,N_5740,N_5558);
or U6471 (N_6471,N_5577,N_5798);
and U6472 (N_6472,N_5574,N_5793);
xnor U6473 (N_6473,N_5890,N_5908);
nand U6474 (N_6474,N_5536,N_5832);
and U6475 (N_6475,N_5705,N_5694);
nand U6476 (N_6476,N_5543,N_5929);
nor U6477 (N_6477,N_5554,N_5883);
and U6478 (N_6478,N_5663,N_5762);
nor U6479 (N_6479,N_5670,N_5572);
nor U6480 (N_6480,N_5882,N_5741);
or U6481 (N_6481,N_5896,N_5841);
nand U6482 (N_6482,N_5621,N_5654);
or U6483 (N_6483,N_5783,N_5822);
and U6484 (N_6484,N_5502,N_5526);
or U6485 (N_6485,N_5908,N_5909);
or U6486 (N_6486,N_5796,N_5816);
and U6487 (N_6487,N_5562,N_5771);
or U6488 (N_6488,N_5603,N_5786);
xnor U6489 (N_6489,N_5789,N_5716);
nor U6490 (N_6490,N_5838,N_5772);
nand U6491 (N_6491,N_5525,N_5944);
nor U6492 (N_6492,N_5921,N_5598);
nand U6493 (N_6493,N_5647,N_5661);
or U6494 (N_6494,N_5583,N_5906);
nand U6495 (N_6495,N_5668,N_5921);
and U6496 (N_6496,N_5640,N_5699);
and U6497 (N_6497,N_5667,N_5787);
nor U6498 (N_6498,N_5534,N_5575);
nand U6499 (N_6499,N_5988,N_5658);
or U6500 (N_6500,N_6234,N_6088);
or U6501 (N_6501,N_6253,N_6276);
and U6502 (N_6502,N_6254,N_6441);
nand U6503 (N_6503,N_6408,N_6446);
and U6504 (N_6504,N_6235,N_6494);
nor U6505 (N_6505,N_6431,N_6221);
nand U6506 (N_6506,N_6171,N_6230);
or U6507 (N_6507,N_6433,N_6351);
nand U6508 (N_6508,N_6135,N_6275);
and U6509 (N_6509,N_6289,N_6498);
nand U6510 (N_6510,N_6092,N_6291);
or U6511 (N_6511,N_6488,N_6232);
and U6512 (N_6512,N_6024,N_6039);
xnor U6513 (N_6513,N_6250,N_6423);
nor U6514 (N_6514,N_6086,N_6213);
nand U6515 (N_6515,N_6200,N_6357);
nor U6516 (N_6516,N_6393,N_6339);
and U6517 (N_6517,N_6182,N_6363);
nor U6518 (N_6518,N_6105,N_6004);
xnor U6519 (N_6519,N_6085,N_6388);
nand U6520 (N_6520,N_6141,N_6185);
nand U6521 (N_6521,N_6391,N_6394);
nor U6522 (N_6522,N_6473,N_6266);
nor U6523 (N_6523,N_6063,N_6440);
and U6524 (N_6524,N_6176,N_6144);
nand U6525 (N_6525,N_6160,N_6152);
nor U6526 (N_6526,N_6075,N_6199);
nand U6527 (N_6527,N_6369,N_6427);
nor U6528 (N_6528,N_6143,N_6018);
or U6529 (N_6529,N_6158,N_6166);
or U6530 (N_6530,N_6150,N_6387);
or U6531 (N_6531,N_6027,N_6132);
or U6532 (N_6532,N_6013,N_6284);
xor U6533 (N_6533,N_6084,N_6303);
xnor U6534 (N_6534,N_6416,N_6207);
and U6535 (N_6535,N_6308,N_6381);
and U6536 (N_6536,N_6231,N_6424);
nand U6537 (N_6537,N_6469,N_6272);
or U6538 (N_6538,N_6102,N_6313);
nor U6539 (N_6539,N_6344,N_6282);
nand U6540 (N_6540,N_6035,N_6153);
nor U6541 (N_6541,N_6455,N_6029);
and U6542 (N_6542,N_6352,N_6002);
xor U6543 (N_6543,N_6019,N_6205);
or U6544 (N_6544,N_6123,N_6090);
and U6545 (N_6545,N_6025,N_6097);
nand U6546 (N_6546,N_6046,N_6398);
and U6547 (N_6547,N_6076,N_6038);
xnor U6548 (N_6548,N_6259,N_6318);
and U6549 (N_6549,N_6120,N_6444);
or U6550 (N_6550,N_6331,N_6103);
xnor U6551 (N_6551,N_6425,N_6479);
and U6552 (N_6552,N_6336,N_6358);
nor U6553 (N_6553,N_6297,N_6225);
nand U6554 (N_6554,N_6093,N_6484);
or U6555 (N_6555,N_6030,N_6380);
nor U6556 (N_6556,N_6285,N_6294);
or U6557 (N_6557,N_6167,N_6386);
nand U6558 (N_6558,N_6443,N_6136);
nand U6559 (N_6559,N_6061,N_6251);
and U6560 (N_6560,N_6055,N_6007);
and U6561 (N_6561,N_6260,N_6212);
nor U6562 (N_6562,N_6091,N_6470);
and U6563 (N_6563,N_6257,N_6390);
nor U6564 (N_6564,N_6264,N_6245);
or U6565 (N_6565,N_6252,N_6345);
and U6566 (N_6566,N_6137,N_6162);
nor U6567 (N_6567,N_6227,N_6379);
xor U6568 (N_6568,N_6215,N_6073);
and U6569 (N_6569,N_6377,N_6273);
nand U6570 (N_6570,N_6319,N_6114);
nand U6571 (N_6571,N_6417,N_6110);
and U6572 (N_6572,N_6006,N_6140);
or U6573 (N_6573,N_6483,N_6321);
nor U6574 (N_6574,N_6109,N_6005);
and U6575 (N_6575,N_6054,N_6128);
and U6576 (N_6576,N_6396,N_6464);
nor U6577 (N_6577,N_6341,N_6405);
xor U6578 (N_6578,N_6311,N_6069);
nand U6579 (N_6579,N_6001,N_6042);
and U6580 (N_6580,N_6392,N_6323);
and U6581 (N_6581,N_6402,N_6228);
nor U6582 (N_6582,N_6467,N_6413);
or U6583 (N_6583,N_6126,N_6249);
and U6584 (N_6584,N_6220,N_6330);
and U6585 (N_6585,N_6170,N_6466);
and U6586 (N_6586,N_6190,N_6178);
nor U6587 (N_6587,N_6223,N_6201);
nand U6588 (N_6588,N_6293,N_6490);
nor U6589 (N_6589,N_6026,N_6139);
and U6590 (N_6590,N_6281,N_6059);
xor U6591 (N_6591,N_6146,N_6365);
and U6592 (N_6592,N_6429,N_6359);
nand U6593 (N_6593,N_6057,N_6422);
nor U6594 (N_6594,N_6395,N_6406);
nor U6595 (N_6595,N_6183,N_6437);
and U6596 (N_6596,N_6499,N_6078);
nor U6597 (N_6597,N_6442,N_6347);
xor U6598 (N_6598,N_6175,N_6439);
nor U6599 (N_6599,N_6216,N_6434);
or U6600 (N_6600,N_6083,N_6372);
or U6601 (N_6601,N_6181,N_6485);
xnor U6602 (N_6602,N_6172,N_6186);
and U6603 (N_6603,N_6236,N_6465);
and U6604 (N_6604,N_6112,N_6173);
and U6605 (N_6605,N_6169,N_6288);
xnor U6606 (N_6606,N_6108,N_6101);
and U6607 (N_6607,N_6348,N_6191);
nor U6608 (N_6608,N_6492,N_6415);
and U6609 (N_6609,N_6229,N_6364);
and U6610 (N_6610,N_6195,N_6463);
nand U6611 (N_6611,N_6335,N_6304);
nor U6612 (N_6612,N_6401,N_6329);
nor U6613 (N_6613,N_6217,N_6487);
nand U6614 (N_6614,N_6326,N_6119);
or U6615 (N_6615,N_6050,N_6298);
or U6616 (N_6616,N_6138,N_6189);
or U6617 (N_6617,N_6246,N_6338);
nand U6618 (N_6618,N_6486,N_6481);
or U6619 (N_6619,N_6077,N_6067);
and U6620 (N_6620,N_6022,N_6051);
and U6621 (N_6621,N_6070,N_6295);
or U6622 (N_6622,N_6023,N_6286);
nand U6623 (N_6623,N_6262,N_6450);
nand U6624 (N_6624,N_6474,N_6130);
and U6625 (N_6625,N_6305,N_6451);
nand U6626 (N_6626,N_6041,N_6476);
and U6627 (N_6627,N_6468,N_6210);
or U6628 (N_6628,N_6320,N_6017);
nor U6629 (N_6629,N_6163,N_6399);
xor U6630 (N_6630,N_6382,N_6371);
nor U6631 (N_6631,N_6087,N_6309);
nor U6632 (N_6632,N_6037,N_6133);
or U6633 (N_6633,N_6362,N_6204);
nor U6634 (N_6634,N_6458,N_6478);
xor U6635 (N_6635,N_6242,N_6271);
and U6636 (N_6636,N_6459,N_6471);
and U6637 (N_6637,N_6021,N_6420);
nand U6638 (N_6638,N_6340,N_6480);
nand U6639 (N_6639,N_6475,N_6403);
xnor U6640 (N_6640,N_6373,N_6278);
or U6641 (N_6641,N_6412,N_6496);
nand U6642 (N_6642,N_6202,N_6145);
and U6643 (N_6643,N_6040,N_6407);
and U6644 (N_6644,N_6003,N_6010);
or U6645 (N_6645,N_6274,N_6317);
or U6646 (N_6646,N_6012,N_6047);
and U6647 (N_6647,N_6325,N_6107);
xnor U6648 (N_6648,N_6461,N_6094);
nor U6649 (N_6649,N_6062,N_6306);
or U6650 (N_6650,N_6244,N_6302);
or U6651 (N_6651,N_6174,N_6277);
or U6652 (N_6652,N_6314,N_6241);
or U6653 (N_6653,N_6065,N_6290);
or U6654 (N_6654,N_6219,N_6310);
nor U6655 (N_6655,N_6375,N_6008);
nor U6656 (N_6656,N_6356,N_6177);
and U6657 (N_6657,N_6360,N_6324);
nand U6658 (N_6658,N_6154,N_6301);
or U6659 (N_6659,N_6389,N_6081);
or U6660 (N_6660,N_6292,N_6280);
nand U6661 (N_6661,N_6203,N_6188);
and U6662 (N_6662,N_6445,N_6454);
and U6663 (N_6663,N_6134,N_6124);
nor U6664 (N_6664,N_6072,N_6238);
nand U6665 (N_6665,N_6196,N_6168);
or U6666 (N_6666,N_6131,N_6098);
nand U6667 (N_6667,N_6009,N_6179);
nand U6668 (N_6668,N_6355,N_6115);
nor U6669 (N_6669,N_6015,N_6247);
nand U6670 (N_6670,N_6327,N_6432);
nor U6671 (N_6671,N_6099,N_6438);
and U6672 (N_6672,N_6267,N_6155);
nor U6673 (N_6673,N_6161,N_6270);
nand U6674 (N_6674,N_6118,N_6095);
nand U6675 (N_6675,N_6187,N_6457);
or U6676 (N_6676,N_6028,N_6343);
or U6677 (N_6677,N_6034,N_6000);
nand U6678 (N_6678,N_6383,N_6261);
and U6679 (N_6679,N_6447,N_6493);
xnor U6680 (N_6680,N_6036,N_6071);
xor U6681 (N_6681,N_6489,N_6049);
or U6682 (N_6682,N_6052,N_6193);
and U6683 (N_6683,N_6453,N_6226);
or U6684 (N_6684,N_6410,N_6349);
or U6685 (N_6685,N_6409,N_6127);
or U6686 (N_6686,N_6222,N_6315);
or U6687 (N_6687,N_6113,N_6361);
or U6688 (N_6688,N_6350,N_6268);
nor U6689 (N_6689,N_6121,N_6332);
and U6690 (N_6690,N_6233,N_6157);
nand U6691 (N_6691,N_6328,N_6125);
nor U6692 (N_6692,N_6016,N_6426);
or U6693 (N_6693,N_6106,N_6370);
and U6694 (N_6694,N_6068,N_6214);
and U6695 (N_6695,N_6064,N_6421);
nor U6696 (N_6696,N_6209,N_6011);
and U6697 (N_6697,N_6248,N_6149);
nand U6698 (N_6698,N_6430,N_6316);
nand U6699 (N_6699,N_6079,N_6384);
and U6700 (N_6700,N_6452,N_6045);
nor U6701 (N_6701,N_6033,N_6449);
and U6702 (N_6702,N_6333,N_6096);
xor U6703 (N_6703,N_6269,N_6020);
nor U6704 (N_6704,N_6197,N_6198);
nand U6705 (N_6705,N_6256,N_6472);
or U6706 (N_6706,N_6299,N_6491);
nor U6707 (N_6707,N_6404,N_6074);
nor U6708 (N_6708,N_6385,N_6100);
nor U6709 (N_6709,N_6116,N_6482);
nand U6710 (N_6710,N_6428,N_6164);
or U6711 (N_6711,N_6296,N_6156);
and U6712 (N_6712,N_6218,N_6044);
and U6713 (N_6713,N_6346,N_6147);
and U6714 (N_6714,N_6436,N_6192);
and U6715 (N_6715,N_6032,N_6184);
nand U6716 (N_6716,N_6056,N_6411);
nand U6717 (N_6717,N_6435,N_6082);
nor U6718 (N_6718,N_6414,N_6374);
nor U6719 (N_6719,N_6368,N_6334);
nand U6720 (N_6720,N_6367,N_6477);
and U6721 (N_6721,N_6497,N_6165);
and U6722 (N_6722,N_6337,N_6448);
nand U6723 (N_6723,N_6208,N_6255);
or U6724 (N_6724,N_6224,N_6495);
or U6725 (N_6725,N_6142,N_6111);
nand U6726 (N_6726,N_6053,N_6400);
nor U6727 (N_6727,N_6151,N_6397);
or U6728 (N_6728,N_6378,N_6265);
xnor U6729 (N_6729,N_6283,N_6300);
xnor U6730 (N_6730,N_6060,N_6117);
nand U6731 (N_6731,N_6287,N_6066);
and U6732 (N_6732,N_6031,N_6243);
nand U6733 (N_6733,N_6419,N_6354);
or U6734 (N_6734,N_6129,N_6258);
and U6735 (N_6735,N_6080,N_6148);
and U6736 (N_6736,N_6376,N_6014);
xnor U6737 (N_6737,N_6342,N_6462);
or U6738 (N_6738,N_6058,N_6211);
xnor U6739 (N_6739,N_6312,N_6159);
and U6740 (N_6740,N_6322,N_6460);
and U6741 (N_6741,N_6366,N_6048);
xor U6742 (N_6742,N_6263,N_6194);
and U6743 (N_6743,N_6104,N_6279);
or U6744 (N_6744,N_6122,N_6240);
nand U6745 (N_6745,N_6206,N_6353);
xnor U6746 (N_6746,N_6307,N_6237);
or U6747 (N_6747,N_6239,N_6456);
and U6748 (N_6748,N_6418,N_6180);
and U6749 (N_6749,N_6043,N_6089);
or U6750 (N_6750,N_6198,N_6377);
and U6751 (N_6751,N_6058,N_6124);
nor U6752 (N_6752,N_6044,N_6144);
and U6753 (N_6753,N_6488,N_6401);
nand U6754 (N_6754,N_6423,N_6204);
and U6755 (N_6755,N_6388,N_6416);
nor U6756 (N_6756,N_6141,N_6393);
and U6757 (N_6757,N_6029,N_6186);
nor U6758 (N_6758,N_6081,N_6006);
and U6759 (N_6759,N_6387,N_6425);
nand U6760 (N_6760,N_6164,N_6041);
nor U6761 (N_6761,N_6318,N_6197);
xnor U6762 (N_6762,N_6377,N_6229);
nor U6763 (N_6763,N_6173,N_6124);
and U6764 (N_6764,N_6238,N_6191);
nor U6765 (N_6765,N_6199,N_6246);
nor U6766 (N_6766,N_6140,N_6227);
nor U6767 (N_6767,N_6205,N_6139);
and U6768 (N_6768,N_6270,N_6166);
nor U6769 (N_6769,N_6346,N_6291);
or U6770 (N_6770,N_6421,N_6066);
nand U6771 (N_6771,N_6333,N_6057);
nor U6772 (N_6772,N_6218,N_6018);
nand U6773 (N_6773,N_6095,N_6377);
xor U6774 (N_6774,N_6064,N_6219);
or U6775 (N_6775,N_6222,N_6272);
nor U6776 (N_6776,N_6249,N_6378);
or U6777 (N_6777,N_6497,N_6345);
nor U6778 (N_6778,N_6178,N_6413);
nand U6779 (N_6779,N_6486,N_6063);
nand U6780 (N_6780,N_6427,N_6118);
and U6781 (N_6781,N_6078,N_6426);
nand U6782 (N_6782,N_6036,N_6149);
nand U6783 (N_6783,N_6209,N_6043);
or U6784 (N_6784,N_6428,N_6372);
and U6785 (N_6785,N_6383,N_6175);
or U6786 (N_6786,N_6147,N_6379);
or U6787 (N_6787,N_6074,N_6236);
nor U6788 (N_6788,N_6167,N_6274);
nand U6789 (N_6789,N_6278,N_6395);
nor U6790 (N_6790,N_6438,N_6153);
xnor U6791 (N_6791,N_6447,N_6465);
nor U6792 (N_6792,N_6286,N_6328);
nand U6793 (N_6793,N_6162,N_6104);
and U6794 (N_6794,N_6374,N_6470);
or U6795 (N_6795,N_6321,N_6403);
nor U6796 (N_6796,N_6263,N_6317);
nand U6797 (N_6797,N_6399,N_6217);
nand U6798 (N_6798,N_6094,N_6057);
and U6799 (N_6799,N_6343,N_6078);
nor U6800 (N_6800,N_6052,N_6196);
and U6801 (N_6801,N_6447,N_6248);
and U6802 (N_6802,N_6346,N_6284);
xor U6803 (N_6803,N_6167,N_6202);
nor U6804 (N_6804,N_6407,N_6218);
or U6805 (N_6805,N_6307,N_6365);
nor U6806 (N_6806,N_6172,N_6111);
or U6807 (N_6807,N_6388,N_6173);
nor U6808 (N_6808,N_6401,N_6354);
nor U6809 (N_6809,N_6332,N_6202);
nand U6810 (N_6810,N_6356,N_6265);
and U6811 (N_6811,N_6189,N_6071);
or U6812 (N_6812,N_6239,N_6369);
or U6813 (N_6813,N_6102,N_6021);
nor U6814 (N_6814,N_6370,N_6364);
and U6815 (N_6815,N_6233,N_6221);
nor U6816 (N_6816,N_6141,N_6447);
and U6817 (N_6817,N_6053,N_6162);
nor U6818 (N_6818,N_6230,N_6040);
or U6819 (N_6819,N_6125,N_6049);
or U6820 (N_6820,N_6032,N_6361);
xnor U6821 (N_6821,N_6493,N_6179);
nor U6822 (N_6822,N_6333,N_6159);
nor U6823 (N_6823,N_6466,N_6235);
nor U6824 (N_6824,N_6193,N_6406);
and U6825 (N_6825,N_6308,N_6061);
or U6826 (N_6826,N_6418,N_6153);
xor U6827 (N_6827,N_6426,N_6222);
or U6828 (N_6828,N_6175,N_6116);
nor U6829 (N_6829,N_6432,N_6160);
or U6830 (N_6830,N_6376,N_6115);
nor U6831 (N_6831,N_6105,N_6119);
nor U6832 (N_6832,N_6174,N_6267);
nor U6833 (N_6833,N_6004,N_6211);
nand U6834 (N_6834,N_6094,N_6306);
and U6835 (N_6835,N_6264,N_6248);
nor U6836 (N_6836,N_6059,N_6326);
nor U6837 (N_6837,N_6328,N_6108);
or U6838 (N_6838,N_6248,N_6361);
nor U6839 (N_6839,N_6103,N_6002);
nand U6840 (N_6840,N_6149,N_6450);
or U6841 (N_6841,N_6384,N_6067);
nand U6842 (N_6842,N_6322,N_6009);
nor U6843 (N_6843,N_6134,N_6389);
and U6844 (N_6844,N_6368,N_6260);
nor U6845 (N_6845,N_6467,N_6376);
and U6846 (N_6846,N_6245,N_6050);
nand U6847 (N_6847,N_6469,N_6359);
nor U6848 (N_6848,N_6022,N_6357);
or U6849 (N_6849,N_6396,N_6460);
nor U6850 (N_6850,N_6437,N_6409);
nand U6851 (N_6851,N_6374,N_6348);
nor U6852 (N_6852,N_6058,N_6463);
nand U6853 (N_6853,N_6333,N_6081);
and U6854 (N_6854,N_6215,N_6273);
and U6855 (N_6855,N_6311,N_6272);
nor U6856 (N_6856,N_6241,N_6067);
or U6857 (N_6857,N_6386,N_6256);
nand U6858 (N_6858,N_6336,N_6302);
and U6859 (N_6859,N_6118,N_6469);
nand U6860 (N_6860,N_6410,N_6191);
or U6861 (N_6861,N_6066,N_6187);
xnor U6862 (N_6862,N_6088,N_6170);
nand U6863 (N_6863,N_6159,N_6292);
nor U6864 (N_6864,N_6001,N_6322);
nand U6865 (N_6865,N_6483,N_6292);
nor U6866 (N_6866,N_6309,N_6070);
nor U6867 (N_6867,N_6218,N_6461);
xor U6868 (N_6868,N_6015,N_6070);
or U6869 (N_6869,N_6496,N_6093);
nand U6870 (N_6870,N_6103,N_6215);
nor U6871 (N_6871,N_6143,N_6474);
or U6872 (N_6872,N_6251,N_6475);
nor U6873 (N_6873,N_6038,N_6315);
nand U6874 (N_6874,N_6092,N_6137);
and U6875 (N_6875,N_6246,N_6313);
nand U6876 (N_6876,N_6455,N_6418);
nand U6877 (N_6877,N_6012,N_6141);
nor U6878 (N_6878,N_6059,N_6198);
and U6879 (N_6879,N_6282,N_6386);
xor U6880 (N_6880,N_6499,N_6113);
xnor U6881 (N_6881,N_6201,N_6125);
nand U6882 (N_6882,N_6252,N_6227);
and U6883 (N_6883,N_6251,N_6115);
and U6884 (N_6884,N_6068,N_6031);
xor U6885 (N_6885,N_6245,N_6275);
or U6886 (N_6886,N_6252,N_6072);
nor U6887 (N_6887,N_6139,N_6213);
and U6888 (N_6888,N_6442,N_6387);
nand U6889 (N_6889,N_6115,N_6391);
nor U6890 (N_6890,N_6083,N_6251);
nand U6891 (N_6891,N_6377,N_6075);
or U6892 (N_6892,N_6406,N_6318);
or U6893 (N_6893,N_6068,N_6370);
nand U6894 (N_6894,N_6046,N_6080);
nor U6895 (N_6895,N_6033,N_6418);
nand U6896 (N_6896,N_6199,N_6340);
xnor U6897 (N_6897,N_6194,N_6407);
nand U6898 (N_6898,N_6395,N_6187);
nor U6899 (N_6899,N_6178,N_6092);
nor U6900 (N_6900,N_6185,N_6097);
nor U6901 (N_6901,N_6133,N_6245);
and U6902 (N_6902,N_6091,N_6019);
or U6903 (N_6903,N_6191,N_6387);
nand U6904 (N_6904,N_6432,N_6170);
xnor U6905 (N_6905,N_6370,N_6358);
xnor U6906 (N_6906,N_6267,N_6468);
and U6907 (N_6907,N_6412,N_6060);
nor U6908 (N_6908,N_6152,N_6027);
xor U6909 (N_6909,N_6482,N_6404);
or U6910 (N_6910,N_6447,N_6464);
or U6911 (N_6911,N_6252,N_6129);
and U6912 (N_6912,N_6018,N_6158);
nand U6913 (N_6913,N_6362,N_6044);
or U6914 (N_6914,N_6064,N_6432);
nand U6915 (N_6915,N_6085,N_6163);
or U6916 (N_6916,N_6198,N_6153);
and U6917 (N_6917,N_6286,N_6192);
or U6918 (N_6918,N_6499,N_6027);
nand U6919 (N_6919,N_6116,N_6311);
or U6920 (N_6920,N_6420,N_6304);
or U6921 (N_6921,N_6070,N_6357);
nor U6922 (N_6922,N_6344,N_6479);
nand U6923 (N_6923,N_6211,N_6427);
and U6924 (N_6924,N_6195,N_6224);
nor U6925 (N_6925,N_6214,N_6476);
nand U6926 (N_6926,N_6016,N_6270);
nand U6927 (N_6927,N_6295,N_6259);
nand U6928 (N_6928,N_6083,N_6467);
nand U6929 (N_6929,N_6478,N_6124);
or U6930 (N_6930,N_6317,N_6369);
xor U6931 (N_6931,N_6368,N_6396);
and U6932 (N_6932,N_6410,N_6202);
nor U6933 (N_6933,N_6025,N_6244);
nor U6934 (N_6934,N_6427,N_6421);
nor U6935 (N_6935,N_6366,N_6261);
nand U6936 (N_6936,N_6045,N_6284);
nand U6937 (N_6937,N_6352,N_6173);
xor U6938 (N_6938,N_6136,N_6472);
nor U6939 (N_6939,N_6403,N_6261);
nor U6940 (N_6940,N_6151,N_6416);
xnor U6941 (N_6941,N_6450,N_6464);
xnor U6942 (N_6942,N_6260,N_6129);
and U6943 (N_6943,N_6094,N_6213);
nand U6944 (N_6944,N_6150,N_6433);
nand U6945 (N_6945,N_6463,N_6305);
nand U6946 (N_6946,N_6389,N_6407);
nand U6947 (N_6947,N_6217,N_6230);
and U6948 (N_6948,N_6115,N_6005);
nand U6949 (N_6949,N_6139,N_6358);
nor U6950 (N_6950,N_6416,N_6136);
or U6951 (N_6951,N_6362,N_6075);
and U6952 (N_6952,N_6147,N_6488);
nand U6953 (N_6953,N_6226,N_6131);
or U6954 (N_6954,N_6079,N_6328);
nor U6955 (N_6955,N_6127,N_6486);
nand U6956 (N_6956,N_6305,N_6254);
or U6957 (N_6957,N_6216,N_6147);
or U6958 (N_6958,N_6261,N_6332);
xor U6959 (N_6959,N_6296,N_6049);
nor U6960 (N_6960,N_6181,N_6007);
xnor U6961 (N_6961,N_6101,N_6081);
nand U6962 (N_6962,N_6281,N_6062);
and U6963 (N_6963,N_6288,N_6447);
and U6964 (N_6964,N_6225,N_6281);
or U6965 (N_6965,N_6398,N_6009);
and U6966 (N_6966,N_6462,N_6497);
nor U6967 (N_6967,N_6433,N_6168);
nand U6968 (N_6968,N_6196,N_6107);
and U6969 (N_6969,N_6437,N_6251);
and U6970 (N_6970,N_6172,N_6364);
or U6971 (N_6971,N_6155,N_6083);
nor U6972 (N_6972,N_6331,N_6100);
nor U6973 (N_6973,N_6326,N_6251);
and U6974 (N_6974,N_6462,N_6193);
nor U6975 (N_6975,N_6292,N_6231);
and U6976 (N_6976,N_6113,N_6339);
and U6977 (N_6977,N_6333,N_6083);
and U6978 (N_6978,N_6089,N_6341);
nand U6979 (N_6979,N_6173,N_6082);
or U6980 (N_6980,N_6044,N_6327);
and U6981 (N_6981,N_6036,N_6073);
xor U6982 (N_6982,N_6494,N_6498);
and U6983 (N_6983,N_6116,N_6330);
nor U6984 (N_6984,N_6168,N_6293);
or U6985 (N_6985,N_6383,N_6130);
or U6986 (N_6986,N_6210,N_6483);
or U6987 (N_6987,N_6398,N_6363);
nor U6988 (N_6988,N_6211,N_6005);
nor U6989 (N_6989,N_6230,N_6423);
and U6990 (N_6990,N_6375,N_6127);
nand U6991 (N_6991,N_6215,N_6387);
nand U6992 (N_6992,N_6138,N_6031);
nand U6993 (N_6993,N_6398,N_6422);
nand U6994 (N_6994,N_6496,N_6017);
or U6995 (N_6995,N_6345,N_6034);
or U6996 (N_6996,N_6168,N_6067);
nand U6997 (N_6997,N_6413,N_6216);
and U6998 (N_6998,N_6401,N_6304);
or U6999 (N_6999,N_6038,N_6473);
and U7000 (N_7000,N_6539,N_6657);
nand U7001 (N_7001,N_6766,N_6541);
nand U7002 (N_7002,N_6614,N_6637);
nand U7003 (N_7003,N_6638,N_6596);
nand U7004 (N_7004,N_6672,N_6502);
and U7005 (N_7005,N_6667,N_6640);
nand U7006 (N_7006,N_6641,N_6671);
and U7007 (N_7007,N_6894,N_6778);
or U7008 (N_7008,N_6974,N_6941);
xor U7009 (N_7009,N_6628,N_6835);
or U7010 (N_7010,N_6837,N_6907);
and U7011 (N_7011,N_6903,N_6720);
nand U7012 (N_7012,N_6562,N_6542);
and U7013 (N_7013,N_6985,N_6955);
or U7014 (N_7014,N_6990,N_6506);
and U7015 (N_7015,N_6743,N_6515);
nor U7016 (N_7016,N_6939,N_6885);
or U7017 (N_7017,N_6962,N_6507);
or U7018 (N_7018,N_6887,N_6533);
xnor U7019 (N_7019,N_6675,N_6775);
or U7020 (N_7020,N_6928,N_6954);
nand U7021 (N_7021,N_6929,N_6861);
and U7022 (N_7022,N_6710,N_6920);
nor U7023 (N_7023,N_6817,N_6748);
and U7024 (N_7024,N_6519,N_6682);
nand U7025 (N_7025,N_6568,N_6664);
nor U7026 (N_7026,N_6845,N_6935);
and U7027 (N_7027,N_6595,N_6613);
nor U7028 (N_7028,N_6970,N_6732);
nand U7029 (N_7029,N_6945,N_6800);
or U7030 (N_7030,N_6727,N_6769);
xor U7031 (N_7031,N_6914,N_6582);
nor U7032 (N_7032,N_6537,N_6911);
and U7033 (N_7033,N_6683,N_6599);
or U7034 (N_7034,N_6785,N_6656);
and U7035 (N_7035,N_6839,N_6740);
or U7036 (N_7036,N_6846,N_6879);
xnor U7037 (N_7037,N_6663,N_6697);
nand U7038 (N_7038,N_6617,N_6632);
and U7039 (N_7039,N_6991,N_6953);
nor U7040 (N_7040,N_6677,N_6755);
or U7041 (N_7041,N_6504,N_6918);
nor U7042 (N_7042,N_6517,N_6650);
or U7043 (N_7043,N_6780,N_6959);
nand U7044 (N_7044,N_6813,N_6698);
nand U7045 (N_7045,N_6610,N_6925);
or U7046 (N_7046,N_6898,N_6500);
nand U7047 (N_7047,N_6699,N_6691);
nor U7048 (N_7048,N_6913,N_6761);
or U7049 (N_7049,N_6888,N_6713);
and U7050 (N_7050,N_6525,N_6685);
nand U7051 (N_7051,N_6708,N_6810);
nor U7052 (N_7052,N_6625,N_6612);
and U7053 (N_7053,N_6790,N_6965);
nand U7054 (N_7054,N_6616,N_6803);
or U7055 (N_7055,N_6739,N_6544);
and U7056 (N_7056,N_6724,N_6892);
and U7057 (N_7057,N_6526,N_6608);
nand U7058 (N_7058,N_6654,N_6828);
and U7059 (N_7059,N_6549,N_6598);
nand U7060 (N_7060,N_6882,N_6702);
nand U7061 (N_7061,N_6771,N_6588);
or U7062 (N_7062,N_6797,N_6633);
nor U7063 (N_7063,N_6681,N_6505);
or U7064 (N_7064,N_6722,N_6923);
xnor U7065 (N_7065,N_6659,N_6872);
nand U7066 (N_7066,N_6591,N_6709);
nor U7067 (N_7067,N_6660,N_6716);
nor U7068 (N_7068,N_6621,N_6733);
or U7069 (N_7069,N_6678,N_6569);
nor U7070 (N_7070,N_6731,N_6574);
nand U7071 (N_7071,N_6714,N_6862);
and U7072 (N_7072,N_6645,N_6866);
and U7073 (N_7073,N_6741,N_6558);
and U7074 (N_7074,N_6876,N_6750);
and U7075 (N_7075,N_6581,N_6982);
xor U7076 (N_7076,N_6503,N_6728);
nand U7077 (N_7077,N_6978,N_6630);
nand U7078 (N_7078,N_6804,N_6662);
nor U7079 (N_7079,N_6852,N_6979);
nand U7080 (N_7080,N_6870,N_6587);
and U7081 (N_7081,N_6551,N_6805);
nor U7082 (N_7082,N_6934,N_6538);
nand U7083 (N_7083,N_6824,N_6980);
or U7084 (N_7084,N_6917,N_6795);
and U7085 (N_7085,N_6942,N_6999);
or U7086 (N_7086,N_6635,N_6791);
and U7087 (N_7087,N_6773,N_6809);
xor U7088 (N_7088,N_6565,N_6704);
or U7089 (N_7089,N_6687,N_6744);
or U7090 (N_7090,N_6912,N_6971);
nand U7091 (N_7091,N_6829,N_6554);
nor U7092 (N_7092,N_6859,N_6585);
xor U7093 (N_7093,N_6513,N_6865);
nor U7094 (N_7094,N_6995,N_6622);
nor U7095 (N_7095,N_6627,N_6665);
or U7096 (N_7096,N_6973,N_6853);
and U7097 (N_7097,N_6547,N_6933);
or U7098 (N_7098,N_6792,N_6840);
xor U7099 (N_7099,N_6871,N_6703);
and U7100 (N_7100,N_6961,N_6512);
and U7101 (N_7101,N_6508,N_6567);
or U7102 (N_7102,N_6666,N_6602);
or U7103 (N_7103,N_6832,N_6956);
or U7104 (N_7104,N_6788,N_6536);
nand U7105 (N_7105,N_6550,N_6717);
and U7106 (N_7106,N_6661,N_6543);
and U7107 (N_7107,N_6523,N_6589);
or U7108 (N_7108,N_6757,N_6793);
and U7109 (N_7109,N_6566,N_6692);
nor U7110 (N_7110,N_6799,N_6629);
nand U7111 (N_7111,N_6777,N_6590);
and U7112 (N_7112,N_6874,N_6904);
xor U7113 (N_7113,N_6900,N_6725);
and U7114 (N_7114,N_6729,N_6963);
xnor U7115 (N_7115,N_6573,N_6895);
xnor U7116 (N_7116,N_6814,N_6509);
nor U7117 (N_7117,N_6700,N_6742);
nor U7118 (N_7118,N_6571,N_6764);
nand U7119 (N_7119,N_6924,N_6735);
and U7120 (N_7120,N_6986,N_6606);
nand U7121 (N_7121,N_6770,N_6592);
and U7122 (N_7122,N_6578,N_6737);
nor U7123 (N_7123,N_6864,N_6715);
and U7124 (N_7124,N_6532,N_6877);
and U7125 (N_7125,N_6851,N_6619);
nand U7126 (N_7126,N_6915,N_6652);
or U7127 (N_7127,N_6639,N_6579);
xor U7128 (N_7128,N_6563,N_6774);
nand U7129 (N_7129,N_6899,N_6931);
nand U7130 (N_7130,N_6674,N_6987);
and U7131 (N_7131,N_6753,N_6712);
and U7132 (N_7132,N_6796,N_6827);
nand U7133 (N_7133,N_6643,N_6968);
and U7134 (N_7134,N_6919,N_6746);
and U7135 (N_7135,N_6561,N_6897);
or U7136 (N_7136,N_6932,N_6760);
nor U7137 (N_7137,N_6552,N_6998);
nor U7138 (N_7138,N_6601,N_6719);
or U7139 (N_7139,N_6734,N_6922);
nand U7140 (N_7140,N_6649,N_6926);
nand U7141 (N_7141,N_6763,N_6531);
and U7142 (N_7142,N_6984,N_6992);
xnor U7143 (N_7143,N_6594,N_6868);
and U7144 (N_7144,N_6891,N_6997);
and U7145 (N_7145,N_6854,N_6684);
xnor U7146 (N_7146,N_6812,N_6946);
nand U7147 (N_7147,N_6584,N_6921);
nand U7148 (N_7148,N_6825,N_6546);
nand U7149 (N_7149,N_6972,N_6875);
nand U7150 (N_7150,N_6723,N_6711);
nor U7151 (N_7151,N_6781,N_6624);
and U7152 (N_7152,N_6988,N_6749);
nor U7153 (N_7153,N_6858,N_6836);
nor U7154 (N_7154,N_6878,N_6943);
nand U7155 (N_7155,N_6593,N_6586);
or U7156 (N_7156,N_6756,N_6981);
or U7157 (N_7157,N_6510,N_6950);
and U7158 (N_7158,N_6758,N_6863);
nand U7159 (N_7159,N_6528,N_6556);
nor U7160 (N_7160,N_6947,N_6553);
xor U7161 (N_7161,N_6860,N_6636);
and U7162 (N_7162,N_6937,N_6522);
xnor U7163 (N_7163,N_6607,N_6842);
and U7164 (N_7164,N_6647,N_6808);
xor U7165 (N_7165,N_6807,N_6576);
or U7166 (N_7166,N_6816,N_6535);
nor U7167 (N_7167,N_6653,N_6881);
nor U7168 (N_7168,N_6841,N_6906);
xor U7169 (N_7169,N_6844,N_6850);
or U7170 (N_7170,N_6767,N_6540);
or U7171 (N_7171,N_6964,N_6938);
and U7172 (N_7172,N_6949,N_6580);
nor U7173 (N_7173,N_6977,N_6655);
xnor U7174 (N_7174,N_6676,N_6747);
nand U7175 (N_7175,N_6768,N_6516);
nand U7176 (N_7176,N_6886,N_6718);
nand U7177 (N_7177,N_6693,N_6967);
xor U7178 (N_7178,N_6905,N_6686);
or U7179 (N_7179,N_6901,N_6694);
or U7180 (N_7180,N_6787,N_6560);
and U7181 (N_7181,N_6529,N_6690);
or U7182 (N_7182,N_6570,N_6884);
nand U7183 (N_7183,N_6557,N_6668);
and U7184 (N_7184,N_6823,N_6801);
nand U7185 (N_7185,N_6501,N_6572);
nand U7186 (N_7186,N_6604,N_6658);
nor U7187 (N_7187,N_6669,N_6811);
nor U7188 (N_7188,N_6615,N_6772);
or U7189 (N_7189,N_6848,N_6646);
xor U7190 (N_7190,N_6524,N_6752);
and U7191 (N_7191,N_6784,N_6521);
nor U7192 (N_7192,N_6944,N_6644);
xor U7193 (N_7193,N_6873,N_6511);
nand U7194 (N_7194,N_6798,N_6957);
or U7195 (N_7195,N_6754,N_6948);
nand U7196 (N_7196,N_6908,N_6555);
nand U7197 (N_7197,N_6815,N_6626);
and U7198 (N_7198,N_6806,N_6966);
or U7199 (N_7199,N_6623,N_6889);
nor U7200 (N_7200,N_6843,N_6820);
and U7201 (N_7201,N_6759,N_6611);
xnor U7202 (N_7202,N_6670,N_6830);
nor U7203 (N_7203,N_6856,N_6518);
or U7204 (N_7204,N_6786,N_6527);
xor U7205 (N_7205,N_6765,N_6969);
and U7206 (N_7206,N_6762,N_6642);
nand U7207 (N_7207,N_6651,N_6680);
and U7208 (N_7208,N_6603,N_6896);
and U7209 (N_7209,N_6930,N_6620);
and U7210 (N_7210,N_6833,N_6618);
and U7211 (N_7211,N_6548,N_6520);
or U7212 (N_7212,N_6559,N_6706);
nand U7213 (N_7213,N_6869,N_6819);
xor U7214 (N_7214,N_6927,N_6634);
and U7215 (N_7215,N_6958,N_6783);
and U7216 (N_7216,N_6631,N_6893);
or U7217 (N_7217,N_6818,N_6802);
nor U7218 (N_7218,N_6940,N_6910);
nand U7219 (N_7219,N_6794,N_6831);
nor U7220 (N_7220,N_6847,N_6721);
xnor U7221 (N_7221,N_6993,N_6855);
or U7222 (N_7222,N_6890,N_6534);
xor U7223 (N_7223,N_6883,N_6600);
or U7224 (N_7224,N_6609,N_6679);
nand U7225 (N_7225,N_6951,N_6960);
nor U7226 (N_7226,N_6564,N_6545);
or U7227 (N_7227,N_6909,N_6857);
or U7228 (N_7228,N_6782,N_6696);
nand U7229 (N_7229,N_6902,N_6705);
nor U7230 (N_7230,N_6838,N_6983);
or U7231 (N_7231,N_6936,N_6776);
nand U7232 (N_7232,N_6689,N_6726);
and U7233 (N_7233,N_6688,N_6577);
xor U7234 (N_7234,N_6673,N_6916);
and U7235 (N_7235,N_6745,N_6880);
and U7236 (N_7236,N_6996,N_6826);
nand U7237 (N_7237,N_6975,N_6849);
nand U7238 (N_7238,N_6605,N_6779);
or U7239 (N_7239,N_6695,N_6994);
nor U7240 (N_7240,N_6976,N_6583);
and U7241 (N_7241,N_6701,N_6821);
nand U7242 (N_7242,N_6834,N_6738);
nor U7243 (N_7243,N_6736,N_6789);
or U7244 (N_7244,N_6648,N_6989);
nor U7245 (N_7245,N_6751,N_6707);
nand U7246 (N_7246,N_6575,N_6952);
or U7247 (N_7247,N_6514,N_6822);
nand U7248 (N_7248,N_6730,N_6597);
or U7249 (N_7249,N_6867,N_6530);
nand U7250 (N_7250,N_6758,N_6526);
nand U7251 (N_7251,N_6658,N_6872);
and U7252 (N_7252,N_6547,N_6921);
or U7253 (N_7253,N_6932,N_6737);
nor U7254 (N_7254,N_6751,N_6590);
or U7255 (N_7255,N_6618,N_6718);
nand U7256 (N_7256,N_6745,N_6628);
nand U7257 (N_7257,N_6887,N_6849);
and U7258 (N_7258,N_6622,N_6787);
or U7259 (N_7259,N_6962,N_6812);
or U7260 (N_7260,N_6511,N_6703);
nand U7261 (N_7261,N_6962,N_6674);
nor U7262 (N_7262,N_6863,N_6955);
and U7263 (N_7263,N_6584,N_6993);
nor U7264 (N_7264,N_6940,N_6777);
or U7265 (N_7265,N_6649,N_6817);
and U7266 (N_7266,N_6733,N_6825);
or U7267 (N_7267,N_6899,N_6701);
nand U7268 (N_7268,N_6592,N_6656);
and U7269 (N_7269,N_6563,N_6550);
nor U7270 (N_7270,N_6715,N_6702);
nor U7271 (N_7271,N_6929,N_6966);
nor U7272 (N_7272,N_6681,N_6574);
nor U7273 (N_7273,N_6639,N_6728);
and U7274 (N_7274,N_6807,N_6737);
or U7275 (N_7275,N_6773,N_6599);
nand U7276 (N_7276,N_6941,N_6666);
and U7277 (N_7277,N_6768,N_6810);
or U7278 (N_7278,N_6620,N_6810);
and U7279 (N_7279,N_6780,N_6910);
nand U7280 (N_7280,N_6501,N_6610);
nand U7281 (N_7281,N_6804,N_6706);
nand U7282 (N_7282,N_6675,N_6791);
or U7283 (N_7283,N_6517,N_6813);
or U7284 (N_7284,N_6706,N_6708);
xor U7285 (N_7285,N_6501,N_6545);
nand U7286 (N_7286,N_6888,N_6779);
nor U7287 (N_7287,N_6925,N_6819);
nor U7288 (N_7288,N_6866,N_6894);
or U7289 (N_7289,N_6737,N_6876);
nor U7290 (N_7290,N_6949,N_6889);
nand U7291 (N_7291,N_6508,N_6543);
or U7292 (N_7292,N_6952,N_6805);
xnor U7293 (N_7293,N_6877,N_6737);
nor U7294 (N_7294,N_6929,N_6814);
nor U7295 (N_7295,N_6695,N_6830);
or U7296 (N_7296,N_6906,N_6724);
nand U7297 (N_7297,N_6628,N_6688);
nand U7298 (N_7298,N_6748,N_6719);
and U7299 (N_7299,N_6946,N_6990);
nor U7300 (N_7300,N_6601,N_6926);
nor U7301 (N_7301,N_6817,N_6529);
xnor U7302 (N_7302,N_6548,N_6868);
nand U7303 (N_7303,N_6733,N_6747);
and U7304 (N_7304,N_6977,N_6503);
xnor U7305 (N_7305,N_6996,N_6580);
nand U7306 (N_7306,N_6748,N_6976);
nor U7307 (N_7307,N_6927,N_6539);
or U7308 (N_7308,N_6543,N_6522);
and U7309 (N_7309,N_6948,N_6666);
xor U7310 (N_7310,N_6976,N_6692);
or U7311 (N_7311,N_6766,N_6754);
nand U7312 (N_7312,N_6867,N_6774);
nand U7313 (N_7313,N_6833,N_6709);
nand U7314 (N_7314,N_6801,N_6968);
nand U7315 (N_7315,N_6880,N_6751);
nor U7316 (N_7316,N_6967,N_6711);
nor U7317 (N_7317,N_6556,N_6855);
or U7318 (N_7318,N_6948,N_6908);
xnor U7319 (N_7319,N_6875,N_6786);
or U7320 (N_7320,N_6761,N_6976);
or U7321 (N_7321,N_6919,N_6856);
and U7322 (N_7322,N_6771,N_6675);
or U7323 (N_7323,N_6706,N_6639);
or U7324 (N_7324,N_6653,N_6758);
and U7325 (N_7325,N_6899,N_6952);
and U7326 (N_7326,N_6565,N_6586);
nand U7327 (N_7327,N_6524,N_6572);
xor U7328 (N_7328,N_6883,N_6760);
or U7329 (N_7329,N_6506,N_6673);
and U7330 (N_7330,N_6823,N_6900);
xor U7331 (N_7331,N_6796,N_6969);
xnor U7332 (N_7332,N_6911,N_6923);
and U7333 (N_7333,N_6954,N_6982);
nor U7334 (N_7334,N_6549,N_6583);
nand U7335 (N_7335,N_6743,N_6691);
or U7336 (N_7336,N_6915,N_6576);
or U7337 (N_7337,N_6541,N_6851);
nor U7338 (N_7338,N_6650,N_6946);
xor U7339 (N_7339,N_6726,N_6951);
nand U7340 (N_7340,N_6751,N_6566);
nand U7341 (N_7341,N_6962,N_6755);
nand U7342 (N_7342,N_6912,N_6569);
nor U7343 (N_7343,N_6502,N_6572);
nor U7344 (N_7344,N_6660,N_6872);
and U7345 (N_7345,N_6742,N_6796);
and U7346 (N_7346,N_6611,N_6931);
and U7347 (N_7347,N_6570,N_6692);
xnor U7348 (N_7348,N_6992,N_6857);
and U7349 (N_7349,N_6956,N_6899);
nand U7350 (N_7350,N_6880,N_6705);
nand U7351 (N_7351,N_6714,N_6680);
or U7352 (N_7352,N_6546,N_6629);
nor U7353 (N_7353,N_6943,N_6816);
and U7354 (N_7354,N_6561,N_6507);
xor U7355 (N_7355,N_6985,N_6505);
xor U7356 (N_7356,N_6552,N_6723);
nand U7357 (N_7357,N_6723,N_6666);
nand U7358 (N_7358,N_6679,N_6861);
or U7359 (N_7359,N_6629,N_6556);
or U7360 (N_7360,N_6645,N_6869);
or U7361 (N_7361,N_6752,N_6789);
or U7362 (N_7362,N_6551,N_6527);
nand U7363 (N_7363,N_6701,N_6568);
or U7364 (N_7364,N_6761,N_6832);
or U7365 (N_7365,N_6753,N_6501);
or U7366 (N_7366,N_6936,N_6749);
or U7367 (N_7367,N_6980,N_6642);
and U7368 (N_7368,N_6591,N_6532);
or U7369 (N_7369,N_6965,N_6985);
and U7370 (N_7370,N_6563,N_6802);
and U7371 (N_7371,N_6844,N_6573);
nand U7372 (N_7372,N_6942,N_6552);
or U7373 (N_7373,N_6844,N_6791);
or U7374 (N_7374,N_6841,N_6887);
or U7375 (N_7375,N_6905,N_6607);
and U7376 (N_7376,N_6942,N_6661);
xor U7377 (N_7377,N_6607,N_6611);
and U7378 (N_7378,N_6996,N_6624);
and U7379 (N_7379,N_6818,N_6966);
nand U7380 (N_7380,N_6849,N_6525);
xor U7381 (N_7381,N_6621,N_6764);
nor U7382 (N_7382,N_6896,N_6723);
nand U7383 (N_7383,N_6992,N_6733);
xor U7384 (N_7384,N_6540,N_6897);
nor U7385 (N_7385,N_6852,N_6777);
and U7386 (N_7386,N_6779,N_6506);
or U7387 (N_7387,N_6922,N_6809);
and U7388 (N_7388,N_6793,N_6658);
nand U7389 (N_7389,N_6862,N_6829);
and U7390 (N_7390,N_6911,N_6649);
and U7391 (N_7391,N_6892,N_6738);
or U7392 (N_7392,N_6973,N_6865);
nor U7393 (N_7393,N_6509,N_6644);
or U7394 (N_7394,N_6550,N_6920);
or U7395 (N_7395,N_6772,N_6654);
or U7396 (N_7396,N_6663,N_6652);
nor U7397 (N_7397,N_6865,N_6559);
or U7398 (N_7398,N_6963,N_6645);
or U7399 (N_7399,N_6537,N_6987);
nand U7400 (N_7400,N_6679,N_6527);
or U7401 (N_7401,N_6595,N_6636);
nand U7402 (N_7402,N_6583,N_6847);
nand U7403 (N_7403,N_6919,N_6719);
nor U7404 (N_7404,N_6924,N_6809);
or U7405 (N_7405,N_6677,N_6820);
or U7406 (N_7406,N_6702,N_6909);
nor U7407 (N_7407,N_6751,N_6827);
nor U7408 (N_7408,N_6637,N_6918);
or U7409 (N_7409,N_6718,N_6640);
or U7410 (N_7410,N_6792,N_6698);
and U7411 (N_7411,N_6916,N_6649);
xor U7412 (N_7412,N_6608,N_6984);
nand U7413 (N_7413,N_6611,N_6708);
or U7414 (N_7414,N_6689,N_6904);
or U7415 (N_7415,N_6723,N_6709);
nand U7416 (N_7416,N_6710,N_6769);
nor U7417 (N_7417,N_6811,N_6826);
nand U7418 (N_7418,N_6654,N_6710);
nor U7419 (N_7419,N_6953,N_6905);
xnor U7420 (N_7420,N_6918,N_6936);
nor U7421 (N_7421,N_6640,N_6857);
or U7422 (N_7422,N_6517,N_6889);
or U7423 (N_7423,N_6853,N_6927);
nand U7424 (N_7424,N_6925,N_6810);
nand U7425 (N_7425,N_6520,N_6517);
or U7426 (N_7426,N_6619,N_6837);
nand U7427 (N_7427,N_6692,N_6516);
or U7428 (N_7428,N_6695,N_6892);
or U7429 (N_7429,N_6650,N_6545);
nor U7430 (N_7430,N_6575,N_6845);
and U7431 (N_7431,N_6742,N_6930);
or U7432 (N_7432,N_6938,N_6781);
or U7433 (N_7433,N_6936,N_6765);
nor U7434 (N_7434,N_6872,N_6852);
nor U7435 (N_7435,N_6835,N_6607);
nand U7436 (N_7436,N_6542,N_6628);
and U7437 (N_7437,N_6659,N_6597);
nor U7438 (N_7438,N_6823,N_6693);
xnor U7439 (N_7439,N_6945,N_6830);
nand U7440 (N_7440,N_6808,N_6541);
or U7441 (N_7441,N_6711,N_6937);
nor U7442 (N_7442,N_6797,N_6877);
or U7443 (N_7443,N_6767,N_6755);
or U7444 (N_7444,N_6541,N_6543);
nor U7445 (N_7445,N_6974,N_6504);
xnor U7446 (N_7446,N_6680,N_6911);
nand U7447 (N_7447,N_6800,N_6578);
nor U7448 (N_7448,N_6633,N_6778);
xnor U7449 (N_7449,N_6736,N_6697);
nor U7450 (N_7450,N_6543,N_6854);
xor U7451 (N_7451,N_6662,N_6836);
nor U7452 (N_7452,N_6514,N_6923);
or U7453 (N_7453,N_6793,N_6766);
nand U7454 (N_7454,N_6676,N_6843);
nand U7455 (N_7455,N_6882,N_6667);
and U7456 (N_7456,N_6700,N_6807);
xnor U7457 (N_7457,N_6715,N_6785);
and U7458 (N_7458,N_6979,N_6942);
xor U7459 (N_7459,N_6680,N_6774);
and U7460 (N_7460,N_6832,N_6579);
and U7461 (N_7461,N_6559,N_6810);
nor U7462 (N_7462,N_6606,N_6763);
xor U7463 (N_7463,N_6563,N_6709);
nor U7464 (N_7464,N_6749,N_6606);
or U7465 (N_7465,N_6636,N_6750);
or U7466 (N_7466,N_6579,N_6835);
or U7467 (N_7467,N_6990,N_6879);
nor U7468 (N_7468,N_6992,N_6777);
xor U7469 (N_7469,N_6714,N_6783);
nor U7470 (N_7470,N_6737,N_6540);
nand U7471 (N_7471,N_6855,N_6946);
or U7472 (N_7472,N_6883,N_6859);
nor U7473 (N_7473,N_6950,N_6944);
and U7474 (N_7474,N_6724,N_6713);
nor U7475 (N_7475,N_6839,N_6922);
nor U7476 (N_7476,N_6583,N_6825);
nand U7477 (N_7477,N_6720,N_6965);
or U7478 (N_7478,N_6778,N_6529);
nor U7479 (N_7479,N_6601,N_6754);
and U7480 (N_7480,N_6639,N_6560);
nor U7481 (N_7481,N_6745,N_6705);
and U7482 (N_7482,N_6586,N_6691);
nand U7483 (N_7483,N_6675,N_6690);
and U7484 (N_7484,N_6605,N_6695);
and U7485 (N_7485,N_6966,N_6833);
xnor U7486 (N_7486,N_6618,N_6905);
and U7487 (N_7487,N_6708,N_6767);
nor U7488 (N_7488,N_6729,N_6576);
nor U7489 (N_7489,N_6538,N_6792);
and U7490 (N_7490,N_6582,N_6724);
or U7491 (N_7491,N_6631,N_6726);
nor U7492 (N_7492,N_6908,N_6893);
or U7493 (N_7493,N_6801,N_6584);
xor U7494 (N_7494,N_6773,N_6525);
and U7495 (N_7495,N_6720,N_6968);
xnor U7496 (N_7496,N_6915,N_6624);
nor U7497 (N_7497,N_6909,N_6820);
or U7498 (N_7498,N_6757,N_6975);
or U7499 (N_7499,N_6557,N_6658);
nor U7500 (N_7500,N_7188,N_7454);
or U7501 (N_7501,N_7385,N_7119);
or U7502 (N_7502,N_7296,N_7475);
nand U7503 (N_7503,N_7068,N_7148);
or U7504 (N_7504,N_7203,N_7184);
nand U7505 (N_7505,N_7223,N_7459);
nand U7506 (N_7506,N_7431,N_7329);
or U7507 (N_7507,N_7001,N_7158);
nand U7508 (N_7508,N_7395,N_7298);
nor U7509 (N_7509,N_7392,N_7266);
nor U7510 (N_7510,N_7433,N_7198);
nand U7511 (N_7511,N_7069,N_7353);
nor U7512 (N_7512,N_7421,N_7348);
and U7513 (N_7513,N_7036,N_7293);
or U7514 (N_7514,N_7383,N_7321);
or U7515 (N_7515,N_7343,N_7129);
and U7516 (N_7516,N_7291,N_7160);
and U7517 (N_7517,N_7281,N_7252);
or U7518 (N_7518,N_7088,N_7074);
nor U7519 (N_7519,N_7403,N_7190);
nand U7520 (N_7520,N_7164,N_7155);
or U7521 (N_7521,N_7081,N_7194);
nand U7522 (N_7522,N_7241,N_7393);
or U7523 (N_7523,N_7378,N_7330);
nor U7524 (N_7524,N_7286,N_7331);
nand U7525 (N_7525,N_7104,N_7031);
and U7526 (N_7526,N_7018,N_7213);
and U7527 (N_7527,N_7206,N_7280);
nor U7528 (N_7528,N_7128,N_7492);
nand U7529 (N_7529,N_7022,N_7046);
and U7530 (N_7530,N_7010,N_7204);
nand U7531 (N_7531,N_7019,N_7245);
nor U7532 (N_7532,N_7217,N_7272);
nor U7533 (N_7533,N_7114,N_7359);
and U7534 (N_7534,N_7028,N_7312);
and U7535 (N_7535,N_7000,N_7465);
or U7536 (N_7536,N_7288,N_7024);
or U7537 (N_7537,N_7029,N_7290);
nor U7538 (N_7538,N_7169,N_7166);
and U7539 (N_7539,N_7450,N_7432);
or U7540 (N_7540,N_7175,N_7186);
nor U7541 (N_7541,N_7411,N_7409);
nor U7542 (N_7542,N_7357,N_7248);
and U7543 (N_7543,N_7285,N_7368);
nor U7544 (N_7544,N_7275,N_7261);
and U7545 (N_7545,N_7082,N_7294);
nand U7546 (N_7546,N_7376,N_7137);
and U7547 (N_7547,N_7373,N_7415);
and U7548 (N_7548,N_7192,N_7308);
nor U7549 (N_7549,N_7416,N_7447);
xor U7550 (N_7550,N_7300,N_7140);
or U7551 (N_7551,N_7159,N_7320);
xor U7552 (N_7552,N_7101,N_7078);
xnor U7553 (N_7553,N_7356,N_7058);
nor U7554 (N_7554,N_7136,N_7344);
nor U7555 (N_7555,N_7438,N_7076);
nand U7556 (N_7556,N_7458,N_7180);
nand U7557 (N_7557,N_7045,N_7236);
xor U7558 (N_7558,N_7048,N_7146);
nand U7559 (N_7559,N_7259,N_7299);
and U7560 (N_7560,N_7407,N_7044);
or U7561 (N_7561,N_7151,N_7077);
xor U7562 (N_7562,N_7485,N_7212);
nand U7563 (N_7563,N_7173,N_7424);
nor U7564 (N_7564,N_7349,N_7242);
and U7565 (N_7565,N_7418,N_7142);
or U7566 (N_7566,N_7215,N_7362);
xnor U7567 (N_7567,N_7319,N_7209);
nand U7568 (N_7568,N_7282,N_7115);
nand U7569 (N_7569,N_7391,N_7276);
nand U7570 (N_7570,N_7253,N_7381);
nand U7571 (N_7571,N_7066,N_7124);
and U7572 (N_7572,N_7480,N_7254);
or U7573 (N_7573,N_7419,N_7020);
xor U7574 (N_7574,N_7205,N_7191);
or U7575 (N_7575,N_7322,N_7352);
and U7576 (N_7576,N_7176,N_7084);
and U7577 (N_7577,N_7455,N_7039);
and U7578 (N_7578,N_7444,N_7310);
nor U7579 (N_7579,N_7038,N_7086);
or U7580 (N_7580,N_7334,N_7149);
or U7581 (N_7581,N_7496,N_7161);
xor U7582 (N_7582,N_7333,N_7139);
nand U7583 (N_7583,N_7478,N_7145);
xnor U7584 (N_7584,N_7013,N_7218);
nor U7585 (N_7585,N_7097,N_7225);
nor U7586 (N_7586,N_7477,N_7179);
nand U7587 (N_7587,N_7273,N_7072);
nor U7588 (N_7588,N_7420,N_7351);
xnor U7589 (N_7589,N_7135,N_7283);
and U7590 (N_7590,N_7345,N_7093);
or U7591 (N_7591,N_7486,N_7240);
and U7592 (N_7592,N_7152,N_7092);
and U7593 (N_7593,N_7441,N_7361);
nand U7594 (N_7594,N_7167,N_7274);
and U7595 (N_7595,N_7462,N_7346);
and U7596 (N_7596,N_7413,N_7055);
and U7597 (N_7597,N_7335,N_7111);
nor U7598 (N_7598,N_7047,N_7228);
and U7599 (N_7599,N_7121,N_7023);
nand U7600 (N_7600,N_7095,N_7439);
or U7601 (N_7601,N_7292,N_7452);
and U7602 (N_7602,N_7182,N_7040);
nor U7603 (N_7603,N_7295,N_7473);
nand U7604 (N_7604,N_7318,N_7263);
and U7605 (N_7605,N_7165,N_7127);
xnor U7606 (N_7606,N_7302,N_7015);
nand U7607 (N_7607,N_7487,N_7289);
nand U7608 (N_7608,N_7436,N_7163);
and U7609 (N_7609,N_7355,N_7340);
or U7610 (N_7610,N_7270,N_7075);
xnor U7611 (N_7611,N_7278,N_7417);
or U7612 (N_7612,N_7109,N_7133);
and U7613 (N_7613,N_7143,N_7265);
and U7614 (N_7614,N_7037,N_7153);
nor U7615 (N_7615,N_7157,N_7277);
or U7616 (N_7616,N_7354,N_7162);
and U7617 (N_7617,N_7434,N_7035);
nand U7618 (N_7618,N_7399,N_7414);
or U7619 (N_7619,N_7271,N_7379);
xnor U7620 (N_7620,N_7112,N_7369);
and U7621 (N_7621,N_7033,N_7249);
or U7622 (N_7622,N_7107,N_7118);
nand U7623 (N_7623,N_7269,N_7233);
or U7624 (N_7624,N_7073,N_7187);
nand U7625 (N_7625,N_7490,N_7126);
or U7626 (N_7626,N_7006,N_7105);
or U7627 (N_7627,N_7460,N_7284);
or U7628 (N_7628,N_7339,N_7117);
nand U7629 (N_7629,N_7375,N_7065);
or U7630 (N_7630,N_7400,N_7017);
or U7631 (N_7631,N_7437,N_7493);
nand U7632 (N_7632,N_7096,N_7472);
nand U7633 (N_7633,N_7260,N_7232);
nand U7634 (N_7634,N_7174,N_7430);
nand U7635 (N_7635,N_7134,N_7138);
nor U7636 (N_7636,N_7262,N_7324);
nor U7637 (N_7637,N_7482,N_7364);
nor U7638 (N_7638,N_7014,N_7476);
nand U7639 (N_7639,N_7484,N_7326);
xor U7640 (N_7640,N_7387,N_7427);
nor U7641 (N_7641,N_7264,N_7305);
xor U7642 (N_7642,N_7085,N_7311);
and U7643 (N_7643,N_7464,N_7398);
nor U7644 (N_7644,N_7440,N_7234);
and U7645 (N_7645,N_7250,N_7062);
or U7646 (N_7646,N_7297,N_7216);
xor U7647 (N_7647,N_7102,N_7230);
nor U7648 (N_7648,N_7094,N_7202);
and U7649 (N_7649,N_7497,N_7199);
and U7650 (N_7650,N_7314,N_7113);
and U7651 (N_7651,N_7374,N_7195);
nand U7652 (N_7652,N_7483,N_7489);
nand U7653 (N_7653,N_7172,N_7193);
or U7654 (N_7654,N_7005,N_7007);
and U7655 (N_7655,N_7309,N_7168);
nor U7656 (N_7656,N_7004,N_7287);
nor U7657 (N_7657,N_7003,N_7200);
nor U7658 (N_7658,N_7422,N_7222);
and U7659 (N_7659,N_7388,N_7238);
nand U7660 (N_7660,N_7426,N_7453);
nand U7661 (N_7661,N_7367,N_7012);
or U7662 (N_7662,N_7246,N_7443);
and U7663 (N_7663,N_7408,N_7057);
xor U7664 (N_7664,N_7214,N_7009);
or U7665 (N_7665,N_7435,N_7061);
nand U7666 (N_7666,N_7389,N_7177);
nor U7667 (N_7667,N_7327,N_7108);
nor U7668 (N_7668,N_7406,N_7323);
and U7669 (N_7669,N_7481,N_7197);
or U7670 (N_7670,N_7103,N_7243);
nand U7671 (N_7671,N_7207,N_7456);
or U7672 (N_7672,N_7042,N_7201);
and U7673 (N_7673,N_7110,N_7171);
and U7674 (N_7674,N_7052,N_7499);
nor U7675 (N_7675,N_7377,N_7116);
nor U7676 (N_7676,N_7067,N_7247);
nor U7677 (N_7677,N_7258,N_7396);
nand U7678 (N_7678,N_7027,N_7231);
or U7679 (N_7679,N_7041,N_7170);
nand U7680 (N_7680,N_7227,N_7196);
nor U7681 (N_7681,N_7123,N_7071);
or U7682 (N_7682,N_7394,N_7423);
and U7683 (N_7683,N_7342,N_7132);
or U7684 (N_7684,N_7008,N_7016);
and U7685 (N_7685,N_7026,N_7050);
or U7686 (N_7686,N_7366,N_7079);
nand U7687 (N_7687,N_7470,N_7156);
nand U7688 (N_7688,N_7498,N_7144);
nand U7689 (N_7689,N_7181,N_7358);
xor U7690 (N_7690,N_7474,N_7446);
nor U7691 (N_7691,N_7428,N_7043);
nand U7692 (N_7692,N_7150,N_7466);
nor U7693 (N_7693,N_7221,N_7063);
nand U7694 (N_7694,N_7030,N_7099);
or U7695 (N_7695,N_7235,N_7060);
nor U7696 (N_7696,N_7316,N_7106);
or U7697 (N_7697,N_7479,N_7380);
and U7698 (N_7698,N_7336,N_7051);
or U7699 (N_7699,N_7468,N_7226);
nor U7700 (N_7700,N_7384,N_7494);
and U7701 (N_7701,N_7087,N_7338);
nand U7702 (N_7702,N_7495,N_7328);
or U7703 (N_7703,N_7341,N_7315);
and U7704 (N_7704,N_7131,N_7491);
nand U7705 (N_7705,N_7224,N_7448);
and U7706 (N_7706,N_7463,N_7365);
nand U7707 (N_7707,N_7429,N_7125);
xnor U7708 (N_7708,N_7091,N_7053);
or U7709 (N_7709,N_7332,N_7021);
xnor U7710 (N_7710,N_7350,N_7467);
nand U7711 (N_7711,N_7154,N_7239);
and U7712 (N_7712,N_7363,N_7056);
nor U7713 (N_7713,N_7451,N_7471);
nor U7714 (N_7714,N_7229,N_7059);
nor U7715 (N_7715,N_7244,N_7268);
xnor U7716 (N_7716,N_7442,N_7313);
nand U7717 (N_7717,N_7301,N_7401);
or U7718 (N_7718,N_7189,N_7461);
nand U7719 (N_7719,N_7210,N_7410);
nor U7720 (N_7720,N_7337,N_7141);
nor U7721 (N_7721,N_7185,N_7080);
nor U7722 (N_7722,N_7412,N_7390);
nor U7723 (N_7723,N_7025,N_7032);
nand U7724 (N_7724,N_7445,N_7070);
or U7725 (N_7725,N_7370,N_7303);
and U7726 (N_7726,N_7402,N_7089);
or U7727 (N_7727,N_7449,N_7317);
nand U7728 (N_7728,N_7279,N_7219);
and U7729 (N_7729,N_7011,N_7090);
nand U7730 (N_7730,N_7372,N_7347);
or U7731 (N_7731,N_7211,N_7267);
and U7732 (N_7732,N_7120,N_7054);
and U7733 (N_7733,N_7130,N_7002);
nand U7734 (N_7734,N_7304,N_7183);
nand U7735 (N_7735,N_7237,N_7425);
or U7736 (N_7736,N_7307,N_7360);
and U7737 (N_7737,N_7034,N_7469);
and U7738 (N_7738,N_7257,N_7122);
or U7739 (N_7739,N_7256,N_7208);
or U7740 (N_7740,N_7382,N_7100);
xor U7741 (N_7741,N_7397,N_7064);
nor U7742 (N_7742,N_7457,N_7306);
nand U7743 (N_7743,N_7049,N_7371);
xnor U7744 (N_7744,N_7405,N_7098);
and U7745 (N_7745,N_7220,N_7083);
nand U7746 (N_7746,N_7147,N_7488);
nor U7747 (N_7747,N_7386,N_7404);
and U7748 (N_7748,N_7255,N_7178);
nand U7749 (N_7749,N_7325,N_7251);
and U7750 (N_7750,N_7422,N_7319);
xnor U7751 (N_7751,N_7007,N_7346);
or U7752 (N_7752,N_7060,N_7222);
nand U7753 (N_7753,N_7178,N_7202);
xor U7754 (N_7754,N_7280,N_7204);
and U7755 (N_7755,N_7447,N_7192);
and U7756 (N_7756,N_7227,N_7014);
nor U7757 (N_7757,N_7410,N_7196);
or U7758 (N_7758,N_7127,N_7219);
nand U7759 (N_7759,N_7361,N_7054);
nor U7760 (N_7760,N_7332,N_7105);
nor U7761 (N_7761,N_7172,N_7180);
or U7762 (N_7762,N_7085,N_7486);
and U7763 (N_7763,N_7455,N_7152);
nand U7764 (N_7764,N_7027,N_7413);
and U7765 (N_7765,N_7308,N_7244);
nand U7766 (N_7766,N_7156,N_7384);
nand U7767 (N_7767,N_7223,N_7238);
nor U7768 (N_7768,N_7458,N_7072);
nand U7769 (N_7769,N_7200,N_7448);
xor U7770 (N_7770,N_7382,N_7116);
or U7771 (N_7771,N_7473,N_7225);
nand U7772 (N_7772,N_7214,N_7347);
xnor U7773 (N_7773,N_7065,N_7183);
or U7774 (N_7774,N_7384,N_7241);
nor U7775 (N_7775,N_7131,N_7143);
or U7776 (N_7776,N_7387,N_7458);
nand U7777 (N_7777,N_7289,N_7008);
nor U7778 (N_7778,N_7336,N_7084);
or U7779 (N_7779,N_7434,N_7233);
and U7780 (N_7780,N_7019,N_7420);
nor U7781 (N_7781,N_7205,N_7100);
nand U7782 (N_7782,N_7099,N_7353);
and U7783 (N_7783,N_7459,N_7328);
and U7784 (N_7784,N_7425,N_7341);
and U7785 (N_7785,N_7253,N_7460);
nand U7786 (N_7786,N_7413,N_7419);
nor U7787 (N_7787,N_7457,N_7189);
or U7788 (N_7788,N_7367,N_7247);
nand U7789 (N_7789,N_7237,N_7274);
nand U7790 (N_7790,N_7425,N_7384);
nor U7791 (N_7791,N_7092,N_7137);
or U7792 (N_7792,N_7359,N_7062);
and U7793 (N_7793,N_7286,N_7041);
nor U7794 (N_7794,N_7426,N_7221);
or U7795 (N_7795,N_7380,N_7493);
or U7796 (N_7796,N_7094,N_7384);
or U7797 (N_7797,N_7073,N_7366);
xnor U7798 (N_7798,N_7143,N_7304);
xnor U7799 (N_7799,N_7449,N_7214);
and U7800 (N_7800,N_7280,N_7319);
nand U7801 (N_7801,N_7303,N_7457);
nand U7802 (N_7802,N_7397,N_7062);
and U7803 (N_7803,N_7367,N_7449);
nor U7804 (N_7804,N_7323,N_7010);
and U7805 (N_7805,N_7353,N_7456);
nand U7806 (N_7806,N_7033,N_7449);
or U7807 (N_7807,N_7295,N_7325);
nor U7808 (N_7808,N_7076,N_7240);
xnor U7809 (N_7809,N_7239,N_7481);
and U7810 (N_7810,N_7398,N_7199);
or U7811 (N_7811,N_7342,N_7453);
and U7812 (N_7812,N_7086,N_7490);
nand U7813 (N_7813,N_7059,N_7123);
nor U7814 (N_7814,N_7311,N_7275);
and U7815 (N_7815,N_7154,N_7455);
and U7816 (N_7816,N_7224,N_7142);
nor U7817 (N_7817,N_7157,N_7334);
xnor U7818 (N_7818,N_7219,N_7360);
nor U7819 (N_7819,N_7435,N_7323);
nand U7820 (N_7820,N_7386,N_7442);
and U7821 (N_7821,N_7055,N_7071);
nand U7822 (N_7822,N_7172,N_7390);
xor U7823 (N_7823,N_7393,N_7037);
nor U7824 (N_7824,N_7339,N_7095);
and U7825 (N_7825,N_7237,N_7124);
and U7826 (N_7826,N_7379,N_7414);
nor U7827 (N_7827,N_7096,N_7259);
and U7828 (N_7828,N_7184,N_7242);
nand U7829 (N_7829,N_7069,N_7088);
nor U7830 (N_7830,N_7392,N_7347);
nor U7831 (N_7831,N_7091,N_7495);
and U7832 (N_7832,N_7103,N_7442);
nor U7833 (N_7833,N_7265,N_7070);
and U7834 (N_7834,N_7290,N_7249);
and U7835 (N_7835,N_7086,N_7253);
nand U7836 (N_7836,N_7321,N_7433);
or U7837 (N_7837,N_7138,N_7193);
nand U7838 (N_7838,N_7465,N_7419);
nor U7839 (N_7839,N_7248,N_7318);
or U7840 (N_7840,N_7497,N_7005);
or U7841 (N_7841,N_7079,N_7437);
or U7842 (N_7842,N_7082,N_7106);
nor U7843 (N_7843,N_7297,N_7401);
nand U7844 (N_7844,N_7215,N_7212);
nor U7845 (N_7845,N_7435,N_7234);
nor U7846 (N_7846,N_7063,N_7486);
nor U7847 (N_7847,N_7250,N_7352);
or U7848 (N_7848,N_7420,N_7025);
nand U7849 (N_7849,N_7456,N_7190);
nand U7850 (N_7850,N_7368,N_7064);
nor U7851 (N_7851,N_7476,N_7342);
and U7852 (N_7852,N_7190,N_7062);
and U7853 (N_7853,N_7429,N_7124);
nor U7854 (N_7854,N_7489,N_7136);
nand U7855 (N_7855,N_7225,N_7484);
nand U7856 (N_7856,N_7486,N_7263);
and U7857 (N_7857,N_7455,N_7356);
xor U7858 (N_7858,N_7200,N_7193);
or U7859 (N_7859,N_7100,N_7448);
nor U7860 (N_7860,N_7092,N_7075);
nand U7861 (N_7861,N_7066,N_7120);
and U7862 (N_7862,N_7241,N_7032);
or U7863 (N_7863,N_7351,N_7025);
and U7864 (N_7864,N_7444,N_7138);
nor U7865 (N_7865,N_7203,N_7476);
nor U7866 (N_7866,N_7495,N_7336);
nand U7867 (N_7867,N_7477,N_7361);
nand U7868 (N_7868,N_7383,N_7483);
xnor U7869 (N_7869,N_7108,N_7040);
nor U7870 (N_7870,N_7344,N_7242);
nor U7871 (N_7871,N_7005,N_7310);
or U7872 (N_7872,N_7024,N_7289);
and U7873 (N_7873,N_7311,N_7297);
xnor U7874 (N_7874,N_7419,N_7297);
or U7875 (N_7875,N_7455,N_7149);
xor U7876 (N_7876,N_7473,N_7113);
nand U7877 (N_7877,N_7380,N_7178);
and U7878 (N_7878,N_7295,N_7407);
and U7879 (N_7879,N_7003,N_7013);
xnor U7880 (N_7880,N_7292,N_7461);
nor U7881 (N_7881,N_7252,N_7009);
or U7882 (N_7882,N_7465,N_7141);
or U7883 (N_7883,N_7410,N_7120);
and U7884 (N_7884,N_7207,N_7401);
or U7885 (N_7885,N_7429,N_7206);
and U7886 (N_7886,N_7010,N_7210);
nand U7887 (N_7887,N_7062,N_7113);
or U7888 (N_7888,N_7134,N_7196);
xor U7889 (N_7889,N_7208,N_7317);
and U7890 (N_7890,N_7305,N_7454);
and U7891 (N_7891,N_7026,N_7114);
nor U7892 (N_7892,N_7211,N_7186);
nor U7893 (N_7893,N_7104,N_7281);
nor U7894 (N_7894,N_7366,N_7458);
or U7895 (N_7895,N_7448,N_7234);
nand U7896 (N_7896,N_7453,N_7102);
or U7897 (N_7897,N_7005,N_7308);
nor U7898 (N_7898,N_7312,N_7114);
nor U7899 (N_7899,N_7085,N_7027);
nand U7900 (N_7900,N_7488,N_7271);
nand U7901 (N_7901,N_7345,N_7173);
nand U7902 (N_7902,N_7253,N_7028);
or U7903 (N_7903,N_7335,N_7163);
or U7904 (N_7904,N_7421,N_7302);
nand U7905 (N_7905,N_7376,N_7231);
and U7906 (N_7906,N_7301,N_7076);
and U7907 (N_7907,N_7098,N_7026);
and U7908 (N_7908,N_7198,N_7399);
and U7909 (N_7909,N_7282,N_7189);
nand U7910 (N_7910,N_7370,N_7235);
nand U7911 (N_7911,N_7245,N_7337);
nor U7912 (N_7912,N_7285,N_7493);
nor U7913 (N_7913,N_7091,N_7151);
and U7914 (N_7914,N_7357,N_7193);
or U7915 (N_7915,N_7385,N_7230);
or U7916 (N_7916,N_7071,N_7419);
nor U7917 (N_7917,N_7284,N_7017);
nand U7918 (N_7918,N_7095,N_7040);
nor U7919 (N_7919,N_7473,N_7186);
or U7920 (N_7920,N_7237,N_7351);
and U7921 (N_7921,N_7323,N_7225);
or U7922 (N_7922,N_7305,N_7288);
nor U7923 (N_7923,N_7260,N_7244);
nand U7924 (N_7924,N_7279,N_7211);
nand U7925 (N_7925,N_7224,N_7093);
or U7926 (N_7926,N_7115,N_7022);
or U7927 (N_7927,N_7068,N_7127);
and U7928 (N_7928,N_7418,N_7331);
nor U7929 (N_7929,N_7320,N_7188);
nand U7930 (N_7930,N_7355,N_7010);
and U7931 (N_7931,N_7381,N_7441);
or U7932 (N_7932,N_7397,N_7270);
xnor U7933 (N_7933,N_7454,N_7358);
or U7934 (N_7934,N_7309,N_7264);
nor U7935 (N_7935,N_7419,N_7401);
xnor U7936 (N_7936,N_7241,N_7115);
nor U7937 (N_7937,N_7000,N_7338);
or U7938 (N_7938,N_7000,N_7137);
or U7939 (N_7939,N_7139,N_7002);
nand U7940 (N_7940,N_7325,N_7173);
or U7941 (N_7941,N_7359,N_7479);
nor U7942 (N_7942,N_7386,N_7182);
and U7943 (N_7943,N_7036,N_7336);
and U7944 (N_7944,N_7294,N_7355);
xnor U7945 (N_7945,N_7230,N_7157);
nor U7946 (N_7946,N_7482,N_7191);
nand U7947 (N_7947,N_7157,N_7301);
or U7948 (N_7948,N_7421,N_7449);
nand U7949 (N_7949,N_7065,N_7451);
and U7950 (N_7950,N_7288,N_7311);
or U7951 (N_7951,N_7045,N_7120);
xnor U7952 (N_7952,N_7029,N_7078);
nor U7953 (N_7953,N_7017,N_7133);
or U7954 (N_7954,N_7399,N_7313);
nor U7955 (N_7955,N_7183,N_7156);
and U7956 (N_7956,N_7381,N_7173);
nor U7957 (N_7957,N_7275,N_7145);
nand U7958 (N_7958,N_7357,N_7295);
nand U7959 (N_7959,N_7057,N_7081);
nand U7960 (N_7960,N_7057,N_7001);
and U7961 (N_7961,N_7396,N_7009);
xnor U7962 (N_7962,N_7288,N_7367);
nand U7963 (N_7963,N_7347,N_7482);
nand U7964 (N_7964,N_7120,N_7299);
xnor U7965 (N_7965,N_7063,N_7195);
and U7966 (N_7966,N_7035,N_7072);
nand U7967 (N_7967,N_7185,N_7120);
xnor U7968 (N_7968,N_7257,N_7221);
and U7969 (N_7969,N_7312,N_7081);
nand U7970 (N_7970,N_7215,N_7365);
nand U7971 (N_7971,N_7269,N_7062);
or U7972 (N_7972,N_7110,N_7324);
nor U7973 (N_7973,N_7109,N_7033);
and U7974 (N_7974,N_7434,N_7368);
or U7975 (N_7975,N_7099,N_7405);
nor U7976 (N_7976,N_7120,N_7191);
and U7977 (N_7977,N_7465,N_7437);
nand U7978 (N_7978,N_7029,N_7270);
nand U7979 (N_7979,N_7212,N_7341);
nor U7980 (N_7980,N_7293,N_7372);
and U7981 (N_7981,N_7106,N_7318);
nor U7982 (N_7982,N_7465,N_7322);
and U7983 (N_7983,N_7196,N_7250);
and U7984 (N_7984,N_7488,N_7333);
and U7985 (N_7985,N_7046,N_7081);
nand U7986 (N_7986,N_7202,N_7231);
xor U7987 (N_7987,N_7140,N_7059);
and U7988 (N_7988,N_7388,N_7007);
xnor U7989 (N_7989,N_7456,N_7104);
nand U7990 (N_7990,N_7444,N_7221);
and U7991 (N_7991,N_7344,N_7025);
nand U7992 (N_7992,N_7037,N_7189);
and U7993 (N_7993,N_7178,N_7347);
nand U7994 (N_7994,N_7157,N_7268);
or U7995 (N_7995,N_7071,N_7146);
and U7996 (N_7996,N_7493,N_7240);
nand U7997 (N_7997,N_7280,N_7431);
and U7998 (N_7998,N_7109,N_7241);
or U7999 (N_7999,N_7088,N_7424);
nand U8000 (N_8000,N_7581,N_7864);
and U8001 (N_8001,N_7522,N_7523);
or U8002 (N_8002,N_7958,N_7559);
nand U8003 (N_8003,N_7704,N_7698);
nand U8004 (N_8004,N_7915,N_7974);
nand U8005 (N_8005,N_7848,N_7754);
and U8006 (N_8006,N_7727,N_7562);
and U8007 (N_8007,N_7926,N_7549);
nor U8008 (N_8008,N_7905,N_7572);
xnor U8009 (N_8009,N_7855,N_7668);
nor U8010 (N_8010,N_7595,N_7837);
nor U8011 (N_8011,N_7953,N_7814);
or U8012 (N_8012,N_7988,N_7710);
nand U8013 (N_8013,N_7952,N_7567);
nand U8014 (N_8014,N_7665,N_7806);
xor U8015 (N_8015,N_7598,N_7870);
or U8016 (N_8016,N_7502,N_7714);
nor U8017 (N_8017,N_7633,N_7943);
or U8018 (N_8018,N_7865,N_7740);
or U8019 (N_8019,N_7722,N_7604);
xnor U8020 (N_8020,N_7690,N_7520);
nand U8021 (N_8021,N_7741,N_7677);
or U8022 (N_8022,N_7532,N_7718);
nor U8023 (N_8023,N_7916,N_7627);
xnor U8024 (N_8024,N_7928,N_7687);
xnor U8025 (N_8025,N_7575,N_7664);
nand U8026 (N_8026,N_7607,N_7553);
and U8027 (N_8027,N_7745,N_7695);
nor U8028 (N_8028,N_7775,N_7582);
xnor U8029 (N_8029,N_7858,N_7666);
nor U8030 (N_8030,N_7646,N_7630);
or U8031 (N_8031,N_7993,N_7786);
xor U8032 (N_8032,N_7977,N_7501);
nand U8033 (N_8033,N_7892,N_7798);
or U8034 (N_8034,N_7500,N_7693);
nand U8035 (N_8035,N_7964,N_7810);
and U8036 (N_8036,N_7876,N_7660);
nor U8037 (N_8037,N_7817,N_7623);
nand U8038 (N_8038,N_7579,N_7732);
or U8039 (N_8039,N_7818,N_7896);
or U8040 (N_8040,N_7984,N_7857);
or U8041 (N_8041,N_7976,N_7600);
nor U8042 (N_8042,N_7563,N_7746);
nor U8043 (N_8043,N_7853,N_7967);
or U8044 (N_8044,N_7531,N_7962);
or U8045 (N_8045,N_7628,N_7925);
nor U8046 (N_8046,N_7783,N_7849);
and U8047 (N_8047,N_7622,N_7577);
nor U8048 (N_8048,N_7791,N_7621);
nand U8049 (N_8049,N_7702,N_7803);
nand U8050 (N_8050,N_7932,N_7947);
xor U8051 (N_8051,N_7635,N_7655);
or U8052 (N_8052,N_7963,N_7766);
and U8053 (N_8053,N_7835,N_7919);
xor U8054 (N_8054,N_7524,N_7752);
xor U8055 (N_8055,N_7744,N_7724);
or U8056 (N_8056,N_7975,N_7779);
xnor U8057 (N_8057,N_7869,N_7739);
and U8058 (N_8058,N_7936,N_7957);
and U8059 (N_8059,N_7878,N_7920);
or U8060 (N_8060,N_7822,N_7797);
nor U8061 (N_8061,N_7640,N_7790);
xnor U8062 (N_8062,N_7770,N_7840);
or U8063 (N_8063,N_7662,N_7641);
or U8064 (N_8064,N_7914,N_7990);
xor U8065 (N_8065,N_7676,N_7513);
nand U8066 (N_8066,N_7960,N_7801);
and U8067 (N_8067,N_7591,N_7830);
xor U8068 (N_8068,N_7565,N_7707);
or U8069 (N_8069,N_7829,N_7514);
nor U8070 (N_8070,N_7902,N_7948);
or U8071 (N_8071,N_7999,N_7648);
or U8072 (N_8072,N_7706,N_7900);
or U8073 (N_8073,N_7804,N_7750);
xnor U8074 (N_8074,N_7881,N_7877);
nand U8075 (N_8075,N_7542,N_7844);
or U8076 (N_8076,N_7923,N_7545);
nand U8077 (N_8077,N_7527,N_7561);
and U8078 (N_8078,N_7645,N_7515);
nor U8079 (N_8079,N_7777,N_7736);
and U8080 (N_8080,N_7670,N_7649);
or U8081 (N_8081,N_7899,N_7634);
or U8082 (N_8082,N_7715,N_7654);
xor U8083 (N_8083,N_7726,N_7592);
nor U8084 (N_8084,N_7965,N_7731);
or U8085 (N_8085,N_7626,N_7541);
nor U8086 (N_8086,N_7728,N_7884);
nor U8087 (N_8087,N_7644,N_7653);
and U8088 (N_8088,N_7788,N_7705);
xnor U8089 (N_8089,N_7929,N_7889);
xor U8090 (N_8090,N_7535,N_7951);
and U8091 (N_8091,N_7934,N_7652);
or U8092 (N_8092,N_7983,N_7605);
and U8093 (N_8093,N_7940,N_7518);
nor U8094 (N_8094,N_7658,N_7753);
nand U8095 (N_8095,N_7872,N_7700);
and U8096 (N_8096,N_7986,N_7898);
or U8097 (N_8097,N_7989,N_7566);
nor U8098 (N_8098,N_7800,N_7911);
nor U8099 (N_8099,N_7765,N_7610);
and U8100 (N_8100,N_7956,N_7525);
nor U8101 (N_8101,N_7908,N_7743);
nor U8102 (N_8102,N_7890,N_7901);
and U8103 (N_8103,N_7576,N_7764);
nor U8104 (N_8104,N_7927,N_7816);
nand U8105 (N_8105,N_7552,N_7650);
nand U8106 (N_8106,N_7767,N_7792);
nand U8107 (N_8107,N_7504,N_7815);
nor U8108 (N_8108,N_7834,N_7760);
nand U8109 (N_8109,N_7587,N_7906);
or U8110 (N_8110,N_7533,N_7509);
nand U8111 (N_8111,N_7987,N_7867);
xnor U8112 (N_8112,N_7820,N_7992);
nor U8113 (N_8113,N_7546,N_7895);
or U8114 (N_8114,N_7709,N_7723);
and U8115 (N_8115,N_7510,N_7680);
nand U8116 (N_8116,N_7871,N_7874);
nor U8117 (N_8117,N_7588,N_7856);
nor U8118 (N_8118,N_7597,N_7773);
nor U8119 (N_8119,N_7508,N_7560);
or U8120 (N_8120,N_7769,N_7969);
nor U8121 (N_8121,N_7671,N_7802);
nor U8122 (N_8122,N_7826,N_7781);
or U8123 (N_8123,N_7517,N_7937);
or U8124 (N_8124,N_7894,N_7618);
nand U8125 (N_8125,N_7910,N_7893);
xor U8126 (N_8126,N_7845,N_7782);
or U8127 (N_8127,N_7512,N_7918);
and U8128 (N_8128,N_7696,N_7719);
nand U8129 (N_8129,N_7970,N_7772);
or U8130 (N_8130,N_7946,N_7912);
nand U8131 (N_8131,N_7536,N_7735);
nand U8132 (N_8132,N_7636,N_7589);
nor U8133 (N_8133,N_7995,N_7538);
nor U8134 (N_8134,N_7998,N_7778);
and U8135 (N_8135,N_7585,N_7882);
and U8136 (N_8136,N_7679,N_7613);
nand U8137 (N_8137,N_7742,N_7991);
or U8138 (N_8138,N_7907,N_7812);
nor U8139 (N_8139,N_7643,N_7609);
nand U8140 (N_8140,N_7819,N_7836);
or U8141 (N_8141,N_7580,N_7843);
or U8142 (N_8142,N_7748,N_7590);
and U8143 (N_8143,N_7860,N_7530);
or U8144 (N_8144,N_7578,N_7716);
xor U8145 (N_8145,N_7651,N_7933);
nand U8146 (N_8146,N_7921,N_7558);
or U8147 (N_8147,N_7528,N_7981);
and U8148 (N_8148,N_7959,N_7673);
xor U8149 (N_8149,N_7663,N_7596);
or U8150 (N_8150,N_7616,N_7697);
or U8151 (N_8151,N_7608,N_7729);
nor U8152 (N_8152,N_7675,N_7885);
or U8153 (N_8153,N_7543,N_7771);
and U8154 (N_8154,N_7672,N_7941);
and U8155 (N_8155,N_7968,N_7584);
nand U8156 (N_8156,N_7712,N_7838);
xnor U8157 (N_8157,N_7711,N_7511);
nand U8158 (N_8158,N_7661,N_7738);
nor U8159 (N_8159,N_7540,N_7720);
nor U8160 (N_8160,N_7821,N_7808);
nor U8161 (N_8161,N_7824,N_7611);
and U8162 (N_8162,N_7931,N_7863);
nor U8163 (N_8163,N_7620,N_7945);
xor U8164 (N_8164,N_7994,N_7631);
xnor U8165 (N_8165,N_7701,N_7691);
or U8166 (N_8166,N_7625,N_7883);
nand U8167 (N_8167,N_7717,N_7859);
and U8168 (N_8168,N_7903,N_7887);
nand U8169 (N_8169,N_7868,N_7725);
nand U8170 (N_8170,N_7564,N_7713);
and U8171 (N_8171,N_7516,N_7688);
or U8172 (N_8172,N_7684,N_7548);
or U8173 (N_8173,N_7573,N_7593);
nor U8174 (N_8174,N_7678,N_7694);
nand U8175 (N_8175,N_7569,N_7796);
and U8176 (N_8176,N_7904,N_7544);
or U8177 (N_8177,N_7852,N_7763);
nor U8178 (N_8178,N_7922,N_7550);
nor U8179 (N_8179,N_7985,N_7632);
nand U8180 (N_8180,N_7734,N_7997);
and U8181 (N_8181,N_7537,N_7539);
or U8182 (N_8182,N_7521,N_7813);
nand U8183 (N_8183,N_7789,N_7833);
xnor U8184 (N_8184,N_7776,N_7954);
nand U8185 (N_8185,N_7659,N_7642);
or U8186 (N_8186,N_7944,N_7917);
nand U8187 (N_8187,N_7950,N_7973);
nor U8188 (N_8188,N_7529,N_7924);
nand U8189 (N_8189,N_7823,N_7612);
xor U8190 (N_8190,N_7554,N_7913);
nor U8191 (N_8191,N_7749,N_7755);
nor U8192 (N_8192,N_7886,N_7614);
and U8193 (N_8193,N_7861,N_7825);
nand U8194 (N_8194,N_7703,N_7692);
nand U8195 (N_8195,N_7751,N_7811);
nor U8196 (N_8196,N_7656,N_7557);
xnor U8197 (N_8197,N_7759,N_7873);
and U8198 (N_8198,N_7846,N_7862);
nand U8199 (N_8199,N_7681,N_7555);
nor U8200 (N_8200,N_7851,N_7888);
or U8201 (N_8201,N_7526,N_7762);
nor U8202 (N_8202,N_7938,N_7571);
or U8203 (N_8203,N_7606,N_7619);
or U8204 (N_8204,N_7949,N_7657);
nand U8205 (N_8205,N_7850,N_7730);
nor U8206 (N_8206,N_7784,N_7547);
and U8207 (N_8207,N_7982,N_7978);
xnor U8208 (N_8208,N_7756,N_7787);
and U8209 (N_8209,N_7629,N_7667);
nand U8210 (N_8210,N_7961,N_7624);
nor U8211 (N_8211,N_7795,N_7601);
or U8212 (N_8212,N_7768,N_7682);
nand U8213 (N_8213,N_7568,N_7930);
and U8214 (N_8214,N_7841,N_7979);
and U8215 (N_8215,N_7747,N_7505);
nand U8216 (N_8216,N_7794,N_7879);
or U8217 (N_8217,N_7737,N_7556);
nand U8218 (N_8218,N_7831,N_7880);
and U8219 (N_8219,N_7689,N_7866);
nand U8220 (N_8220,N_7971,N_7551);
nand U8221 (N_8221,N_7955,N_7503);
nor U8222 (N_8222,N_7854,N_7980);
or U8223 (N_8223,N_7839,N_7875);
xor U8224 (N_8224,N_7807,N_7583);
xor U8225 (N_8225,N_7785,N_7647);
or U8226 (N_8226,N_7683,N_7721);
nand U8227 (N_8227,N_7996,N_7793);
nor U8228 (N_8228,N_7674,N_7897);
nand U8229 (N_8229,N_7699,N_7669);
nand U8230 (N_8230,N_7708,N_7832);
and U8231 (N_8231,N_7594,N_7780);
and U8232 (N_8232,N_7686,N_7939);
nor U8233 (N_8233,N_7615,N_7966);
nor U8234 (N_8234,N_7617,N_7847);
xnor U8235 (N_8235,N_7828,N_7506);
xor U8236 (N_8236,N_7935,N_7972);
nand U8237 (N_8237,N_7842,N_7638);
or U8238 (N_8238,N_7799,N_7519);
nand U8239 (N_8239,N_7809,N_7827);
or U8240 (N_8240,N_7574,N_7758);
xnor U8241 (N_8241,N_7757,N_7602);
xor U8242 (N_8242,N_7637,N_7586);
and U8243 (N_8243,N_7909,N_7599);
nand U8244 (N_8244,N_7942,N_7603);
xor U8245 (N_8245,N_7685,N_7507);
nand U8246 (N_8246,N_7534,N_7570);
nand U8247 (N_8247,N_7761,N_7639);
nand U8248 (N_8248,N_7891,N_7733);
or U8249 (N_8249,N_7805,N_7774);
nor U8250 (N_8250,N_7783,N_7691);
nand U8251 (N_8251,N_7903,N_7602);
nand U8252 (N_8252,N_7927,N_7618);
nor U8253 (N_8253,N_7746,N_7884);
and U8254 (N_8254,N_7853,N_7607);
nor U8255 (N_8255,N_7574,N_7891);
nor U8256 (N_8256,N_7821,N_7560);
nand U8257 (N_8257,N_7664,N_7987);
nand U8258 (N_8258,N_7576,N_7743);
and U8259 (N_8259,N_7704,N_7694);
xnor U8260 (N_8260,N_7931,N_7954);
or U8261 (N_8261,N_7713,N_7682);
nand U8262 (N_8262,N_7886,N_7597);
and U8263 (N_8263,N_7605,N_7681);
or U8264 (N_8264,N_7723,N_7649);
nand U8265 (N_8265,N_7801,N_7698);
nand U8266 (N_8266,N_7798,N_7914);
or U8267 (N_8267,N_7975,N_7946);
or U8268 (N_8268,N_7589,N_7567);
nand U8269 (N_8269,N_7954,N_7956);
or U8270 (N_8270,N_7718,N_7581);
or U8271 (N_8271,N_7597,N_7803);
and U8272 (N_8272,N_7576,N_7607);
or U8273 (N_8273,N_7989,N_7696);
nand U8274 (N_8274,N_7514,N_7602);
nand U8275 (N_8275,N_7946,N_7799);
nor U8276 (N_8276,N_7805,N_7529);
nand U8277 (N_8277,N_7885,N_7868);
xor U8278 (N_8278,N_7689,N_7554);
nor U8279 (N_8279,N_7902,N_7936);
nand U8280 (N_8280,N_7660,N_7561);
nand U8281 (N_8281,N_7898,N_7706);
nor U8282 (N_8282,N_7757,N_7611);
and U8283 (N_8283,N_7952,N_7629);
and U8284 (N_8284,N_7578,N_7537);
nor U8285 (N_8285,N_7758,N_7837);
and U8286 (N_8286,N_7855,N_7978);
or U8287 (N_8287,N_7795,N_7513);
nor U8288 (N_8288,N_7873,N_7920);
nand U8289 (N_8289,N_7921,N_7630);
and U8290 (N_8290,N_7719,N_7978);
or U8291 (N_8291,N_7846,N_7832);
xnor U8292 (N_8292,N_7511,N_7523);
nor U8293 (N_8293,N_7563,N_7884);
and U8294 (N_8294,N_7732,N_7568);
or U8295 (N_8295,N_7915,N_7630);
nor U8296 (N_8296,N_7720,N_7668);
nor U8297 (N_8297,N_7733,N_7554);
nand U8298 (N_8298,N_7745,N_7703);
nand U8299 (N_8299,N_7614,N_7918);
xnor U8300 (N_8300,N_7905,N_7894);
or U8301 (N_8301,N_7948,N_7763);
or U8302 (N_8302,N_7973,N_7857);
nand U8303 (N_8303,N_7917,N_7784);
nand U8304 (N_8304,N_7831,N_7604);
xnor U8305 (N_8305,N_7692,N_7996);
nand U8306 (N_8306,N_7748,N_7670);
nor U8307 (N_8307,N_7720,N_7744);
nor U8308 (N_8308,N_7831,N_7853);
nand U8309 (N_8309,N_7535,N_7762);
and U8310 (N_8310,N_7591,N_7839);
xnor U8311 (N_8311,N_7520,N_7724);
xnor U8312 (N_8312,N_7816,N_7579);
or U8313 (N_8313,N_7648,N_7914);
xnor U8314 (N_8314,N_7899,N_7645);
nor U8315 (N_8315,N_7853,N_7617);
or U8316 (N_8316,N_7711,N_7831);
or U8317 (N_8317,N_7507,N_7694);
nand U8318 (N_8318,N_7922,N_7688);
or U8319 (N_8319,N_7532,N_7617);
and U8320 (N_8320,N_7676,N_7873);
xor U8321 (N_8321,N_7973,N_7853);
xor U8322 (N_8322,N_7814,N_7519);
xnor U8323 (N_8323,N_7894,N_7763);
and U8324 (N_8324,N_7891,N_7916);
or U8325 (N_8325,N_7787,N_7595);
and U8326 (N_8326,N_7646,N_7726);
or U8327 (N_8327,N_7720,N_7872);
nor U8328 (N_8328,N_7828,N_7884);
nor U8329 (N_8329,N_7941,N_7777);
nor U8330 (N_8330,N_7961,N_7998);
xnor U8331 (N_8331,N_7679,N_7835);
or U8332 (N_8332,N_7851,N_7913);
and U8333 (N_8333,N_7872,N_7525);
nor U8334 (N_8334,N_7957,N_7831);
nand U8335 (N_8335,N_7606,N_7640);
nor U8336 (N_8336,N_7748,N_7725);
xnor U8337 (N_8337,N_7617,N_7552);
and U8338 (N_8338,N_7875,N_7735);
and U8339 (N_8339,N_7769,N_7794);
nor U8340 (N_8340,N_7845,N_7921);
or U8341 (N_8341,N_7850,N_7999);
nand U8342 (N_8342,N_7703,N_7922);
xnor U8343 (N_8343,N_7930,N_7536);
or U8344 (N_8344,N_7897,N_7597);
or U8345 (N_8345,N_7675,N_7898);
nor U8346 (N_8346,N_7998,N_7569);
nor U8347 (N_8347,N_7674,N_7821);
and U8348 (N_8348,N_7906,N_7778);
nand U8349 (N_8349,N_7853,N_7923);
nand U8350 (N_8350,N_7554,N_7954);
and U8351 (N_8351,N_7808,N_7624);
nand U8352 (N_8352,N_7813,N_7583);
nand U8353 (N_8353,N_7755,N_7702);
xnor U8354 (N_8354,N_7647,N_7883);
nand U8355 (N_8355,N_7602,N_7744);
or U8356 (N_8356,N_7804,N_7504);
and U8357 (N_8357,N_7739,N_7908);
or U8358 (N_8358,N_7702,N_7757);
nand U8359 (N_8359,N_7680,N_7885);
nor U8360 (N_8360,N_7888,N_7987);
and U8361 (N_8361,N_7844,N_7580);
nand U8362 (N_8362,N_7506,N_7972);
and U8363 (N_8363,N_7717,N_7624);
xnor U8364 (N_8364,N_7711,N_7774);
nand U8365 (N_8365,N_7792,N_7556);
and U8366 (N_8366,N_7808,N_7943);
and U8367 (N_8367,N_7700,N_7579);
and U8368 (N_8368,N_7984,N_7800);
xnor U8369 (N_8369,N_7798,N_7620);
nand U8370 (N_8370,N_7954,N_7960);
and U8371 (N_8371,N_7696,N_7632);
nand U8372 (N_8372,N_7830,N_7700);
or U8373 (N_8373,N_7669,N_7719);
or U8374 (N_8374,N_7664,N_7512);
nor U8375 (N_8375,N_7740,N_7655);
nand U8376 (N_8376,N_7513,N_7697);
or U8377 (N_8377,N_7511,N_7996);
nand U8378 (N_8378,N_7524,N_7643);
or U8379 (N_8379,N_7608,N_7534);
and U8380 (N_8380,N_7972,N_7554);
nor U8381 (N_8381,N_7787,N_7727);
or U8382 (N_8382,N_7741,N_7854);
xnor U8383 (N_8383,N_7739,N_7890);
nand U8384 (N_8384,N_7809,N_7585);
nor U8385 (N_8385,N_7587,N_7840);
and U8386 (N_8386,N_7830,N_7733);
nand U8387 (N_8387,N_7575,N_7573);
and U8388 (N_8388,N_7937,N_7816);
nand U8389 (N_8389,N_7558,N_7851);
nand U8390 (N_8390,N_7623,N_7896);
nand U8391 (N_8391,N_7848,N_7677);
or U8392 (N_8392,N_7676,N_7919);
or U8393 (N_8393,N_7839,N_7555);
nand U8394 (N_8394,N_7992,N_7989);
or U8395 (N_8395,N_7845,N_7586);
or U8396 (N_8396,N_7833,N_7535);
nor U8397 (N_8397,N_7559,N_7571);
nand U8398 (N_8398,N_7870,N_7604);
and U8399 (N_8399,N_7884,N_7705);
or U8400 (N_8400,N_7952,N_7687);
or U8401 (N_8401,N_7931,N_7586);
xor U8402 (N_8402,N_7779,N_7829);
and U8403 (N_8403,N_7681,N_7686);
nand U8404 (N_8404,N_7780,N_7721);
nand U8405 (N_8405,N_7921,N_7958);
nor U8406 (N_8406,N_7943,N_7792);
nor U8407 (N_8407,N_7743,N_7769);
nand U8408 (N_8408,N_7622,N_7991);
xor U8409 (N_8409,N_7778,N_7773);
and U8410 (N_8410,N_7813,N_7959);
nor U8411 (N_8411,N_7562,N_7745);
nand U8412 (N_8412,N_7735,N_7758);
nand U8413 (N_8413,N_7508,N_7904);
and U8414 (N_8414,N_7907,N_7688);
nand U8415 (N_8415,N_7611,N_7500);
nor U8416 (N_8416,N_7582,N_7923);
and U8417 (N_8417,N_7834,N_7856);
and U8418 (N_8418,N_7586,N_7973);
nor U8419 (N_8419,N_7852,N_7902);
and U8420 (N_8420,N_7513,N_7698);
nor U8421 (N_8421,N_7523,N_7662);
and U8422 (N_8422,N_7950,N_7607);
nor U8423 (N_8423,N_7737,N_7667);
nor U8424 (N_8424,N_7825,N_7902);
and U8425 (N_8425,N_7915,N_7759);
nand U8426 (N_8426,N_7736,N_7602);
nand U8427 (N_8427,N_7505,N_7525);
nand U8428 (N_8428,N_7798,N_7941);
and U8429 (N_8429,N_7958,N_7950);
and U8430 (N_8430,N_7626,N_7946);
or U8431 (N_8431,N_7618,N_7906);
nor U8432 (N_8432,N_7751,N_7800);
and U8433 (N_8433,N_7866,N_7531);
xor U8434 (N_8434,N_7589,N_7910);
nand U8435 (N_8435,N_7850,N_7907);
and U8436 (N_8436,N_7670,N_7709);
and U8437 (N_8437,N_7809,N_7837);
xnor U8438 (N_8438,N_7800,N_7899);
and U8439 (N_8439,N_7986,N_7912);
nand U8440 (N_8440,N_7896,N_7825);
nor U8441 (N_8441,N_7910,N_7565);
xor U8442 (N_8442,N_7549,N_7930);
or U8443 (N_8443,N_7709,N_7645);
nand U8444 (N_8444,N_7810,N_7892);
and U8445 (N_8445,N_7986,N_7556);
nand U8446 (N_8446,N_7985,N_7818);
nor U8447 (N_8447,N_7720,N_7984);
nand U8448 (N_8448,N_7967,N_7929);
and U8449 (N_8449,N_7866,N_7623);
or U8450 (N_8450,N_7797,N_7978);
or U8451 (N_8451,N_7875,N_7963);
nor U8452 (N_8452,N_7517,N_7660);
nor U8453 (N_8453,N_7873,N_7610);
and U8454 (N_8454,N_7566,N_7939);
or U8455 (N_8455,N_7584,N_7867);
xnor U8456 (N_8456,N_7817,N_7737);
nand U8457 (N_8457,N_7597,N_7810);
and U8458 (N_8458,N_7910,N_7632);
or U8459 (N_8459,N_7758,N_7965);
and U8460 (N_8460,N_7908,N_7902);
or U8461 (N_8461,N_7598,N_7690);
and U8462 (N_8462,N_7616,N_7860);
nor U8463 (N_8463,N_7754,N_7830);
nor U8464 (N_8464,N_7787,N_7826);
nor U8465 (N_8465,N_7823,N_7731);
nand U8466 (N_8466,N_7965,N_7547);
nor U8467 (N_8467,N_7718,N_7987);
and U8468 (N_8468,N_7825,N_7640);
nand U8469 (N_8469,N_7932,N_7548);
nand U8470 (N_8470,N_7986,N_7758);
or U8471 (N_8471,N_7867,N_7828);
xor U8472 (N_8472,N_7749,N_7679);
nand U8473 (N_8473,N_7898,N_7935);
and U8474 (N_8474,N_7635,N_7564);
nor U8475 (N_8475,N_7726,N_7811);
nand U8476 (N_8476,N_7518,N_7767);
or U8477 (N_8477,N_7775,N_7691);
nor U8478 (N_8478,N_7685,N_7857);
and U8479 (N_8479,N_7914,N_7986);
nor U8480 (N_8480,N_7526,N_7733);
nand U8481 (N_8481,N_7618,N_7834);
and U8482 (N_8482,N_7972,N_7749);
or U8483 (N_8483,N_7854,N_7845);
nand U8484 (N_8484,N_7918,N_7866);
nor U8485 (N_8485,N_7912,N_7611);
nor U8486 (N_8486,N_7730,N_7764);
nor U8487 (N_8487,N_7617,N_7800);
or U8488 (N_8488,N_7980,N_7976);
and U8489 (N_8489,N_7504,N_7794);
or U8490 (N_8490,N_7985,N_7643);
xor U8491 (N_8491,N_7620,N_7745);
xor U8492 (N_8492,N_7859,N_7794);
xor U8493 (N_8493,N_7846,N_7576);
xor U8494 (N_8494,N_7975,N_7835);
nor U8495 (N_8495,N_7659,N_7681);
nor U8496 (N_8496,N_7777,N_7649);
and U8497 (N_8497,N_7941,N_7943);
nand U8498 (N_8498,N_7846,N_7724);
xor U8499 (N_8499,N_7631,N_7521);
or U8500 (N_8500,N_8411,N_8010);
nor U8501 (N_8501,N_8427,N_8110);
and U8502 (N_8502,N_8087,N_8280);
and U8503 (N_8503,N_8467,N_8476);
and U8504 (N_8504,N_8256,N_8288);
or U8505 (N_8505,N_8132,N_8369);
or U8506 (N_8506,N_8305,N_8154);
nor U8507 (N_8507,N_8205,N_8005);
nand U8508 (N_8508,N_8294,N_8174);
nor U8509 (N_8509,N_8223,N_8416);
nor U8510 (N_8510,N_8080,N_8171);
xnor U8511 (N_8511,N_8477,N_8108);
and U8512 (N_8512,N_8357,N_8035);
and U8513 (N_8513,N_8073,N_8295);
or U8514 (N_8514,N_8189,N_8095);
nand U8515 (N_8515,N_8359,N_8198);
nor U8516 (N_8516,N_8157,N_8133);
nand U8517 (N_8517,N_8315,N_8193);
or U8518 (N_8518,N_8128,N_8203);
nand U8519 (N_8519,N_8377,N_8019);
and U8520 (N_8520,N_8362,N_8141);
nor U8521 (N_8521,N_8286,N_8471);
nand U8522 (N_8522,N_8025,N_8221);
or U8523 (N_8523,N_8121,N_8227);
xnor U8524 (N_8524,N_8301,N_8097);
nor U8525 (N_8525,N_8155,N_8066);
or U8526 (N_8526,N_8351,N_8045);
nand U8527 (N_8527,N_8389,N_8451);
nor U8528 (N_8528,N_8465,N_8468);
or U8529 (N_8529,N_8074,N_8418);
nor U8530 (N_8530,N_8163,N_8378);
nor U8531 (N_8531,N_8214,N_8493);
or U8532 (N_8532,N_8094,N_8494);
nor U8533 (N_8533,N_8404,N_8370);
nor U8534 (N_8534,N_8313,N_8423);
or U8535 (N_8535,N_8446,N_8492);
and U8536 (N_8536,N_8440,N_8491);
nor U8537 (N_8537,N_8081,N_8020);
nor U8538 (N_8538,N_8324,N_8405);
nor U8539 (N_8539,N_8173,N_8320);
or U8540 (N_8540,N_8103,N_8085);
xor U8541 (N_8541,N_8233,N_8188);
nand U8542 (N_8542,N_8147,N_8015);
nor U8543 (N_8543,N_8435,N_8044);
or U8544 (N_8544,N_8258,N_8250);
xor U8545 (N_8545,N_8031,N_8486);
and U8546 (N_8546,N_8199,N_8244);
or U8547 (N_8547,N_8116,N_8177);
and U8548 (N_8548,N_8145,N_8499);
or U8549 (N_8549,N_8225,N_8292);
or U8550 (N_8550,N_8026,N_8265);
or U8551 (N_8551,N_8410,N_8114);
or U8552 (N_8552,N_8488,N_8356);
nor U8553 (N_8553,N_8249,N_8375);
and U8554 (N_8554,N_8234,N_8284);
and U8555 (N_8555,N_8072,N_8376);
xnor U8556 (N_8556,N_8119,N_8136);
nand U8557 (N_8557,N_8075,N_8212);
and U8558 (N_8558,N_8328,N_8152);
and U8559 (N_8559,N_8325,N_8253);
and U8560 (N_8560,N_8187,N_8299);
and U8561 (N_8561,N_8176,N_8064);
nor U8562 (N_8562,N_8402,N_8118);
nand U8563 (N_8563,N_8135,N_8282);
or U8564 (N_8564,N_8470,N_8243);
and U8565 (N_8565,N_8083,N_8002);
nand U8566 (N_8566,N_8323,N_8086);
or U8567 (N_8567,N_8478,N_8429);
and U8568 (N_8568,N_8395,N_8390);
nor U8569 (N_8569,N_8159,N_8428);
or U8570 (N_8570,N_8436,N_8140);
or U8571 (N_8571,N_8424,N_8481);
and U8572 (N_8572,N_8007,N_8175);
or U8573 (N_8573,N_8455,N_8460);
or U8574 (N_8574,N_8151,N_8146);
nand U8575 (N_8575,N_8371,N_8077);
nand U8576 (N_8576,N_8222,N_8268);
or U8577 (N_8577,N_8398,N_8247);
or U8578 (N_8578,N_8421,N_8303);
or U8579 (N_8579,N_8049,N_8437);
and U8580 (N_8580,N_8215,N_8425);
nand U8581 (N_8581,N_8270,N_8207);
xnor U8582 (N_8582,N_8041,N_8358);
nor U8583 (N_8583,N_8373,N_8281);
or U8584 (N_8584,N_8084,N_8403);
nand U8585 (N_8585,N_8091,N_8224);
and U8586 (N_8586,N_8172,N_8480);
and U8587 (N_8587,N_8329,N_8442);
and U8588 (N_8588,N_8150,N_8192);
and U8589 (N_8589,N_8431,N_8191);
and U8590 (N_8590,N_8257,N_8479);
nor U8591 (N_8591,N_8238,N_8381);
nand U8592 (N_8592,N_8104,N_8184);
and U8593 (N_8593,N_8003,N_8266);
nand U8594 (N_8594,N_8498,N_8018);
or U8595 (N_8595,N_8346,N_8228);
and U8596 (N_8596,N_8453,N_8209);
or U8597 (N_8597,N_8400,N_8229);
nor U8598 (N_8598,N_8165,N_8012);
and U8599 (N_8599,N_8076,N_8226);
nand U8600 (N_8600,N_8106,N_8495);
nor U8601 (N_8601,N_8466,N_8269);
and U8602 (N_8602,N_8245,N_8113);
or U8603 (N_8603,N_8053,N_8261);
and U8604 (N_8604,N_8321,N_8319);
and U8605 (N_8605,N_8100,N_8006);
and U8606 (N_8606,N_8298,N_8332);
nor U8607 (N_8607,N_8186,N_8485);
xnor U8608 (N_8608,N_8160,N_8289);
and U8609 (N_8609,N_8040,N_8211);
xor U8610 (N_8610,N_8343,N_8052);
nand U8611 (N_8611,N_8341,N_8048);
and U8612 (N_8612,N_8058,N_8069);
xor U8613 (N_8613,N_8120,N_8099);
and U8614 (N_8614,N_8017,N_8237);
nand U8615 (N_8615,N_8393,N_8038);
nor U8616 (N_8616,N_8456,N_8216);
nor U8617 (N_8617,N_8070,N_8318);
nor U8618 (N_8618,N_8008,N_8326);
nor U8619 (N_8619,N_8050,N_8392);
nor U8620 (N_8620,N_8422,N_8056);
nor U8621 (N_8621,N_8409,N_8461);
and U8622 (N_8622,N_8380,N_8408);
and U8623 (N_8623,N_8415,N_8065);
nor U8624 (N_8624,N_8349,N_8401);
nand U8625 (N_8625,N_8129,N_8430);
and U8626 (N_8626,N_8279,N_8014);
and U8627 (N_8627,N_8230,N_8296);
and U8628 (N_8628,N_8235,N_8213);
xnor U8629 (N_8629,N_8454,N_8028);
or U8630 (N_8630,N_8021,N_8051);
nand U8631 (N_8631,N_8219,N_8004);
and U8632 (N_8632,N_8178,N_8383);
and U8633 (N_8633,N_8490,N_8023);
or U8634 (N_8634,N_8310,N_8208);
or U8635 (N_8635,N_8354,N_8122);
nand U8636 (N_8636,N_8361,N_8475);
nor U8637 (N_8637,N_8293,N_8267);
or U8638 (N_8638,N_8197,N_8316);
and U8639 (N_8639,N_8090,N_8201);
xor U8640 (N_8640,N_8300,N_8054);
nor U8641 (N_8641,N_8444,N_8032);
or U8642 (N_8642,N_8312,N_8259);
nor U8643 (N_8643,N_8275,N_8263);
and U8644 (N_8644,N_8042,N_8413);
nor U8645 (N_8645,N_8452,N_8030);
or U8646 (N_8646,N_8384,N_8331);
and U8647 (N_8647,N_8092,N_8079);
or U8648 (N_8648,N_8335,N_8483);
nor U8649 (N_8649,N_8196,N_8181);
nand U8650 (N_8650,N_8443,N_8387);
xnor U8651 (N_8651,N_8338,N_8170);
or U8652 (N_8652,N_8285,N_8182);
xnor U8653 (N_8653,N_8134,N_8434);
nand U8654 (N_8654,N_8127,N_8399);
nor U8655 (N_8655,N_8412,N_8448);
xor U8656 (N_8656,N_8333,N_8102);
or U8657 (N_8657,N_8304,N_8447);
nand U8658 (N_8658,N_8123,N_8394);
and U8659 (N_8659,N_8462,N_8089);
nor U8660 (N_8660,N_8334,N_8126);
nor U8661 (N_8661,N_8016,N_8449);
and U8662 (N_8662,N_8439,N_8445);
nor U8663 (N_8663,N_8314,N_8148);
nor U8664 (N_8664,N_8469,N_8397);
xnor U8665 (N_8665,N_8463,N_8242);
xnor U8666 (N_8666,N_8464,N_8330);
or U8667 (N_8667,N_8363,N_8240);
nor U8668 (N_8668,N_8153,N_8364);
or U8669 (N_8669,N_8098,N_8185);
and U8670 (N_8670,N_8396,N_8027);
or U8671 (N_8671,N_8302,N_8391);
or U8672 (N_8672,N_8450,N_8009);
nand U8673 (N_8673,N_8039,N_8047);
or U8674 (N_8674,N_8386,N_8220);
and U8675 (N_8675,N_8183,N_8365);
nand U8676 (N_8676,N_8034,N_8179);
nor U8677 (N_8677,N_8327,N_8071);
nor U8678 (N_8678,N_8271,N_8291);
and U8679 (N_8679,N_8414,N_8000);
and U8680 (N_8680,N_8082,N_8441);
nand U8681 (N_8681,N_8496,N_8372);
nand U8682 (N_8682,N_8057,N_8117);
and U8683 (N_8683,N_8037,N_8283);
nor U8684 (N_8684,N_8149,N_8278);
nor U8685 (N_8685,N_8060,N_8360);
and U8686 (N_8686,N_8489,N_8474);
nor U8687 (N_8687,N_8317,N_8180);
nand U8688 (N_8688,N_8239,N_8385);
nand U8689 (N_8689,N_8206,N_8264);
nor U8690 (N_8690,N_8236,N_8011);
and U8691 (N_8691,N_8407,N_8347);
xor U8692 (N_8692,N_8043,N_8307);
or U8693 (N_8693,N_8033,N_8022);
xnor U8694 (N_8694,N_8482,N_8487);
xnor U8695 (N_8695,N_8130,N_8204);
nor U8696 (N_8696,N_8210,N_8139);
or U8697 (N_8697,N_8344,N_8067);
or U8698 (N_8698,N_8366,N_8277);
or U8699 (N_8699,N_8059,N_8459);
xor U8700 (N_8700,N_8231,N_8190);
nor U8701 (N_8701,N_8308,N_8194);
and U8702 (N_8702,N_8306,N_8156);
and U8703 (N_8703,N_8339,N_8246);
nand U8704 (N_8704,N_8337,N_8202);
xnor U8705 (N_8705,N_8232,N_8001);
and U8706 (N_8706,N_8260,N_8368);
xor U8707 (N_8707,N_8311,N_8274);
and U8708 (N_8708,N_8144,N_8168);
nand U8709 (N_8709,N_8309,N_8426);
nor U8710 (N_8710,N_8112,N_8162);
and U8711 (N_8711,N_8367,N_8379);
nand U8712 (N_8712,N_8169,N_8167);
nor U8713 (N_8713,N_8458,N_8124);
or U8714 (N_8714,N_8350,N_8107);
xnor U8715 (N_8715,N_8109,N_8115);
nor U8716 (N_8716,N_8420,N_8195);
nand U8717 (N_8717,N_8273,N_8484);
or U8718 (N_8718,N_8096,N_8241);
nand U8719 (N_8719,N_8125,N_8322);
and U8720 (N_8720,N_8158,N_8248);
or U8721 (N_8721,N_8088,N_8336);
nor U8722 (N_8722,N_8252,N_8438);
or U8723 (N_8723,N_8164,N_8143);
xnor U8724 (N_8724,N_8348,N_8353);
nor U8725 (N_8725,N_8374,N_8200);
nor U8726 (N_8726,N_8078,N_8254);
and U8727 (N_8727,N_8472,N_8024);
and U8728 (N_8728,N_8217,N_8101);
and U8729 (N_8729,N_8068,N_8287);
and U8730 (N_8730,N_8093,N_8013);
nand U8731 (N_8731,N_8111,N_8161);
nor U8732 (N_8732,N_8262,N_8406);
nor U8733 (N_8733,N_8457,N_8382);
nor U8734 (N_8734,N_8417,N_8473);
nor U8735 (N_8735,N_8345,N_8388);
and U8736 (N_8736,N_8272,N_8131);
nand U8737 (N_8737,N_8251,N_8297);
nor U8738 (N_8738,N_8036,N_8340);
nor U8739 (N_8739,N_8355,N_8055);
nor U8740 (N_8740,N_8352,N_8029);
xnor U8741 (N_8741,N_8419,N_8218);
and U8742 (N_8742,N_8137,N_8166);
and U8743 (N_8743,N_8276,N_8342);
nor U8744 (N_8744,N_8142,N_8432);
and U8745 (N_8745,N_8063,N_8046);
nand U8746 (N_8746,N_8497,N_8255);
or U8747 (N_8747,N_8433,N_8138);
nand U8748 (N_8748,N_8061,N_8290);
or U8749 (N_8749,N_8105,N_8062);
and U8750 (N_8750,N_8227,N_8127);
nor U8751 (N_8751,N_8236,N_8366);
xnor U8752 (N_8752,N_8263,N_8049);
or U8753 (N_8753,N_8186,N_8228);
and U8754 (N_8754,N_8172,N_8349);
and U8755 (N_8755,N_8461,N_8172);
nor U8756 (N_8756,N_8389,N_8316);
or U8757 (N_8757,N_8454,N_8155);
nor U8758 (N_8758,N_8429,N_8252);
nand U8759 (N_8759,N_8042,N_8473);
nand U8760 (N_8760,N_8412,N_8115);
or U8761 (N_8761,N_8094,N_8411);
nand U8762 (N_8762,N_8120,N_8322);
or U8763 (N_8763,N_8354,N_8485);
and U8764 (N_8764,N_8127,N_8366);
nor U8765 (N_8765,N_8123,N_8160);
and U8766 (N_8766,N_8442,N_8223);
or U8767 (N_8767,N_8295,N_8052);
nand U8768 (N_8768,N_8166,N_8380);
or U8769 (N_8769,N_8335,N_8048);
and U8770 (N_8770,N_8270,N_8045);
or U8771 (N_8771,N_8030,N_8157);
or U8772 (N_8772,N_8224,N_8406);
or U8773 (N_8773,N_8071,N_8481);
xor U8774 (N_8774,N_8066,N_8148);
nand U8775 (N_8775,N_8175,N_8379);
nand U8776 (N_8776,N_8442,N_8440);
and U8777 (N_8777,N_8136,N_8135);
xnor U8778 (N_8778,N_8099,N_8490);
nand U8779 (N_8779,N_8075,N_8301);
nor U8780 (N_8780,N_8077,N_8404);
or U8781 (N_8781,N_8129,N_8429);
nand U8782 (N_8782,N_8310,N_8387);
or U8783 (N_8783,N_8298,N_8389);
and U8784 (N_8784,N_8094,N_8258);
xnor U8785 (N_8785,N_8171,N_8274);
nand U8786 (N_8786,N_8167,N_8247);
nand U8787 (N_8787,N_8241,N_8184);
nand U8788 (N_8788,N_8403,N_8007);
or U8789 (N_8789,N_8222,N_8331);
nor U8790 (N_8790,N_8446,N_8132);
nor U8791 (N_8791,N_8251,N_8053);
nor U8792 (N_8792,N_8363,N_8436);
nor U8793 (N_8793,N_8090,N_8337);
and U8794 (N_8794,N_8137,N_8231);
or U8795 (N_8795,N_8285,N_8206);
and U8796 (N_8796,N_8449,N_8273);
nand U8797 (N_8797,N_8190,N_8451);
xor U8798 (N_8798,N_8177,N_8497);
nor U8799 (N_8799,N_8137,N_8356);
nor U8800 (N_8800,N_8028,N_8033);
nand U8801 (N_8801,N_8234,N_8275);
nor U8802 (N_8802,N_8189,N_8367);
and U8803 (N_8803,N_8201,N_8478);
and U8804 (N_8804,N_8276,N_8328);
nand U8805 (N_8805,N_8065,N_8401);
or U8806 (N_8806,N_8141,N_8118);
and U8807 (N_8807,N_8066,N_8071);
nor U8808 (N_8808,N_8290,N_8268);
or U8809 (N_8809,N_8385,N_8477);
nor U8810 (N_8810,N_8329,N_8275);
or U8811 (N_8811,N_8195,N_8317);
nor U8812 (N_8812,N_8298,N_8427);
nor U8813 (N_8813,N_8231,N_8315);
nor U8814 (N_8814,N_8487,N_8253);
xor U8815 (N_8815,N_8113,N_8277);
nand U8816 (N_8816,N_8148,N_8126);
xor U8817 (N_8817,N_8091,N_8250);
nor U8818 (N_8818,N_8051,N_8093);
or U8819 (N_8819,N_8182,N_8495);
nor U8820 (N_8820,N_8354,N_8059);
or U8821 (N_8821,N_8423,N_8284);
xnor U8822 (N_8822,N_8448,N_8000);
and U8823 (N_8823,N_8401,N_8037);
or U8824 (N_8824,N_8051,N_8023);
xnor U8825 (N_8825,N_8431,N_8128);
or U8826 (N_8826,N_8095,N_8274);
or U8827 (N_8827,N_8325,N_8475);
nor U8828 (N_8828,N_8202,N_8445);
nand U8829 (N_8829,N_8387,N_8405);
xnor U8830 (N_8830,N_8361,N_8480);
and U8831 (N_8831,N_8469,N_8389);
xnor U8832 (N_8832,N_8263,N_8406);
xnor U8833 (N_8833,N_8141,N_8116);
nor U8834 (N_8834,N_8206,N_8472);
nand U8835 (N_8835,N_8459,N_8466);
nand U8836 (N_8836,N_8371,N_8069);
and U8837 (N_8837,N_8318,N_8022);
or U8838 (N_8838,N_8280,N_8093);
and U8839 (N_8839,N_8464,N_8413);
nand U8840 (N_8840,N_8097,N_8008);
or U8841 (N_8841,N_8141,N_8185);
nand U8842 (N_8842,N_8332,N_8385);
nand U8843 (N_8843,N_8314,N_8294);
and U8844 (N_8844,N_8124,N_8464);
nand U8845 (N_8845,N_8439,N_8129);
nor U8846 (N_8846,N_8119,N_8304);
nand U8847 (N_8847,N_8077,N_8000);
nand U8848 (N_8848,N_8395,N_8113);
and U8849 (N_8849,N_8204,N_8470);
nor U8850 (N_8850,N_8064,N_8110);
xor U8851 (N_8851,N_8234,N_8248);
xnor U8852 (N_8852,N_8384,N_8313);
nand U8853 (N_8853,N_8084,N_8145);
nand U8854 (N_8854,N_8213,N_8128);
and U8855 (N_8855,N_8102,N_8274);
and U8856 (N_8856,N_8046,N_8499);
or U8857 (N_8857,N_8205,N_8478);
and U8858 (N_8858,N_8206,N_8464);
nor U8859 (N_8859,N_8150,N_8263);
or U8860 (N_8860,N_8497,N_8295);
or U8861 (N_8861,N_8226,N_8462);
and U8862 (N_8862,N_8380,N_8285);
nor U8863 (N_8863,N_8270,N_8358);
nor U8864 (N_8864,N_8325,N_8450);
or U8865 (N_8865,N_8361,N_8466);
nand U8866 (N_8866,N_8061,N_8136);
nor U8867 (N_8867,N_8061,N_8013);
nor U8868 (N_8868,N_8408,N_8170);
xor U8869 (N_8869,N_8019,N_8065);
and U8870 (N_8870,N_8055,N_8018);
and U8871 (N_8871,N_8307,N_8128);
and U8872 (N_8872,N_8259,N_8005);
nor U8873 (N_8873,N_8461,N_8052);
nor U8874 (N_8874,N_8149,N_8469);
and U8875 (N_8875,N_8468,N_8249);
and U8876 (N_8876,N_8101,N_8037);
and U8877 (N_8877,N_8221,N_8253);
or U8878 (N_8878,N_8006,N_8286);
and U8879 (N_8879,N_8428,N_8002);
nand U8880 (N_8880,N_8024,N_8351);
and U8881 (N_8881,N_8080,N_8211);
or U8882 (N_8882,N_8072,N_8379);
nor U8883 (N_8883,N_8298,N_8262);
nand U8884 (N_8884,N_8150,N_8080);
and U8885 (N_8885,N_8206,N_8383);
and U8886 (N_8886,N_8429,N_8198);
or U8887 (N_8887,N_8083,N_8474);
xor U8888 (N_8888,N_8449,N_8337);
nand U8889 (N_8889,N_8276,N_8289);
nor U8890 (N_8890,N_8243,N_8355);
nor U8891 (N_8891,N_8053,N_8036);
and U8892 (N_8892,N_8213,N_8188);
nand U8893 (N_8893,N_8329,N_8465);
or U8894 (N_8894,N_8255,N_8368);
nand U8895 (N_8895,N_8115,N_8205);
and U8896 (N_8896,N_8464,N_8195);
and U8897 (N_8897,N_8017,N_8000);
and U8898 (N_8898,N_8446,N_8016);
nor U8899 (N_8899,N_8213,N_8240);
and U8900 (N_8900,N_8371,N_8448);
nor U8901 (N_8901,N_8345,N_8173);
or U8902 (N_8902,N_8368,N_8476);
and U8903 (N_8903,N_8315,N_8115);
xnor U8904 (N_8904,N_8369,N_8309);
nor U8905 (N_8905,N_8196,N_8287);
nor U8906 (N_8906,N_8460,N_8305);
or U8907 (N_8907,N_8228,N_8379);
or U8908 (N_8908,N_8348,N_8330);
and U8909 (N_8909,N_8352,N_8421);
nor U8910 (N_8910,N_8220,N_8259);
and U8911 (N_8911,N_8183,N_8095);
xor U8912 (N_8912,N_8420,N_8135);
and U8913 (N_8913,N_8109,N_8407);
and U8914 (N_8914,N_8451,N_8061);
and U8915 (N_8915,N_8300,N_8442);
and U8916 (N_8916,N_8271,N_8092);
or U8917 (N_8917,N_8377,N_8172);
nand U8918 (N_8918,N_8437,N_8499);
xor U8919 (N_8919,N_8066,N_8370);
and U8920 (N_8920,N_8183,N_8473);
or U8921 (N_8921,N_8399,N_8210);
and U8922 (N_8922,N_8386,N_8438);
and U8923 (N_8923,N_8021,N_8004);
nor U8924 (N_8924,N_8139,N_8248);
and U8925 (N_8925,N_8282,N_8162);
nand U8926 (N_8926,N_8436,N_8261);
and U8927 (N_8927,N_8068,N_8307);
and U8928 (N_8928,N_8005,N_8322);
and U8929 (N_8929,N_8409,N_8318);
and U8930 (N_8930,N_8175,N_8414);
nor U8931 (N_8931,N_8405,N_8105);
or U8932 (N_8932,N_8186,N_8022);
or U8933 (N_8933,N_8497,N_8344);
or U8934 (N_8934,N_8050,N_8131);
nand U8935 (N_8935,N_8293,N_8490);
or U8936 (N_8936,N_8267,N_8250);
or U8937 (N_8937,N_8409,N_8298);
nor U8938 (N_8938,N_8246,N_8048);
and U8939 (N_8939,N_8457,N_8126);
xnor U8940 (N_8940,N_8290,N_8043);
nor U8941 (N_8941,N_8496,N_8330);
nor U8942 (N_8942,N_8176,N_8346);
xor U8943 (N_8943,N_8401,N_8440);
xnor U8944 (N_8944,N_8351,N_8145);
nand U8945 (N_8945,N_8408,N_8441);
nor U8946 (N_8946,N_8399,N_8244);
xnor U8947 (N_8947,N_8453,N_8153);
or U8948 (N_8948,N_8442,N_8475);
or U8949 (N_8949,N_8170,N_8013);
and U8950 (N_8950,N_8444,N_8294);
or U8951 (N_8951,N_8017,N_8416);
xor U8952 (N_8952,N_8108,N_8379);
nand U8953 (N_8953,N_8099,N_8329);
or U8954 (N_8954,N_8221,N_8266);
nand U8955 (N_8955,N_8271,N_8494);
xor U8956 (N_8956,N_8137,N_8095);
nand U8957 (N_8957,N_8149,N_8498);
nor U8958 (N_8958,N_8029,N_8415);
nand U8959 (N_8959,N_8264,N_8466);
nor U8960 (N_8960,N_8388,N_8107);
nand U8961 (N_8961,N_8362,N_8338);
and U8962 (N_8962,N_8386,N_8029);
nor U8963 (N_8963,N_8390,N_8207);
and U8964 (N_8964,N_8397,N_8479);
or U8965 (N_8965,N_8392,N_8240);
nand U8966 (N_8966,N_8453,N_8369);
nor U8967 (N_8967,N_8027,N_8467);
xor U8968 (N_8968,N_8117,N_8476);
nand U8969 (N_8969,N_8345,N_8366);
and U8970 (N_8970,N_8358,N_8330);
or U8971 (N_8971,N_8060,N_8207);
nand U8972 (N_8972,N_8268,N_8301);
nand U8973 (N_8973,N_8308,N_8321);
or U8974 (N_8974,N_8398,N_8159);
and U8975 (N_8975,N_8273,N_8091);
or U8976 (N_8976,N_8108,N_8132);
or U8977 (N_8977,N_8025,N_8155);
and U8978 (N_8978,N_8179,N_8035);
and U8979 (N_8979,N_8001,N_8439);
or U8980 (N_8980,N_8492,N_8230);
and U8981 (N_8981,N_8245,N_8373);
or U8982 (N_8982,N_8216,N_8343);
nor U8983 (N_8983,N_8440,N_8236);
xnor U8984 (N_8984,N_8094,N_8409);
nand U8985 (N_8985,N_8488,N_8408);
and U8986 (N_8986,N_8062,N_8295);
nor U8987 (N_8987,N_8108,N_8462);
and U8988 (N_8988,N_8279,N_8153);
nand U8989 (N_8989,N_8247,N_8043);
nor U8990 (N_8990,N_8036,N_8486);
nand U8991 (N_8991,N_8047,N_8426);
and U8992 (N_8992,N_8075,N_8190);
nor U8993 (N_8993,N_8280,N_8253);
or U8994 (N_8994,N_8224,N_8192);
nand U8995 (N_8995,N_8117,N_8322);
nand U8996 (N_8996,N_8035,N_8165);
nor U8997 (N_8997,N_8481,N_8094);
and U8998 (N_8998,N_8188,N_8306);
xor U8999 (N_8999,N_8335,N_8365);
or U9000 (N_9000,N_8713,N_8741);
and U9001 (N_9001,N_8745,N_8712);
nor U9002 (N_9002,N_8677,N_8669);
xnor U9003 (N_9003,N_8815,N_8884);
nor U9004 (N_9004,N_8701,N_8634);
and U9005 (N_9005,N_8670,N_8936);
nand U9006 (N_9006,N_8934,N_8557);
or U9007 (N_9007,N_8740,N_8552);
nand U9008 (N_9008,N_8590,N_8940);
xor U9009 (N_9009,N_8807,N_8734);
nand U9010 (N_9010,N_8766,N_8641);
or U9011 (N_9011,N_8796,N_8563);
or U9012 (N_9012,N_8919,N_8653);
nand U9013 (N_9013,N_8850,N_8719);
and U9014 (N_9014,N_8503,N_8793);
nand U9015 (N_9015,N_8820,N_8879);
nand U9016 (N_9016,N_8671,N_8823);
or U9017 (N_9017,N_8529,N_8862);
nor U9018 (N_9018,N_8939,N_8863);
and U9019 (N_9019,N_8517,N_8831);
nor U9020 (N_9020,N_8658,N_8895);
or U9021 (N_9021,N_8759,N_8500);
nand U9022 (N_9022,N_8958,N_8989);
or U9023 (N_9023,N_8644,N_8646);
and U9024 (N_9024,N_8867,N_8572);
nand U9025 (N_9025,N_8767,N_8636);
and U9026 (N_9026,N_8853,N_8900);
nor U9027 (N_9027,N_8847,N_8663);
or U9028 (N_9028,N_8645,N_8979);
and U9029 (N_9029,N_8525,N_8684);
or U9030 (N_9030,N_8717,N_8893);
xor U9031 (N_9031,N_8542,N_8627);
and U9032 (N_9032,N_8654,N_8660);
and U9033 (N_9033,N_8642,N_8956);
nand U9034 (N_9034,N_8891,N_8533);
or U9035 (N_9035,N_8686,N_8812);
nand U9036 (N_9036,N_8649,N_8571);
nor U9037 (N_9037,N_8960,N_8833);
and U9038 (N_9038,N_8518,N_8507);
nor U9039 (N_9039,N_8547,N_8966);
or U9040 (N_9040,N_8926,N_8846);
nand U9041 (N_9041,N_8816,N_8953);
and U9042 (N_9042,N_8886,N_8744);
nor U9043 (N_9043,N_8664,N_8996);
and U9044 (N_9044,N_8675,N_8651);
and U9045 (N_9045,N_8769,N_8785);
and U9046 (N_9046,N_8594,N_8791);
and U9047 (N_9047,N_8625,N_8944);
nand U9048 (N_9048,N_8530,N_8802);
nor U9049 (N_9049,N_8808,N_8839);
and U9050 (N_9050,N_8779,N_8822);
or U9051 (N_9051,N_8694,N_8856);
xor U9052 (N_9052,N_8790,N_8591);
or U9053 (N_9053,N_8898,N_8986);
or U9054 (N_9054,N_8993,N_8509);
nor U9055 (N_9055,N_8848,N_8697);
nor U9056 (N_9056,N_8849,N_8782);
and U9057 (N_9057,N_8809,N_8558);
nand U9058 (N_9058,N_8760,N_8826);
or U9059 (N_9059,N_8994,N_8723);
and U9060 (N_9060,N_8623,N_8585);
and U9061 (N_9061,N_8976,N_8764);
nor U9062 (N_9062,N_8883,N_8611);
or U9063 (N_9063,N_8549,N_8511);
nor U9064 (N_9064,N_8655,N_8523);
xnor U9065 (N_9065,N_8521,N_8567);
nand U9066 (N_9066,N_8681,N_8730);
nor U9067 (N_9067,N_8845,N_8855);
or U9068 (N_9068,N_8505,N_8544);
and U9069 (N_9069,N_8817,N_8914);
nand U9070 (N_9070,N_8582,N_8922);
nor U9071 (N_9071,N_8588,N_8874);
nor U9072 (N_9072,N_8532,N_8749);
and U9073 (N_9073,N_8595,N_8650);
nand U9074 (N_9074,N_8616,N_8871);
and U9075 (N_9075,N_8576,N_8931);
nand U9076 (N_9076,N_8661,N_8955);
xnor U9077 (N_9077,N_8710,N_8562);
xnor U9078 (N_9078,N_8805,N_8535);
nor U9079 (N_9079,N_8774,N_8763);
and U9080 (N_9080,N_8548,N_8668);
nand U9081 (N_9081,N_8672,N_8860);
nor U9082 (N_9082,N_8758,N_8673);
nand U9083 (N_9083,N_8689,N_8602);
and U9084 (N_9084,N_8925,N_8866);
or U9085 (N_9085,N_8693,N_8735);
or U9086 (N_9086,N_8937,N_8910);
and U9087 (N_9087,N_8890,N_8827);
nand U9088 (N_9088,N_8948,N_8695);
nand U9089 (N_9089,N_8980,N_8584);
nand U9090 (N_9090,N_8656,N_8972);
and U9091 (N_9091,N_8998,N_8825);
xnor U9092 (N_9092,N_8707,N_8913);
or U9093 (N_9093,N_8528,N_8869);
nand U9094 (N_9094,N_8516,N_8539);
or U9095 (N_9095,N_8633,N_8514);
nand U9096 (N_9096,N_8703,N_8501);
or U9097 (N_9097,N_8512,N_8872);
and U9098 (N_9098,N_8965,N_8714);
or U9099 (N_9099,N_8810,N_8959);
and U9100 (N_9100,N_8834,N_8698);
and U9101 (N_9101,N_8792,N_8708);
nand U9102 (N_9102,N_8962,N_8909);
nor U9103 (N_9103,N_8924,N_8918);
nand U9104 (N_9104,N_8750,N_8773);
or U9105 (N_9105,N_8941,N_8865);
xnor U9106 (N_9106,N_8852,N_8731);
nand U9107 (N_9107,N_8752,N_8702);
and U9108 (N_9108,N_8945,N_8566);
nand U9109 (N_9109,N_8737,N_8682);
and U9110 (N_9110,N_8970,N_8711);
and U9111 (N_9111,N_8604,N_8508);
and U9112 (N_9112,N_8699,N_8772);
nor U9113 (N_9113,N_8967,N_8836);
xnor U9114 (N_9114,N_8929,N_8899);
nand U9115 (N_9115,N_8643,N_8932);
nor U9116 (N_9116,N_8841,N_8538);
or U9117 (N_9117,N_8587,N_8605);
nand U9118 (N_9118,N_8685,N_8575);
or U9119 (N_9119,N_8902,N_8504);
nand U9120 (N_9120,N_8506,N_8840);
nor U9121 (N_9121,N_8519,N_8678);
xnor U9122 (N_9122,N_8999,N_8596);
nand U9123 (N_9123,N_8640,N_8531);
nand U9124 (N_9124,N_8803,N_8720);
nor U9125 (N_9125,N_8964,N_8901);
or U9126 (N_9126,N_8923,N_8709);
nor U9127 (N_9127,N_8515,N_8739);
or U9128 (N_9128,N_8592,N_8727);
and U9129 (N_9129,N_8811,N_8800);
nand U9130 (N_9130,N_8502,N_8553);
or U9131 (N_9131,N_8513,N_8554);
or U9132 (N_9132,N_8639,N_8835);
nand U9133 (N_9133,N_8832,N_8888);
or U9134 (N_9134,N_8635,N_8599);
or U9135 (N_9135,N_8543,N_8838);
nor U9136 (N_9136,N_8534,N_8700);
or U9137 (N_9137,N_8804,N_8947);
or U9138 (N_9138,N_8814,N_8565);
nand U9139 (N_9139,N_8747,N_8935);
xor U9140 (N_9140,N_8706,N_8729);
nand U9141 (N_9141,N_8968,N_8778);
or U9142 (N_9142,N_8921,N_8662);
or U9143 (N_9143,N_8632,N_8877);
and U9144 (N_9144,N_8927,N_8854);
and U9145 (N_9145,N_8715,N_8622);
xor U9146 (N_9146,N_8577,N_8928);
and U9147 (N_9147,N_8736,N_8875);
or U9148 (N_9148,N_8679,N_8917);
and U9149 (N_9149,N_8579,N_8786);
xor U9150 (N_9150,N_8732,N_8560);
nand U9151 (N_9151,N_8615,N_8780);
nand U9152 (N_9152,N_8873,N_8526);
nor U9153 (N_9153,N_8768,N_8789);
nor U9154 (N_9154,N_8783,N_8995);
and U9155 (N_9155,N_8683,N_8600);
nand U9156 (N_9156,N_8775,N_8894);
and U9157 (N_9157,N_8943,N_8889);
or U9158 (N_9158,N_8905,N_8522);
nor U9159 (N_9159,N_8788,N_8546);
nand U9160 (N_9160,N_8527,N_8844);
or U9161 (N_9161,N_8957,N_8969);
and U9162 (N_9162,N_8665,N_8536);
nand U9163 (N_9163,N_8716,N_8887);
and U9164 (N_9164,N_8620,N_8950);
xnor U9165 (N_9165,N_8537,N_8991);
and U9166 (N_9166,N_8907,N_8801);
or U9167 (N_9167,N_8568,N_8601);
nor U9168 (N_9168,N_8743,N_8906);
nor U9169 (N_9169,N_8981,N_8837);
nand U9170 (N_9170,N_8946,N_8510);
or U9171 (N_9171,N_8988,N_8586);
and U9172 (N_9172,N_8770,N_8718);
or U9173 (N_9173,N_8762,N_8608);
and U9174 (N_9174,N_8676,N_8961);
and U9175 (N_9175,N_8692,N_8753);
and U9176 (N_9176,N_8722,N_8621);
nor U9177 (N_9177,N_8593,N_8912);
xor U9178 (N_9178,N_8550,N_8896);
nor U9179 (N_9179,N_8859,N_8541);
nand U9180 (N_9180,N_8583,N_8569);
nor U9181 (N_9181,N_8614,N_8892);
xnor U9182 (N_9182,N_8761,N_8674);
nand U9183 (N_9183,N_8637,N_8626);
nor U9184 (N_9184,N_8757,N_8612);
and U9185 (N_9185,N_8657,N_8659);
or U9186 (N_9186,N_8581,N_8933);
and U9187 (N_9187,N_8580,N_8971);
nor U9188 (N_9188,N_8748,N_8911);
or U9189 (N_9189,N_8798,N_8992);
or U9190 (N_9190,N_8619,N_8952);
nor U9191 (N_9191,N_8705,N_8806);
nor U9192 (N_9192,N_8648,N_8987);
and U9193 (N_9193,N_8742,N_8843);
or U9194 (N_9194,N_8573,N_8666);
and U9195 (N_9195,N_8578,N_8696);
xor U9196 (N_9196,N_8771,N_8880);
nand U9197 (N_9197,N_8618,N_8667);
nand U9198 (N_9198,N_8861,N_8813);
and U9199 (N_9199,N_8828,N_8631);
or U9200 (N_9200,N_8606,N_8830);
or U9201 (N_9201,N_8977,N_8545);
or U9202 (N_9202,N_8876,N_8897);
xor U9203 (N_9203,N_8975,N_8857);
nor U9204 (N_9204,N_8795,N_8603);
and U9205 (N_9205,N_8551,N_8638);
and U9206 (N_9206,N_8870,N_8610);
nor U9207 (N_9207,N_8652,N_8756);
and U9208 (N_9208,N_8690,N_8738);
or U9209 (N_9209,N_8751,N_8915);
nor U9210 (N_9210,N_8597,N_8868);
xor U9211 (N_9211,N_8574,N_8559);
and U9212 (N_9212,N_8725,N_8824);
xnor U9213 (N_9213,N_8985,N_8754);
or U9214 (N_9214,N_8777,N_8647);
and U9215 (N_9215,N_8842,N_8797);
and U9216 (N_9216,N_8949,N_8916);
nand U9217 (N_9217,N_8990,N_8903);
and U9218 (N_9218,N_8556,N_8881);
and U9219 (N_9219,N_8726,N_8555);
nand U9220 (N_9220,N_8570,N_8878);
nor U9221 (N_9221,N_8818,N_8520);
nand U9222 (N_9222,N_8942,N_8983);
nand U9223 (N_9223,N_8963,N_8617);
nor U9224 (N_9224,N_8561,N_8904);
nor U9225 (N_9225,N_8628,N_8733);
nor U9226 (N_9226,N_8864,N_8938);
and U9227 (N_9227,N_8630,N_8858);
and U9228 (N_9228,N_8784,N_8589);
nand U9229 (N_9229,N_8564,N_8704);
and U9230 (N_9230,N_8984,N_8908);
nor U9231 (N_9231,N_8680,N_8920);
or U9232 (N_9232,N_8746,N_8721);
nor U9233 (N_9233,N_8728,N_8540);
nand U9234 (N_9234,N_8982,N_8821);
nand U9235 (N_9235,N_8930,N_8688);
nand U9236 (N_9236,N_8794,N_8624);
nor U9237 (N_9237,N_8951,N_8978);
and U9238 (N_9238,N_8787,N_8724);
nor U9239 (N_9239,N_8829,N_8974);
or U9240 (N_9240,N_8776,N_8781);
nand U9241 (N_9241,N_8613,N_8885);
and U9242 (N_9242,N_8882,N_8954);
xnor U9243 (N_9243,N_8629,N_8691);
and U9244 (N_9244,N_8997,N_8765);
and U9245 (N_9245,N_8609,N_8687);
or U9246 (N_9246,N_8524,N_8598);
nand U9247 (N_9247,N_8973,N_8607);
nor U9248 (N_9248,N_8799,N_8851);
and U9249 (N_9249,N_8755,N_8819);
nor U9250 (N_9250,N_8697,N_8585);
nand U9251 (N_9251,N_8598,N_8567);
nor U9252 (N_9252,N_8617,N_8978);
or U9253 (N_9253,N_8688,N_8744);
nand U9254 (N_9254,N_8785,N_8815);
nand U9255 (N_9255,N_8580,N_8956);
nor U9256 (N_9256,N_8630,N_8870);
and U9257 (N_9257,N_8568,N_8919);
xor U9258 (N_9258,N_8730,N_8866);
nand U9259 (N_9259,N_8827,N_8929);
xor U9260 (N_9260,N_8838,N_8538);
or U9261 (N_9261,N_8934,N_8789);
or U9262 (N_9262,N_8765,N_8590);
xnor U9263 (N_9263,N_8600,N_8674);
and U9264 (N_9264,N_8576,N_8901);
nor U9265 (N_9265,N_8519,N_8717);
and U9266 (N_9266,N_8729,N_8788);
or U9267 (N_9267,N_8718,N_8753);
xor U9268 (N_9268,N_8940,N_8744);
or U9269 (N_9269,N_8808,N_8971);
nor U9270 (N_9270,N_8526,N_8977);
and U9271 (N_9271,N_8737,N_8907);
and U9272 (N_9272,N_8812,N_8616);
or U9273 (N_9273,N_8816,N_8598);
nor U9274 (N_9274,N_8519,N_8584);
and U9275 (N_9275,N_8703,N_8899);
or U9276 (N_9276,N_8610,N_8594);
and U9277 (N_9277,N_8910,N_8524);
or U9278 (N_9278,N_8839,N_8746);
or U9279 (N_9279,N_8970,N_8808);
nand U9280 (N_9280,N_8978,N_8804);
nand U9281 (N_9281,N_8671,N_8613);
or U9282 (N_9282,N_8583,N_8980);
nand U9283 (N_9283,N_8770,N_8813);
or U9284 (N_9284,N_8577,N_8818);
nand U9285 (N_9285,N_8811,N_8970);
nor U9286 (N_9286,N_8705,N_8863);
and U9287 (N_9287,N_8823,N_8802);
or U9288 (N_9288,N_8629,N_8926);
xor U9289 (N_9289,N_8540,N_8680);
nor U9290 (N_9290,N_8933,N_8562);
nor U9291 (N_9291,N_8593,N_8872);
or U9292 (N_9292,N_8855,N_8817);
and U9293 (N_9293,N_8756,N_8806);
or U9294 (N_9294,N_8661,N_8993);
and U9295 (N_9295,N_8645,N_8855);
or U9296 (N_9296,N_8698,N_8934);
nand U9297 (N_9297,N_8860,N_8524);
and U9298 (N_9298,N_8512,N_8772);
xnor U9299 (N_9299,N_8855,N_8529);
xor U9300 (N_9300,N_8882,N_8567);
nor U9301 (N_9301,N_8730,N_8638);
or U9302 (N_9302,N_8886,N_8735);
and U9303 (N_9303,N_8627,N_8708);
nor U9304 (N_9304,N_8611,N_8727);
and U9305 (N_9305,N_8541,N_8852);
or U9306 (N_9306,N_8829,N_8916);
nand U9307 (N_9307,N_8665,N_8980);
or U9308 (N_9308,N_8533,N_8963);
nand U9309 (N_9309,N_8962,N_8576);
or U9310 (N_9310,N_8523,N_8825);
and U9311 (N_9311,N_8829,N_8984);
and U9312 (N_9312,N_8708,N_8943);
nand U9313 (N_9313,N_8618,N_8732);
or U9314 (N_9314,N_8768,N_8835);
nand U9315 (N_9315,N_8914,N_8537);
nor U9316 (N_9316,N_8823,N_8781);
nor U9317 (N_9317,N_8875,N_8688);
nor U9318 (N_9318,N_8620,N_8630);
xor U9319 (N_9319,N_8623,N_8995);
or U9320 (N_9320,N_8729,N_8941);
nor U9321 (N_9321,N_8788,N_8961);
nor U9322 (N_9322,N_8758,N_8692);
and U9323 (N_9323,N_8693,N_8821);
nand U9324 (N_9324,N_8730,N_8805);
nor U9325 (N_9325,N_8926,N_8792);
nand U9326 (N_9326,N_8659,N_8985);
xnor U9327 (N_9327,N_8925,N_8606);
nor U9328 (N_9328,N_8793,N_8734);
xnor U9329 (N_9329,N_8701,N_8542);
nand U9330 (N_9330,N_8759,N_8832);
or U9331 (N_9331,N_8699,N_8658);
and U9332 (N_9332,N_8905,N_8949);
nor U9333 (N_9333,N_8518,N_8888);
or U9334 (N_9334,N_8642,N_8859);
and U9335 (N_9335,N_8595,N_8581);
nand U9336 (N_9336,N_8867,N_8528);
or U9337 (N_9337,N_8959,N_8833);
nand U9338 (N_9338,N_8517,N_8846);
nor U9339 (N_9339,N_8566,N_8580);
or U9340 (N_9340,N_8701,N_8915);
nor U9341 (N_9341,N_8807,N_8601);
or U9342 (N_9342,N_8573,N_8872);
nand U9343 (N_9343,N_8748,N_8566);
nand U9344 (N_9344,N_8771,N_8842);
and U9345 (N_9345,N_8948,N_8757);
and U9346 (N_9346,N_8957,N_8772);
nand U9347 (N_9347,N_8603,N_8529);
nand U9348 (N_9348,N_8854,N_8532);
or U9349 (N_9349,N_8974,N_8836);
nor U9350 (N_9350,N_8511,N_8729);
nand U9351 (N_9351,N_8542,N_8858);
and U9352 (N_9352,N_8994,N_8737);
and U9353 (N_9353,N_8813,N_8752);
nor U9354 (N_9354,N_8566,N_8899);
nor U9355 (N_9355,N_8630,N_8788);
and U9356 (N_9356,N_8542,N_8965);
and U9357 (N_9357,N_8705,N_8787);
nor U9358 (N_9358,N_8677,N_8962);
nor U9359 (N_9359,N_8950,N_8597);
nand U9360 (N_9360,N_8530,N_8963);
or U9361 (N_9361,N_8896,N_8892);
and U9362 (N_9362,N_8974,N_8874);
and U9363 (N_9363,N_8800,N_8832);
nand U9364 (N_9364,N_8668,N_8522);
nor U9365 (N_9365,N_8522,N_8821);
nor U9366 (N_9366,N_8671,N_8790);
xor U9367 (N_9367,N_8586,N_8741);
and U9368 (N_9368,N_8619,N_8796);
xor U9369 (N_9369,N_8691,N_8770);
xor U9370 (N_9370,N_8973,N_8613);
and U9371 (N_9371,N_8612,N_8551);
or U9372 (N_9372,N_8671,N_8795);
or U9373 (N_9373,N_8637,N_8595);
and U9374 (N_9374,N_8844,N_8827);
nor U9375 (N_9375,N_8700,N_8655);
and U9376 (N_9376,N_8631,N_8523);
and U9377 (N_9377,N_8663,N_8952);
nor U9378 (N_9378,N_8845,N_8674);
or U9379 (N_9379,N_8761,N_8586);
nand U9380 (N_9380,N_8956,N_8661);
nand U9381 (N_9381,N_8539,N_8838);
and U9382 (N_9382,N_8619,N_8630);
and U9383 (N_9383,N_8992,N_8523);
nand U9384 (N_9384,N_8849,N_8718);
nor U9385 (N_9385,N_8781,N_8991);
and U9386 (N_9386,N_8909,N_8810);
and U9387 (N_9387,N_8728,N_8870);
nand U9388 (N_9388,N_8565,N_8507);
nor U9389 (N_9389,N_8958,N_8776);
nand U9390 (N_9390,N_8745,N_8703);
and U9391 (N_9391,N_8714,N_8981);
nor U9392 (N_9392,N_8608,N_8621);
or U9393 (N_9393,N_8911,N_8761);
nand U9394 (N_9394,N_8946,N_8922);
nor U9395 (N_9395,N_8851,N_8856);
nand U9396 (N_9396,N_8792,N_8888);
nor U9397 (N_9397,N_8687,N_8755);
nor U9398 (N_9398,N_8921,N_8611);
nor U9399 (N_9399,N_8709,N_8800);
nand U9400 (N_9400,N_8769,N_8715);
nand U9401 (N_9401,N_8604,N_8876);
nor U9402 (N_9402,N_8526,N_8938);
xor U9403 (N_9403,N_8729,N_8553);
nor U9404 (N_9404,N_8614,N_8782);
or U9405 (N_9405,N_8722,N_8767);
nand U9406 (N_9406,N_8674,N_8742);
nor U9407 (N_9407,N_8677,N_8837);
and U9408 (N_9408,N_8651,N_8614);
or U9409 (N_9409,N_8903,N_8696);
or U9410 (N_9410,N_8709,N_8767);
and U9411 (N_9411,N_8991,N_8840);
xnor U9412 (N_9412,N_8884,N_8773);
xor U9413 (N_9413,N_8976,N_8584);
or U9414 (N_9414,N_8783,N_8843);
nor U9415 (N_9415,N_8607,N_8989);
or U9416 (N_9416,N_8520,N_8564);
nand U9417 (N_9417,N_8880,N_8720);
or U9418 (N_9418,N_8997,N_8933);
nand U9419 (N_9419,N_8597,N_8535);
nand U9420 (N_9420,N_8659,N_8629);
and U9421 (N_9421,N_8964,N_8811);
or U9422 (N_9422,N_8886,N_8665);
and U9423 (N_9423,N_8670,N_8981);
or U9424 (N_9424,N_8869,N_8778);
and U9425 (N_9425,N_8829,N_8857);
nor U9426 (N_9426,N_8642,N_8988);
xnor U9427 (N_9427,N_8987,N_8503);
and U9428 (N_9428,N_8970,N_8906);
xor U9429 (N_9429,N_8548,N_8703);
or U9430 (N_9430,N_8587,N_8935);
and U9431 (N_9431,N_8824,N_8897);
and U9432 (N_9432,N_8908,N_8589);
or U9433 (N_9433,N_8579,N_8794);
xnor U9434 (N_9434,N_8967,N_8691);
and U9435 (N_9435,N_8580,N_8946);
and U9436 (N_9436,N_8911,N_8535);
nor U9437 (N_9437,N_8710,N_8906);
nand U9438 (N_9438,N_8593,N_8932);
and U9439 (N_9439,N_8634,N_8683);
nor U9440 (N_9440,N_8549,N_8763);
nor U9441 (N_9441,N_8689,N_8953);
and U9442 (N_9442,N_8829,N_8520);
and U9443 (N_9443,N_8685,N_8567);
or U9444 (N_9444,N_8944,N_8910);
nand U9445 (N_9445,N_8840,N_8629);
or U9446 (N_9446,N_8582,N_8529);
nor U9447 (N_9447,N_8529,N_8863);
or U9448 (N_9448,N_8914,N_8915);
nor U9449 (N_9449,N_8788,N_8507);
or U9450 (N_9450,N_8821,N_8531);
or U9451 (N_9451,N_8956,N_8927);
nand U9452 (N_9452,N_8936,N_8586);
nor U9453 (N_9453,N_8672,N_8615);
nand U9454 (N_9454,N_8961,N_8988);
nor U9455 (N_9455,N_8970,N_8706);
nor U9456 (N_9456,N_8750,N_8732);
nor U9457 (N_9457,N_8568,N_8818);
and U9458 (N_9458,N_8523,N_8641);
nand U9459 (N_9459,N_8866,N_8971);
and U9460 (N_9460,N_8571,N_8617);
xor U9461 (N_9461,N_8648,N_8534);
nand U9462 (N_9462,N_8710,N_8634);
or U9463 (N_9463,N_8689,N_8599);
nor U9464 (N_9464,N_8946,N_8863);
nor U9465 (N_9465,N_8606,N_8904);
nor U9466 (N_9466,N_8658,N_8634);
or U9467 (N_9467,N_8743,N_8981);
xor U9468 (N_9468,N_8777,N_8609);
nand U9469 (N_9469,N_8661,N_8978);
nor U9470 (N_9470,N_8631,N_8590);
and U9471 (N_9471,N_8778,N_8928);
or U9472 (N_9472,N_8800,N_8944);
nor U9473 (N_9473,N_8558,N_8680);
and U9474 (N_9474,N_8813,N_8881);
or U9475 (N_9475,N_8829,N_8991);
or U9476 (N_9476,N_8918,N_8727);
xor U9477 (N_9477,N_8555,N_8851);
or U9478 (N_9478,N_8942,N_8576);
and U9479 (N_9479,N_8636,N_8590);
or U9480 (N_9480,N_8618,N_8876);
nand U9481 (N_9481,N_8648,N_8551);
nor U9482 (N_9482,N_8661,N_8848);
nor U9483 (N_9483,N_8884,N_8806);
and U9484 (N_9484,N_8537,N_8986);
nand U9485 (N_9485,N_8779,N_8849);
nand U9486 (N_9486,N_8606,N_8696);
nand U9487 (N_9487,N_8950,N_8665);
and U9488 (N_9488,N_8755,N_8704);
xnor U9489 (N_9489,N_8781,N_8932);
nand U9490 (N_9490,N_8956,N_8522);
nor U9491 (N_9491,N_8684,N_8992);
nor U9492 (N_9492,N_8702,N_8537);
and U9493 (N_9493,N_8853,N_8687);
xor U9494 (N_9494,N_8799,N_8906);
nand U9495 (N_9495,N_8575,N_8921);
xor U9496 (N_9496,N_8798,N_8768);
and U9497 (N_9497,N_8829,N_8738);
nand U9498 (N_9498,N_8600,N_8790);
or U9499 (N_9499,N_8502,N_8524);
or U9500 (N_9500,N_9410,N_9021);
or U9501 (N_9501,N_9222,N_9221);
nand U9502 (N_9502,N_9292,N_9071);
nor U9503 (N_9503,N_9412,N_9261);
and U9504 (N_9504,N_9102,N_9141);
nand U9505 (N_9505,N_9086,N_9123);
nand U9506 (N_9506,N_9143,N_9247);
nand U9507 (N_9507,N_9002,N_9263);
and U9508 (N_9508,N_9054,N_9363);
and U9509 (N_9509,N_9415,N_9219);
or U9510 (N_9510,N_9194,N_9444);
nand U9511 (N_9511,N_9160,N_9290);
and U9512 (N_9512,N_9182,N_9385);
and U9513 (N_9513,N_9231,N_9214);
or U9514 (N_9514,N_9293,N_9358);
and U9515 (N_9515,N_9027,N_9210);
xnor U9516 (N_9516,N_9333,N_9316);
nand U9517 (N_9517,N_9116,N_9060);
xnor U9518 (N_9518,N_9327,N_9236);
and U9519 (N_9519,N_9050,N_9268);
nand U9520 (N_9520,N_9201,N_9284);
nor U9521 (N_9521,N_9381,N_9346);
or U9522 (N_9522,N_9245,N_9131);
xor U9523 (N_9523,N_9049,N_9379);
nor U9524 (N_9524,N_9092,N_9438);
nand U9525 (N_9525,N_9421,N_9373);
or U9526 (N_9526,N_9476,N_9249);
and U9527 (N_9527,N_9258,N_9097);
nand U9528 (N_9528,N_9202,N_9163);
and U9529 (N_9529,N_9224,N_9463);
nor U9530 (N_9530,N_9154,N_9350);
nand U9531 (N_9531,N_9165,N_9023);
and U9532 (N_9532,N_9398,N_9034);
nand U9533 (N_9533,N_9462,N_9341);
nor U9534 (N_9534,N_9191,N_9348);
nand U9535 (N_9535,N_9349,N_9260);
nor U9536 (N_9536,N_9129,N_9195);
xnor U9537 (N_9537,N_9483,N_9240);
nand U9538 (N_9538,N_9397,N_9389);
nor U9539 (N_9539,N_9101,N_9057);
and U9540 (N_9540,N_9081,N_9113);
xnor U9541 (N_9541,N_9220,N_9144);
nand U9542 (N_9542,N_9134,N_9303);
or U9543 (N_9543,N_9487,N_9099);
nand U9544 (N_9544,N_9045,N_9416);
and U9545 (N_9545,N_9190,N_9361);
and U9546 (N_9546,N_9048,N_9169);
or U9547 (N_9547,N_9419,N_9271);
and U9548 (N_9548,N_9153,N_9337);
nand U9549 (N_9549,N_9365,N_9390);
and U9550 (N_9550,N_9152,N_9436);
xor U9551 (N_9551,N_9184,N_9321);
or U9552 (N_9552,N_9461,N_9331);
or U9553 (N_9553,N_9145,N_9037);
or U9554 (N_9554,N_9380,N_9474);
and U9555 (N_9555,N_9176,N_9353);
or U9556 (N_9556,N_9432,N_9198);
or U9557 (N_9557,N_9109,N_9022);
xnor U9558 (N_9558,N_9400,N_9253);
and U9559 (N_9559,N_9157,N_9428);
nand U9560 (N_9560,N_9019,N_9264);
nand U9561 (N_9561,N_9124,N_9304);
and U9562 (N_9562,N_9082,N_9283);
and U9563 (N_9563,N_9059,N_9417);
and U9564 (N_9564,N_9025,N_9107);
nor U9565 (N_9565,N_9007,N_9492);
or U9566 (N_9566,N_9375,N_9180);
xor U9567 (N_9567,N_9014,N_9368);
nand U9568 (N_9568,N_9056,N_9067);
xor U9569 (N_9569,N_9068,N_9323);
xor U9570 (N_9570,N_9382,N_9174);
or U9571 (N_9571,N_9020,N_9343);
nand U9572 (N_9572,N_9424,N_9026);
nand U9573 (N_9573,N_9013,N_9089);
and U9574 (N_9574,N_9105,N_9139);
nor U9575 (N_9575,N_9356,N_9427);
nor U9576 (N_9576,N_9093,N_9238);
or U9577 (N_9577,N_9171,N_9120);
nand U9578 (N_9578,N_9326,N_9429);
nand U9579 (N_9579,N_9032,N_9499);
nand U9580 (N_9580,N_9062,N_9309);
xnor U9581 (N_9581,N_9008,N_9423);
nand U9582 (N_9582,N_9345,N_9396);
nand U9583 (N_9583,N_9447,N_9076);
nor U9584 (N_9584,N_9005,N_9012);
and U9585 (N_9585,N_9469,N_9334);
nor U9586 (N_9586,N_9192,N_9016);
or U9587 (N_9587,N_9112,N_9272);
or U9588 (N_9588,N_9282,N_9243);
nand U9589 (N_9589,N_9278,N_9497);
xnor U9590 (N_9590,N_9445,N_9015);
nand U9591 (N_9591,N_9362,N_9186);
xnor U9592 (N_9592,N_9401,N_9246);
xor U9593 (N_9593,N_9480,N_9471);
nand U9594 (N_9594,N_9308,N_9472);
or U9595 (N_9595,N_9226,N_9262);
or U9596 (N_9596,N_9332,N_9166);
or U9597 (N_9597,N_9460,N_9248);
nor U9598 (N_9598,N_9473,N_9302);
or U9599 (N_9599,N_9030,N_9420);
and U9600 (N_9600,N_9065,N_9108);
nand U9601 (N_9601,N_9074,N_9273);
and U9602 (N_9602,N_9127,N_9149);
nor U9603 (N_9603,N_9399,N_9244);
or U9604 (N_9604,N_9147,N_9205);
and U9605 (N_9605,N_9442,N_9256);
nor U9606 (N_9606,N_9465,N_9208);
nor U9607 (N_9607,N_9150,N_9087);
or U9608 (N_9608,N_9235,N_9212);
xor U9609 (N_9609,N_9041,N_9291);
nand U9610 (N_9610,N_9320,N_9374);
and U9611 (N_9611,N_9018,N_9435);
and U9612 (N_9612,N_9338,N_9259);
and U9613 (N_9613,N_9162,N_9265);
or U9614 (N_9614,N_9223,N_9126);
nand U9615 (N_9615,N_9340,N_9464);
or U9616 (N_9616,N_9342,N_9252);
and U9617 (N_9617,N_9161,N_9458);
nor U9618 (N_9618,N_9498,N_9151);
or U9619 (N_9619,N_9364,N_9075);
nor U9620 (N_9620,N_9009,N_9117);
and U9621 (N_9621,N_9122,N_9482);
and U9622 (N_9622,N_9029,N_9354);
nor U9623 (N_9623,N_9204,N_9178);
nor U9624 (N_9624,N_9481,N_9392);
nand U9625 (N_9625,N_9197,N_9359);
xor U9626 (N_9626,N_9006,N_9280);
nand U9627 (N_9627,N_9010,N_9215);
or U9628 (N_9628,N_9307,N_9310);
xor U9629 (N_9629,N_9237,N_9360);
xor U9630 (N_9630,N_9218,N_9175);
or U9631 (N_9631,N_9227,N_9241);
xor U9632 (N_9632,N_9386,N_9043);
and U9633 (N_9633,N_9287,N_9207);
nand U9634 (N_9634,N_9485,N_9179);
and U9635 (N_9635,N_9267,N_9489);
nand U9636 (N_9636,N_9046,N_9403);
or U9637 (N_9637,N_9233,N_9311);
xor U9638 (N_9638,N_9196,N_9185);
and U9639 (N_9639,N_9314,N_9189);
nand U9640 (N_9640,N_9078,N_9090);
or U9641 (N_9641,N_9443,N_9004);
and U9642 (N_9642,N_9437,N_9156);
and U9643 (N_9643,N_9251,N_9325);
or U9644 (N_9644,N_9275,N_9077);
nor U9645 (N_9645,N_9404,N_9330);
or U9646 (N_9646,N_9211,N_9477);
xor U9647 (N_9647,N_9328,N_9494);
nor U9648 (N_9648,N_9072,N_9199);
nor U9649 (N_9649,N_9322,N_9384);
or U9650 (N_9650,N_9305,N_9234);
and U9651 (N_9651,N_9301,N_9289);
or U9652 (N_9652,N_9387,N_9193);
nor U9653 (N_9653,N_9270,N_9490);
and U9654 (N_9654,N_9335,N_9430);
nand U9655 (N_9655,N_9414,N_9459);
or U9656 (N_9656,N_9170,N_9257);
and U9657 (N_9657,N_9003,N_9047);
and U9658 (N_9658,N_9319,N_9033);
or U9659 (N_9659,N_9313,N_9426);
or U9660 (N_9660,N_9213,N_9266);
nand U9661 (N_9661,N_9425,N_9298);
nor U9662 (N_9662,N_9052,N_9355);
nor U9663 (N_9663,N_9225,N_9281);
nor U9664 (N_9664,N_9091,N_9111);
and U9665 (N_9665,N_9017,N_9155);
xor U9666 (N_9666,N_9409,N_9312);
or U9667 (N_9667,N_9230,N_9453);
nor U9668 (N_9668,N_9133,N_9066);
nand U9669 (N_9669,N_9285,N_9434);
nand U9670 (N_9670,N_9168,N_9055);
or U9671 (N_9671,N_9394,N_9457);
xor U9672 (N_9672,N_9255,N_9376);
or U9673 (N_9673,N_9402,N_9115);
xor U9674 (N_9674,N_9254,N_9058);
nand U9675 (N_9675,N_9391,N_9393);
nand U9676 (N_9676,N_9164,N_9318);
and U9677 (N_9677,N_9172,N_9377);
or U9678 (N_9678,N_9486,N_9061);
xor U9679 (N_9679,N_9095,N_9466);
nor U9680 (N_9680,N_9200,N_9142);
nor U9681 (N_9681,N_9339,N_9096);
and U9682 (N_9682,N_9135,N_9063);
nand U9683 (N_9683,N_9118,N_9452);
and U9684 (N_9684,N_9036,N_9478);
and U9685 (N_9685,N_9069,N_9229);
nor U9686 (N_9686,N_9294,N_9378);
nor U9687 (N_9687,N_9408,N_9468);
xnor U9688 (N_9688,N_9084,N_9479);
and U9689 (N_9689,N_9455,N_9159);
or U9690 (N_9690,N_9232,N_9274);
or U9691 (N_9691,N_9035,N_9028);
and U9692 (N_9692,N_9053,N_9228);
nand U9693 (N_9693,N_9418,N_9119);
and U9694 (N_9694,N_9173,N_9146);
or U9695 (N_9695,N_9406,N_9446);
nor U9696 (N_9696,N_9366,N_9306);
nor U9697 (N_9697,N_9440,N_9299);
or U9698 (N_9698,N_9357,N_9411);
and U9699 (N_9699,N_9024,N_9070);
or U9700 (N_9700,N_9085,N_9079);
xnor U9701 (N_9701,N_9125,N_9422);
nor U9702 (N_9702,N_9106,N_9140);
nand U9703 (N_9703,N_9039,N_9203);
nand U9704 (N_9704,N_9369,N_9080);
or U9705 (N_9705,N_9040,N_9395);
or U9706 (N_9706,N_9297,N_9137);
xor U9707 (N_9707,N_9098,N_9000);
nor U9708 (N_9708,N_9051,N_9295);
nand U9709 (N_9709,N_9044,N_9148);
or U9710 (N_9710,N_9110,N_9372);
nor U9711 (N_9711,N_9493,N_9324);
or U9712 (N_9712,N_9104,N_9488);
or U9713 (N_9713,N_9276,N_9431);
nand U9714 (N_9714,N_9183,N_9042);
or U9715 (N_9715,N_9250,N_9296);
or U9716 (N_9716,N_9467,N_9064);
nor U9717 (N_9717,N_9371,N_9484);
nand U9718 (N_9718,N_9288,N_9239);
nand U9719 (N_9719,N_9495,N_9470);
or U9720 (N_9720,N_9405,N_9279);
nor U9721 (N_9721,N_9088,N_9351);
or U9722 (N_9722,N_9031,N_9001);
and U9723 (N_9723,N_9491,N_9352);
nand U9724 (N_9724,N_9475,N_9128);
nor U9725 (N_9725,N_9011,N_9413);
nor U9726 (N_9726,N_9269,N_9187);
xnor U9727 (N_9727,N_9209,N_9433);
nor U9728 (N_9728,N_9456,N_9094);
nand U9729 (N_9729,N_9450,N_9407);
or U9730 (N_9730,N_9103,N_9100);
nand U9731 (N_9731,N_9188,N_9130);
and U9732 (N_9732,N_9336,N_9242);
nor U9733 (N_9733,N_9344,N_9300);
or U9734 (N_9734,N_9114,N_9181);
or U9735 (N_9735,N_9038,N_9286);
and U9736 (N_9736,N_9121,N_9073);
or U9737 (N_9737,N_9167,N_9138);
xor U9738 (N_9738,N_9451,N_9136);
or U9739 (N_9739,N_9388,N_9448);
nand U9740 (N_9740,N_9206,N_9216);
and U9741 (N_9741,N_9383,N_9329);
nand U9742 (N_9742,N_9277,N_9454);
nand U9743 (N_9743,N_9317,N_9439);
or U9744 (N_9744,N_9347,N_9132);
nor U9745 (N_9745,N_9370,N_9315);
nand U9746 (N_9746,N_9177,N_9367);
nor U9747 (N_9747,N_9496,N_9441);
and U9748 (N_9748,N_9449,N_9217);
xnor U9749 (N_9749,N_9158,N_9083);
and U9750 (N_9750,N_9024,N_9237);
and U9751 (N_9751,N_9094,N_9041);
or U9752 (N_9752,N_9289,N_9494);
nand U9753 (N_9753,N_9343,N_9450);
or U9754 (N_9754,N_9089,N_9285);
or U9755 (N_9755,N_9468,N_9011);
nand U9756 (N_9756,N_9281,N_9084);
nand U9757 (N_9757,N_9088,N_9444);
nand U9758 (N_9758,N_9305,N_9299);
or U9759 (N_9759,N_9185,N_9267);
or U9760 (N_9760,N_9073,N_9000);
and U9761 (N_9761,N_9460,N_9446);
or U9762 (N_9762,N_9053,N_9058);
and U9763 (N_9763,N_9311,N_9218);
or U9764 (N_9764,N_9257,N_9271);
nor U9765 (N_9765,N_9011,N_9046);
and U9766 (N_9766,N_9097,N_9205);
and U9767 (N_9767,N_9075,N_9254);
and U9768 (N_9768,N_9383,N_9463);
nor U9769 (N_9769,N_9005,N_9299);
or U9770 (N_9770,N_9232,N_9070);
nor U9771 (N_9771,N_9094,N_9406);
or U9772 (N_9772,N_9306,N_9181);
nor U9773 (N_9773,N_9373,N_9096);
nor U9774 (N_9774,N_9327,N_9468);
nand U9775 (N_9775,N_9304,N_9178);
nand U9776 (N_9776,N_9309,N_9202);
nand U9777 (N_9777,N_9340,N_9469);
nand U9778 (N_9778,N_9350,N_9281);
and U9779 (N_9779,N_9171,N_9360);
or U9780 (N_9780,N_9237,N_9182);
nor U9781 (N_9781,N_9459,N_9038);
nor U9782 (N_9782,N_9114,N_9250);
or U9783 (N_9783,N_9249,N_9305);
xnor U9784 (N_9784,N_9284,N_9383);
nor U9785 (N_9785,N_9276,N_9237);
or U9786 (N_9786,N_9023,N_9017);
or U9787 (N_9787,N_9284,N_9341);
or U9788 (N_9788,N_9357,N_9369);
nand U9789 (N_9789,N_9410,N_9220);
and U9790 (N_9790,N_9310,N_9485);
xor U9791 (N_9791,N_9222,N_9106);
nand U9792 (N_9792,N_9196,N_9394);
xnor U9793 (N_9793,N_9079,N_9020);
and U9794 (N_9794,N_9387,N_9239);
nand U9795 (N_9795,N_9149,N_9441);
nand U9796 (N_9796,N_9461,N_9371);
nand U9797 (N_9797,N_9253,N_9029);
nand U9798 (N_9798,N_9101,N_9444);
nand U9799 (N_9799,N_9233,N_9437);
nor U9800 (N_9800,N_9366,N_9312);
nor U9801 (N_9801,N_9259,N_9185);
nor U9802 (N_9802,N_9096,N_9126);
nor U9803 (N_9803,N_9436,N_9297);
or U9804 (N_9804,N_9231,N_9091);
nor U9805 (N_9805,N_9367,N_9448);
or U9806 (N_9806,N_9219,N_9006);
and U9807 (N_9807,N_9116,N_9054);
nor U9808 (N_9808,N_9283,N_9431);
nor U9809 (N_9809,N_9361,N_9469);
or U9810 (N_9810,N_9025,N_9204);
or U9811 (N_9811,N_9495,N_9472);
and U9812 (N_9812,N_9369,N_9464);
nor U9813 (N_9813,N_9105,N_9402);
nor U9814 (N_9814,N_9177,N_9390);
or U9815 (N_9815,N_9282,N_9345);
xor U9816 (N_9816,N_9463,N_9160);
or U9817 (N_9817,N_9211,N_9483);
xnor U9818 (N_9818,N_9144,N_9430);
nor U9819 (N_9819,N_9468,N_9433);
or U9820 (N_9820,N_9461,N_9394);
and U9821 (N_9821,N_9401,N_9410);
and U9822 (N_9822,N_9193,N_9163);
nand U9823 (N_9823,N_9107,N_9110);
or U9824 (N_9824,N_9219,N_9498);
or U9825 (N_9825,N_9373,N_9356);
nand U9826 (N_9826,N_9184,N_9403);
or U9827 (N_9827,N_9434,N_9457);
nor U9828 (N_9828,N_9202,N_9115);
xor U9829 (N_9829,N_9108,N_9473);
nor U9830 (N_9830,N_9389,N_9187);
and U9831 (N_9831,N_9246,N_9462);
nor U9832 (N_9832,N_9123,N_9379);
nor U9833 (N_9833,N_9452,N_9146);
or U9834 (N_9834,N_9025,N_9496);
or U9835 (N_9835,N_9169,N_9249);
nor U9836 (N_9836,N_9328,N_9426);
or U9837 (N_9837,N_9311,N_9031);
and U9838 (N_9838,N_9148,N_9038);
nand U9839 (N_9839,N_9067,N_9299);
xnor U9840 (N_9840,N_9183,N_9409);
xnor U9841 (N_9841,N_9225,N_9452);
and U9842 (N_9842,N_9418,N_9166);
or U9843 (N_9843,N_9344,N_9247);
nor U9844 (N_9844,N_9072,N_9036);
or U9845 (N_9845,N_9316,N_9321);
xnor U9846 (N_9846,N_9368,N_9366);
nand U9847 (N_9847,N_9364,N_9369);
or U9848 (N_9848,N_9324,N_9067);
xor U9849 (N_9849,N_9142,N_9198);
nand U9850 (N_9850,N_9478,N_9291);
nor U9851 (N_9851,N_9242,N_9174);
or U9852 (N_9852,N_9043,N_9442);
nand U9853 (N_9853,N_9251,N_9039);
xor U9854 (N_9854,N_9247,N_9308);
nand U9855 (N_9855,N_9476,N_9193);
and U9856 (N_9856,N_9327,N_9008);
nand U9857 (N_9857,N_9424,N_9180);
nand U9858 (N_9858,N_9424,N_9041);
and U9859 (N_9859,N_9392,N_9308);
xnor U9860 (N_9860,N_9443,N_9045);
or U9861 (N_9861,N_9176,N_9225);
and U9862 (N_9862,N_9242,N_9493);
or U9863 (N_9863,N_9237,N_9391);
nand U9864 (N_9864,N_9079,N_9431);
and U9865 (N_9865,N_9168,N_9275);
xnor U9866 (N_9866,N_9413,N_9053);
and U9867 (N_9867,N_9188,N_9338);
nor U9868 (N_9868,N_9233,N_9469);
nand U9869 (N_9869,N_9435,N_9458);
and U9870 (N_9870,N_9327,N_9422);
nor U9871 (N_9871,N_9099,N_9245);
nand U9872 (N_9872,N_9408,N_9498);
nand U9873 (N_9873,N_9063,N_9380);
and U9874 (N_9874,N_9164,N_9220);
xnor U9875 (N_9875,N_9300,N_9447);
nand U9876 (N_9876,N_9256,N_9338);
nor U9877 (N_9877,N_9410,N_9222);
nor U9878 (N_9878,N_9213,N_9339);
nand U9879 (N_9879,N_9086,N_9021);
and U9880 (N_9880,N_9314,N_9045);
xnor U9881 (N_9881,N_9314,N_9403);
nand U9882 (N_9882,N_9196,N_9416);
and U9883 (N_9883,N_9034,N_9386);
nand U9884 (N_9884,N_9089,N_9316);
and U9885 (N_9885,N_9037,N_9263);
and U9886 (N_9886,N_9186,N_9073);
and U9887 (N_9887,N_9052,N_9009);
or U9888 (N_9888,N_9307,N_9444);
and U9889 (N_9889,N_9159,N_9304);
nor U9890 (N_9890,N_9438,N_9025);
nand U9891 (N_9891,N_9345,N_9288);
xor U9892 (N_9892,N_9186,N_9145);
and U9893 (N_9893,N_9336,N_9371);
nand U9894 (N_9894,N_9063,N_9461);
nand U9895 (N_9895,N_9051,N_9403);
nor U9896 (N_9896,N_9486,N_9152);
and U9897 (N_9897,N_9488,N_9498);
nor U9898 (N_9898,N_9169,N_9084);
and U9899 (N_9899,N_9246,N_9077);
nand U9900 (N_9900,N_9099,N_9289);
or U9901 (N_9901,N_9168,N_9450);
and U9902 (N_9902,N_9148,N_9380);
or U9903 (N_9903,N_9310,N_9096);
nor U9904 (N_9904,N_9394,N_9216);
xnor U9905 (N_9905,N_9181,N_9164);
or U9906 (N_9906,N_9022,N_9207);
nor U9907 (N_9907,N_9277,N_9332);
and U9908 (N_9908,N_9353,N_9027);
nand U9909 (N_9909,N_9280,N_9128);
nand U9910 (N_9910,N_9020,N_9286);
and U9911 (N_9911,N_9426,N_9343);
nor U9912 (N_9912,N_9148,N_9008);
or U9913 (N_9913,N_9058,N_9217);
xor U9914 (N_9914,N_9459,N_9312);
or U9915 (N_9915,N_9259,N_9018);
nand U9916 (N_9916,N_9430,N_9410);
or U9917 (N_9917,N_9231,N_9333);
nor U9918 (N_9918,N_9050,N_9223);
nor U9919 (N_9919,N_9475,N_9046);
nor U9920 (N_9920,N_9080,N_9372);
xnor U9921 (N_9921,N_9188,N_9302);
nor U9922 (N_9922,N_9451,N_9356);
nand U9923 (N_9923,N_9253,N_9474);
and U9924 (N_9924,N_9255,N_9134);
or U9925 (N_9925,N_9042,N_9191);
or U9926 (N_9926,N_9180,N_9444);
nand U9927 (N_9927,N_9473,N_9076);
nor U9928 (N_9928,N_9361,N_9300);
and U9929 (N_9929,N_9418,N_9149);
xor U9930 (N_9930,N_9259,N_9178);
nand U9931 (N_9931,N_9318,N_9243);
or U9932 (N_9932,N_9188,N_9462);
nor U9933 (N_9933,N_9278,N_9480);
nor U9934 (N_9934,N_9406,N_9219);
nand U9935 (N_9935,N_9482,N_9303);
nor U9936 (N_9936,N_9158,N_9141);
and U9937 (N_9937,N_9455,N_9340);
and U9938 (N_9938,N_9433,N_9281);
and U9939 (N_9939,N_9398,N_9343);
or U9940 (N_9940,N_9068,N_9415);
nor U9941 (N_9941,N_9234,N_9353);
nor U9942 (N_9942,N_9322,N_9334);
or U9943 (N_9943,N_9498,N_9263);
nand U9944 (N_9944,N_9295,N_9268);
or U9945 (N_9945,N_9497,N_9155);
nand U9946 (N_9946,N_9424,N_9152);
or U9947 (N_9947,N_9487,N_9477);
nor U9948 (N_9948,N_9157,N_9029);
and U9949 (N_9949,N_9394,N_9044);
nor U9950 (N_9950,N_9103,N_9210);
and U9951 (N_9951,N_9166,N_9093);
nor U9952 (N_9952,N_9147,N_9080);
or U9953 (N_9953,N_9053,N_9154);
nand U9954 (N_9954,N_9248,N_9264);
nand U9955 (N_9955,N_9231,N_9235);
nand U9956 (N_9956,N_9026,N_9043);
and U9957 (N_9957,N_9100,N_9456);
and U9958 (N_9958,N_9213,N_9168);
nor U9959 (N_9959,N_9352,N_9203);
or U9960 (N_9960,N_9054,N_9337);
nor U9961 (N_9961,N_9277,N_9007);
and U9962 (N_9962,N_9393,N_9283);
and U9963 (N_9963,N_9456,N_9365);
and U9964 (N_9964,N_9132,N_9326);
and U9965 (N_9965,N_9355,N_9071);
nand U9966 (N_9966,N_9433,N_9479);
or U9967 (N_9967,N_9348,N_9164);
nand U9968 (N_9968,N_9477,N_9106);
nand U9969 (N_9969,N_9422,N_9041);
nand U9970 (N_9970,N_9383,N_9398);
xor U9971 (N_9971,N_9331,N_9237);
xor U9972 (N_9972,N_9170,N_9237);
nand U9973 (N_9973,N_9182,N_9153);
nand U9974 (N_9974,N_9410,N_9203);
nor U9975 (N_9975,N_9169,N_9081);
and U9976 (N_9976,N_9354,N_9230);
xor U9977 (N_9977,N_9383,N_9048);
or U9978 (N_9978,N_9260,N_9434);
or U9979 (N_9979,N_9049,N_9238);
nor U9980 (N_9980,N_9298,N_9311);
nand U9981 (N_9981,N_9348,N_9022);
nor U9982 (N_9982,N_9091,N_9246);
nor U9983 (N_9983,N_9418,N_9392);
nand U9984 (N_9984,N_9234,N_9241);
nor U9985 (N_9985,N_9428,N_9425);
nor U9986 (N_9986,N_9099,N_9394);
nor U9987 (N_9987,N_9146,N_9073);
nand U9988 (N_9988,N_9000,N_9167);
or U9989 (N_9989,N_9241,N_9402);
nor U9990 (N_9990,N_9196,N_9186);
and U9991 (N_9991,N_9491,N_9412);
nor U9992 (N_9992,N_9115,N_9055);
nor U9993 (N_9993,N_9282,N_9154);
or U9994 (N_9994,N_9148,N_9075);
nand U9995 (N_9995,N_9099,N_9443);
nand U9996 (N_9996,N_9050,N_9432);
or U9997 (N_9997,N_9250,N_9406);
or U9998 (N_9998,N_9156,N_9042);
nor U9999 (N_9999,N_9110,N_9484);
nand UO_0 (O_0,N_9691,N_9790);
xor UO_1 (O_1,N_9880,N_9764);
nand UO_2 (O_2,N_9536,N_9916);
or UO_3 (O_3,N_9861,N_9506);
or UO_4 (O_4,N_9918,N_9785);
and UO_5 (O_5,N_9595,N_9558);
xor UO_6 (O_6,N_9737,N_9721);
and UO_7 (O_7,N_9652,N_9728);
or UO_8 (O_8,N_9964,N_9634);
and UO_9 (O_9,N_9935,N_9948);
or UO_10 (O_10,N_9954,N_9925);
and UO_11 (O_11,N_9600,N_9692);
and UO_12 (O_12,N_9674,N_9503);
nor UO_13 (O_13,N_9718,N_9646);
nor UO_14 (O_14,N_9505,N_9519);
and UO_15 (O_15,N_9981,N_9758);
nand UO_16 (O_16,N_9798,N_9965);
nor UO_17 (O_17,N_9654,N_9883);
or UO_18 (O_18,N_9770,N_9601);
and UO_19 (O_19,N_9663,N_9852);
or UO_20 (O_20,N_9914,N_9507);
nand UO_21 (O_21,N_9958,N_9650);
nor UO_22 (O_22,N_9768,N_9618);
and UO_23 (O_23,N_9690,N_9651);
nor UO_24 (O_24,N_9774,N_9734);
or UO_25 (O_25,N_9990,N_9963);
nor UO_26 (O_26,N_9816,N_9658);
xor UO_27 (O_27,N_9730,N_9851);
nand UO_28 (O_28,N_9573,N_9788);
nand UO_29 (O_29,N_9738,N_9942);
or UO_30 (O_30,N_9677,N_9629);
xor UO_31 (O_31,N_9742,N_9806);
and UO_32 (O_32,N_9619,N_9800);
or UO_33 (O_33,N_9676,N_9797);
and UO_34 (O_34,N_9864,N_9946);
xnor UO_35 (O_35,N_9613,N_9858);
nand UO_36 (O_36,N_9833,N_9775);
and UO_37 (O_37,N_9823,N_9602);
xor UO_38 (O_38,N_9560,N_9894);
nor UO_39 (O_39,N_9756,N_9989);
or UO_40 (O_40,N_9675,N_9678);
nand UO_41 (O_41,N_9923,N_9520);
nor UO_42 (O_42,N_9594,N_9992);
or UO_43 (O_43,N_9943,N_9753);
or UO_44 (O_44,N_9897,N_9735);
or UO_45 (O_45,N_9604,N_9726);
and UO_46 (O_46,N_9926,N_9615);
nor UO_47 (O_47,N_9696,N_9898);
nand UO_48 (O_48,N_9695,N_9588);
xnor UO_49 (O_49,N_9781,N_9644);
nor UO_50 (O_50,N_9875,N_9809);
and UO_51 (O_51,N_9521,N_9599);
nor UO_52 (O_52,N_9638,N_9952);
xor UO_53 (O_53,N_9722,N_9666);
nand UO_54 (O_54,N_9636,N_9553);
and UO_55 (O_55,N_9708,N_9821);
and UO_56 (O_56,N_9596,N_9986);
nand UO_57 (O_57,N_9642,N_9856);
nand UO_58 (O_58,N_9955,N_9540);
nand UO_59 (O_59,N_9870,N_9834);
nor UO_60 (O_60,N_9524,N_9847);
and UO_61 (O_61,N_9713,N_9578);
nand UO_62 (O_62,N_9773,N_9882);
or UO_63 (O_63,N_9569,N_9736);
and UO_64 (O_64,N_9777,N_9538);
and UO_65 (O_65,N_9866,N_9577);
xnor UO_66 (O_66,N_9912,N_9513);
nor UO_67 (O_67,N_9716,N_9939);
and UO_68 (O_68,N_9749,N_9702);
xor UO_69 (O_69,N_9687,N_9759);
and UO_70 (O_70,N_9732,N_9717);
nor UO_71 (O_71,N_9757,N_9628);
and UO_72 (O_72,N_9525,N_9705);
and UO_73 (O_73,N_9610,N_9917);
or UO_74 (O_74,N_9671,N_9924);
or UO_75 (O_75,N_9731,N_9932);
nand UO_76 (O_76,N_9526,N_9820);
nor UO_77 (O_77,N_9913,N_9899);
nand UO_78 (O_78,N_9900,N_9996);
or UO_79 (O_79,N_9714,N_9684);
nor UO_80 (O_80,N_9543,N_9751);
nand UO_81 (O_81,N_9984,N_9665);
nor UO_82 (O_82,N_9745,N_9761);
xor UO_83 (O_83,N_9985,N_9804);
nand UO_84 (O_84,N_9968,N_9941);
nand UO_85 (O_85,N_9853,N_9871);
nand UO_86 (O_86,N_9973,N_9793);
or UO_87 (O_87,N_9822,N_9700);
xnor UO_88 (O_88,N_9607,N_9814);
or UO_89 (O_89,N_9789,N_9533);
nor UO_90 (O_90,N_9576,N_9639);
nor UO_91 (O_91,N_9621,N_9575);
nor UO_92 (O_92,N_9827,N_9509);
and UO_93 (O_93,N_9672,N_9906);
or UO_94 (O_94,N_9921,N_9617);
or UO_95 (O_95,N_9859,N_9582);
and UO_96 (O_96,N_9763,N_9528);
and UO_97 (O_97,N_9787,N_9508);
or UO_98 (O_98,N_9872,N_9635);
or UO_99 (O_99,N_9655,N_9517);
nor UO_100 (O_100,N_9938,N_9562);
and UO_101 (O_101,N_9530,N_9895);
and UO_102 (O_102,N_9704,N_9739);
xor UO_103 (O_103,N_9776,N_9896);
or UO_104 (O_104,N_9873,N_9534);
xnor UO_105 (O_105,N_9659,N_9572);
nand UO_106 (O_106,N_9679,N_9893);
or UO_107 (O_107,N_9541,N_9727);
xor UO_108 (O_108,N_9555,N_9546);
or UO_109 (O_109,N_9720,N_9614);
nand UO_110 (O_110,N_9584,N_9699);
xnor UO_111 (O_111,N_9750,N_9854);
and UO_112 (O_112,N_9840,N_9826);
xnor UO_113 (O_113,N_9624,N_9991);
nand UO_114 (O_114,N_9987,N_9755);
or UO_115 (O_115,N_9598,N_9792);
nand UO_116 (O_116,N_9979,N_9648);
and UO_117 (O_117,N_9529,N_9901);
nand UO_118 (O_118,N_9567,N_9885);
nand UO_119 (O_119,N_9828,N_9623);
or UO_120 (O_120,N_9746,N_9590);
or UO_121 (O_121,N_9850,N_9725);
nand UO_122 (O_122,N_9778,N_9929);
nand UO_123 (O_123,N_9910,N_9904);
or UO_124 (O_124,N_9664,N_9733);
nor UO_125 (O_125,N_9998,N_9796);
nor UO_126 (O_126,N_9835,N_9620);
and UO_127 (O_127,N_9608,N_9802);
and UO_128 (O_128,N_9510,N_9518);
and UO_129 (O_129,N_9633,N_9951);
and UO_130 (O_130,N_9504,N_9581);
nor UO_131 (O_131,N_9765,N_9817);
and UO_132 (O_132,N_9724,N_9995);
and UO_133 (O_133,N_9927,N_9782);
and UO_134 (O_134,N_9640,N_9762);
nor UO_135 (O_135,N_9551,N_9891);
and UO_136 (O_136,N_9975,N_9824);
and UO_137 (O_137,N_9589,N_9501);
nor UO_138 (O_138,N_9974,N_9579);
nand UO_139 (O_139,N_9668,N_9825);
nand UO_140 (O_140,N_9686,N_9626);
or UO_141 (O_141,N_9653,N_9813);
and UO_142 (O_142,N_9689,N_9863);
nor UO_143 (O_143,N_9953,N_9832);
or UO_144 (O_144,N_9911,N_9632);
nor UO_145 (O_145,N_9741,N_9630);
nand UO_146 (O_146,N_9516,N_9922);
nor UO_147 (O_147,N_9849,N_9808);
and UO_148 (O_148,N_9846,N_9673);
and UO_149 (O_149,N_9645,N_9947);
nor UO_150 (O_150,N_9845,N_9747);
xnor UO_151 (O_151,N_9881,N_9969);
nand UO_152 (O_152,N_9580,N_9961);
nand UO_153 (O_153,N_9616,N_9637);
and UO_154 (O_154,N_9934,N_9748);
and UO_155 (O_155,N_9933,N_9656);
nor UO_156 (O_156,N_9593,N_9962);
or UO_157 (O_157,N_9869,N_9527);
nor UO_158 (O_158,N_9545,N_9936);
nand UO_159 (O_159,N_9815,N_9694);
and UO_160 (O_160,N_9643,N_9627);
and UO_161 (O_161,N_9878,N_9683);
nor UO_162 (O_162,N_9994,N_9799);
and UO_163 (O_163,N_9783,N_9556);
nand UO_164 (O_164,N_9769,N_9950);
nor UO_165 (O_165,N_9886,N_9919);
and UO_166 (O_166,N_9554,N_9848);
or UO_167 (O_167,N_9549,N_9937);
nor UO_168 (O_168,N_9535,N_9930);
or UO_169 (O_169,N_9574,N_9522);
xnor UO_170 (O_170,N_9729,N_9795);
nor UO_171 (O_171,N_9818,N_9592);
nand UO_172 (O_172,N_9537,N_9597);
xnor UO_173 (O_173,N_9585,N_9945);
and UO_174 (O_174,N_9843,N_9752);
or UO_175 (O_175,N_9928,N_9903);
nor UO_176 (O_176,N_9523,N_9908);
nor UO_177 (O_177,N_9772,N_9966);
nor UO_178 (O_178,N_9810,N_9997);
and UO_179 (O_179,N_9819,N_9844);
or UO_180 (O_180,N_9876,N_9669);
nor UO_181 (O_181,N_9801,N_9548);
nand UO_182 (O_182,N_9662,N_9612);
nor UO_183 (O_183,N_9547,N_9740);
or UO_184 (O_184,N_9557,N_9559);
or UO_185 (O_185,N_9682,N_9681);
nand UO_186 (O_186,N_9707,N_9649);
and UO_187 (O_187,N_9887,N_9879);
nand UO_188 (O_188,N_9905,N_9542);
xor UO_189 (O_189,N_9657,N_9855);
and UO_190 (O_190,N_9931,N_9957);
nand UO_191 (O_191,N_9571,N_9760);
and UO_192 (O_192,N_9811,N_9712);
and UO_193 (O_193,N_9940,N_9701);
or UO_194 (O_194,N_9983,N_9999);
and UO_195 (O_195,N_9971,N_9976);
or UO_196 (O_196,N_9711,N_9862);
and UO_197 (O_197,N_9715,N_9703);
xnor UO_198 (O_198,N_9583,N_9564);
nand UO_199 (O_199,N_9902,N_9511);
or UO_200 (O_200,N_9641,N_9680);
and UO_201 (O_201,N_9874,N_9515);
nor UO_202 (O_202,N_9920,N_9867);
or UO_203 (O_203,N_9693,N_9888);
or UO_204 (O_204,N_9550,N_9803);
and UO_205 (O_205,N_9842,N_9709);
nor UO_206 (O_206,N_9531,N_9754);
and UO_207 (O_207,N_9944,N_9982);
xor UO_208 (O_208,N_9967,N_9514);
or UO_209 (O_209,N_9631,N_9697);
nand UO_210 (O_210,N_9606,N_9771);
nand UO_211 (O_211,N_9830,N_9909);
nor UO_212 (O_212,N_9780,N_9977);
nand UO_213 (O_213,N_9865,N_9685);
or UO_214 (O_214,N_9988,N_9960);
and UO_215 (O_215,N_9892,N_9609);
and UO_216 (O_216,N_9622,N_9544);
nand UO_217 (O_217,N_9868,N_9719);
nand UO_218 (O_218,N_9698,N_9647);
nor UO_219 (O_219,N_9836,N_9603);
or UO_220 (O_220,N_9744,N_9670);
and UO_221 (O_221,N_9784,N_9563);
xnor UO_222 (O_222,N_9794,N_9660);
or UO_223 (O_223,N_9889,N_9625);
nor UO_224 (O_224,N_9532,N_9706);
nor UO_225 (O_225,N_9552,N_9884);
nand UO_226 (O_226,N_9959,N_9956);
nand UO_227 (O_227,N_9831,N_9829);
nand UO_228 (O_228,N_9841,N_9972);
nor UO_229 (O_229,N_9838,N_9907);
or UO_230 (O_230,N_9539,N_9766);
and UO_231 (O_231,N_9605,N_9860);
nand UO_232 (O_232,N_9586,N_9993);
nand UO_233 (O_233,N_9566,N_9779);
nor UO_234 (O_234,N_9743,N_9970);
nor UO_235 (O_235,N_9767,N_9502);
or UO_236 (O_236,N_9667,N_9791);
nor UO_237 (O_237,N_9568,N_9839);
or UO_238 (O_238,N_9565,N_9591);
nand UO_239 (O_239,N_9890,N_9980);
and UO_240 (O_240,N_9661,N_9500);
xnor UO_241 (O_241,N_9837,N_9570);
and UO_242 (O_242,N_9915,N_9561);
nand UO_243 (O_243,N_9807,N_9611);
nand UO_244 (O_244,N_9857,N_9812);
nand UO_245 (O_245,N_9512,N_9710);
or UO_246 (O_246,N_9877,N_9786);
and UO_247 (O_247,N_9949,N_9805);
nor UO_248 (O_248,N_9723,N_9978);
nor UO_249 (O_249,N_9688,N_9587);
nand UO_250 (O_250,N_9580,N_9792);
nand UO_251 (O_251,N_9508,N_9629);
nor UO_252 (O_252,N_9527,N_9938);
xor UO_253 (O_253,N_9594,N_9884);
and UO_254 (O_254,N_9740,N_9888);
and UO_255 (O_255,N_9903,N_9924);
xnor UO_256 (O_256,N_9865,N_9959);
or UO_257 (O_257,N_9585,N_9524);
and UO_258 (O_258,N_9943,N_9859);
nand UO_259 (O_259,N_9691,N_9997);
or UO_260 (O_260,N_9674,N_9952);
or UO_261 (O_261,N_9560,N_9601);
nor UO_262 (O_262,N_9840,N_9646);
or UO_263 (O_263,N_9518,N_9852);
nor UO_264 (O_264,N_9785,N_9500);
xnor UO_265 (O_265,N_9646,N_9865);
and UO_266 (O_266,N_9620,N_9860);
xor UO_267 (O_267,N_9651,N_9968);
or UO_268 (O_268,N_9947,N_9928);
nor UO_269 (O_269,N_9874,N_9736);
or UO_270 (O_270,N_9658,N_9695);
or UO_271 (O_271,N_9737,N_9802);
xor UO_272 (O_272,N_9687,N_9603);
or UO_273 (O_273,N_9664,N_9946);
or UO_274 (O_274,N_9920,N_9727);
xnor UO_275 (O_275,N_9978,N_9709);
and UO_276 (O_276,N_9938,N_9720);
and UO_277 (O_277,N_9670,N_9608);
nor UO_278 (O_278,N_9546,N_9988);
nand UO_279 (O_279,N_9650,N_9603);
nand UO_280 (O_280,N_9852,N_9505);
nand UO_281 (O_281,N_9537,N_9703);
nand UO_282 (O_282,N_9792,N_9660);
nor UO_283 (O_283,N_9519,N_9767);
nor UO_284 (O_284,N_9897,N_9578);
and UO_285 (O_285,N_9590,N_9891);
and UO_286 (O_286,N_9700,N_9703);
and UO_287 (O_287,N_9634,N_9540);
nand UO_288 (O_288,N_9755,N_9650);
or UO_289 (O_289,N_9684,N_9529);
nor UO_290 (O_290,N_9817,N_9566);
nand UO_291 (O_291,N_9833,N_9849);
nor UO_292 (O_292,N_9990,N_9782);
nor UO_293 (O_293,N_9626,N_9801);
and UO_294 (O_294,N_9591,N_9880);
or UO_295 (O_295,N_9736,N_9888);
nor UO_296 (O_296,N_9999,N_9656);
nor UO_297 (O_297,N_9763,N_9735);
nor UO_298 (O_298,N_9874,N_9945);
or UO_299 (O_299,N_9817,N_9543);
nor UO_300 (O_300,N_9850,N_9590);
nor UO_301 (O_301,N_9541,N_9692);
and UO_302 (O_302,N_9502,N_9705);
or UO_303 (O_303,N_9973,N_9615);
xor UO_304 (O_304,N_9671,N_9898);
or UO_305 (O_305,N_9765,N_9912);
xnor UO_306 (O_306,N_9543,N_9564);
nand UO_307 (O_307,N_9743,N_9967);
xor UO_308 (O_308,N_9634,N_9733);
nor UO_309 (O_309,N_9668,N_9889);
nand UO_310 (O_310,N_9616,N_9765);
and UO_311 (O_311,N_9870,N_9825);
nand UO_312 (O_312,N_9553,N_9766);
xnor UO_313 (O_313,N_9615,N_9724);
nand UO_314 (O_314,N_9819,N_9875);
xor UO_315 (O_315,N_9950,N_9614);
and UO_316 (O_316,N_9921,N_9904);
nand UO_317 (O_317,N_9935,N_9616);
xor UO_318 (O_318,N_9976,N_9562);
nand UO_319 (O_319,N_9699,N_9803);
nand UO_320 (O_320,N_9982,N_9820);
and UO_321 (O_321,N_9603,N_9575);
nand UO_322 (O_322,N_9581,N_9798);
nand UO_323 (O_323,N_9983,N_9535);
nand UO_324 (O_324,N_9811,N_9573);
or UO_325 (O_325,N_9823,N_9506);
nor UO_326 (O_326,N_9881,N_9541);
and UO_327 (O_327,N_9978,N_9546);
or UO_328 (O_328,N_9661,N_9633);
nor UO_329 (O_329,N_9579,N_9926);
or UO_330 (O_330,N_9928,N_9753);
nand UO_331 (O_331,N_9934,N_9690);
and UO_332 (O_332,N_9939,N_9764);
nor UO_333 (O_333,N_9676,N_9528);
nand UO_334 (O_334,N_9554,N_9569);
and UO_335 (O_335,N_9708,N_9950);
and UO_336 (O_336,N_9509,N_9807);
nand UO_337 (O_337,N_9552,N_9587);
nor UO_338 (O_338,N_9912,N_9525);
or UO_339 (O_339,N_9880,N_9697);
xor UO_340 (O_340,N_9677,N_9573);
nor UO_341 (O_341,N_9637,N_9631);
nand UO_342 (O_342,N_9941,N_9987);
xnor UO_343 (O_343,N_9884,N_9783);
nor UO_344 (O_344,N_9764,N_9741);
xor UO_345 (O_345,N_9576,N_9571);
and UO_346 (O_346,N_9944,N_9805);
or UO_347 (O_347,N_9753,N_9782);
nand UO_348 (O_348,N_9850,N_9828);
and UO_349 (O_349,N_9992,N_9549);
nand UO_350 (O_350,N_9737,N_9647);
and UO_351 (O_351,N_9890,N_9807);
or UO_352 (O_352,N_9634,N_9557);
nand UO_353 (O_353,N_9506,N_9684);
xor UO_354 (O_354,N_9556,N_9903);
nor UO_355 (O_355,N_9524,N_9808);
and UO_356 (O_356,N_9550,N_9759);
or UO_357 (O_357,N_9718,N_9581);
nand UO_358 (O_358,N_9702,N_9874);
and UO_359 (O_359,N_9651,N_9563);
nand UO_360 (O_360,N_9942,N_9602);
nand UO_361 (O_361,N_9665,N_9668);
or UO_362 (O_362,N_9813,N_9693);
nor UO_363 (O_363,N_9979,N_9679);
or UO_364 (O_364,N_9961,N_9876);
and UO_365 (O_365,N_9900,N_9756);
xnor UO_366 (O_366,N_9639,N_9563);
nor UO_367 (O_367,N_9956,N_9921);
nor UO_368 (O_368,N_9816,N_9676);
nor UO_369 (O_369,N_9874,N_9537);
nand UO_370 (O_370,N_9826,N_9954);
nor UO_371 (O_371,N_9507,N_9536);
nor UO_372 (O_372,N_9993,N_9843);
and UO_373 (O_373,N_9692,N_9552);
nand UO_374 (O_374,N_9835,N_9654);
nor UO_375 (O_375,N_9504,N_9735);
and UO_376 (O_376,N_9598,N_9553);
or UO_377 (O_377,N_9869,N_9935);
nand UO_378 (O_378,N_9774,N_9909);
nand UO_379 (O_379,N_9601,N_9636);
and UO_380 (O_380,N_9919,N_9684);
or UO_381 (O_381,N_9752,N_9602);
and UO_382 (O_382,N_9684,N_9584);
nor UO_383 (O_383,N_9643,N_9820);
nor UO_384 (O_384,N_9897,N_9755);
or UO_385 (O_385,N_9841,N_9760);
or UO_386 (O_386,N_9756,N_9842);
xnor UO_387 (O_387,N_9877,N_9967);
and UO_388 (O_388,N_9852,N_9651);
and UO_389 (O_389,N_9924,N_9900);
and UO_390 (O_390,N_9699,N_9816);
or UO_391 (O_391,N_9561,N_9542);
or UO_392 (O_392,N_9733,N_9736);
nand UO_393 (O_393,N_9631,N_9732);
or UO_394 (O_394,N_9558,N_9996);
nor UO_395 (O_395,N_9639,N_9906);
nand UO_396 (O_396,N_9738,N_9847);
nor UO_397 (O_397,N_9996,N_9910);
nor UO_398 (O_398,N_9633,N_9997);
nor UO_399 (O_399,N_9764,N_9726);
nand UO_400 (O_400,N_9849,N_9688);
or UO_401 (O_401,N_9537,N_9673);
and UO_402 (O_402,N_9807,N_9765);
or UO_403 (O_403,N_9640,N_9876);
nand UO_404 (O_404,N_9952,N_9749);
nor UO_405 (O_405,N_9949,N_9536);
nand UO_406 (O_406,N_9699,N_9724);
nand UO_407 (O_407,N_9772,N_9919);
nor UO_408 (O_408,N_9586,N_9631);
nand UO_409 (O_409,N_9980,N_9663);
xnor UO_410 (O_410,N_9562,N_9748);
nor UO_411 (O_411,N_9600,N_9710);
or UO_412 (O_412,N_9846,N_9916);
and UO_413 (O_413,N_9516,N_9680);
or UO_414 (O_414,N_9749,N_9816);
nor UO_415 (O_415,N_9718,N_9789);
and UO_416 (O_416,N_9634,N_9629);
nor UO_417 (O_417,N_9704,N_9973);
or UO_418 (O_418,N_9580,N_9753);
or UO_419 (O_419,N_9887,N_9595);
and UO_420 (O_420,N_9611,N_9867);
xnor UO_421 (O_421,N_9678,N_9890);
nor UO_422 (O_422,N_9635,N_9550);
or UO_423 (O_423,N_9660,N_9520);
and UO_424 (O_424,N_9523,N_9796);
and UO_425 (O_425,N_9765,N_9963);
nor UO_426 (O_426,N_9523,N_9924);
nand UO_427 (O_427,N_9938,N_9534);
nor UO_428 (O_428,N_9729,N_9637);
nor UO_429 (O_429,N_9792,N_9870);
or UO_430 (O_430,N_9712,N_9603);
nor UO_431 (O_431,N_9597,N_9744);
or UO_432 (O_432,N_9529,N_9564);
nand UO_433 (O_433,N_9671,N_9674);
or UO_434 (O_434,N_9688,N_9623);
and UO_435 (O_435,N_9850,N_9561);
nand UO_436 (O_436,N_9676,N_9786);
nor UO_437 (O_437,N_9598,N_9502);
nor UO_438 (O_438,N_9635,N_9541);
nand UO_439 (O_439,N_9601,N_9924);
or UO_440 (O_440,N_9632,N_9719);
and UO_441 (O_441,N_9992,N_9697);
and UO_442 (O_442,N_9800,N_9548);
and UO_443 (O_443,N_9668,N_9902);
and UO_444 (O_444,N_9689,N_9796);
xnor UO_445 (O_445,N_9924,N_9514);
or UO_446 (O_446,N_9687,N_9989);
nand UO_447 (O_447,N_9538,N_9652);
or UO_448 (O_448,N_9618,N_9640);
nor UO_449 (O_449,N_9517,N_9979);
nand UO_450 (O_450,N_9989,N_9697);
xnor UO_451 (O_451,N_9941,N_9922);
or UO_452 (O_452,N_9804,N_9991);
nand UO_453 (O_453,N_9512,N_9644);
nand UO_454 (O_454,N_9818,N_9707);
and UO_455 (O_455,N_9579,N_9691);
nor UO_456 (O_456,N_9538,N_9645);
xnor UO_457 (O_457,N_9793,N_9913);
nand UO_458 (O_458,N_9674,N_9650);
or UO_459 (O_459,N_9880,N_9643);
and UO_460 (O_460,N_9991,N_9786);
and UO_461 (O_461,N_9772,N_9949);
nand UO_462 (O_462,N_9686,N_9815);
nor UO_463 (O_463,N_9674,N_9958);
and UO_464 (O_464,N_9563,N_9994);
nor UO_465 (O_465,N_9868,N_9675);
nor UO_466 (O_466,N_9976,N_9869);
or UO_467 (O_467,N_9890,N_9977);
nand UO_468 (O_468,N_9741,N_9607);
nand UO_469 (O_469,N_9905,N_9912);
and UO_470 (O_470,N_9777,N_9669);
or UO_471 (O_471,N_9571,N_9657);
nand UO_472 (O_472,N_9780,N_9572);
xor UO_473 (O_473,N_9961,N_9627);
nor UO_474 (O_474,N_9994,N_9820);
nand UO_475 (O_475,N_9530,N_9866);
nand UO_476 (O_476,N_9812,N_9952);
nand UO_477 (O_477,N_9837,N_9651);
and UO_478 (O_478,N_9713,N_9536);
nor UO_479 (O_479,N_9521,N_9765);
and UO_480 (O_480,N_9536,N_9819);
nor UO_481 (O_481,N_9677,N_9798);
nand UO_482 (O_482,N_9962,N_9552);
or UO_483 (O_483,N_9684,N_9634);
and UO_484 (O_484,N_9559,N_9931);
nand UO_485 (O_485,N_9966,N_9917);
nand UO_486 (O_486,N_9580,N_9938);
nor UO_487 (O_487,N_9529,N_9820);
nand UO_488 (O_488,N_9729,N_9960);
nand UO_489 (O_489,N_9984,N_9805);
and UO_490 (O_490,N_9639,N_9764);
nand UO_491 (O_491,N_9982,N_9712);
and UO_492 (O_492,N_9762,N_9562);
and UO_493 (O_493,N_9587,N_9511);
nor UO_494 (O_494,N_9844,N_9575);
and UO_495 (O_495,N_9840,N_9889);
nand UO_496 (O_496,N_9792,N_9505);
or UO_497 (O_497,N_9969,N_9882);
nand UO_498 (O_498,N_9956,N_9840);
nand UO_499 (O_499,N_9727,N_9995);
nor UO_500 (O_500,N_9789,N_9665);
nor UO_501 (O_501,N_9988,N_9936);
nand UO_502 (O_502,N_9590,N_9975);
or UO_503 (O_503,N_9788,N_9975);
and UO_504 (O_504,N_9998,N_9818);
or UO_505 (O_505,N_9915,N_9720);
nor UO_506 (O_506,N_9988,N_9836);
or UO_507 (O_507,N_9798,N_9800);
and UO_508 (O_508,N_9507,N_9732);
or UO_509 (O_509,N_9591,N_9950);
and UO_510 (O_510,N_9809,N_9938);
or UO_511 (O_511,N_9872,N_9660);
nand UO_512 (O_512,N_9838,N_9596);
nand UO_513 (O_513,N_9914,N_9939);
and UO_514 (O_514,N_9554,N_9517);
and UO_515 (O_515,N_9630,N_9904);
or UO_516 (O_516,N_9850,N_9720);
or UO_517 (O_517,N_9892,N_9698);
nor UO_518 (O_518,N_9813,N_9601);
nand UO_519 (O_519,N_9512,N_9770);
and UO_520 (O_520,N_9582,N_9938);
nand UO_521 (O_521,N_9961,N_9858);
or UO_522 (O_522,N_9723,N_9543);
and UO_523 (O_523,N_9660,N_9557);
nor UO_524 (O_524,N_9763,N_9750);
and UO_525 (O_525,N_9938,N_9553);
nand UO_526 (O_526,N_9915,N_9710);
or UO_527 (O_527,N_9600,N_9956);
nand UO_528 (O_528,N_9682,N_9708);
nor UO_529 (O_529,N_9571,N_9549);
and UO_530 (O_530,N_9786,N_9578);
xor UO_531 (O_531,N_9848,N_9815);
xnor UO_532 (O_532,N_9856,N_9503);
nand UO_533 (O_533,N_9590,N_9829);
nor UO_534 (O_534,N_9707,N_9704);
nand UO_535 (O_535,N_9720,N_9784);
and UO_536 (O_536,N_9817,N_9602);
nand UO_537 (O_537,N_9568,N_9586);
or UO_538 (O_538,N_9833,N_9767);
nor UO_539 (O_539,N_9514,N_9758);
nand UO_540 (O_540,N_9554,N_9633);
nand UO_541 (O_541,N_9791,N_9760);
and UO_542 (O_542,N_9770,N_9768);
nand UO_543 (O_543,N_9829,N_9571);
or UO_544 (O_544,N_9805,N_9923);
nor UO_545 (O_545,N_9669,N_9506);
or UO_546 (O_546,N_9645,N_9898);
nor UO_547 (O_547,N_9862,N_9800);
or UO_548 (O_548,N_9597,N_9677);
or UO_549 (O_549,N_9991,N_9923);
or UO_550 (O_550,N_9600,N_9581);
and UO_551 (O_551,N_9919,N_9604);
xnor UO_552 (O_552,N_9739,N_9904);
nor UO_553 (O_553,N_9527,N_9777);
nand UO_554 (O_554,N_9544,N_9550);
xor UO_555 (O_555,N_9818,N_9883);
nand UO_556 (O_556,N_9902,N_9784);
and UO_557 (O_557,N_9698,N_9957);
nand UO_558 (O_558,N_9659,N_9925);
and UO_559 (O_559,N_9966,N_9854);
xnor UO_560 (O_560,N_9539,N_9743);
or UO_561 (O_561,N_9607,N_9893);
or UO_562 (O_562,N_9846,N_9821);
nor UO_563 (O_563,N_9537,N_9814);
xnor UO_564 (O_564,N_9985,N_9740);
or UO_565 (O_565,N_9696,N_9530);
and UO_566 (O_566,N_9688,N_9780);
and UO_567 (O_567,N_9822,N_9726);
or UO_568 (O_568,N_9537,N_9644);
or UO_569 (O_569,N_9782,N_9969);
nand UO_570 (O_570,N_9789,N_9707);
nand UO_571 (O_571,N_9745,N_9755);
xnor UO_572 (O_572,N_9578,N_9763);
nand UO_573 (O_573,N_9720,N_9577);
nand UO_574 (O_574,N_9587,N_9797);
or UO_575 (O_575,N_9760,N_9620);
nand UO_576 (O_576,N_9551,N_9696);
nor UO_577 (O_577,N_9566,N_9717);
nor UO_578 (O_578,N_9997,N_9679);
nor UO_579 (O_579,N_9945,N_9914);
nand UO_580 (O_580,N_9895,N_9701);
nand UO_581 (O_581,N_9598,N_9809);
nor UO_582 (O_582,N_9556,N_9904);
or UO_583 (O_583,N_9578,N_9599);
nand UO_584 (O_584,N_9694,N_9762);
and UO_585 (O_585,N_9661,N_9742);
and UO_586 (O_586,N_9875,N_9665);
nand UO_587 (O_587,N_9890,N_9636);
or UO_588 (O_588,N_9904,N_9636);
and UO_589 (O_589,N_9651,N_9746);
nand UO_590 (O_590,N_9885,N_9792);
nor UO_591 (O_591,N_9909,N_9855);
or UO_592 (O_592,N_9574,N_9920);
nor UO_593 (O_593,N_9642,N_9555);
nor UO_594 (O_594,N_9719,N_9833);
and UO_595 (O_595,N_9541,N_9709);
or UO_596 (O_596,N_9916,N_9502);
nor UO_597 (O_597,N_9516,N_9539);
xor UO_598 (O_598,N_9826,N_9589);
xor UO_599 (O_599,N_9844,N_9715);
or UO_600 (O_600,N_9838,N_9712);
or UO_601 (O_601,N_9831,N_9855);
or UO_602 (O_602,N_9784,N_9726);
xor UO_603 (O_603,N_9667,N_9592);
or UO_604 (O_604,N_9811,N_9707);
and UO_605 (O_605,N_9842,N_9566);
nor UO_606 (O_606,N_9816,N_9640);
nand UO_607 (O_607,N_9812,N_9938);
nor UO_608 (O_608,N_9807,N_9575);
nor UO_609 (O_609,N_9918,N_9777);
nor UO_610 (O_610,N_9936,N_9770);
nand UO_611 (O_611,N_9620,N_9693);
or UO_612 (O_612,N_9500,N_9659);
or UO_613 (O_613,N_9807,N_9948);
xnor UO_614 (O_614,N_9595,N_9943);
nand UO_615 (O_615,N_9765,N_9655);
and UO_616 (O_616,N_9717,N_9844);
xor UO_617 (O_617,N_9638,N_9759);
nand UO_618 (O_618,N_9647,N_9988);
or UO_619 (O_619,N_9933,N_9546);
or UO_620 (O_620,N_9730,N_9913);
nand UO_621 (O_621,N_9742,N_9693);
nor UO_622 (O_622,N_9854,N_9853);
and UO_623 (O_623,N_9636,N_9618);
and UO_624 (O_624,N_9638,N_9772);
and UO_625 (O_625,N_9651,N_9762);
nand UO_626 (O_626,N_9604,N_9692);
and UO_627 (O_627,N_9734,N_9633);
or UO_628 (O_628,N_9749,N_9761);
xnor UO_629 (O_629,N_9525,N_9502);
nand UO_630 (O_630,N_9933,N_9523);
nand UO_631 (O_631,N_9800,N_9832);
or UO_632 (O_632,N_9985,N_9850);
nand UO_633 (O_633,N_9960,N_9520);
nor UO_634 (O_634,N_9956,N_9807);
xor UO_635 (O_635,N_9566,N_9536);
and UO_636 (O_636,N_9707,N_9653);
nand UO_637 (O_637,N_9742,N_9776);
nor UO_638 (O_638,N_9578,N_9916);
or UO_639 (O_639,N_9750,N_9848);
nor UO_640 (O_640,N_9815,N_9927);
and UO_641 (O_641,N_9827,N_9823);
xor UO_642 (O_642,N_9856,N_9936);
nor UO_643 (O_643,N_9668,N_9583);
or UO_644 (O_644,N_9541,N_9894);
nor UO_645 (O_645,N_9565,N_9699);
nand UO_646 (O_646,N_9879,N_9678);
nand UO_647 (O_647,N_9609,N_9902);
or UO_648 (O_648,N_9754,N_9654);
or UO_649 (O_649,N_9560,N_9544);
nor UO_650 (O_650,N_9982,N_9667);
and UO_651 (O_651,N_9792,N_9851);
xnor UO_652 (O_652,N_9988,N_9642);
nor UO_653 (O_653,N_9938,N_9551);
nand UO_654 (O_654,N_9655,N_9568);
xnor UO_655 (O_655,N_9539,N_9824);
and UO_656 (O_656,N_9689,N_9584);
nand UO_657 (O_657,N_9766,N_9667);
or UO_658 (O_658,N_9694,N_9657);
nand UO_659 (O_659,N_9704,N_9784);
nor UO_660 (O_660,N_9569,N_9771);
and UO_661 (O_661,N_9597,N_9709);
nor UO_662 (O_662,N_9693,N_9529);
nor UO_663 (O_663,N_9605,N_9697);
and UO_664 (O_664,N_9871,N_9741);
and UO_665 (O_665,N_9600,N_9514);
and UO_666 (O_666,N_9628,N_9855);
xnor UO_667 (O_667,N_9646,N_9557);
and UO_668 (O_668,N_9683,N_9719);
xnor UO_669 (O_669,N_9683,N_9692);
and UO_670 (O_670,N_9605,N_9515);
or UO_671 (O_671,N_9512,N_9731);
nand UO_672 (O_672,N_9768,N_9686);
and UO_673 (O_673,N_9890,N_9915);
nand UO_674 (O_674,N_9804,N_9590);
and UO_675 (O_675,N_9905,N_9522);
nand UO_676 (O_676,N_9972,N_9756);
nor UO_677 (O_677,N_9903,N_9670);
or UO_678 (O_678,N_9666,N_9993);
nand UO_679 (O_679,N_9936,N_9787);
nand UO_680 (O_680,N_9791,N_9552);
nand UO_681 (O_681,N_9533,N_9764);
xor UO_682 (O_682,N_9915,N_9788);
or UO_683 (O_683,N_9929,N_9504);
and UO_684 (O_684,N_9612,N_9764);
and UO_685 (O_685,N_9755,N_9791);
nand UO_686 (O_686,N_9859,N_9818);
or UO_687 (O_687,N_9806,N_9870);
or UO_688 (O_688,N_9646,N_9963);
and UO_689 (O_689,N_9909,N_9744);
xor UO_690 (O_690,N_9863,N_9676);
nor UO_691 (O_691,N_9612,N_9689);
nor UO_692 (O_692,N_9827,N_9714);
nand UO_693 (O_693,N_9810,N_9969);
or UO_694 (O_694,N_9943,N_9790);
nand UO_695 (O_695,N_9980,N_9692);
nand UO_696 (O_696,N_9577,N_9882);
nand UO_697 (O_697,N_9555,N_9680);
nor UO_698 (O_698,N_9876,N_9818);
and UO_699 (O_699,N_9876,N_9858);
xnor UO_700 (O_700,N_9972,N_9801);
xor UO_701 (O_701,N_9970,N_9609);
nor UO_702 (O_702,N_9997,N_9965);
and UO_703 (O_703,N_9639,N_9537);
nand UO_704 (O_704,N_9932,N_9971);
nor UO_705 (O_705,N_9564,N_9961);
and UO_706 (O_706,N_9567,N_9925);
nor UO_707 (O_707,N_9880,N_9859);
nand UO_708 (O_708,N_9952,N_9944);
and UO_709 (O_709,N_9704,N_9512);
nand UO_710 (O_710,N_9735,N_9600);
nor UO_711 (O_711,N_9808,N_9681);
xnor UO_712 (O_712,N_9910,N_9870);
xor UO_713 (O_713,N_9772,N_9876);
and UO_714 (O_714,N_9549,N_9865);
or UO_715 (O_715,N_9948,N_9882);
and UO_716 (O_716,N_9527,N_9982);
nand UO_717 (O_717,N_9524,N_9872);
nor UO_718 (O_718,N_9912,N_9838);
or UO_719 (O_719,N_9735,N_9754);
xor UO_720 (O_720,N_9925,N_9851);
nor UO_721 (O_721,N_9862,N_9827);
nor UO_722 (O_722,N_9834,N_9930);
or UO_723 (O_723,N_9793,N_9565);
nor UO_724 (O_724,N_9863,N_9964);
nor UO_725 (O_725,N_9746,N_9827);
nor UO_726 (O_726,N_9827,N_9986);
nand UO_727 (O_727,N_9521,N_9625);
nand UO_728 (O_728,N_9800,N_9781);
nor UO_729 (O_729,N_9583,N_9694);
nand UO_730 (O_730,N_9523,N_9558);
xor UO_731 (O_731,N_9915,N_9882);
and UO_732 (O_732,N_9658,N_9591);
and UO_733 (O_733,N_9524,N_9795);
nor UO_734 (O_734,N_9845,N_9848);
and UO_735 (O_735,N_9982,N_9932);
nand UO_736 (O_736,N_9959,N_9762);
nor UO_737 (O_737,N_9934,N_9618);
nand UO_738 (O_738,N_9891,N_9902);
and UO_739 (O_739,N_9618,N_9782);
and UO_740 (O_740,N_9556,N_9717);
or UO_741 (O_741,N_9758,N_9921);
nand UO_742 (O_742,N_9559,N_9674);
xor UO_743 (O_743,N_9987,N_9994);
and UO_744 (O_744,N_9953,N_9699);
and UO_745 (O_745,N_9715,N_9916);
nor UO_746 (O_746,N_9657,N_9919);
nor UO_747 (O_747,N_9947,N_9879);
or UO_748 (O_748,N_9634,N_9594);
nor UO_749 (O_749,N_9610,N_9527);
or UO_750 (O_750,N_9602,N_9793);
and UO_751 (O_751,N_9837,N_9967);
nor UO_752 (O_752,N_9877,N_9913);
or UO_753 (O_753,N_9895,N_9874);
and UO_754 (O_754,N_9631,N_9861);
nand UO_755 (O_755,N_9971,N_9680);
and UO_756 (O_756,N_9633,N_9568);
or UO_757 (O_757,N_9851,N_9596);
and UO_758 (O_758,N_9662,N_9706);
nand UO_759 (O_759,N_9774,N_9881);
and UO_760 (O_760,N_9902,N_9760);
or UO_761 (O_761,N_9668,N_9714);
and UO_762 (O_762,N_9667,N_9705);
nand UO_763 (O_763,N_9521,N_9856);
or UO_764 (O_764,N_9616,N_9982);
xor UO_765 (O_765,N_9929,N_9529);
or UO_766 (O_766,N_9657,N_9962);
and UO_767 (O_767,N_9565,N_9736);
nor UO_768 (O_768,N_9549,N_9851);
and UO_769 (O_769,N_9990,N_9815);
nor UO_770 (O_770,N_9953,N_9564);
nand UO_771 (O_771,N_9784,N_9941);
and UO_772 (O_772,N_9881,N_9903);
nand UO_773 (O_773,N_9552,N_9867);
and UO_774 (O_774,N_9999,N_9978);
nor UO_775 (O_775,N_9599,N_9509);
or UO_776 (O_776,N_9640,N_9842);
xnor UO_777 (O_777,N_9824,N_9699);
or UO_778 (O_778,N_9602,N_9686);
or UO_779 (O_779,N_9797,N_9582);
nand UO_780 (O_780,N_9680,N_9545);
nor UO_781 (O_781,N_9957,N_9994);
xnor UO_782 (O_782,N_9628,N_9533);
xor UO_783 (O_783,N_9996,N_9618);
or UO_784 (O_784,N_9682,N_9559);
or UO_785 (O_785,N_9760,N_9510);
nand UO_786 (O_786,N_9736,N_9926);
or UO_787 (O_787,N_9883,N_9771);
nand UO_788 (O_788,N_9946,N_9942);
and UO_789 (O_789,N_9805,N_9649);
or UO_790 (O_790,N_9659,N_9626);
xor UO_791 (O_791,N_9579,N_9673);
and UO_792 (O_792,N_9975,N_9760);
xor UO_793 (O_793,N_9824,N_9648);
or UO_794 (O_794,N_9977,N_9599);
nand UO_795 (O_795,N_9558,N_9734);
or UO_796 (O_796,N_9700,N_9569);
or UO_797 (O_797,N_9953,N_9694);
and UO_798 (O_798,N_9874,N_9609);
nand UO_799 (O_799,N_9509,N_9536);
or UO_800 (O_800,N_9666,N_9933);
or UO_801 (O_801,N_9558,N_9727);
and UO_802 (O_802,N_9897,N_9766);
and UO_803 (O_803,N_9677,N_9679);
nor UO_804 (O_804,N_9642,N_9818);
and UO_805 (O_805,N_9554,N_9990);
or UO_806 (O_806,N_9946,N_9779);
nand UO_807 (O_807,N_9859,N_9897);
and UO_808 (O_808,N_9575,N_9938);
and UO_809 (O_809,N_9945,N_9581);
or UO_810 (O_810,N_9687,N_9868);
nor UO_811 (O_811,N_9902,N_9959);
or UO_812 (O_812,N_9614,N_9547);
or UO_813 (O_813,N_9958,N_9972);
or UO_814 (O_814,N_9744,N_9854);
or UO_815 (O_815,N_9541,N_9982);
nand UO_816 (O_816,N_9646,N_9666);
nor UO_817 (O_817,N_9847,N_9777);
nand UO_818 (O_818,N_9984,N_9973);
xnor UO_819 (O_819,N_9604,N_9599);
or UO_820 (O_820,N_9985,N_9747);
and UO_821 (O_821,N_9970,N_9826);
and UO_822 (O_822,N_9870,N_9615);
nor UO_823 (O_823,N_9587,N_9703);
nand UO_824 (O_824,N_9756,N_9983);
xnor UO_825 (O_825,N_9533,N_9620);
nand UO_826 (O_826,N_9711,N_9544);
and UO_827 (O_827,N_9776,N_9667);
and UO_828 (O_828,N_9550,N_9586);
and UO_829 (O_829,N_9518,N_9823);
xor UO_830 (O_830,N_9503,N_9989);
and UO_831 (O_831,N_9557,N_9562);
xor UO_832 (O_832,N_9939,N_9748);
nor UO_833 (O_833,N_9578,N_9844);
nor UO_834 (O_834,N_9889,N_9500);
and UO_835 (O_835,N_9649,N_9968);
nand UO_836 (O_836,N_9952,N_9903);
nor UO_837 (O_837,N_9687,N_9611);
and UO_838 (O_838,N_9570,N_9848);
or UO_839 (O_839,N_9605,N_9910);
nor UO_840 (O_840,N_9867,N_9753);
or UO_841 (O_841,N_9545,N_9786);
and UO_842 (O_842,N_9580,N_9769);
xnor UO_843 (O_843,N_9742,N_9851);
or UO_844 (O_844,N_9693,N_9988);
nor UO_845 (O_845,N_9772,N_9503);
nand UO_846 (O_846,N_9673,N_9826);
and UO_847 (O_847,N_9748,N_9570);
xor UO_848 (O_848,N_9993,N_9587);
or UO_849 (O_849,N_9562,N_9626);
or UO_850 (O_850,N_9790,N_9692);
nand UO_851 (O_851,N_9814,N_9544);
or UO_852 (O_852,N_9551,N_9576);
nor UO_853 (O_853,N_9620,N_9689);
nand UO_854 (O_854,N_9546,N_9788);
nor UO_855 (O_855,N_9830,N_9531);
xnor UO_856 (O_856,N_9845,N_9741);
or UO_857 (O_857,N_9623,N_9820);
and UO_858 (O_858,N_9579,N_9829);
nand UO_859 (O_859,N_9950,N_9735);
and UO_860 (O_860,N_9672,N_9961);
or UO_861 (O_861,N_9804,N_9951);
and UO_862 (O_862,N_9993,N_9782);
or UO_863 (O_863,N_9594,N_9506);
nand UO_864 (O_864,N_9905,N_9788);
and UO_865 (O_865,N_9635,N_9525);
and UO_866 (O_866,N_9891,N_9898);
xnor UO_867 (O_867,N_9537,N_9865);
nand UO_868 (O_868,N_9614,N_9647);
and UO_869 (O_869,N_9679,N_9675);
nand UO_870 (O_870,N_9725,N_9715);
and UO_871 (O_871,N_9723,N_9561);
nor UO_872 (O_872,N_9689,N_9506);
nand UO_873 (O_873,N_9733,N_9972);
and UO_874 (O_874,N_9953,N_9884);
nand UO_875 (O_875,N_9630,N_9918);
nor UO_876 (O_876,N_9765,N_9781);
nand UO_877 (O_877,N_9552,N_9974);
nor UO_878 (O_878,N_9738,N_9880);
nor UO_879 (O_879,N_9721,N_9869);
or UO_880 (O_880,N_9515,N_9655);
and UO_881 (O_881,N_9982,N_9887);
nor UO_882 (O_882,N_9747,N_9852);
nand UO_883 (O_883,N_9510,N_9959);
nor UO_884 (O_884,N_9613,N_9567);
xnor UO_885 (O_885,N_9598,N_9802);
nand UO_886 (O_886,N_9969,N_9857);
nor UO_887 (O_887,N_9846,N_9503);
nand UO_888 (O_888,N_9554,N_9741);
nand UO_889 (O_889,N_9664,N_9529);
nor UO_890 (O_890,N_9990,N_9544);
and UO_891 (O_891,N_9696,N_9549);
or UO_892 (O_892,N_9513,N_9801);
and UO_893 (O_893,N_9743,N_9535);
or UO_894 (O_894,N_9705,N_9845);
or UO_895 (O_895,N_9609,N_9840);
and UO_896 (O_896,N_9697,N_9996);
nor UO_897 (O_897,N_9823,N_9979);
xor UO_898 (O_898,N_9981,N_9883);
and UO_899 (O_899,N_9519,N_9619);
nor UO_900 (O_900,N_9610,N_9924);
or UO_901 (O_901,N_9813,N_9735);
and UO_902 (O_902,N_9754,N_9527);
nand UO_903 (O_903,N_9992,N_9956);
xor UO_904 (O_904,N_9786,N_9815);
or UO_905 (O_905,N_9511,N_9940);
nor UO_906 (O_906,N_9813,N_9622);
nand UO_907 (O_907,N_9870,N_9805);
or UO_908 (O_908,N_9996,N_9908);
nor UO_909 (O_909,N_9679,N_9734);
xnor UO_910 (O_910,N_9716,N_9707);
and UO_911 (O_911,N_9922,N_9697);
nand UO_912 (O_912,N_9522,N_9908);
or UO_913 (O_913,N_9958,N_9635);
or UO_914 (O_914,N_9990,N_9789);
nand UO_915 (O_915,N_9570,N_9511);
xnor UO_916 (O_916,N_9934,N_9593);
and UO_917 (O_917,N_9582,N_9887);
nand UO_918 (O_918,N_9561,N_9801);
nand UO_919 (O_919,N_9797,N_9717);
and UO_920 (O_920,N_9848,N_9715);
nand UO_921 (O_921,N_9954,N_9832);
and UO_922 (O_922,N_9920,N_9530);
or UO_923 (O_923,N_9545,N_9730);
nor UO_924 (O_924,N_9694,N_9549);
or UO_925 (O_925,N_9757,N_9968);
xor UO_926 (O_926,N_9569,N_9893);
or UO_927 (O_927,N_9956,N_9649);
nand UO_928 (O_928,N_9934,N_9631);
or UO_929 (O_929,N_9526,N_9601);
nor UO_930 (O_930,N_9968,N_9673);
and UO_931 (O_931,N_9540,N_9524);
or UO_932 (O_932,N_9741,N_9603);
nand UO_933 (O_933,N_9742,N_9927);
and UO_934 (O_934,N_9505,N_9594);
xnor UO_935 (O_935,N_9881,N_9990);
or UO_936 (O_936,N_9503,N_9512);
nand UO_937 (O_937,N_9752,N_9716);
nand UO_938 (O_938,N_9756,N_9720);
nand UO_939 (O_939,N_9527,N_9925);
or UO_940 (O_940,N_9621,N_9928);
xor UO_941 (O_941,N_9955,N_9749);
and UO_942 (O_942,N_9842,N_9504);
or UO_943 (O_943,N_9531,N_9953);
nor UO_944 (O_944,N_9956,N_9847);
nand UO_945 (O_945,N_9642,N_9937);
nor UO_946 (O_946,N_9810,N_9521);
and UO_947 (O_947,N_9846,N_9777);
nand UO_948 (O_948,N_9776,N_9904);
nand UO_949 (O_949,N_9775,N_9539);
nand UO_950 (O_950,N_9797,N_9563);
and UO_951 (O_951,N_9944,N_9832);
nand UO_952 (O_952,N_9827,N_9589);
and UO_953 (O_953,N_9997,N_9745);
xnor UO_954 (O_954,N_9917,N_9579);
nand UO_955 (O_955,N_9998,N_9903);
or UO_956 (O_956,N_9871,N_9860);
and UO_957 (O_957,N_9898,N_9692);
nand UO_958 (O_958,N_9535,N_9826);
or UO_959 (O_959,N_9931,N_9517);
xor UO_960 (O_960,N_9568,N_9604);
or UO_961 (O_961,N_9709,N_9974);
and UO_962 (O_962,N_9543,N_9567);
nor UO_963 (O_963,N_9927,N_9981);
nor UO_964 (O_964,N_9593,N_9900);
nand UO_965 (O_965,N_9686,N_9996);
and UO_966 (O_966,N_9759,N_9586);
nor UO_967 (O_967,N_9608,N_9937);
nor UO_968 (O_968,N_9902,N_9909);
or UO_969 (O_969,N_9875,N_9870);
and UO_970 (O_970,N_9874,N_9892);
nor UO_971 (O_971,N_9522,N_9625);
nand UO_972 (O_972,N_9811,N_9737);
and UO_973 (O_973,N_9593,N_9681);
nor UO_974 (O_974,N_9814,N_9806);
and UO_975 (O_975,N_9755,N_9812);
nand UO_976 (O_976,N_9929,N_9604);
xnor UO_977 (O_977,N_9527,N_9965);
nor UO_978 (O_978,N_9671,N_9774);
nor UO_979 (O_979,N_9985,N_9913);
and UO_980 (O_980,N_9845,N_9988);
nand UO_981 (O_981,N_9932,N_9760);
or UO_982 (O_982,N_9704,N_9940);
nand UO_983 (O_983,N_9929,N_9530);
nor UO_984 (O_984,N_9792,N_9760);
or UO_985 (O_985,N_9877,N_9928);
nor UO_986 (O_986,N_9538,N_9814);
nor UO_987 (O_987,N_9591,N_9613);
nand UO_988 (O_988,N_9959,N_9625);
or UO_989 (O_989,N_9611,N_9662);
nor UO_990 (O_990,N_9687,N_9948);
nand UO_991 (O_991,N_9798,N_9671);
and UO_992 (O_992,N_9624,N_9576);
or UO_993 (O_993,N_9611,N_9587);
nand UO_994 (O_994,N_9517,N_9977);
nor UO_995 (O_995,N_9518,N_9906);
and UO_996 (O_996,N_9786,N_9971);
xnor UO_997 (O_997,N_9797,N_9610);
or UO_998 (O_998,N_9500,N_9980);
and UO_999 (O_999,N_9914,N_9643);
and UO_1000 (O_1000,N_9869,N_9785);
nand UO_1001 (O_1001,N_9525,N_9748);
or UO_1002 (O_1002,N_9813,N_9938);
or UO_1003 (O_1003,N_9589,N_9742);
xor UO_1004 (O_1004,N_9797,N_9753);
or UO_1005 (O_1005,N_9937,N_9657);
or UO_1006 (O_1006,N_9985,N_9853);
xnor UO_1007 (O_1007,N_9719,N_9802);
nand UO_1008 (O_1008,N_9863,N_9835);
nor UO_1009 (O_1009,N_9813,N_9990);
and UO_1010 (O_1010,N_9906,N_9965);
and UO_1011 (O_1011,N_9733,N_9536);
nand UO_1012 (O_1012,N_9609,N_9740);
nor UO_1013 (O_1013,N_9905,N_9690);
nor UO_1014 (O_1014,N_9874,N_9953);
or UO_1015 (O_1015,N_9862,N_9730);
nor UO_1016 (O_1016,N_9974,N_9567);
or UO_1017 (O_1017,N_9717,N_9571);
and UO_1018 (O_1018,N_9578,N_9737);
and UO_1019 (O_1019,N_9686,N_9862);
or UO_1020 (O_1020,N_9753,N_9704);
nor UO_1021 (O_1021,N_9958,N_9670);
nand UO_1022 (O_1022,N_9800,N_9769);
nand UO_1023 (O_1023,N_9844,N_9671);
nand UO_1024 (O_1024,N_9806,N_9699);
xnor UO_1025 (O_1025,N_9793,N_9681);
nor UO_1026 (O_1026,N_9688,N_9701);
xnor UO_1027 (O_1027,N_9787,N_9563);
nor UO_1028 (O_1028,N_9636,N_9611);
xor UO_1029 (O_1029,N_9674,N_9835);
nor UO_1030 (O_1030,N_9961,N_9928);
and UO_1031 (O_1031,N_9514,N_9869);
nor UO_1032 (O_1032,N_9873,N_9613);
nor UO_1033 (O_1033,N_9948,N_9776);
nand UO_1034 (O_1034,N_9568,N_9557);
and UO_1035 (O_1035,N_9811,N_9823);
and UO_1036 (O_1036,N_9651,N_9867);
and UO_1037 (O_1037,N_9537,N_9851);
nor UO_1038 (O_1038,N_9506,N_9648);
nor UO_1039 (O_1039,N_9854,N_9701);
nand UO_1040 (O_1040,N_9936,N_9719);
or UO_1041 (O_1041,N_9806,N_9731);
and UO_1042 (O_1042,N_9867,N_9838);
nor UO_1043 (O_1043,N_9809,N_9737);
nor UO_1044 (O_1044,N_9955,N_9826);
and UO_1045 (O_1045,N_9788,N_9801);
xnor UO_1046 (O_1046,N_9621,N_9601);
or UO_1047 (O_1047,N_9526,N_9980);
and UO_1048 (O_1048,N_9686,N_9901);
or UO_1049 (O_1049,N_9629,N_9626);
nor UO_1050 (O_1050,N_9608,N_9847);
nor UO_1051 (O_1051,N_9977,N_9953);
nor UO_1052 (O_1052,N_9895,N_9841);
nor UO_1053 (O_1053,N_9959,N_9991);
nor UO_1054 (O_1054,N_9785,N_9595);
nor UO_1055 (O_1055,N_9890,N_9715);
nand UO_1056 (O_1056,N_9797,N_9611);
xnor UO_1057 (O_1057,N_9657,N_9774);
or UO_1058 (O_1058,N_9736,N_9930);
nand UO_1059 (O_1059,N_9701,N_9982);
nand UO_1060 (O_1060,N_9745,N_9513);
nor UO_1061 (O_1061,N_9988,N_9886);
and UO_1062 (O_1062,N_9949,N_9595);
or UO_1063 (O_1063,N_9882,N_9820);
nand UO_1064 (O_1064,N_9890,N_9991);
nand UO_1065 (O_1065,N_9939,N_9741);
and UO_1066 (O_1066,N_9868,N_9505);
nand UO_1067 (O_1067,N_9534,N_9995);
nor UO_1068 (O_1068,N_9854,N_9755);
nor UO_1069 (O_1069,N_9948,N_9850);
nand UO_1070 (O_1070,N_9957,N_9521);
or UO_1071 (O_1071,N_9532,N_9967);
nor UO_1072 (O_1072,N_9848,N_9844);
and UO_1073 (O_1073,N_9878,N_9897);
nand UO_1074 (O_1074,N_9575,N_9602);
nand UO_1075 (O_1075,N_9740,N_9522);
or UO_1076 (O_1076,N_9957,N_9742);
and UO_1077 (O_1077,N_9544,N_9539);
nand UO_1078 (O_1078,N_9791,N_9863);
or UO_1079 (O_1079,N_9712,N_9920);
xnor UO_1080 (O_1080,N_9627,N_9635);
or UO_1081 (O_1081,N_9915,N_9682);
xnor UO_1082 (O_1082,N_9609,N_9851);
and UO_1083 (O_1083,N_9888,N_9979);
and UO_1084 (O_1084,N_9594,N_9626);
nand UO_1085 (O_1085,N_9814,N_9736);
nand UO_1086 (O_1086,N_9820,N_9743);
nand UO_1087 (O_1087,N_9656,N_9664);
nand UO_1088 (O_1088,N_9939,N_9713);
and UO_1089 (O_1089,N_9977,N_9706);
or UO_1090 (O_1090,N_9699,N_9548);
and UO_1091 (O_1091,N_9645,N_9570);
nor UO_1092 (O_1092,N_9551,N_9769);
nand UO_1093 (O_1093,N_9885,N_9983);
or UO_1094 (O_1094,N_9670,N_9717);
nand UO_1095 (O_1095,N_9790,N_9836);
and UO_1096 (O_1096,N_9834,N_9820);
and UO_1097 (O_1097,N_9834,N_9945);
or UO_1098 (O_1098,N_9830,N_9839);
and UO_1099 (O_1099,N_9759,N_9804);
nor UO_1100 (O_1100,N_9618,N_9916);
and UO_1101 (O_1101,N_9614,N_9680);
nand UO_1102 (O_1102,N_9782,N_9615);
nand UO_1103 (O_1103,N_9904,N_9860);
xor UO_1104 (O_1104,N_9894,N_9652);
or UO_1105 (O_1105,N_9977,N_9685);
and UO_1106 (O_1106,N_9903,N_9849);
xor UO_1107 (O_1107,N_9720,N_9695);
and UO_1108 (O_1108,N_9803,N_9514);
or UO_1109 (O_1109,N_9534,N_9867);
or UO_1110 (O_1110,N_9692,N_9767);
nand UO_1111 (O_1111,N_9934,N_9851);
nand UO_1112 (O_1112,N_9895,N_9807);
nor UO_1113 (O_1113,N_9789,N_9586);
nand UO_1114 (O_1114,N_9827,N_9572);
xnor UO_1115 (O_1115,N_9636,N_9596);
and UO_1116 (O_1116,N_9511,N_9694);
or UO_1117 (O_1117,N_9689,N_9631);
or UO_1118 (O_1118,N_9820,N_9749);
and UO_1119 (O_1119,N_9830,N_9738);
or UO_1120 (O_1120,N_9542,N_9776);
nand UO_1121 (O_1121,N_9703,N_9741);
nor UO_1122 (O_1122,N_9910,N_9926);
or UO_1123 (O_1123,N_9891,N_9932);
xor UO_1124 (O_1124,N_9820,N_9906);
xor UO_1125 (O_1125,N_9745,N_9822);
or UO_1126 (O_1126,N_9551,N_9559);
and UO_1127 (O_1127,N_9908,N_9639);
or UO_1128 (O_1128,N_9588,N_9850);
and UO_1129 (O_1129,N_9830,N_9686);
nor UO_1130 (O_1130,N_9753,N_9653);
or UO_1131 (O_1131,N_9818,N_9760);
or UO_1132 (O_1132,N_9951,N_9517);
and UO_1133 (O_1133,N_9552,N_9680);
nor UO_1134 (O_1134,N_9661,N_9673);
xor UO_1135 (O_1135,N_9530,N_9584);
nor UO_1136 (O_1136,N_9771,N_9554);
nand UO_1137 (O_1137,N_9702,N_9586);
nor UO_1138 (O_1138,N_9804,N_9953);
xnor UO_1139 (O_1139,N_9575,N_9842);
and UO_1140 (O_1140,N_9737,N_9774);
or UO_1141 (O_1141,N_9955,N_9630);
xnor UO_1142 (O_1142,N_9681,N_9712);
xnor UO_1143 (O_1143,N_9947,N_9566);
and UO_1144 (O_1144,N_9839,N_9869);
and UO_1145 (O_1145,N_9946,N_9829);
or UO_1146 (O_1146,N_9933,N_9908);
or UO_1147 (O_1147,N_9610,N_9656);
nor UO_1148 (O_1148,N_9645,N_9607);
or UO_1149 (O_1149,N_9603,N_9916);
and UO_1150 (O_1150,N_9883,N_9802);
nand UO_1151 (O_1151,N_9925,N_9640);
nand UO_1152 (O_1152,N_9913,N_9706);
nor UO_1153 (O_1153,N_9531,N_9743);
xor UO_1154 (O_1154,N_9973,N_9541);
nand UO_1155 (O_1155,N_9701,N_9740);
or UO_1156 (O_1156,N_9772,N_9932);
and UO_1157 (O_1157,N_9722,N_9891);
or UO_1158 (O_1158,N_9567,N_9832);
and UO_1159 (O_1159,N_9666,N_9667);
nor UO_1160 (O_1160,N_9702,N_9895);
nand UO_1161 (O_1161,N_9962,N_9524);
xnor UO_1162 (O_1162,N_9952,N_9748);
and UO_1163 (O_1163,N_9814,N_9726);
or UO_1164 (O_1164,N_9772,N_9827);
and UO_1165 (O_1165,N_9722,N_9836);
or UO_1166 (O_1166,N_9831,N_9974);
or UO_1167 (O_1167,N_9636,N_9875);
and UO_1168 (O_1168,N_9589,N_9949);
nand UO_1169 (O_1169,N_9972,N_9630);
xor UO_1170 (O_1170,N_9725,N_9726);
nor UO_1171 (O_1171,N_9652,N_9571);
nand UO_1172 (O_1172,N_9536,N_9825);
nor UO_1173 (O_1173,N_9839,N_9712);
nand UO_1174 (O_1174,N_9709,N_9786);
nand UO_1175 (O_1175,N_9629,N_9984);
nor UO_1176 (O_1176,N_9555,N_9969);
nand UO_1177 (O_1177,N_9839,N_9780);
nand UO_1178 (O_1178,N_9918,N_9553);
nor UO_1179 (O_1179,N_9730,N_9541);
or UO_1180 (O_1180,N_9969,N_9961);
or UO_1181 (O_1181,N_9838,N_9776);
nand UO_1182 (O_1182,N_9635,N_9924);
nor UO_1183 (O_1183,N_9532,N_9675);
nor UO_1184 (O_1184,N_9611,N_9574);
nor UO_1185 (O_1185,N_9710,N_9648);
xnor UO_1186 (O_1186,N_9757,N_9865);
and UO_1187 (O_1187,N_9862,N_9660);
nand UO_1188 (O_1188,N_9545,N_9892);
and UO_1189 (O_1189,N_9527,N_9930);
xor UO_1190 (O_1190,N_9641,N_9787);
nand UO_1191 (O_1191,N_9661,N_9639);
xor UO_1192 (O_1192,N_9872,N_9621);
or UO_1193 (O_1193,N_9994,N_9871);
nand UO_1194 (O_1194,N_9874,N_9844);
and UO_1195 (O_1195,N_9947,N_9773);
and UO_1196 (O_1196,N_9992,N_9706);
nand UO_1197 (O_1197,N_9527,N_9595);
and UO_1198 (O_1198,N_9589,N_9722);
nor UO_1199 (O_1199,N_9803,N_9671);
xnor UO_1200 (O_1200,N_9925,N_9829);
nand UO_1201 (O_1201,N_9549,N_9631);
nand UO_1202 (O_1202,N_9640,N_9949);
nor UO_1203 (O_1203,N_9643,N_9989);
and UO_1204 (O_1204,N_9863,N_9741);
nand UO_1205 (O_1205,N_9764,N_9813);
or UO_1206 (O_1206,N_9557,N_9812);
and UO_1207 (O_1207,N_9798,N_9730);
nor UO_1208 (O_1208,N_9601,N_9656);
xnor UO_1209 (O_1209,N_9739,N_9567);
or UO_1210 (O_1210,N_9557,N_9608);
and UO_1211 (O_1211,N_9975,N_9671);
nand UO_1212 (O_1212,N_9799,N_9610);
nor UO_1213 (O_1213,N_9550,N_9578);
nor UO_1214 (O_1214,N_9542,N_9721);
nand UO_1215 (O_1215,N_9751,N_9517);
nor UO_1216 (O_1216,N_9553,N_9948);
nand UO_1217 (O_1217,N_9799,N_9922);
or UO_1218 (O_1218,N_9748,N_9699);
nor UO_1219 (O_1219,N_9825,N_9666);
or UO_1220 (O_1220,N_9744,N_9607);
and UO_1221 (O_1221,N_9631,N_9834);
and UO_1222 (O_1222,N_9991,N_9879);
and UO_1223 (O_1223,N_9541,N_9923);
or UO_1224 (O_1224,N_9642,N_9752);
or UO_1225 (O_1225,N_9556,N_9706);
nand UO_1226 (O_1226,N_9562,N_9830);
xnor UO_1227 (O_1227,N_9850,N_9741);
xor UO_1228 (O_1228,N_9604,N_9909);
or UO_1229 (O_1229,N_9643,N_9692);
nor UO_1230 (O_1230,N_9979,N_9632);
nand UO_1231 (O_1231,N_9818,N_9567);
and UO_1232 (O_1232,N_9726,N_9910);
nor UO_1233 (O_1233,N_9907,N_9878);
or UO_1234 (O_1234,N_9635,N_9912);
and UO_1235 (O_1235,N_9683,N_9646);
or UO_1236 (O_1236,N_9599,N_9737);
nand UO_1237 (O_1237,N_9815,N_9814);
nand UO_1238 (O_1238,N_9640,N_9516);
or UO_1239 (O_1239,N_9646,N_9700);
xor UO_1240 (O_1240,N_9869,N_9532);
nor UO_1241 (O_1241,N_9551,N_9647);
and UO_1242 (O_1242,N_9980,N_9934);
nand UO_1243 (O_1243,N_9724,N_9656);
nor UO_1244 (O_1244,N_9667,N_9656);
and UO_1245 (O_1245,N_9827,N_9608);
or UO_1246 (O_1246,N_9593,N_9945);
nor UO_1247 (O_1247,N_9844,N_9958);
and UO_1248 (O_1248,N_9743,N_9951);
nor UO_1249 (O_1249,N_9640,N_9955);
nand UO_1250 (O_1250,N_9720,N_9889);
nand UO_1251 (O_1251,N_9679,N_9973);
nor UO_1252 (O_1252,N_9577,N_9719);
nor UO_1253 (O_1253,N_9800,N_9529);
nand UO_1254 (O_1254,N_9693,N_9548);
nor UO_1255 (O_1255,N_9739,N_9657);
or UO_1256 (O_1256,N_9526,N_9806);
and UO_1257 (O_1257,N_9694,N_9814);
and UO_1258 (O_1258,N_9986,N_9864);
and UO_1259 (O_1259,N_9516,N_9653);
or UO_1260 (O_1260,N_9672,N_9849);
nor UO_1261 (O_1261,N_9842,N_9571);
or UO_1262 (O_1262,N_9727,N_9988);
and UO_1263 (O_1263,N_9775,N_9679);
nand UO_1264 (O_1264,N_9741,N_9689);
xor UO_1265 (O_1265,N_9791,N_9622);
and UO_1266 (O_1266,N_9721,N_9953);
nor UO_1267 (O_1267,N_9728,N_9913);
or UO_1268 (O_1268,N_9875,N_9592);
nand UO_1269 (O_1269,N_9685,N_9764);
nand UO_1270 (O_1270,N_9773,N_9819);
and UO_1271 (O_1271,N_9657,N_9643);
nor UO_1272 (O_1272,N_9690,N_9632);
nand UO_1273 (O_1273,N_9821,N_9908);
and UO_1274 (O_1274,N_9636,N_9546);
and UO_1275 (O_1275,N_9536,N_9739);
or UO_1276 (O_1276,N_9697,N_9868);
or UO_1277 (O_1277,N_9559,N_9807);
nand UO_1278 (O_1278,N_9765,N_9589);
xnor UO_1279 (O_1279,N_9846,N_9568);
nor UO_1280 (O_1280,N_9880,N_9622);
or UO_1281 (O_1281,N_9763,N_9806);
nor UO_1282 (O_1282,N_9726,N_9667);
nand UO_1283 (O_1283,N_9817,N_9943);
nor UO_1284 (O_1284,N_9599,N_9827);
and UO_1285 (O_1285,N_9675,N_9518);
nor UO_1286 (O_1286,N_9813,N_9529);
and UO_1287 (O_1287,N_9751,N_9682);
nor UO_1288 (O_1288,N_9715,N_9884);
nand UO_1289 (O_1289,N_9896,N_9786);
and UO_1290 (O_1290,N_9997,N_9945);
or UO_1291 (O_1291,N_9775,N_9924);
nor UO_1292 (O_1292,N_9844,N_9905);
nor UO_1293 (O_1293,N_9878,N_9708);
nor UO_1294 (O_1294,N_9840,N_9891);
nor UO_1295 (O_1295,N_9980,N_9621);
or UO_1296 (O_1296,N_9754,N_9551);
nor UO_1297 (O_1297,N_9869,N_9696);
and UO_1298 (O_1298,N_9671,N_9813);
nor UO_1299 (O_1299,N_9982,N_9846);
xnor UO_1300 (O_1300,N_9912,N_9601);
and UO_1301 (O_1301,N_9654,N_9778);
nor UO_1302 (O_1302,N_9893,N_9568);
or UO_1303 (O_1303,N_9953,N_9800);
nand UO_1304 (O_1304,N_9683,N_9998);
and UO_1305 (O_1305,N_9566,N_9772);
or UO_1306 (O_1306,N_9746,N_9616);
and UO_1307 (O_1307,N_9693,N_9596);
or UO_1308 (O_1308,N_9734,N_9818);
and UO_1309 (O_1309,N_9503,N_9750);
nor UO_1310 (O_1310,N_9824,N_9767);
nand UO_1311 (O_1311,N_9508,N_9522);
and UO_1312 (O_1312,N_9539,N_9918);
nand UO_1313 (O_1313,N_9560,N_9905);
and UO_1314 (O_1314,N_9818,N_9800);
nor UO_1315 (O_1315,N_9999,N_9904);
nor UO_1316 (O_1316,N_9683,N_9909);
nor UO_1317 (O_1317,N_9614,N_9501);
nand UO_1318 (O_1318,N_9665,N_9903);
xnor UO_1319 (O_1319,N_9841,N_9723);
or UO_1320 (O_1320,N_9791,N_9794);
nand UO_1321 (O_1321,N_9704,N_9909);
nand UO_1322 (O_1322,N_9926,N_9845);
nand UO_1323 (O_1323,N_9951,N_9704);
nor UO_1324 (O_1324,N_9726,N_9666);
nand UO_1325 (O_1325,N_9580,N_9904);
nor UO_1326 (O_1326,N_9911,N_9635);
nand UO_1327 (O_1327,N_9694,N_9940);
nor UO_1328 (O_1328,N_9521,N_9790);
nand UO_1329 (O_1329,N_9958,N_9520);
and UO_1330 (O_1330,N_9902,N_9716);
and UO_1331 (O_1331,N_9982,N_9719);
xnor UO_1332 (O_1332,N_9637,N_9861);
and UO_1333 (O_1333,N_9788,N_9860);
xnor UO_1334 (O_1334,N_9501,N_9686);
or UO_1335 (O_1335,N_9877,N_9937);
or UO_1336 (O_1336,N_9700,N_9594);
xnor UO_1337 (O_1337,N_9720,N_9885);
and UO_1338 (O_1338,N_9854,N_9535);
nor UO_1339 (O_1339,N_9897,N_9780);
and UO_1340 (O_1340,N_9507,N_9940);
xnor UO_1341 (O_1341,N_9901,N_9728);
xnor UO_1342 (O_1342,N_9791,N_9541);
or UO_1343 (O_1343,N_9887,N_9961);
nor UO_1344 (O_1344,N_9846,N_9528);
nand UO_1345 (O_1345,N_9570,N_9651);
nand UO_1346 (O_1346,N_9801,N_9926);
or UO_1347 (O_1347,N_9625,N_9780);
nor UO_1348 (O_1348,N_9917,N_9899);
or UO_1349 (O_1349,N_9610,N_9954);
nor UO_1350 (O_1350,N_9772,N_9757);
nor UO_1351 (O_1351,N_9652,N_9822);
or UO_1352 (O_1352,N_9861,N_9657);
xor UO_1353 (O_1353,N_9595,N_9689);
nand UO_1354 (O_1354,N_9873,N_9655);
or UO_1355 (O_1355,N_9574,N_9704);
nand UO_1356 (O_1356,N_9564,N_9784);
nor UO_1357 (O_1357,N_9953,N_9770);
nand UO_1358 (O_1358,N_9787,N_9707);
nand UO_1359 (O_1359,N_9566,N_9719);
nor UO_1360 (O_1360,N_9924,N_9763);
nand UO_1361 (O_1361,N_9636,N_9688);
and UO_1362 (O_1362,N_9508,N_9819);
nand UO_1363 (O_1363,N_9964,N_9696);
nor UO_1364 (O_1364,N_9742,N_9850);
nor UO_1365 (O_1365,N_9774,N_9726);
nor UO_1366 (O_1366,N_9914,N_9692);
or UO_1367 (O_1367,N_9594,N_9989);
nor UO_1368 (O_1368,N_9968,N_9510);
xnor UO_1369 (O_1369,N_9502,N_9768);
or UO_1370 (O_1370,N_9734,N_9981);
xor UO_1371 (O_1371,N_9524,N_9990);
or UO_1372 (O_1372,N_9961,N_9842);
nand UO_1373 (O_1373,N_9579,N_9521);
or UO_1374 (O_1374,N_9527,N_9584);
nor UO_1375 (O_1375,N_9614,N_9873);
nor UO_1376 (O_1376,N_9501,N_9806);
nand UO_1377 (O_1377,N_9971,N_9728);
xor UO_1378 (O_1378,N_9831,N_9735);
or UO_1379 (O_1379,N_9533,N_9864);
nor UO_1380 (O_1380,N_9526,N_9554);
nor UO_1381 (O_1381,N_9513,N_9860);
or UO_1382 (O_1382,N_9983,N_9746);
xnor UO_1383 (O_1383,N_9700,N_9797);
or UO_1384 (O_1384,N_9548,N_9536);
nor UO_1385 (O_1385,N_9609,N_9518);
and UO_1386 (O_1386,N_9933,N_9958);
or UO_1387 (O_1387,N_9895,N_9849);
or UO_1388 (O_1388,N_9683,N_9742);
or UO_1389 (O_1389,N_9994,N_9622);
xor UO_1390 (O_1390,N_9969,N_9745);
or UO_1391 (O_1391,N_9647,N_9825);
xnor UO_1392 (O_1392,N_9926,N_9844);
and UO_1393 (O_1393,N_9773,N_9543);
or UO_1394 (O_1394,N_9928,N_9662);
nand UO_1395 (O_1395,N_9673,N_9769);
nor UO_1396 (O_1396,N_9605,N_9553);
nor UO_1397 (O_1397,N_9864,N_9920);
or UO_1398 (O_1398,N_9657,N_9577);
nand UO_1399 (O_1399,N_9839,N_9600);
nor UO_1400 (O_1400,N_9927,N_9727);
nand UO_1401 (O_1401,N_9768,N_9923);
nand UO_1402 (O_1402,N_9686,N_9891);
nor UO_1403 (O_1403,N_9678,N_9952);
and UO_1404 (O_1404,N_9561,N_9835);
nand UO_1405 (O_1405,N_9561,N_9820);
nor UO_1406 (O_1406,N_9920,N_9517);
nand UO_1407 (O_1407,N_9948,N_9813);
xor UO_1408 (O_1408,N_9984,N_9581);
and UO_1409 (O_1409,N_9691,N_9736);
or UO_1410 (O_1410,N_9686,N_9687);
nor UO_1411 (O_1411,N_9535,N_9655);
nand UO_1412 (O_1412,N_9997,N_9820);
or UO_1413 (O_1413,N_9903,N_9859);
nand UO_1414 (O_1414,N_9746,N_9821);
nor UO_1415 (O_1415,N_9510,N_9800);
or UO_1416 (O_1416,N_9992,N_9729);
or UO_1417 (O_1417,N_9677,N_9733);
nand UO_1418 (O_1418,N_9689,N_9640);
nand UO_1419 (O_1419,N_9684,N_9630);
nand UO_1420 (O_1420,N_9701,N_9598);
nor UO_1421 (O_1421,N_9762,N_9622);
or UO_1422 (O_1422,N_9947,N_9872);
nand UO_1423 (O_1423,N_9944,N_9807);
and UO_1424 (O_1424,N_9954,N_9550);
or UO_1425 (O_1425,N_9813,N_9957);
or UO_1426 (O_1426,N_9630,N_9541);
and UO_1427 (O_1427,N_9866,N_9820);
and UO_1428 (O_1428,N_9866,N_9603);
nor UO_1429 (O_1429,N_9506,N_9695);
nor UO_1430 (O_1430,N_9965,N_9737);
nand UO_1431 (O_1431,N_9619,N_9838);
nand UO_1432 (O_1432,N_9594,N_9767);
xnor UO_1433 (O_1433,N_9669,N_9632);
and UO_1434 (O_1434,N_9794,N_9551);
or UO_1435 (O_1435,N_9701,N_9621);
and UO_1436 (O_1436,N_9914,N_9510);
or UO_1437 (O_1437,N_9834,N_9965);
nand UO_1438 (O_1438,N_9589,N_9580);
nand UO_1439 (O_1439,N_9577,N_9716);
nand UO_1440 (O_1440,N_9601,N_9795);
nand UO_1441 (O_1441,N_9979,N_9856);
nor UO_1442 (O_1442,N_9700,N_9740);
xnor UO_1443 (O_1443,N_9592,N_9764);
xnor UO_1444 (O_1444,N_9553,N_9524);
nor UO_1445 (O_1445,N_9658,N_9869);
or UO_1446 (O_1446,N_9836,N_9921);
nor UO_1447 (O_1447,N_9725,N_9984);
nand UO_1448 (O_1448,N_9838,N_9594);
xor UO_1449 (O_1449,N_9933,N_9507);
nor UO_1450 (O_1450,N_9617,N_9623);
xor UO_1451 (O_1451,N_9674,N_9676);
nand UO_1452 (O_1452,N_9841,N_9592);
and UO_1453 (O_1453,N_9571,N_9950);
or UO_1454 (O_1454,N_9843,N_9865);
and UO_1455 (O_1455,N_9609,N_9770);
nor UO_1456 (O_1456,N_9530,N_9550);
xnor UO_1457 (O_1457,N_9672,N_9620);
nor UO_1458 (O_1458,N_9676,N_9977);
nand UO_1459 (O_1459,N_9699,N_9509);
nor UO_1460 (O_1460,N_9678,N_9916);
nand UO_1461 (O_1461,N_9723,N_9599);
nor UO_1462 (O_1462,N_9992,N_9819);
and UO_1463 (O_1463,N_9572,N_9536);
or UO_1464 (O_1464,N_9908,N_9846);
or UO_1465 (O_1465,N_9503,N_9771);
and UO_1466 (O_1466,N_9592,N_9616);
xnor UO_1467 (O_1467,N_9562,N_9685);
nand UO_1468 (O_1468,N_9538,N_9805);
and UO_1469 (O_1469,N_9788,N_9914);
and UO_1470 (O_1470,N_9624,N_9982);
nand UO_1471 (O_1471,N_9843,N_9717);
and UO_1472 (O_1472,N_9596,N_9624);
nor UO_1473 (O_1473,N_9958,N_9680);
nor UO_1474 (O_1474,N_9671,N_9782);
nor UO_1475 (O_1475,N_9598,N_9684);
and UO_1476 (O_1476,N_9638,N_9565);
and UO_1477 (O_1477,N_9722,N_9627);
nand UO_1478 (O_1478,N_9830,N_9883);
nand UO_1479 (O_1479,N_9925,N_9788);
or UO_1480 (O_1480,N_9981,N_9541);
or UO_1481 (O_1481,N_9842,N_9997);
and UO_1482 (O_1482,N_9975,N_9589);
nor UO_1483 (O_1483,N_9506,N_9935);
nand UO_1484 (O_1484,N_9771,N_9795);
xor UO_1485 (O_1485,N_9953,N_9824);
or UO_1486 (O_1486,N_9710,N_9637);
and UO_1487 (O_1487,N_9592,N_9655);
xnor UO_1488 (O_1488,N_9578,N_9758);
nor UO_1489 (O_1489,N_9923,N_9875);
nand UO_1490 (O_1490,N_9526,N_9568);
nand UO_1491 (O_1491,N_9676,N_9517);
xnor UO_1492 (O_1492,N_9983,N_9972);
nor UO_1493 (O_1493,N_9619,N_9557);
nor UO_1494 (O_1494,N_9642,N_9838);
or UO_1495 (O_1495,N_9752,N_9988);
nor UO_1496 (O_1496,N_9848,N_9720);
and UO_1497 (O_1497,N_9820,N_9500);
or UO_1498 (O_1498,N_9578,N_9746);
nor UO_1499 (O_1499,N_9855,N_9745);
endmodule