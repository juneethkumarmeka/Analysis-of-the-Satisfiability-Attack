module basic_1000_10000_1500_5_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_74,In_24);
or U1 (N_1,In_244,In_921);
nand U2 (N_2,In_770,In_29);
nand U3 (N_3,In_796,In_146);
and U4 (N_4,In_601,In_654);
nor U5 (N_5,In_482,In_132);
nor U6 (N_6,In_268,In_498);
or U7 (N_7,In_936,In_975);
xnor U8 (N_8,In_254,In_42);
nor U9 (N_9,In_791,In_327);
or U10 (N_10,In_978,In_869);
or U11 (N_11,In_790,In_675);
nor U12 (N_12,In_465,In_308);
or U13 (N_13,In_958,In_925);
or U14 (N_14,In_585,In_863);
and U15 (N_15,In_350,In_200);
or U16 (N_16,In_34,In_281);
nor U17 (N_17,In_807,In_597);
and U18 (N_18,In_1,In_611);
nand U19 (N_19,In_426,In_462);
nand U20 (N_20,In_195,In_660);
nor U21 (N_21,In_859,In_325);
and U22 (N_22,In_184,In_739);
or U23 (N_23,In_445,In_589);
or U24 (N_24,In_673,In_207);
and U25 (N_25,In_539,In_942);
nor U26 (N_26,In_416,In_726);
nor U27 (N_27,In_917,In_9);
or U28 (N_28,In_624,In_14);
nand U29 (N_29,In_775,In_222);
nand U30 (N_30,In_75,In_950);
and U31 (N_31,In_372,In_121);
xnor U32 (N_32,In_534,In_348);
and U33 (N_33,In_748,In_696);
and U34 (N_34,In_178,In_733);
nand U35 (N_35,In_532,In_377);
nand U36 (N_36,In_605,In_334);
nand U37 (N_37,In_530,In_866);
nor U38 (N_38,In_162,In_158);
or U39 (N_39,In_315,In_930);
nand U40 (N_40,In_272,In_213);
nand U41 (N_41,In_376,In_5);
or U42 (N_42,In_509,In_995);
nor U43 (N_43,In_179,In_880);
nor U44 (N_44,In_744,In_289);
and U45 (N_45,In_900,In_641);
nand U46 (N_46,In_494,In_669);
nand U47 (N_47,In_999,In_485);
and U48 (N_48,In_257,In_461);
or U49 (N_49,In_570,In_64);
and U50 (N_50,In_353,In_398);
and U51 (N_51,In_145,In_36);
nand U52 (N_52,In_864,In_747);
or U53 (N_53,In_568,In_356);
or U54 (N_54,In_810,In_837);
and U55 (N_55,In_766,In_43);
and U56 (N_56,In_778,In_983);
or U57 (N_57,In_715,In_799);
or U58 (N_58,In_932,In_609);
or U59 (N_59,In_6,In_365);
nor U60 (N_60,In_151,In_390);
nand U61 (N_61,In_188,In_111);
nand U62 (N_62,In_663,In_940);
nor U63 (N_63,In_813,In_844);
nand U64 (N_64,In_709,In_408);
nand U65 (N_65,In_223,In_202);
or U66 (N_66,In_0,In_99);
and U67 (N_67,In_683,In_58);
and U68 (N_68,In_206,In_724);
and U69 (N_69,In_19,In_467);
nand U70 (N_70,In_584,In_655);
and U71 (N_71,In_374,In_944);
and U72 (N_72,In_172,In_452);
or U73 (N_73,In_962,In_569);
or U74 (N_74,In_631,In_169);
or U75 (N_75,In_407,In_340);
or U76 (N_76,In_537,In_805);
or U77 (N_77,In_551,In_642);
nor U78 (N_78,In_522,In_681);
and U79 (N_79,In_313,In_309);
nand U80 (N_80,In_66,In_126);
or U81 (N_81,In_41,In_263);
nand U82 (N_82,In_989,In_514);
or U83 (N_83,In_571,In_598);
and U84 (N_84,In_862,In_720);
or U85 (N_85,In_895,In_933);
or U86 (N_86,In_171,In_753);
xor U87 (N_87,In_127,In_705);
or U88 (N_88,In_783,In_959);
nand U89 (N_89,In_897,In_302);
nand U90 (N_90,In_752,In_803);
and U91 (N_91,In_544,In_430);
or U92 (N_92,In_203,In_163);
nor U93 (N_93,In_596,In_891);
nand U94 (N_94,In_706,In_231);
nor U95 (N_95,In_758,In_938);
nor U96 (N_96,In_118,In_4);
or U97 (N_97,In_931,In_314);
and U98 (N_98,In_690,In_361);
nand U99 (N_99,In_299,In_84);
nor U100 (N_100,In_435,In_428);
nand U101 (N_101,In_582,In_830);
nand U102 (N_102,In_650,In_890);
nor U103 (N_103,In_627,In_502);
or U104 (N_104,In_347,In_533);
nand U105 (N_105,In_541,In_155);
nand U106 (N_106,In_639,In_243);
nor U107 (N_107,In_772,In_852);
nor U108 (N_108,In_458,In_67);
nand U109 (N_109,In_335,In_848);
nand U110 (N_110,In_241,In_554);
and U111 (N_111,In_996,In_303);
nand U112 (N_112,In_625,In_985);
or U113 (N_113,In_964,In_849);
nand U114 (N_114,In_405,In_117);
or U115 (N_115,In_635,In_73);
nor U116 (N_116,In_89,In_481);
and U117 (N_117,In_516,In_550);
nand U118 (N_118,In_246,In_547);
or U119 (N_119,In_702,In_275);
or U120 (N_120,In_828,In_364);
nand U121 (N_121,In_682,In_496);
nand U122 (N_122,In_908,In_501);
nand U123 (N_123,In_62,In_271);
nand U124 (N_124,In_298,In_52);
and U125 (N_125,In_90,In_761);
or U126 (N_126,In_977,In_59);
and U127 (N_127,In_618,In_45);
nor U128 (N_128,In_578,In_283);
nand U129 (N_129,In_523,In_60);
nor U130 (N_130,In_746,In_500);
nor U131 (N_131,In_559,In_220);
nand U132 (N_132,In_26,In_451);
nand U133 (N_133,In_258,In_998);
nor U134 (N_134,In_168,In_529);
nand U135 (N_135,In_124,In_901);
nand U136 (N_136,In_37,In_285);
nand U137 (N_137,In_731,In_785);
and U138 (N_138,In_765,In_489);
and U139 (N_139,In_97,In_540);
or U140 (N_140,In_741,In_344);
and U141 (N_141,In_366,In_28);
nor U142 (N_142,In_906,In_535);
nor U143 (N_143,In_883,In_719);
nor U144 (N_144,In_227,In_615);
or U145 (N_145,In_665,In_87);
nand U146 (N_146,In_10,In_905);
nand U147 (N_147,In_245,In_191);
and U148 (N_148,In_924,In_961);
nand U149 (N_149,In_763,In_580);
nor U150 (N_150,In_339,In_256);
nor U151 (N_151,In_881,In_531);
nand U152 (N_152,In_72,In_410);
nand U153 (N_153,In_575,In_175);
nand U154 (N_154,In_923,In_929);
nor U155 (N_155,In_769,In_488);
nor U156 (N_156,In_525,In_479);
and U157 (N_157,In_898,In_692);
or U158 (N_158,In_331,In_513);
nand U159 (N_159,In_504,In_518);
nor U160 (N_160,In_926,In_240);
or U161 (N_161,In_307,In_588);
nand U162 (N_162,In_974,In_873);
and U163 (N_163,In_728,In_219);
nand U164 (N_164,In_2,In_16);
nand U165 (N_165,In_745,In_76);
nand U166 (N_166,In_602,In_809);
or U167 (N_167,In_952,In_459);
nand U168 (N_168,In_198,In_18);
or U169 (N_169,In_499,In_899);
and U170 (N_170,In_468,In_210);
or U171 (N_171,In_177,In_716);
xor U172 (N_172,In_484,In_608);
nor U173 (N_173,In_316,In_301);
nor U174 (N_174,In_406,In_341);
nand U175 (N_175,In_469,In_507);
and U176 (N_176,In_816,In_556);
or U177 (N_177,In_422,In_135);
and U178 (N_178,In_510,In_209);
nand U179 (N_179,In_868,In_980);
nor U180 (N_180,In_7,In_528);
nor U181 (N_181,In_282,In_878);
or U182 (N_182,In_599,In_388);
nor U183 (N_183,In_427,In_782);
or U184 (N_184,In_194,In_110);
nand U185 (N_185,In_438,In_463);
nor U186 (N_186,In_704,In_131);
and U187 (N_187,In_987,In_822);
nand U188 (N_188,In_708,In_320);
and U189 (N_189,In_557,In_512);
nand U190 (N_190,In_969,In_23);
nand U191 (N_191,In_35,In_700);
or U192 (N_192,In_71,In_576);
nand U193 (N_193,In_330,In_511);
nand U194 (N_194,In_332,In_919);
nand U195 (N_195,In_208,In_367);
nor U196 (N_196,In_261,In_199);
or U197 (N_197,In_600,In_317);
or U198 (N_198,In_993,In_833);
or U199 (N_199,In_647,In_225);
and U200 (N_200,In_113,In_968);
or U201 (N_201,In_79,In_238);
and U202 (N_202,In_216,In_221);
nor U203 (N_203,In_234,In_779);
or U204 (N_204,In_735,In_278);
nor U205 (N_205,In_904,In_288);
nor U206 (N_206,In_856,In_536);
nand U207 (N_207,In_907,In_319);
nor U208 (N_208,In_885,In_290);
or U209 (N_209,In_617,In_424);
nor U210 (N_210,In_235,In_842);
or U211 (N_211,In_143,In_957);
or U212 (N_212,In_889,In_338);
or U213 (N_213,In_487,In_586);
and U214 (N_214,In_986,In_835);
or U215 (N_215,In_888,In_399);
nand U216 (N_216,In_149,In_214);
or U217 (N_217,In_723,In_976);
or U218 (N_218,In_108,In_693);
nor U219 (N_219,In_343,In_820);
nor U220 (N_220,In_935,In_773);
xor U221 (N_221,In_734,In_871);
nand U222 (N_222,In_251,In_774);
and U223 (N_223,In_280,In_928);
nand U224 (N_224,In_248,In_230);
nor U225 (N_225,In_561,In_699);
nor U226 (N_226,In_371,In_381);
or U227 (N_227,In_98,In_657);
and U228 (N_228,In_363,In_167);
nor U229 (N_229,In_345,In_797);
and U230 (N_230,In_130,In_493);
and U231 (N_231,In_818,In_483);
and U232 (N_232,In_53,In_100);
and U233 (N_233,In_260,In_232);
or U234 (N_234,In_953,In_215);
nor U235 (N_235,In_159,In_182);
nand U236 (N_236,In_471,In_827);
nor U237 (N_237,In_3,In_106);
nand U238 (N_238,In_437,In_141);
and U239 (N_239,In_357,In_689);
nor U240 (N_240,In_284,In_565);
and U241 (N_241,In_250,In_292);
nor U242 (N_242,In_277,In_579);
nand U243 (N_243,In_712,In_259);
and U244 (N_244,In_725,In_606);
nor U245 (N_245,In_922,In_492);
nand U246 (N_246,In_140,In_156);
nand U247 (N_247,In_454,In_337);
nor U248 (N_248,In_619,In_610);
and U249 (N_249,In_701,In_780);
nor U250 (N_250,In_57,In_306);
or U251 (N_251,In_33,In_434);
nor U252 (N_252,In_270,In_144);
nor U253 (N_253,In_638,In_527);
or U254 (N_254,In_722,In_679);
nor U255 (N_255,In_125,In_391);
or U256 (N_256,In_31,In_517);
nor U257 (N_257,In_808,In_264);
and U258 (N_258,In_94,In_300);
nor U259 (N_259,In_400,In_413);
or U260 (N_260,In_46,In_109);
or U261 (N_261,In_738,In_756);
and U262 (N_262,In_825,In_911);
or U263 (N_263,In_373,In_562);
nor U264 (N_264,In_448,In_170);
nand U265 (N_265,In_414,In_651);
nand U266 (N_266,In_841,In_814);
nand U267 (N_267,In_912,In_560);
or U268 (N_268,In_992,In_949);
nand U269 (N_269,In_328,In_927);
nand U270 (N_270,In_604,In_133);
nand U271 (N_271,In_242,In_186);
nor U272 (N_272,In_392,In_247);
or U273 (N_273,In_322,In_860);
nand U274 (N_274,In_433,In_380);
nand U275 (N_275,In_55,In_351);
and U276 (N_276,In_581,In_920);
nand U277 (N_277,In_896,In_553);
nor U278 (N_278,In_193,In_233);
or U279 (N_279,In_239,In_211);
or U280 (N_280,In_368,In_526);
or U281 (N_281,In_838,In_83);
or U282 (N_282,In_902,In_453);
or U283 (N_283,In_92,In_174);
or U284 (N_284,In_662,In_443);
or U285 (N_285,In_710,In_587);
or U286 (N_286,In_629,In_616);
or U287 (N_287,In_595,In_287);
or U288 (N_288,In_44,In_154);
nand U289 (N_289,In_887,In_508);
nor U290 (N_290,In_872,In_115);
and U291 (N_291,In_362,In_486);
or U292 (N_292,In_592,In_691);
nor U293 (N_293,In_966,In_382);
nor U294 (N_294,In_524,In_449);
and U295 (N_295,In_685,In_764);
nand U296 (N_296,In_676,In_730);
or U297 (N_297,In_718,In_442);
nor U298 (N_298,In_909,In_265);
nor U299 (N_299,In_103,In_670);
nor U300 (N_300,In_793,In_678);
and U301 (N_301,In_776,In_160);
and U302 (N_302,In_48,In_369);
and U303 (N_303,In_123,In_274);
and U304 (N_304,In_142,In_861);
nor U305 (N_305,In_988,In_804);
nand U306 (N_306,In_945,In_972);
and U307 (N_307,In_326,In_736);
and U308 (N_308,In_321,In_80);
nor U309 (N_309,In_914,In_189);
xor U310 (N_310,In_947,In_183);
nor U311 (N_311,In_549,In_114);
and U312 (N_312,In_680,In_455);
nor U313 (N_313,In_632,In_794);
or U314 (N_314,In_379,In_760);
or U315 (N_315,In_768,In_583);
nor U316 (N_316,In_505,In_879);
and U317 (N_317,In_994,In_661);
or U318 (N_318,In_946,In_387);
nor U319 (N_319,In_354,In_164);
and U320 (N_320,In_874,In_555);
nand U321 (N_321,In_875,In_310);
and U322 (N_322,In_751,In_478);
nand U323 (N_323,In_847,In_714);
nor U324 (N_324,In_754,In_82);
nor U325 (N_325,In_312,In_865);
nand U326 (N_326,In_294,In_395);
and U327 (N_327,In_684,In_777);
and U328 (N_328,In_477,In_346);
nand U329 (N_329,In_68,In_711);
or U330 (N_330,In_892,In_107);
or U331 (N_331,In_677,In_291);
and U332 (N_332,In_358,In_150);
or U333 (N_333,In_333,In_717);
nor U334 (N_334,In_205,In_971);
nor U335 (N_335,In_614,In_824);
or U336 (N_336,In_843,In_423);
or U337 (N_337,In_954,In_836);
and U338 (N_338,In_137,In_474);
nor U339 (N_339,In_948,In_686);
nand U340 (N_340,In_538,In_104);
nor U341 (N_341,In_762,In_249);
nand U342 (N_342,In_666,In_17);
nor U343 (N_343,In_378,In_286);
and U344 (N_344,In_336,In_846);
nor U345 (N_345,In_27,In_564);
and U346 (N_346,In_419,In_939);
nor U347 (N_347,In_394,In_593);
and U348 (N_348,In_577,In_749);
nor U349 (N_349,In_558,In_91);
and U350 (N_350,In_991,In_129);
nor U351 (N_351,In_147,In_963);
or U352 (N_352,In_607,In_475);
or U353 (N_353,In_798,In_276);
nor U354 (N_354,In_196,In_645);
or U355 (N_355,In_21,In_411);
nor U356 (N_356,In_819,In_727);
nor U357 (N_357,In_855,In_884);
or U358 (N_358,In_542,In_732);
nor U359 (N_359,In_755,In_834);
nand U360 (N_360,In_77,In_273);
nor U361 (N_361,In_653,In_152);
and U362 (N_362,In_648,In_429);
or U363 (N_363,In_687,In_913);
or U364 (N_364,In_603,In_789);
and U365 (N_365,In_476,In_737);
nor U366 (N_366,In_12,In_829);
or U367 (N_367,In_296,In_444);
or U368 (N_368,In_165,In_65);
or U369 (N_369,In_224,In_743);
or U370 (N_370,In_412,In_323);
nand U371 (N_371,In_421,In_491);
or U372 (N_372,In_187,In_86);
nor U373 (N_373,In_566,In_457);
xor U374 (N_374,In_311,In_418);
or U375 (N_375,In_674,In_456);
nor U376 (N_376,In_401,In_503);
and U377 (N_377,In_646,In_695);
nor U378 (N_378,In_39,In_11);
nor U379 (N_379,In_965,In_51);
nand U380 (N_380,In_546,In_101);
nand U381 (N_381,In_56,In_594);
nor U382 (N_382,In_973,In_63);
nor U383 (N_383,In_229,In_415);
nand U384 (N_384,In_870,In_817);
or U385 (N_385,In_441,In_882);
nand U386 (N_386,In_185,In_573);
and U387 (N_387,In_979,In_590);
or U388 (N_388,In_329,In_397);
nor U389 (N_389,In_318,In_664);
and U390 (N_390,In_621,In_886);
and U391 (N_391,In_385,In_955);
nand U392 (N_392,In_786,In_236);
or U393 (N_393,In_703,In_800);
nand U394 (N_394,In_652,In_40);
nand U395 (N_395,In_237,In_876);
nor U396 (N_396,In_937,In_61);
or U397 (N_397,In_409,In_383);
and U398 (N_398,In_759,In_567);
and U399 (N_399,In_612,In_792);
nand U400 (N_400,In_845,In_497);
nand U401 (N_401,In_370,In_102);
xor U402 (N_402,In_173,In_440);
and U403 (N_403,In_93,In_269);
nor U404 (N_404,In_105,In_49);
nand U405 (N_405,In_644,In_630);
or U406 (N_406,In_697,In_192);
and U407 (N_407,In_47,In_78);
and U408 (N_408,In_688,In_802);
and U409 (N_409,In_548,In_352);
nor U410 (N_410,In_20,In_349);
or U411 (N_411,In_88,In_495);
and U412 (N_412,In_212,In_795);
nor U413 (N_413,In_671,In_267);
and U414 (N_414,In_490,In_622);
nor U415 (N_415,In_997,In_226);
or U416 (N_416,In_519,In_915);
or U417 (N_417,In_543,In_181);
or U418 (N_418,In_506,In_50);
nor U419 (N_419,In_420,In_355);
nor U420 (N_420,In_815,In_729);
nand U421 (N_421,In_81,In_204);
and U422 (N_422,In_941,In_771);
or U423 (N_423,In_255,In_404);
xor U424 (N_424,In_956,In_324);
nor U425 (N_425,In_877,In_831);
or U426 (N_426,In_806,In_436);
nor U427 (N_427,In_649,In_572);
or U428 (N_428,In_470,In_659);
or U429 (N_429,In_116,In_910);
nand U430 (N_430,In_628,In_95);
nor U431 (N_431,In_640,In_396);
nand U432 (N_432,In_417,In_894);
nand U433 (N_433,In_384,In_473);
or U434 (N_434,In_180,In_134);
and U435 (N_435,In_713,In_136);
nor U436 (N_436,In_552,In_13);
nand U437 (N_437,In_197,In_8);
or U438 (N_438,In_857,In_858);
nor U439 (N_439,In_228,In_432);
nand U440 (N_440,In_960,In_851);
and U441 (N_441,In_25,In_967);
and U442 (N_442,In_812,In_757);
nor U443 (N_443,In_982,In_984);
or U444 (N_444,In_636,In_112);
and U445 (N_445,In_360,In_425);
or U446 (N_446,In_721,In_943);
nand U447 (N_447,In_811,In_637);
nor U448 (N_448,In_990,In_217);
or U449 (N_449,In_262,In_821);
or U450 (N_450,In_15,In_672);
nand U451 (N_451,In_431,In_30);
and U452 (N_452,In_801,In_297);
nand U453 (N_453,In_69,In_120);
or U454 (N_454,In_403,In_279);
or U455 (N_455,In_788,In_970);
nor U456 (N_456,In_840,In_439);
and U457 (N_457,In_153,In_839);
nor U458 (N_458,In_591,In_460);
nand U459 (N_459,In_157,In_450);
and U460 (N_460,In_375,In_643);
or U461 (N_461,In_359,In_853);
and U462 (N_462,In_613,In_295);
nor U463 (N_463,In_342,In_201);
and U464 (N_464,In_626,In_466);
and U465 (N_465,In_266,In_750);
nand U466 (N_466,In_176,In_823);
and U467 (N_467,In_464,In_658);
nor U468 (N_468,In_480,In_520);
nor U469 (N_469,In_96,In_694);
nor U470 (N_470,In_668,In_867);
or U471 (N_471,In_667,In_918);
and U472 (N_472,In_122,In_515);
nor U473 (N_473,In_138,In_563);
nand U474 (N_474,In_981,In_826);
nand U475 (N_475,In_656,In_707);
nand U476 (N_476,In_166,In_893);
nand U477 (N_477,In_70,In_545);
nand U478 (N_478,In_218,In_767);
nor U479 (N_479,In_393,In_389);
nand U480 (N_480,In_787,In_934);
xor U481 (N_481,In_916,In_850);
or U482 (N_482,In_740,In_22);
nor U483 (N_483,In_620,In_742);
and U484 (N_484,In_139,In_903);
nand U485 (N_485,In_623,In_634);
nand U486 (N_486,In_574,In_521);
nor U487 (N_487,In_781,In_832);
nand U488 (N_488,In_293,In_386);
nand U489 (N_489,In_85,In_253);
or U490 (N_490,In_446,In_472);
or U491 (N_491,In_304,In_119);
nor U492 (N_492,In_951,In_148);
nand U493 (N_493,In_54,In_161);
or U494 (N_494,In_402,In_128);
nor U495 (N_495,In_698,In_38);
and U496 (N_496,In_784,In_633);
and U497 (N_497,In_190,In_854);
nor U498 (N_498,In_305,In_252);
and U499 (N_499,In_447,In_32);
and U500 (N_500,In_180,In_578);
nand U501 (N_501,In_341,In_891);
or U502 (N_502,In_812,In_67);
or U503 (N_503,In_10,In_629);
nor U504 (N_504,In_480,In_970);
nand U505 (N_505,In_389,In_947);
nor U506 (N_506,In_322,In_817);
and U507 (N_507,In_644,In_768);
nor U508 (N_508,In_452,In_993);
nand U509 (N_509,In_971,In_632);
or U510 (N_510,In_539,In_148);
and U511 (N_511,In_295,In_153);
or U512 (N_512,In_398,In_878);
nand U513 (N_513,In_100,In_219);
nand U514 (N_514,In_897,In_298);
nor U515 (N_515,In_535,In_461);
and U516 (N_516,In_10,In_676);
nand U517 (N_517,In_886,In_625);
nor U518 (N_518,In_836,In_488);
and U519 (N_519,In_815,In_928);
nand U520 (N_520,In_947,In_6);
nor U521 (N_521,In_959,In_206);
or U522 (N_522,In_746,In_445);
nor U523 (N_523,In_825,In_532);
and U524 (N_524,In_697,In_590);
and U525 (N_525,In_128,In_432);
nand U526 (N_526,In_529,In_806);
and U527 (N_527,In_263,In_510);
and U528 (N_528,In_248,In_961);
nor U529 (N_529,In_353,In_73);
or U530 (N_530,In_17,In_522);
nor U531 (N_531,In_232,In_452);
nor U532 (N_532,In_691,In_87);
nor U533 (N_533,In_843,In_397);
and U534 (N_534,In_270,In_896);
and U535 (N_535,In_572,In_265);
or U536 (N_536,In_752,In_47);
or U537 (N_537,In_561,In_123);
nand U538 (N_538,In_726,In_81);
or U539 (N_539,In_625,In_37);
and U540 (N_540,In_492,In_337);
nor U541 (N_541,In_474,In_781);
nand U542 (N_542,In_617,In_901);
or U543 (N_543,In_885,In_787);
nand U544 (N_544,In_110,In_920);
nand U545 (N_545,In_127,In_44);
nor U546 (N_546,In_648,In_66);
nand U547 (N_547,In_113,In_925);
or U548 (N_548,In_88,In_666);
and U549 (N_549,In_982,In_323);
nor U550 (N_550,In_583,In_951);
nand U551 (N_551,In_579,In_264);
or U552 (N_552,In_351,In_928);
nor U553 (N_553,In_641,In_680);
nand U554 (N_554,In_44,In_862);
or U555 (N_555,In_202,In_446);
nand U556 (N_556,In_182,In_283);
and U557 (N_557,In_835,In_154);
or U558 (N_558,In_607,In_963);
nor U559 (N_559,In_345,In_424);
nand U560 (N_560,In_609,In_117);
nor U561 (N_561,In_52,In_451);
and U562 (N_562,In_595,In_76);
nand U563 (N_563,In_168,In_566);
or U564 (N_564,In_346,In_576);
nand U565 (N_565,In_883,In_196);
nand U566 (N_566,In_138,In_259);
or U567 (N_567,In_730,In_675);
or U568 (N_568,In_545,In_858);
nor U569 (N_569,In_48,In_256);
nor U570 (N_570,In_696,In_587);
nor U571 (N_571,In_283,In_833);
or U572 (N_572,In_771,In_826);
nor U573 (N_573,In_93,In_987);
and U574 (N_574,In_196,In_847);
and U575 (N_575,In_851,In_695);
and U576 (N_576,In_655,In_339);
and U577 (N_577,In_490,In_186);
and U578 (N_578,In_860,In_650);
nand U579 (N_579,In_354,In_831);
nand U580 (N_580,In_396,In_764);
and U581 (N_581,In_932,In_460);
nand U582 (N_582,In_642,In_751);
nand U583 (N_583,In_817,In_511);
and U584 (N_584,In_204,In_371);
nor U585 (N_585,In_917,In_612);
and U586 (N_586,In_79,In_104);
nand U587 (N_587,In_800,In_854);
and U588 (N_588,In_186,In_163);
and U589 (N_589,In_773,In_440);
and U590 (N_590,In_203,In_767);
nand U591 (N_591,In_315,In_293);
and U592 (N_592,In_520,In_503);
nand U593 (N_593,In_201,In_105);
nand U594 (N_594,In_927,In_447);
or U595 (N_595,In_297,In_18);
nand U596 (N_596,In_965,In_693);
nand U597 (N_597,In_219,In_228);
nand U598 (N_598,In_16,In_40);
nand U599 (N_599,In_184,In_325);
or U600 (N_600,In_443,In_234);
nor U601 (N_601,In_213,In_948);
and U602 (N_602,In_597,In_71);
and U603 (N_603,In_980,In_555);
and U604 (N_604,In_63,In_578);
or U605 (N_605,In_108,In_249);
nor U606 (N_606,In_561,In_197);
or U607 (N_607,In_934,In_47);
xnor U608 (N_608,In_882,In_159);
nor U609 (N_609,In_527,In_968);
nand U610 (N_610,In_301,In_997);
nor U611 (N_611,In_348,In_250);
and U612 (N_612,In_794,In_697);
and U613 (N_613,In_790,In_74);
nor U614 (N_614,In_240,In_604);
and U615 (N_615,In_789,In_495);
xnor U616 (N_616,In_642,In_480);
nor U617 (N_617,In_874,In_905);
nor U618 (N_618,In_601,In_380);
nor U619 (N_619,In_600,In_25);
or U620 (N_620,In_291,In_640);
or U621 (N_621,In_40,In_585);
or U622 (N_622,In_444,In_343);
nand U623 (N_623,In_153,In_327);
and U624 (N_624,In_252,In_736);
or U625 (N_625,In_413,In_228);
nand U626 (N_626,In_443,In_240);
or U627 (N_627,In_539,In_187);
or U628 (N_628,In_797,In_834);
nor U629 (N_629,In_127,In_375);
nor U630 (N_630,In_76,In_441);
and U631 (N_631,In_944,In_265);
and U632 (N_632,In_357,In_535);
nor U633 (N_633,In_960,In_965);
nand U634 (N_634,In_966,In_817);
and U635 (N_635,In_384,In_968);
nor U636 (N_636,In_223,In_335);
or U637 (N_637,In_664,In_502);
nand U638 (N_638,In_336,In_726);
nor U639 (N_639,In_84,In_55);
or U640 (N_640,In_189,In_905);
nand U641 (N_641,In_186,In_245);
nor U642 (N_642,In_35,In_385);
or U643 (N_643,In_355,In_532);
nor U644 (N_644,In_211,In_950);
nor U645 (N_645,In_904,In_955);
and U646 (N_646,In_685,In_260);
and U647 (N_647,In_130,In_435);
nor U648 (N_648,In_706,In_818);
nand U649 (N_649,In_889,In_526);
nand U650 (N_650,In_556,In_452);
and U651 (N_651,In_362,In_216);
nor U652 (N_652,In_379,In_713);
nor U653 (N_653,In_8,In_244);
or U654 (N_654,In_322,In_410);
nor U655 (N_655,In_344,In_698);
nand U656 (N_656,In_362,In_570);
nand U657 (N_657,In_899,In_514);
nand U658 (N_658,In_861,In_740);
nand U659 (N_659,In_947,In_295);
and U660 (N_660,In_826,In_790);
xor U661 (N_661,In_746,In_460);
nor U662 (N_662,In_6,In_481);
nor U663 (N_663,In_777,In_627);
or U664 (N_664,In_991,In_10);
nand U665 (N_665,In_212,In_921);
or U666 (N_666,In_405,In_129);
nand U667 (N_667,In_400,In_824);
nor U668 (N_668,In_649,In_938);
xor U669 (N_669,In_421,In_241);
nor U670 (N_670,In_445,In_856);
nor U671 (N_671,In_595,In_707);
or U672 (N_672,In_71,In_51);
nor U673 (N_673,In_383,In_478);
nand U674 (N_674,In_849,In_668);
nor U675 (N_675,In_65,In_12);
or U676 (N_676,In_689,In_382);
or U677 (N_677,In_996,In_212);
or U678 (N_678,In_820,In_854);
nor U679 (N_679,In_749,In_149);
nand U680 (N_680,In_271,In_728);
nor U681 (N_681,In_778,In_493);
and U682 (N_682,In_738,In_425);
nand U683 (N_683,In_854,In_397);
nor U684 (N_684,In_395,In_679);
nor U685 (N_685,In_128,In_707);
nor U686 (N_686,In_22,In_57);
or U687 (N_687,In_76,In_41);
nor U688 (N_688,In_639,In_747);
nand U689 (N_689,In_814,In_363);
nor U690 (N_690,In_175,In_856);
nand U691 (N_691,In_486,In_922);
nand U692 (N_692,In_553,In_131);
or U693 (N_693,In_836,In_710);
nor U694 (N_694,In_901,In_583);
nor U695 (N_695,In_714,In_320);
or U696 (N_696,In_43,In_331);
and U697 (N_697,In_261,In_141);
nor U698 (N_698,In_571,In_958);
nor U699 (N_699,In_659,In_103);
nor U700 (N_700,In_973,In_349);
and U701 (N_701,In_129,In_250);
and U702 (N_702,In_654,In_534);
nor U703 (N_703,In_19,In_970);
or U704 (N_704,In_334,In_856);
nand U705 (N_705,In_921,In_951);
and U706 (N_706,In_750,In_226);
nand U707 (N_707,In_999,In_131);
and U708 (N_708,In_876,In_758);
or U709 (N_709,In_495,In_84);
nand U710 (N_710,In_72,In_832);
nor U711 (N_711,In_732,In_599);
nand U712 (N_712,In_278,In_7);
nand U713 (N_713,In_113,In_32);
or U714 (N_714,In_240,In_316);
nand U715 (N_715,In_928,In_701);
and U716 (N_716,In_208,In_657);
nand U717 (N_717,In_768,In_435);
nand U718 (N_718,In_689,In_7);
nand U719 (N_719,In_26,In_349);
and U720 (N_720,In_19,In_141);
and U721 (N_721,In_308,In_530);
nor U722 (N_722,In_50,In_164);
or U723 (N_723,In_377,In_500);
and U724 (N_724,In_213,In_869);
nand U725 (N_725,In_275,In_465);
nand U726 (N_726,In_205,In_199);
xor U727 (N_727,In_254,In_664);
and U728 (N_728,In_481,In_174);
nor U729 (N_729,In_834,In_214);
or U730 (N_730,In_595,In_779);
nor U731 (N_731,In_448,In_787);
and U732 (N_732,In_701,In_793);
or U733 (N_733,In_294,In_19);
nor U734 (N_734,In_860,In_878);
or U735 (N_735,In_648,In_514);
nand U736 (N_736,In_871,In_469);
nor U737 (N_737,In_676,In_918);
nor U738 (N_738,In_848,In_684);
and U739 (N_739,In_481,In_187);
nand U740 (N_740,In_662,In_122);
and U741 (N_741,In_902,In_77);
nor U742 (N_742,In_571,In_166);
nand U743 (N_743,In_544,In_384);
nor U744 (N_744,In_801,In_153);
nor U745 (N_745,In_781,In_986);
nand U746 (N_746,In_761,In_488);
nor U747 (N_747,In_982,In_506);
nor U748 (N_748,In_97,In_506);
nand U749 (N_749,In_757,In_139);
nand U750 (N_750,In_268,In_943);
nor U751 (N_751,In_971,In_614);
or U752 (N_752,In_173,In_298);
nor U753 (N_753,In_870,In_932);
nor U754 (N_754,In_513,In_411);
nand U755 (N_755,In_339,In_752);
nand U756 (N_756,In_736,In_595);
nand U757 (N_757,In_969,In_795);
nor U758 (N_758,In_543,In_245);
and U759 (N_759,In_779,In_542);
nor U760 (N_760,In_329,In_584);
and U761 (N_761,In_217,In_736);
and U762 (N_762,In_772,In_692);
nand U763 (N_763,In_810,In_402);
nand U764 (N_764,In_210,In_972);
nand U765 (N_765,In_338,In_457);
nand U766 (N_766,In_658,In_474);
nand U767 (N_767,In_220,In_807);
and U768 (N_768,In_765,In_450);
and U769 (N_769,In_787,In_654);
nor U770 (N_770,In_123,In_256);
and U771 (N_771,In_267,In_771);
or U772 (N_772,In_680,In_685);
or U773 (N_773,In_293,In_371);
nand U774 (N_774,In_36,In_97);
and U775 (N_775,In_714,In_849);
nor U776 (N_776,In_483,In_846);
nor U777 (N_777,In_506,In_188);
nor U778 (N_778,In_38,In_933);
or U779 (N_779,In_307,In_868);
nor U780 (N_780,In_820,In_448);
nand U781 (N_781,In_208,In_608);
and U782 (N_782,In_849,In_211);
nor U783 (N_783,In_837,In_539);
and U784 (N_784,In_782,In_204);
nor U785 (N_785,In_279,In_235);
or U786 (N_786,In_460,In_56);
nand U787 (N_787,In_618,In_885);
nand U788 (N_788,In_709,In_47);
nand U789 (N_789,In_469,In_64);
nor U790 (N_790,In_260,In_255);
or U791 (N_791,In_736,In_37);
nor U792 (N_792,In_778,In_107);
nor U793 (N_793,In_406,In_605);
and U794 (N_794,In_890,In_319);
nand U795 (N_795,In_589,In_394);
or U796 (N_796,In_507,In_24);
and U797 (N_797,In_805,In_669);
nor U798 (N_798,In_850,In_363);
or U799 (N_799,In_420,In_308);
or U800 (N_800,In_378,In_525);
and U801 (N_801,In_984,In_69);
nand U802 (N_802,In_449,In_7);
nand U803 (N_803,In_111,In_705);
and U804 (N_804,In_695,In_973);
nor U805 (N_805,In_301,In_855);
nor U806 (N_806,In_565,In_148);
nor U807 (N_807,In_53,In_327);
or U808 (N_808,In_888,In_112);
or U809 (N_809,In_755,In_780);
nor U810 (N_810,In_106,In_575);
or U811 (N_811,In_227,In_105);
nor U812 (N_812,In_388,In_560);
or U813 (N_813,In_754,In_11);
nand U814 (N_814,In_103,In_68);
and U815 (N_815,In_465,In_24);
nor U816 (N_816,In_350,In_322);
nor U817 (N_817,In_729,In_505);
nand U818 (N_818,In_845,In_729);
or U819 (N_819,In_946,In_198);
or U820 (N_820,In_2,In_151);
nor U821 (N_821,In_271,In_279);
and U822 (N_822,In_222,In_30);
nor U823 (N_823,In_206,In_613);
nand U824 (N_824,In_900,In_116);
or U825 (N_825,In_862,In_750);
nand U826 (N_826,In_136,In_606);
xor U827 (N_827,In_157,In_64);
nand U828 (N_828,In_159,In_223);
nor U829 (N_829,In_296,In_760);
nor U830 (N_830,In_432,In_250);
nand U831 (N_831,In_11,In_811);
or U832 (N_832,In_291,In_979);
and U833 (N_833,In_794,In_373);
nand U834 (N_834,In_605,In_830);
nand U835 (N_835,In_845,In_701);
and U836 (N_836,In_622,In_949);
nor U837 (N_837,In_76,In_888);
nand U838 (N_838,In_665,In_607);
and U839 (N_839,In_31,In_529);
or U840 (N_840,In_98,In_591);
and U841 (N_841,In_293,In_260);
or U842 (N_842,In_448,In_452);
nand U843 (N_843,In_337,In_548);
and U844 (N_844,In_539,In_839);
and U845 (N_845,In_499,In_271);
nand U846 (N_846,In_820,In_67);
nand U847 (N_847,In_14,In_68);
nand U848 (N_848,In_348,In_167);
nand U849 (N_849,In_401,In_114);
nor U850 (N_850,In_488,In_94);
nand U851 (N_851,In_485,In_827);
nand U852 (N_852,In_378,In_188);
nand U853 (N_853,In_47,In_18);
or U854 (N_854,In_875,In_791);
and U855 (N_855,In_795,In_699);
and U856 (N_856,In_607,In_915);
nor U857 (N_857,In_231,In_579);
or U858 (N_858,In_839,In_249);
and U859 (N_859,In_725,In_644);
nand U860 (N_860,In_280,In_20);
nor U861 (N_861,In_796,In_568);
nand U862 (N_862,In_639,In_857);
or U863 (N_863,In_814,In_526);
or U864 (N_864,In_863,In_638);
nand U865 (N_865,In_97,In_887);
nor U866 (N_866,In_945,In_340);
nand U867 (N_867,In_301,In_86);
or U868 (N_868,In_186,In_372);
nand U869 (N_869,In_634,In_254);
and U870 (N_870,In_378,In_147);
nand U871 (N_871,In_605,In_817);
nand U872 (N_872,In_79,In_856);
nor U873 (N_873,In_917,In_251);
nor U874 (N_874,In_351,In_647);
nand U875 (N_875,In_632,In_159);
or U876 (N_876,In_696,In_40);
and U877 (N_877,In_675,In_802);
or U878 (N_878,In_166,In_370);
or U879 (N_879,In_562,In_767);
and U880 (N_880,In_282,In_595);
nor U881 (N_881,In_566,In_871);
and U882 (N_882,In_863,In_932);
or U883 (N_883,In_285,In_846);
nor U884 (N_884,In_989,In_125);
nand U885 (N_885,In_41,In_423);
and U886 (N_886,In_453,In_833);
nand U887 (N_887,In_520,In_4);
nor U888 (N_888,In_685,In_236);
nor U889 (N_889,In_478,In_56);
and U890 (N_890,In_756,In_289);
or U891 (N_891,In_388,In_362);
or U892 (N_892,In_322,In_656);
or U893 (N_893,In_78,In_687);
nor U894 (N_894,In_813,In_625);
nor U895 (N_895,In_552,In_9);
nor U896 (N_896,In_170,In_419);
and U897 (N_897,In_642,In_942);
nor U898 (N_898,In_690,In_541);
nand U899 (N_899,In_572,In_496);
and U900 (N_900,In_195,In_883);
nor U901 (N_901,In_381,In_582);
nor U902 (N_902,In_501,In_112);
or U903 (N_903,In_0,In_378);
nor U904 (N_904,In_778,In_137);
or U905 (N_905,In_417,In_400);
nor U906 (N_906,In_463,In_325);
nand U907 (N_907,In_841,In_356);
nor U908 (N_908,In_830,In_663);
nand U909 (N_909,In_444,In_971);
nor U910 (N_910,In_708,In_274);
nand U911 (N_911,In_308,In_666);
nand U912 (N_912,In_842,In_107);
nand U913 (N_913,In_402,In_848);
nand U914 (N_914,In_444,In_158);
nand U915 (N_915,In_887,In_155);
nor U916 (N_916,In_22,In_348);
nand U917 (N_917,In_987,In_862);
or U918 (N_918,In_774,In_347);
nor U919 (N_919,In_117,In_738);
and U920 (N_920,In_543,In_708);
and U921 (N_921,In_937,In_884);
nand U922 (N_922,In_670,In_478);
nand U923 (N_923,In_636,In_913);
and U924 (N_924,In_175,In_189);
nand U925 (N_925,In_309,In_267);
and U926 (N_926,In_863,In_572);
and U927 (N_927,In_754,In_322);
nor U928 (N_928,In_178,In_804);
and U929 (N_929,In_110,In_863);
or U930 (N_930,In_888,In_606);
nor U931 (N_931,In_94,In_675);
nor U932 (N_932,In_467,In_362);
nor U933 (N_933,In_825,In_645);
or U934 (N_934,In_981,In_576);
and U935 (N_935,In_133,In_785);
or U936 (N_936,In_8,In_774);
and U937 (N_937,In_840,In_997);
or U938 (N_938,In_992,In_540);
nor U939 (N_939,In_905,In_665);
and U940 (N_940,In_563,In_308);
and U941 (N_941,In_983,In_185);
nor U942 (N_942,In_876,In_78);
or U943 (N_943,In_740,In_50);
nand U944 (N_944,In_896,In_195);
and U945 (N_945,In_401,In_585);
nor U946 (N_946,In_807,In_588);
nand U947 (N_947,In_433,In_407);
nor U948 (N_948,In_844,In_479);
nor U949 (N_949,In_890,In_540);
nand U950 (N_950,In_54,In_243);
or U951 (N_951,In_790,In_679);
and U952 (N_952,In_930,In_469);
nand U953 (N_953,In_625,In_435);
and U954 (N_954,In_990,In_589);
or U955 (N_955,In_326,In_359);
or U956 (N_956,In_126,In_933);
nand U957 (N_957,In_774,In_726);
or U958 (N_958,In_181,In_565);
nand U959 (N_959,In_463,In_171);
nand U960 (N_960,In_476,In_856);
or U961 (N_961,In_452,In_578);
nor U962 (N_962,In_604,In_746);
nand U963 (N_963,In_334,In_414);
nand U964 (N_964,In_893,In_16);
nor U965 (N_965,In_254,In_258);
nand U966 (N_966,In_634,In_108);
nand U967 (N_967,In_849,In_289);
or U968 (N_968,In_110,In_689);
and U969 (N_969,In_884,In_704);
nand U970 (N_970,In_507,In_962);
or U971 (N_971,In_674,In_950);
nor U972 (N_972,In_419,In_672);
nand U973 (N_973,In_527,In_352);
nor U974 (N_974,In_413,In_930);
nand U975 (N_975,In_739,In_415);
or U976 (N_976,In_972,In_297);
nand U977 (N_977,In_5,In_286);
nand U978 (N_978,In_788,In_833);
nor U979 (N_979,In_665,In_546);
nor U980 (N_980,In_823,In_15);
or U981 (N_981,In_923,In_38);
or U982 (N_982,In_226,In_795);
and U983 (N_983,In_298,In_799);
xor U984 (N_984,In_43,In_144);
nor U985 (N_985,In_870,In_894);
or U986 (N_986,In_713,In_683);
or U987 (N_987,In_106,In_974);
or U988 (N_988,In_79,In_718);
nand U989 (N_989,In_560,In_593);
nor U990 (N_990,In_545,In_578);
nor U991 (N_991,In_991,In_303);
nor U992 (N_992,In_44,In_355);
and U993 (N_993,In_763,In_124);
nand U994 (N_994,In_624,In_227);
or U995 (N_995,In_314,In_541);
nor U996 (N_996,In_517,In_345);
and U997 (N_997,In_87,In_482);
nand U998 (N_998,In_90,In_150);
nor U999 (N_999,In_0,In_716);
nor U1000 (N_1000,In_60,In_731);
nor U1001 (N_1001,In_869,In_486);
nor U1002 (N_1002,In_998,In_640);
nor U1003 (N_1003,In_554,In_565);
and U1004 (N_1004,In_395,In_629);
and U1005 (N_1005,In_531,In_301);
nand U1006 (N_1006,In_942,In_392);
or U1007 (N_1007,In_167,In_559);
nand U1008 (N_1008,In_530,In_659);
and U1009 (N_1009,In_176,In_199);
nor U1010 (N_1010,In_277,In_108);
nand U1011 (N_1011,In_630,In_53);
nor U1012 (N_1012,In_474,In_924);
nand U1013 (N_1013,In_457,In_581);
and U1014 (N_1014,In_932,In_413);
nor U1015 (N_1015,In_854,In_172);
or U1016 (N_1016,In_648,In_477);
and U1017 (N_1017,In_540,In_917);
nand U1018 (N_1018,In_442,In_554);
and U1019 (N_1019,In_293,In_937);
nand U1020 (N_1020,In_222,In_1);
nor U1021 (N_1021,In_368,In_67);
nor U1022 (N_1022,In_432,In_827);
nor U1023 (N_1023,In_240,In_402);
nand U1024 (N_1024,In_858,In_569);
nand U1025 (N_1025,In_485,In_944);
or U1026 (N_1026,In_909,In_214);
nand U1027 (N_1027,In_440,In_291);
nor U1028 (N_1028,In_436,In_761);
nand U1029 (N_1029,In_967,In_73);
xnor U1030 (N_1030,In_879,In_786);
nor U1031 (N_1031,In_77,In_338);
or U1032 (N_1032,In_670,In_291);
nand U1033 (N_1033,In_658,In_429);
and U1034 (N_1034,In_871,In_106);
and U1035 (N_1035,In_245,In_885);
nor U1036 (N_1036,In_478,In_270);
nand U1037 (N_1037,In_39,In_411);
nand U1038 (N_1038,In_852,In_534);
nand U1039 (N_1039,In_993,In_375);
or U1040 (N_1040,In_213,In_694);
nor U1041 (N_1041,In_393,In_733);
and U1042 (N_1042,In_388,In_58);
and U1043 (N_1043,In_343,In_548);
or U1044 (N_1044,In_291,In_406);
or U1045 (N_1045,In_66,In_917);
nor U1046 (N_1046,In_50,In_334);
nand U1047 (N_1047,In_563,In_141);
nor U1048 (N_1048,In_323,In_656);
and U1049 (N_1049,In_105,In_236);
nand U1050 (N_1050,In_401,In_50);
and U1051 (N_1051,In_354,In_342);
and U1052 (N_1052,In_87,In_305);
nand U1053 (N_1053,In_661,In_918);
or U1054 (N_1054,In_676,In_493);
or U1055 (N_1055,In_556,In_885);
or U1056 (N_1056,In_686,In_158);
and U1057 (N_1057,In_543,In_150);
or U1058 (N_1058,In_908,In_858);
nand U1059 (N_1059,In_602,In_287);
nand U1060 (N_1060,In_466,In_826);
or U1061 (N_1061,In_623,In_691);
nor U1062 (N_1062,In_403,In_146);
or U1063 (N_1063,In_207,In_208);
and U1064 (N_1064,In_160,In_755);
or U1065 (N_1065,In_630,In_880);
nor U1066 (N_1066,In_521,In_889);
or U1067 (N_1067,In_441,In_423);
and U1068 (N_1068,In_82,In_259);
or U1069 (N_1069,In_414,In_462);
or U1070 (N_1070,In_615,In_823);
nor U1071 (N_1071,In_681,In_367);
and U1072 (N_1072,In_933,In_496);
nor U1073 (N_1073,In_376,In_664);
or U1074 (N_1074,In_675,In_804);
nand U1075 (N_1075,In_786,In_38);
or U1076 (N_1076,In_369,In_141);
and U1077 (N_1077,In_973,In_149);
and U1078 (N_1078,In_803,In_266);
or U1079 (N_1079,In_78,In_314);
nand U1080 (N_1080,In_572,In_105);
nor U1081 (N_1081,In_508,In_673);
and U1082 (N_1082,In_798,In_283);
or U1083 (N_1083,In_499,In_953);
or U1084 (N_1084,In_582,In_552);
and U1085 (N_1085,In_700,In_327);
nor U1086 (N_1086,In_819,In_423);
nor U1087 (N_1087,In_770,In_776);
or U1088 (N_1088,In_657,In_574);
nand U1089 (N_1089,In_101,In_318);
nand U1090 (N_1090,In_597,In_579);
and U1091 (N_1091,In_758,In_840);
nand U1092 (N_1092,In_323,In_485);
and U1093 (N_1093,In_589,In_363);
nand U1094 (N_1094,In_213,In_351);
or U1095 (N_1095,In_794,In_949);
or U1096 (N_1096,In_445,In_704);
nand U1097 (N_1097,In_972,In_741);
or U1098 (N_1098,In_807,In_26);
and U1099 (N_1099,In_622,In_113);
and U1100 (N_1100,In_927,In_158);
or U1101 (N_1101,In_211,In_866);
or U1102 (N_1102,In_386,In_962);
or U1103 (N_1103,In_75,In_103);
or U1104 (N_1104,In_905,In_155);
nand U1105 (N_1105,In_844,In_671);
nor U1106 (N_1106,In_925,In_620);
nand U1107 (N_1107,In_773,In_916);
or U1108 (N_1108,In_643,In_478);
and U1109 (N_1109,In_672,In_406);
nor U1110 (N_1110,In_853,In_79);
nand U1111 (N_1111,In_625,In_372);
nand U1112 (N_1112,In_144,In_367);
nor U1113 (N_1113,In_313,In_318);
nand U1114 (N_1114,In_90,In_707);
or U1115 (N_1115,In_774,In_182);
nor U1116 (N_1116,In_260,In_344);
nand U1117 (N_1117,In_570,In_689);
or U1118 (N_1118,In_124,In_918);
and U1119 (N_1119,In_895,In_833);
or U1120 (N_1120,In_861,In_431);
and U1121 (N_1121,In_112,In_385);
nand U1122 (N_1122,In_800,In_303);
and U1123 (N_1123,In_433,In_726);
or U1124 (N_1124,In_844,In_840);
nand U1125 (N_1125,In_88,In_860);
and U1126 (N_1126,In_855,In_746);
or U1127 (N_1127,In_620,In_561);
and U1128 (N_1128,In_94,In_762);
and U1129 (N_1129,In_598,In_338);
nor U1130 (N_1130,In_851,In_509);
nand U1131 (N_1131,In_368,In_953);
nor U1132 (N_1132,In_532,In_289);
and U1133 (N_1133,In_352,In_281);
and U1134 (N_1134,In_232,In_794);
and U1135 (N_1135,In_309,In_693);
nand U1136 (N_1136,In_420,In_494);
and U1137 (N_1137,In_751,In_270);
and U1138 (N_1138,In_901,In_119);
nand U1139 (N_1139,In_50,In_538);
nand U1140 (N_1140,In_649,In_826);
and U1141 (N_1141,In_447,In_490);
and U1142 (N_1142,In_731,In_739);
or U1143 (N_1143,In_510,In_189);
and U1144 (N_1144,In_799,In_113);
and U1145 (N_1145,In_893,In_269);
nor U1146 (N_1146,In_917,In_522);
nor U1147 (N_1147,In_291,In_510);
nor U1148 (N_1148,In_866,In_885);
nand U1149 (N_1149,In_830,In_214);
nand U1150 (N_1150,In_430,In_341);
and U1151 (N_1151,In_160,In_907);
xor U1152 (N_1152,In_370,In_201);
nor U1153 (N_1153,In_604,In_964);
nor U1154 (N_1154,In_239,In_636);
nor U1155 (N_1155,In_480,In_569);
and U1156 (N_1156,In_561,In_977);
nand U1157 (N_1157,In_355,In_450);
or U1158 (N_1158,In_71,In_96);
nand U1159 (N_1159,In_76,In_269);
and U1160 (N_1160,In_209,In_425);
nor U1161 (N_1161,In_907,In_209);
and U1162 (N_1162,In_562,In_169);
or U1163 (N_1163,In_696,In_102);
and U1164 (N_1164,In_391,In_858);
and U1165 (N_1165,In_332,In_660);
nor U1166 (N_1166,In_629,In_657);
or U1167 (N_1167,In_840,In_84);
and U1168 (N_1168,In_152,In_760);
and U1169 (N_1169,In_466,In_943);
nand U1170 (N_1170,In_382,In_408);
nand U1171 (N_1171,In_769,In_14);
and U1172 (N_1172,In_948,In_982);
nand U1173 (N_1173,In_215,In_481);
or U1174 (N_1174,In_350,In_158);
nand U1175 (N_1175,In_581,In_578);
and U1176 (N_1176,In_764,In_431);
or U1177 (N_1177,In_614,In_656);
and U1178 (N_1178,In_736,In_409);
nor U1179 (N_1179,In_392,In_386);
and U1180 (N_1180,In_978,In_996);
nand U1181 (N_1181,In_868,In_34);
nand U1182 (N_1182,In_554,In_701);
nand U1183 (N_1183,In_559,In_63);
xnor U1184 (N_1184,In_529,In_776);
nand U1185 (N_1185,In_476,In_110);
nand U1186 (N_1186,In_274,In_158);
nor U1187 (N_1187,In_794,In_222);
and U1188 (N_1188,In_787,In_194);
and U1189 (N_1189,In_318,In_881);
nand U1190 (N_1190,In_62,In_467);
nand U1191 (N_1191,In_22,In_589);
nand U1192 (N_1192,In_460,In_145);
or U1193 (N_1193,In_51,In_800);
and U1194 (N_1194,In_723,In_968);
nand U1195 (N_1195,In_938,In_380);
and U1196 (N_1196,In_271,In_754);
or U1197 (N_1197,In_235,In_294);
xor U1198 (N_1198,In_504,In_53);
nand U1199 (N_1199,In_902,In_219);
nor U1200 (N_1200,In_997,In_817);
and U1201 (N_1201,In_680,In_904);
or U1202 (N_1202,In_870,In_536);
nor U1203 (N_1203,In_17,In_598);
or U1204 (N_1204,In_641,In_198);
nand U1205 (N_1205,In_54,In_110);
nand U1206 (N_1206,In_108,In_244);
or U1207 (N_1207,In_267,In_886);
or U1208 (N_1208,In_428,In_726);
and U1209 (N_1209,In_223,In_811);
nand U1210 (N_1210,In_678,In_830);
or U1211 (N_1211,In_890,In_796);
nand U1212 (N_1212,In_649,In_46);
nand U1213 (N_1213,In_822,In_260);
nor U1214 (N_1214,In_969,In_683);
nand U1215 (N_1215,In_450,In_304);
nor U1216 (N_1216,In_114,In_445);
nor U1217 (N_1217,In_907,In_455);
nor U1218 (N_1218,In_473,In_882);
nor U1219 (N_1219,In_233,In_809);
or U1220 (N_1220,In_96,In_182);
nand U1221 (N_1221,In_256,In_433);
or U1222 (N_1222,In_557,In_789);
and U1223 (N_1223,In_536,In_474);
or U1224 (N_1224,In_313,In_332);
nor U1225 (N_1225,In_792,In_257);
nor U1226 (N_1226,In_332,In_1);
or U1227 (N_1227,In_839,In_713);
nor U1228 (N_1228,In_619,In_92);
nand U1229 (N_1229,In_199,In_311);
nand U1230 (N_1230,In_201,In_337);
or U1231 (N_1231,In_799,In_251);
nor U1232 (N_1232,In_691,In_650);
and U1233 (N_1233,In_396,In_883);
or U1234 (N_1234,In_197,In_641);
nand U1235 (N_1235,In_240,In_771);
nor U1236 (N_1236,In_655,In_343);
and U1237 (N_1237,In_643,In_543);
and U1238 (N_1238,In_742,In_881);
nand U1239 (N_1239,In_783,In_944);
nor U1240 (N_1240,In_39,In_896);
xor U1241 (N_1241,In_159,In_155);
nand U1242 (N_1242,In_52,In_323);
nor U1243 (N_1243,In_135,In_512);
nand U1244 (N_1244,In_863,In_453);
or U1245 (N_1245,In_188,In_372);
nand U1246 (N_1246,In_695,In_882);
nand U1247 (N_1247,In_283,In_256);
and U1248 (N_1248,In_758,In_0);
and U1249 (N_1249,In_946,In_722);
nand U1250 (N_1250,In_356,In_911);
or U1251 (N_1251,In_980,In_405);
nand U1252 (N_1252,In_495,In_328);
or U1253 (N_1253,In_889,In_746);
or U1254 (N_1254,In_646,In_717);
and U1255 (N_1255,In_62,In_807);
and U1256 (N_1256,In_471,In_213);
nor U1257 (N_1257,In_898,In_644);
or U1258 (N_1258,In_803,In_180);
nor U1259 (N_1259,In_711,In_837);
and U1260 (N_1260,In_317,In_459);
nand U1261 (N_1261,In_755,In_646);
nand U1262 (N_1262,In_266,In_799);
nor U1263 (N_1263,In_670,In_854);
and U1264 (N_1264,In_274,In_593);
or U1265 (N_1265,In_784,In_752);
or U1266 (N_1266,In_234,In_507);
nor U1267 (N_1267,In_122,In_812);
nand U1268 (N_1268,In_450,In_629);
or U1269 (N_1269,In_45,In_310);
or U1270 (N_1270,In_453,In_634);
and U1271 (N_1271,In_604,In_736);
or U1272 (N_1272,In_214,In_291);
or U1273 (N_1273,In_435,In_177);
nand U1274 (N_1274,In_678,In_348);
or U1275 (N_1275,In_109,In_695);
or U1276 (N_1276,In_44,In_599);
nor U1277 (N_1277,In_358,In_58);
nor U1278 (N_1278,In_29,In_894);
nand U1279 (N_1279,In_159,In_405);
nor U1280 (N_1280,In_681,In_442);
nor U1281 (N_1281,In_841,In_469);
or U1282 (N_1282,In_191,In_332);
and U1283 (N_1283,In_64,In_252);
or U1284 (N_1284,In_651,In_759);
nor U1285 (N_1285,In_186,In_177);
nor U1286 (N_1286,In_964,In_350);
nor U1287 (N_1287,In_642,In_985);
or U1288 (N_1288,In_25,In_51);
nand U1289 (N_1289,In_90,In_311);
and U1290 (N_1290,In_633,In_929);
or U1291 (N_1291,In_103,In_125);
or U1292 (N_1292,In_526,In_342);
nor U1293 (N_1293,In_392,In_360);
and U1294 (N_1294,In_171,In_912);
nor U1295 (N_1295,In_131,In_143);
nand U1296 (N_1296,In_242,In_659);
and U1297 (N_1297,In_284,In_952);
nor U1298 (N_1298,In_943,In_122);
nand U1299 (N_1299,In_121,In_972);
or U1300 (N_1300,In_152,In_945);
or U1301 (N_1301,In_321,In_189);
nor U1302 (N_1302,In_597,In_305);
xor U1303 (N_1303,In_925,In_668);
and U1304 (N_1304,In_824,In_316);
nor U1305 (N_1305,In_91,In_974);
nor U1306 (N_1306,In_247,In_836);
nand U1307 (N_1307,In_829,In_324);
nor U1308 (N_1308,In_236,In_584);
nor U1309 (N_1309,In_24,In_877);
or U1310 (N_1310,In_186,In_662);
or U1311 (N_1311,In_149,In_660);
nor U1312 (N_1312,In_681,In_166);
nand U1313 (N_1313,In_565,In_977);
or U1314 (N_1314,In_3,In_481);
and U1315 (N_1315,In_525,In_824);
and U1316 (N_1316,In_44,In_142);
nor U1317 (N_1317,In_674,In_52);
nor U1318 (N_1318,In_328,In_446);
nand U1319 (N_1319,In_94,In_645);
xor U1320 (N_1320,In_643,In_228);
nor U1321 (N_1321,In_150,In_652);
or U1322 (N_1322,In_999,In_55);
nand U1323 (N_1323,In_930,In_374);
and U1324 (N_1324,In_103,In_274);
nor U1325 (N_1325,In_36,In_84);
and U1326 (N_1326,In_110,In_136);
nand U1327 (N_1327,In_632,In_564);
or U1328 (N_1328,In_641,In_552);
nor U1329 (N_1329,In_893,In_939);
nand U1330 (N_1330,In_992,In_188);
nand U1331 (N_1331,In_472,In_51);
nor U1332 (N_1332,In_1,In_988);
or U1333 (N_1333,In_806,In_486);
or U1334 (N_1334,In_193,In_600);
nand U1335 (N_1335,In_67,In_911);
nor U1336 (N_1336,In_175,In_592);
nor U1337 (N_1337,In_278,In_598);
nor U1338 (N_1338,In_469,In_72);
nand U1339 (N_1339,In_552,In_313);
nand U1340 (N_1340,In_110,In_178);
nor U1341 (N_1341,In_753,In_488);
or U1342 (N_1342,In_331,In_913);
nor U1343 (N_1343,In_171,In_855);
nor U1344 (N_1344,In_413,In_601);
and U1345 (N_1345,In_56,In_461);
and U1346 (N_1346,In_4,In_493);
and U1347 (N_1347,In_226,In_520);
or U1348 (N_1348,In_358,In_763);
and U1349 (N_1349,In_920,In_573);
or U1350 (N_1350,In_316,In_237);
nor U1351 (N_1351,In_437,In_413);
nor U1352 (N_1352,In_765,In_159);
nor U1353 (N_1353,In_718,In_169);
nor U1354 (N_1354,In_582,In_615);
and U1355 (N_1355,In_358,In_45);
nor U1356 (N_1356,In_964,In_732);
nor U1357 (N_1357,In_570,In_660);
and U1358 (N_1358,In_97,In_563);
and U1359 (N_1359,In_90,In_709);
or U1360 (N_1360,In_830,In_886);
or U1361 (N_1361,In_939,In_682);
nor U1362 (N_1362,In_867,In_704);
xnor U1363 (N_1363,In_686,In_225);
nor U1364 (N_1364,In_975,In_457);
and U1365 (N_1365,In_823,In_909);
nand U1366 (N_1366,In_101,In_652);
and U1367 (N_1367,In_663,In_2);
or U1368 (N_1368,In_559,In_953);
and U1369 (N_1369,In_373,In_287);
and U1370 (N_1370,In_569,In_209);
nand U1371 (N_1371,In_278,In_901);
or U1372 (N_1372,In_538,In_748);
nor U1373 (N_1373,In_753,In_211);
nor U1374 (N_1374,In_821,In_134);
nand U1375 (N_1375,In_564,In_15);
nand U1376 (N_1376,In_699,In_112);
nor U1377 (N_1377,In_752,In_486);
nand U1378 (N_1378,In_661,In_38);
and U1379 (N_1379,In_693,In_520);
nand U1380 (N_1380,In_939,In_82);
or U1381 (N_1381,In_964,In_494);
or U1382 (N_1382,In_685,In_914);
and U1383 (N_1383,In_419,In_575);
and U1384 (N_1384,In_360,In_940);
or U1385 (N_1385,In_53,In_355);
nor U1386 (N_1386,In_200,In_626);
nand U1387 (N_1387,In_727,In_738);
nor U1388 (N_1388,In_612,In_190);
nor U1389 (N_1389,In_607,In_787);
nor U1390 (N_1390,In_925,In_67);
xnor U1391 (N_1391,In_879,In_609);
nand U1392 (N_1392,In_690,In_429);
or U1393 (N_1393,In_259,In_186);
or U1394 (N_1394,In_388,In_506);
nor U1395 (N_1395,In_168,In_99);
nor U1396 (N_1396,In_51,In_419);
nand U1397 (N_1397,In_696,In_13);
or U1398 (N_1398,In_263,In_699);
nor U1399 (N_1399,In_374,In_787);
or U1400 (N_1400,In_672,In_738);
or U1401 (N_1401,In_264,In_183);
or U1402 (N_1402,In_395,In_571);
or U1403 (N_1403,In_721,In_824);
or U1404 (N_1404,In_731,In_280);
nor U1405 (N_1405,In_130,In_439);
or U1406 (N_1406,In_104,In_491);
and U1407 (N_1407,In_203,In_634);
nand U1408 (N_1408,In_722,In_346);
nand U1409 (N_1409,In_363,In_935);
and U1410 (N_1410,In_831,In_33);
nor U1411 (N_1411,In_560,In_863);
nor U1412 (N_1412,In_494,In_4);
nor U1413 (N_1413,In_469,In_837);
and U1414 (N_1414,In_512,In_60);
nand U1415 (N_1415,In_251,In_163);
nand U1416 (N_1416,In_183,In_944);
nor U1417 (N_1417,In_214,In_550);
and U1418 (N_1418,In_926,In_719);
nor U1419 (N_1419,In_246,In_516);
nor U1420 (N_1420,In_901,In_205);
or U1421 (N_1421,In_353,In_259);
and U1422 (N_1422,In_24,In_314);
or U1423 (N_1423,In_995,In_890);
or U1424 (N_1424,In_703,In_276);
nand U1425 (N_1425,In_800,In_265);
nand U1426 (N_1426,In_994,In_114);
or U1427 (N_1427,In_23,In_195);
and U1428 (N_1428,In_113,In_15);
and U1429 (N_1429,In_357,In_622);
nand U1430 (N_1430,In_225,In_479);
and U1431 (N_1431,In_206,In_673);
nand U1432 (N_1432,In_809,In_497);
nor U1433 (N_1433,In_325,In_58);
nor U1434 (N_1434,In_784,In_114);
nand U1435 (N_1435,In_638,In_510);
nor U1436 (N_1436,In_69,In_264);
or U1437 (N_1437,In_726,In_125);
nand U1438 (N_1438,In_621,In_801);
nor U1439 (N_1439,In_690,In_156);
or U1440 (N_1440,In_863,In_237);
nor U1441 (N_1441,In_625,In_388);
or U1442 (N_1442,In_786,In_608);
and U1443 (N_1443,In_993,In_215);
or U1444 (N_1444,In_142,In_222);
or U1445 (N_1445,In_496,In_694);
nand U1446 (N_1446,In_835,In_475);
or U1447 (N_1447,In_606,In_83);
and U1448 (N_1448,In_144,In_363);
nor U1449 (N_1449,In_693,In_536);
nor U1450 (N_1450,In_115,In_578);
nand U1451 (N_1451,In_862,In_365);
or U1452 (N_1452,In_27,In_425);
nor U1453 (N_1453,In_535,In_632);
and U1454 (N_1454,In_976,In_396);
nand U1455 (N_1455,In_7,In_77);
or U1456 (N_1456,In_507,In_75);
nor U1457 (N_1457,In_317,In_164);
nor U1458 (N_1458,In_849,In_191);
and U1459 (N_1459,In_728,In_915);
nand U1460 (N_1460,In_188,In_832);
xor U1461 (N_1461,In_124,In_794);
nor U1462 (N_1462,In_626,In_68);
and U1463 (N_1463,In_882,In_431);
or U1464 (N_1464,In_489,In_711);
and U1465 (N_1465,In_490,In_963);
nand U1466 (N_1466,In_538,In_457);
nor U1467 (N_1467,In_308,In_107);
nor U1468 (N_1468,In_680,In_560);
nand U1469 (N_1469,In_232,In_400);
nand U1470 (N_1470,In_456,In_852);
nand U1471 (N_1471,In_236,In_565);
or U1472 (N_1472,In_983,In_483);
nand U1473 (N_1473,In_641,In_154);
nor U1474 (N_1474,In_111,In_716);
nor U1475 (N_1475,In_680,In_440);
nand U1476 (N_1476,In_531,In_109);
nand U1477 (N_1477,In_921,In_726);
nor U1478 (N_1478,In_259,In_362);
nand U1479 (N_1479,In_794,In_95);
or U1480 (N_1480,In_948,In_647);
and U1481 (N_1481,In_841,In_11);
and U1482 (N_1482,In_196,In_518);
xor U1483 (N_1483,In_342,In_360);
or U1484 (N_1484,In_196,In_198);
nand U1485 (N_1485,In_257,In_729);
or U1486 (N_1486,In_793,In_689);
nor U1487 (N_1487,In_938,In_696);
or U1488 (N_1488,In_721,In_851);
nand U1489 (N_1489,In_381,In_11);
nand U1490 (N_1490,In_212,In_70);
nor U1491 (N_1491,In_529,In_769);
or U1492 (N_1492,In_858,In_208);
nand U1493 (N_1493,In_461,In_262);
and U1494 (N_1494,In_390,In_171);
nor U1495 (N_1495,In_411,In_487);
and U1496 (N_1496,In_194,In_825);
xor U1497 (N_1497,In_425,In_24);
and U1498 (N_1498,In_603,In_794);
and U1499 (N_1499,In_713,In_236);
or U1500 (N_1500,In_454,In_988);
nand U1501 (N_1501,In_536,In_607);
or U1502 (N_1502,In_86,In_855);
nand U1503 (N_1503,In_269,In_616);
or U1504 (N_1504,In_868,In_6);
and U1505 (N_1505,In_474,In_243);
or U1506 (N_1506,In_783,In_570);
and U1507 (N_1507,In_269,In_519);
nand U1508 (N_1508,In_921,In_822);
or U1509 (N_1509,In_597,In_178);
or U1510 (N_1510,In_797,In_420);
nor U1511 (N_1511,In_696,In_111);
or U1512 (N_1512,In_52,In_620);
nor U1513 (N_1513,In_487,In_936);
nand U1514 (N_1514,In_155,In_675);
or U1515 (N_1515,In_704,In_70);
or U1516 (N_1516,In_743,In_87);
nor U1517 (N_1517,In_455,In_18);
nor U1518 (N_1518,In_963,In_728);
and U1519 (N_1519,In_635,In_843);
nor U1520 (N_1520,In_846,In_826);
nor U1521 (N_1521,In_171,In_112);
and U1522 (N_1522,In_452,In_371);
nor U1523 (N_1523,In_64,In_25);
xor U1524 (N_1524,In_171,In_109);
and U1525 (N_1525,In_392,In_152);
nand U1526 (N_1526,In_720,In_104);
nor U1527 (N_1527,In_55,In_221);
or U1528 (N_1528,In_797,In_107);
or U1529 (N_1529,In_757,In_67);
or U1530 (N_1530,In_184,In_321);
and U1531 (N_1531,In_199,In_265);
and U1532 (N_1532,In_286,In_431);
or U1533 (N_1533,In_283,In_925);
nand U1534 (N_1534,In_750,In_763);
nor U1535 (N_1535,In_433,In_385);
nor U1536 (N_1536,In_968,In_89);
nor U1537 (N_1537,In_994,In_91);
and U1538 (N_1538,In_454,In_300);
nand U1539 (N_1539,In_185,In_434);
or U1540 (N_1540,In_910,In_588);
or U1541 (N_1541,In_267,In_167);
nand U1542 (N_1542,In_294,In_277);
nor U1543 (N_1543,In_801,In_95);
or U1544 (N_1544,In_429,In_247);
nand U1545 (N_1545,In_683,In_682);
nor U1546 (N_1546,In_870,In_228);
nor U1547 (N_1547,In_93,In_407);
and U1548 (N_1548,In_148,In_8);
nor U1549 (N_1549,In_945,In_636);
nand U1550 (N_1550,In_174,In_310);
nor U1551 (N_1551,In_925,In_335);
and U1552 (N_1552,In_327,In_933);
or U1553 (N_1553,In_327,In_275);
and U1554 (N_1554,In_559,In_40);
nand U1555 (N_1555,In_79,In_226);
nand U1556 (N_1556,In_349,In_204);
nor U1557 (N_1557,In_2,In_44);
or U1558 (N_1558,In_547,In_368);
nand U1559 (N_1559,In_775,In_333);
nand U1560 (N_1560,In_167,In_161);
nor U1561 (N_1561,In_691,In_699);
nor U1562 (N_1562,In_738,In_72);
nor U1563 (N_1563,In_835,In_862);
and U1564 (N_1564,In_906,In_416);
and U1565 (N_1565,In_423,In_138);
xnor U1566 (N_1566,In_60,In_349);
and U1567 (N_1567,In_698,In_996);
and U1568 (N_1568,In_949,In_54);
and U1569 (N_1569,In_300,In_774);
or U1570 (N_1570,In_434,In_972);
and U1571 (N_1571,In_505,In_801);
nor U1572 (N_1572,In_168,In_152);
nand U1573 (N_1573,In_175,In_385);
nor U1574 (N_1574,In_807,In_642);
or U1575 (N_1575,In_832,In_984);
and U1576 (N_1576,In_36,In_880);
or U1577 (N_1577,In_181,In_182);
nor U1578 (N_1578,In_165,In_690);
or U1579 (N_1579,In_660,In_553);
nor U1580 (N_1580,In_763,In_478);
and U1581 (N_1581,In_957,In_860);
and U1582 (N_1582,In_410,In_56);
nor U1583 (N_1583,In_833,In_45);
and U1584 (N_1584,In_468,In_203);
and U1585 (N_1585,In_232,In_206);
and U1586 (N_1586,In_645,In_817);
nand U1587 (N_1587,In_593,In_474);
nor U1588 (N_1588,In_944,In_977);
nor U1589 (N_1589,In_432,In_176);
nor U1590 (N_1590,In_510,In_775);
nand U1591 (N_1591,In_947,In_96);
or U1592 (N_1592,In_368,In_566);
and U1593 (N_1593,In_774,In_464);
nand U1594 (N_1594,In_880,In_982);
nand U1595 (N_1595,In_118,In_549);
or U1596 (N_1596,In_447,In_489);
nand U1597 (N_1597,In_213,In_302);
nand U1598 (N_1598,In_234,In_812);
nor U1599 (N_1599,In_199,In_180);
nor U1600 (N_1600,In_654,In_741);
nand U1601 (N_1601,In_296,In_403);
or U1602 (N_1602,In_770,In_959);
nor U1603 (N_1603,In_474,In_283);
nand U1604 (N_1604,In_713,In_1);
or U1605 (N_1605,In_931,In_599);
or U1606 (N_1606,In_546,In_269);
nand U1607 (N_1607,In_109,In_970);
nor U1608 (N_1608,In_751,In_144);
nand U1609 (N_1609,In_168,In_762);
or U1610 (N_1610,In_247,In_246);
nor U1611 (N_1611,In_161,In_173);
nor U1612 (N_1612,In_706,In_285);
nand U1613 (N_1613,In_342,In_610);
or U1614 (N_1614,In_712,In_292);
nand U1615 (N_1615,In_770,In_958);
nand U1616 (N_1616,In_744,In_114);
nor U1617 (N_1617,In_514,In_832);
nand U1618 (N_1618,In_340,In_540);
or U1619 (N_1619,In_802,In_750);
or U1620 (N_1620,In_355,In_757);
nor U1621 (N_1621,In_134,In_861);
or U1622 (N_1622,In_596,In_835);
and U1623 (N_1623,In_375,In_251);
nand U1624 (N_1624,In_433,In_251);
nor U1625 (N_1625,In_574,In_635);
or U1626 (N_1626,In_18,In_99);
and U1627 (N_1627,In_567,In_214);
nand U1628 (N_1628,In_273,In_30);
and U1629 (N_1629,In_850,In_865);
nor U1630 (N_1630,In_853,In_829);
and U1631 (N_1631,In_391,In_365);
and U1632 (N_1632,In_504,In_696);
nor U1633 (N_1633,In_935,In_640);
or U1634 (N_1634,In_707,In_449);
nand U1635 (N_1635,In_59,In_465);
nand U1636 (N_1636,In_584,In_114);
nor U1637 (N_1637,In_900,In_361);
and U1638 (N_1638,In_506,In_380);
and U1639 (N_1639,In_40,In_842);
and U1640 (N_1640,In_669,In_735);
nor U1641 (N_1641,In_236,In_446);
xor U1642 (N_1642,In_751,In_957);
nand U1643 (N_1643,In_576,In_44);
or U1644 (N_1644,In_685,In_944);
nand U1645 (N_1645,In_766,In_827);
nand U1646 (N_1646,In_192,In_909);
or U1647 (N_1647,In_802,In_440);
xor U1648 (N_1648,In_275,In_786);
nand U1649 (N_1649,In_346,In_383);
and U1650 (N_1650,In_149,In_932);
nand U1651 (N_1651,In_582,In_1);
nand U1652 (N_1652,In_448,In_891);
xnor U1653 (N_1653,In_610,In_521);
nor U1654 (N_1654,In_165,In_835);
nand U1655 (N_1655,In_863,In_976);
and U1656 (N_1656,In_376,In_249);
nor U1657 (N_1657,In_267,In_441);
nor U1658 (N_1658,In_527,In_749);
nor U1659 (N_1659,In_762,In_402);
nor U1660 (N_1660,In_292,In_199);
and U1661 (N_1661,In_251,In_116);
or U1662 (N_1662,In_886,In_799);
or U1663 (N_1663,In_524,In_549);
and U1664 (N_1664,In_697,In_191);
and U1665 (N_1665,In_101,In_506);
nor U1666 (N_1666,In_771,In_60);
or U1667 (N_1667,In_459,In_721);
and U1668 (N_1668,In_828,In_675);
and U1669 (N_1669,In_219,In_190);
or U1670 (N_1670,In_83,In_873);
or U1671 (N_1671,In_770,In_364);
nand U1672 (N_1672,In_770,In_707);
nand U1673 (N_1673,In_780,In_757);
or U1674 (N_1674,In_864,In_866);
nor U1675 (N_1675,In_911,In_974);
nor U1676 (N_1676,In_394,In_453);
or U1677 (N_1677,In_411,In_344);
and U1678 (N_1678,In_250,In_411);
or U1679 (N_1679,In_138,In_150);
and U1680 (N_1680,In_61,In_439);
nand U1681 (N_1681,In_786,In_767);
or U1682 (N_1682,In_982,In_607);
and U1683 (N_1683,In_30,In_719);
and U1684 (N_1684,In_466,In_338);
and U1685 (N_1685,In_407,In_289);
nand U1686 (N_1686,In_703,In_899);
nor U1687 (N_1687,In_393,In_420);
nand U1688 (N_1688,In_924,In_635);
nor U1689 (N_1689,In_10,In_744);
nor U1690 (N_1690,In_676,In_491);
nor U1691 (N_1691,In_965,In_399);
nand U1692 (N_1692,In_390,In_355);
nor U1693 (N_1693,In_574,In_794);
nand U1694 (N_1694,In_307,In_578);
nand U1695 (N_1695,In_204,In_656);
nor U1696 (N_1696,In_158,In_368);
nor U1697 (N_1697,In_387,In_532);
xor U1698 (N_1698,In_619,In_771);
and U1699 (N_1699,In_897,In_824);
nor U1700 (N_1700,In_627,In_99);
or U1701 (N_1701,In_425,In_337);
and U1702 (N_1702,In_813,In_176);
or U1703 (N_1703,In_802,In_614);
nor U1704 (N_1704,In_402,In_937);
nand U1705 (N_1705,In_432,In_434);
nor U1706 (N_1706,In_36,In_219);
or U1707 (N_1707,In_349,In_614);
nor U1708 (N_1708,In_575,In_9);
and U1709 (N_1709,In_224,In_315);
or U1710 (N_1710,In_456,In_221);
and U1711 (N_1711,In_969,In_882);
or U1712 (N_1712,In_899,In_93);
and U1713 (N_1713,In_85,In_169);
nand U1714 (N_1714,In_794,In_423);
nand U1715 (N_1715,In_226,In_669);
nor U1716 (N_1716,In_90,In_708);
nand U1717 (N_1717,In_945,In_263);
and U1718 (N_1718,In_904,In_84);
nor U1719 (N_1719,In_658,In_789);
or U1720 (N_1720,In_905,In_646);
or U1721 (N_1721,In_423,In_874);
nor U1722 (N_1722,In_1,In_967);
nor U1723 (N_1723,In_221,In_97);
nand U1724 (N_1724,In_749,In_758);
or U1725 (N_1725,In_836,In_855);
nor U1726 (N_1726,In_981,In_697);
or U1727 (N_1727,In_449,In_309);
and U1728 (N_1728,In_806,In_815);
nand U1729 (N_1729,In_425,In_147);
nor U1730 (N_1730,In_952,In_405);
or U1731 (N_1731,In_60,In_49);
nand U1732 (N_1732,In_212,In_740);
nor U1733 (N_1733,In_142,In_475);
xor U1734 (N_1734,In_627,In_799);
nand U1735 (N_1735,In_717,In_782);
nand U1736 (N_1736,In_876,In_925);
nor U1737 (N_1737,In_818,In_405);
or U1738 (N_1738,In_664,In_244);
and U1739 (N_1739,In_341,In_342);
and U1740 (N_1740,In_973,In_413);
and U1741 (N_1741,In_590,In_38);
and U1742 (N_1742,In_510,In_57);
or U1743 (N_1743,In_127,In_46);
and U1744 (N_1744,In_942,In_755);
nand U1745 (N_1745,In_563,In_844);
or U1746 (N_1746,In_624,In_237);
nor U1747 (N_1747,In_980,In_495);
nand U1748 (N_1748,In_9,In_693);
or U1749 (N_1749,In_778,In_293);
or U1750 (N_1750,In_600,In_41);
nand U1751 (N_1751,In_762,In_260);
or U1752 (N_1752,In_959,In_418);
or U1753 (N_1753,In_255,In_279);
or U1754 (N_1754,In_730,In_22);
nor U1755 (N_1755,In_72,In_23);
nor U1756 (N_1756,In_236,In_753);
or U1757 (N_1757,In_813,In_916);
and U1758 (N_1758,In_419,In_944);
and U1759 (N_1759,In_811,In_333);
nor U1760 (N_1760,In_451,In_368);
and U1761 (N_1761,In_830,In_999);
nand U1762 (N_1762,In_480,In_888);
or U1763 (N_1763,In_657,In_363);
or U1764 (N_1764,In_492,In_465);
nand U1765 (N_1765,In_820,In_341);
nor U1766 (N_1766,In_170,In_582);
and U1767 (N_1767,In_853,In_404);
and U1768 (N_1768,In_95,In_854);
nor U1769 (N_1769,In_686,In_496);
or U1770 (N_1770,In_139,In_547);
nand U1771 (N_1771,In_887,In_634);
nand U1772 (N_1772,In_782,In_741);
nor U1773 (N_1773,In_586,In_879);
nor U1774 (N_1774,In_911,In_837);
or U1775 (N_1775,In_412,In_922);
and U1776 (N_1776,In_125,In_295);
or U1777 (N_1777,In_9,In_967);
or U1778 (N_1778,In_344,In_815);
nand U1779 (N_1779,In_31,In_899);
or U1780 (N_1780,In_576,In_36);
and U1781 (N_1781,In_863,In_292);
and U1782 (N_1782,In_436,In_501);
or U1783 (N_1783,In_941,In_73);
and U1784 (N_1784,In_747,In_115);
or U1785 (N_1785,In_764,In_15);
nor U1786 (N_1786,In_719,In_24);
or U1787 (N_1787,In_432,In_237);
nand U1788 (N_1788,In_556,In_664);
nor U1789 (N_1789,In_538,In_834);
and U1790 (N_1790,In_405,In_492);
or U1791 (N_1791,In_385,In_409);
nor U1792 (N_1792,In_110,In_613);
or U1793 (N_1793,In_458,In_963);
xor U1794 (N_1794,In_140,In_718);
nand U1795 (N_1795,In_767,In_773);
xor U1796 (N_1796,In_553,In_133);
and U1797 (N_1797,In_412,In_168);
nor U1798 (N_1798,In_193,In_709);
and U1799 (N_1799,In_622,In_668);
and U1800 (N_1800,In_252,In_872);
nand U1801 (N_1801,In_108,In_166);
nor U1802 (N_1802,In_49,In_158);
nor U1803 (N_1803,In_409,In_850);
nand U1804 (N_1804,In_828,In_773);
or U1805 (N_1805,In_867,In_475);
or U1806 (N_1806,In_685,In_61);
nand U1807 (N_1807,In_276,In_241);
and U1808 (N_1808,In_780,In_689);
or U1809 (N_1809,In_536,In_809);
and U1810 (N_1810,In_821,In_37);
and U1811 (N_1811,In_213,In_388);
or U1812 (N_1812,In_358,In_360);
nor U1813 (N_1813,In_322,In_26);
nand U1814 (N_1814,In_551,In_731);
nand U1815 (N_1815,In_888,In_15);
nand U1816 (N_1816,In_226,In_676);
nand U1817 (N_1817,In_531,In_303);
and U1818 (N_1818,In_321,In_225);
nand U1819 (N_1819,In_859,In_932);
nor U1820 (N_1820,In_530,In_252);
nor U1821 (N_1821,In_665,In_681);
nor U1822 (N_1822,In_269,In_439);
nand U1823 (N_1823,In_181,In_183);
nand U1824 (N_1824,In_0,In_205);
and U1825 (N_1825,In_550,In_683);
nor U1826 (N_1826,In_739,In_46);
nand U1827 (N_1827,In_661,In_356);
and U1828 (N_1828,In_216,In_327);
and U1829 (N_1829,In_516,In_397);
or U1830 (N_1830,In_290,In_453);
nand U1831 (N_1831,In_309,In_280);
nor U1832 (N_1832,In_592,In_603);
nor U1833 (N_1833,In_695,In_402);
nand U1834 (N_1834,In_191,In_409);
nor U1835 (N_1835,In_270,In_891);
and U1836 (N_1836,In_252,In_478);
and U1837 (N_1837,In_322,In_665);
nor U1838 (N_1838,In_208,In_180);
and U1839 (N_1839,In_684,In_529);
and U1840 (N_1840,In_700,In_884);
nor U1841 (N_1841,In_282,In_883);
nand U1842 (N_1842,In_943,In_738);
and U1843 (N_1843,In_207,In_819);
and U1844 (N_1844,In_870,In_727);
nand U1845 (N_1845,In_594,In_442);
nand U1846 (N_1846,In_82,In_599);
nor U1847 (N_1847,In_331,In_127);
nand U1848 (N_1848,In_375,In_288);
nor U1849 (N_1849,In_58,In_895);
or U1850 (N_1850,In_738,In_930);
or U1851 (N_1851,In_935,In_168);
and U1852 (N_1852,In_405,In_191);
or U1853 (N_1853,In_563,In_242);
and U1854 (N_1854,In_734,In_454);
nand U1855 (N_1855,In_340,In_609);
nor U1856 (N_1856,In_922,In_236);
nand U1857 (N_1857,In_410,In_852);
and U1858 (N_1858,In_905,In_269);
nor U1859 (N_1859,In_325,In_459);
and U1860 (N_1860,In_812,In_64);
or U1861 (N_1861,In_55,In_915);
or U1862 (N_1862,In_38,In_906);
or U1863 (N_1863,In_212,In_222);
nand U1864 (N_1864,In_359,In_272);
or U1865 (N_1865,In_549,In_453);
or U1866 (N_1866,In_949,In_442);
nor U1867 (N_1867,In_745,In_342);
nand U1868 (N_1868,In_260,In_245);
nor U1869 (N_1869,In_657,In_53);
or U1870 (N_1870,In_123,In_651);
or U1871 (N_1871,In_300,In_236);
or U1872 (N_1872,In_8,In_876);
or U1873 (N_1873,In_649,In_588);
or U1874 (N_1874,In_196,In_550);
or U1875 (N_1875,In_773,In_732);
and U1876 (N_1876,In_475,In_78);
or U1877 (N_1877,In_823,In_234);
nand U1878 (N_1878,In_462,In_642);
nor U1879 (N_1879,In_436,In_836);
nor U1880 (N_1880,In_494,In_763);
nor U1881 (N_1881,In_462,In_630);
and U1882 (N_1882,In_792,In_749);
nand U1883 (N_1883,In_463,In_348);
or U1884 (N_1884,In_303,In_904);
and U1885 (N_1885,In_668,In_721);
and U1886 (N_1886,In_872,In_201);
and U1887 (N_1887,In_803,In_735);
nand U1888 (N_1888,In_542,In_31);
or U1889 (N_1889,In_593,In_254);
or U1890 (N_1890,In_368,In_61);
nand U1891 (N_1891,In_515,In_507);
nor U1892 (N_1892,In_35,In_300);
or U1893 (N_1893,In_333,In_595);
nand U1894 (N_1894,In_661,In_268);
nor U1895 (N_1895,In_675,In_972);
nor U1896 (N_1896,In_542,In_824);
nand U1897 (N_1897,In_249,In_870);
or U1898 (N_1898,In_943,In_291);
nand U1899 (N_1899,In_55,In_453);
nor U1900 (N_1900,In_463,In_549);
or U1901 (N_1901,In_463,In_77);
or U1902 (N_1902,In_375,In_119);
nand U1903 (N_1903,In_787,In_686);
and U1904 (N_1904,In_651,In_72);
or U1905 (N_1905,In_119,In_217);
or U1906 (N_1906,In_310,In_315);
nor U1907 (N_1907,In_475,In_889);
nand U1908 (N_1908,In_596,In_640);
xnor U1909 (N_1909,In_607,In_453);
nor U1910 (N_1910,In_90,In_105);
or U1911 (N_1911,In_784,In_43);
nor U1912 (N_1912,In_544,In_614);
nor U1913 (N_1913,In_976,In_721);
and U1914 (N_1914,In_906,In_956);
and U1915 (N_1915,In_962,In_984);
nor U1916 (N_1916,In_918,In_394);
or U1917 (N_1917,In_764,In_577);
or U1918 (N_1918,In_397,In_370);
nor U1919 (N_1919,In_593,In_478);
or U1920 (N_1920,In_327,In_592);
nor U1921 (N_1921,In_851,In_304);
nand U1922 (N_1922,In_967,In_643);
or U1923 (N_1923,In_948,In_759);
nor U1924 (N_1924,In_334,In_262);
nor U1925 (N_1925,In_855,In_354);
nor U1926 (N_1926,In_960,In_705);
or U1927 (N_1927,In_107,In_497);
or U1928 (N_1928,In_242,In_354);
and U1929 (N_1929,In_96,In_733);
nand U1930 (N_1930,In_204,In_255);
nand U1931 (N_1931,In_25,In_326);
nand U1932 (N_1932,In_709,In_972);
nor U1933 (N_1933,In_333,In_466);
nor U1934 (N_1934,In_592,In_335);
nand U1935 (N_1935,In_41,In_448);
and U1936 (N_1936,In_784,In_773);
and U1937 (N_1937,In_413,In_818);
or U1938 (N_1938,In_614,In_255);
nor U1939 (N_1939,In_839,In_715);
nor U1940 (N_1940,In_65,In_156);
nand U1941 (N_1941,In_743,In_995);
or U1942 (N_1942,In_606,In_389);
nand U1943 (N_1943,In_386,In_614);
and U1944 (N_1944,In_772,In_497);
or U1945 (N_1945,In_510,In_984);
and U1946 (N_1946,In_828,In_263);
nor U1947 (N_1947,In_439,In_751);
and U1948 (N_1948,In_945,In_350);
or U1949 (N_1949,In_994,In_475);
or U1950 (N_1950,In_405,In_296);
nand U1951 (N_1951,In_626,In_480);
nand U1952 (N_1952,In_147,In_43);
and U1953 (N_1953,In_652,In_887);
and U1954 (N_1954,In_3,In_782);
or U1955 (N_1955,In_613,In_911);
xnor U1956 (N_1956,In_22,In_23);
nand U1957 (N_1957,In_867,In_852);
nor U1958 (N_1958,In_294,In_572);
and U1959 (N_1959,In_814,In_124);
and U1960 (N_1960,In_489,In_160);
nor U1961 (N_1961,In_760,In_800);
nand U1962 (N_1962,In_711,In_464);
nand U1963 (N_1963,In_80,In_331);
nand U1964 (N_1964,In_117,In_342);
and U1965 (N_1965,In_22,In_881);
or U1966 (N_1966,In_709,In_197);
nand U1967 (N_1967,In_608,In_280);
or U1968 (N_1968,In_388,In_4);
or U1969 (N_1969,In_884,In_397);
nand U1970 (N_1970,In_190,In_802);
or U1971 (N_1971,In_598,In_793);
or U1972 (N_1972,In_840,In_196);
nor U1973 (N_1973,In_853,In_464);
and U1974 (N_1974,In_555,In_783);
and U1975 (N_1975,In_802,In_981);
or U1976 (N_1976,In_462,In_951);
nor U1977 (N_1977,In_815,In_713);
and U1978 (N_1978,In_106,In_963);
nor U1979 (N_1979,In_389,In_379);
or U1980 (N_1980,In_648,In_554);
nor U1981 (N_1981,In_653,In_196);
and U1982 (N_1982,In_636,In_161);
nand U1983 (N_1983,In_421,In_114);
or U1984 (N_1984,In_911,In_405);
and U1985 (N_1985,In_45,In_48);
and U1986 (N_1986,In_570,In_163);
nor U1987 (N_1987,In_354,In_439);
nor U1988 (N_1988,In_709,In_649);
nand U1989 (N_1989,In_726,In_92);
or U1990 (N_1990,In_197,In_568);
nor U1991 (N_1991,In_855,In_393);
nand U1992 (N_1992,In_15,In_922);
nor U1993 (N_1993,In_346,In_480);
nor U1994 (N_1994,In_452,In_276);
nand U1995 (N_1995,In_745,In_528);
or U1996 (N_1996,In_420,In_328);
and U1997 (N_1997,In_392,In_764);
or U1998 (N_1998,In_740,In_182);
nor U1999 (N_1999,In_604,In_481);
nor U2000 (N_2000,N_1233,N_1074);
or U2001 (N_2001,N_1031,N_1001);
or U2002 (N_2002,N_648,N_952);
or U2003 (N_2003,N_692,N_91);
or U2004 (N_2004,N_1399,N_1280);
nand U2005 (N_2005,N_75,N_1323);
nand U2006 (N_2006,N_611,N_12);
or U2007 (N_2007,N_118,N_1558);
and U2008 (N_2008,N_745,N_921);
nor U2009 (N_2009,N_869,N_1746);
and U2010 (N_2010,N_136,N_1624);
or U2011 (N_2011,N_553,N_749);
nand U2012 (N_2012,N_899,N_1146);
or U2013 (N_2013,N_1204,N_7);
or U2014 (N_2014,N_284,N_432);
nor U2015 (N_2015,N_659,N_1852);
or U2016 (N_2016,N_768,N_199);
or U2017 (N_2017,N_1125,N_86);
or U2018 (N_2018,N_1467,N_951);
and U2019 (N_2019,N_1457,N_1231);
nand U2020 (N_2020,N_1207,N_1798);
nor U2021 (N_2021,N_841,N_57);
nor U2022 (N_2022,N_273,N_1637);
or U2023 (N_2023,N_891,N_1550);
nor U2024 (N_2024,N_558,N_1082);
nand U2025 (N_2025,N_218,N_1754);
nor U2026 (N_2026,N_664,N_1839);
nor U2027 (N_2027,N_998,N_303);
nor U2028 (N_2028,N_1854,N_783);
nor U2029 (N_2029,N_819,N_446);
and U2030 (N_2030,N_120,N_1608);
or U2031 (N_2031,N_409,N_366);
or U2032 (N_2032,N_777,N_95);
nor U2033 (N_2033,N_1153,N_1017);
nand U2034 (N_2034,N_438,N_593);
or U2035 (N_2035,N_1961,N_1616);
nand U2036 (N_2036,N_333,N_1236);
nor U2037 (N_2037,N_50,N_1592);
and U2038 (N_2038,N_309,N_1142);
nand U2039 (N_2039,N_197,N_1588);
nor U2040 (N_2040,N_954,N_536);
or U2041 (N_2041,N_1325,N_1032);
nor U2042 (N_2042,N_1685,N_272);
nor U2043 (N_2043,N_792,N_1516);
xnor U2044 (N_2044,N_1393,N_299);
nand U2045 (N_2045,N_762,N_4);
or U2046 (N_2046,N_658,N_669);
nand U2047 (N_2047,N_1450,N_1473);
or U2048 (N_2048,N_565,N_349);
and U2049 (N_2049,N_1828,N_1098);
nor U2050 (N_2050,N_425,N_936);
nand U2051 (N_2051,N_1010,N_1361);
or U2052 (N_2052,N_494,N_1617);
nor U2053 (N_2053,N_958,N_256);
nor U2054 (N_2054,N_401,N_1070);
or U2055 (N_2055,N_1799,N_1573);
nor U2056 (N_2056,N_101,N_149);
nor U2057 (N_2057,N_719,N_1876);
and U2058 (N_2058,N_380,N_1477);
nor U2059 (N_2059,N_627,N_1108);
nor U2060 (N_2060,N_205,N_1865);
and U2061 (N_2061,N_329,N_962);
nand U2062 (N_2062,N_1003,N_1537);
nand U2063 (N_2063,N_571,N_595);
nor U2064 (N_2064,N_18,N_1829);
or U2065 (N_2065,N_1981,N_532);
or U2066 (N_2066,N_1226,N_377);
and U2067 (N_2067,N_1715,N_1520);
nor U2068 (N_2068,N_235,N_867);
nor U2069 (N_2069,N_1980,N_1000);
nand U2070 (N_2070,N_1175,N_1733);
or U2071 (N_2071,N_1436,N_112);
nor U2072 (N_2072,N_142,N_1814);
and U2073 (N_2073,N_392,N_1205);
nor U2074 (N_2074,N_105,N_29);
nor U2075 (N_2075,N_1111,N_1760);
nand U2076 (N_2076,N_1122,N_1986);
and U2077 (N_2077,N_297,N_448);
nor U2078 (N_2078,N_816,N_1210);
nand U2079 (N_2079,N_96,N_1044);
nor U2080 (N_2080,N_1970,N_73);
nor U2081 (N_2081,N_64,N_1194);
nand U2082 (N_2082,N_1405,N_798);
or U2083 (N_2083,N_1818,N_1651);
nand U2084 (N_2084,N_422,N_430);
and U2085 (N_2085,N_797,N_516);
nand U2086 (N_2086,N_300,N_1306);
or U2087 (N_2087,N_471,N_524);
nor U2088 (N_2088,N_1109,N_382);
and U2089 (N_2089,N_594,N_323);
nor U2090 (N_2090,N_1193,N_1340);
nor U2091 (N_2091,N_296,N_1638);
nand U2092 (N_2092,N_1895,N_770);
nand U2093 (N_2093,N_42,N_772);
or U2094 (N_2094,N_561,N_132);
and U2095 (N_2095,N_855,N_1305);
and U2096 (N_2096,N_193,N_1565);
nand U2097 (N_2097,N_1392,N_1902);
nand U2098 (N_2098,N_625,N_647);
nand U2099 (N_2099,N_356,N_201);
or U2100 (N_2100,N_1162,N_367);
nand U2101 (N_2101,N_252,N_1297);
and U2102 (N_2102,N_1947,N_599);
nor U2103 (N_2103,N_1525,N_321);
and U2104 (N_2104,N_1052,N_1);
and U2105 (N_2105,N_181,N_937);
or U2106 (N_2106,N_383,N_1159);
nor U2107 (N_2107,N_906,N_884);
nor U2108 (N_2108,N_1374,N_1335);
or U2109 (N_2109,N_1315,N_1078);
or U2110 (N_2110,N_874,N_589);
nand U2111 (N_2111,N_1647,N_742);
and U2112 (N_2112,N_1282,N_165);
or U2113 (N_2113,N_932,N_945);
and U2114 (N_2114,N_1502,N_51);
and U2115 (N_2115,N_262,N_959);
and U2116 (N_2116,N_693,N_600);
nand U2117 (N_2117,N_172,N_1290);
or U2118 (N_2118,N_925,N_1882);
nor U2119 (N_2119,N_387,N_144);
or U2120 (N_2120,N_102,N_1932);
nor U2121 (N_2121,N_1948,N_280);
and U2122 (N_2122,N_1061,N_702);
or U2123 (N_2123,N_1443,N_452);
or U2124 (N_2124,N_1698,N_1751);
or U2125 (N_2125,N_501,N_1889);
nor U2126 (N_2126,N_1339,N_766);
and U2127 (N_2127,N_705,N_1632);
nor U2128 (N_2128,N_90,N_621);
or U2129 (N_2129,N_98,N_1807);
nand U2130 (N_2130,N_89,N_1049);
nand U2131 (N_2131,N_1256,N_1939);
nand U2132 (N_2132,N_944,N_1904);
nor U2133 (N_2133,N_93,N_228);
or U2134 (N_2134,N_1154,N_1777);
nand U2135 (N_2135,N_1776,N_721);
nor U2136 (N_2136,N_601,N_1300);
nand U2137 (N_2137,N_365,N_288);
or U2138 (N_2138,N_1999,N_439);
nand U2139 (N_2139,N_1097,N_580);
or U2140 (N_2140,N_68,N_1806);
xnor U2141 (N_2141,N_1303,N_1195);
nand U2142 (N_2142,N_1934,N_1984);
nand U2143 (N_2143,N_1844,N_1090);
nor U2144 (N_2144,N_750,N_755);
nor U2145 (N_2145,N_794,N_1433);
and U2146 (N_2146,N_1164,N_110);
nand U2147 (N_2147,N_618,N_1182);
nand U2148 (N_2148,N_1873,N_1222);
and U2149 (N_2149,N_576,N_332);
or U2150 (N_2150,N_191,N_1042);
nor U2151 (N_2151,N_930,N_1350);
nor U2152 (N_2152,N_1369,N_1650);
or U2153 (N_2153,N_1148,N_258);
and U2154 (N_2154,N_1134,N_390);
nand U2155 (N_2155,N_700,N_24);
nor U2156 (N_2156,N_1772,N_718);
and U2157 (N_2157,N_1228,N_1230);
nor U2158 (N_2158,N_904,N_1302);
nand U2159 (N_2159,N_623,N_1783);
nor U2160 (N_2160,N_1587,N_1495);
nand U2161 (N_2161,N_963,N_1756);
and U2162 (N_2162,N_1121,N_1428);
and U2163 (N_2163,N_374,N_735);
nor U2164 (N_2164,N_973,N_1219);
or U2165 (N_2165,N_699,N_1454);
and U2166 (N_2166,N_863,N_982);
and U2167 (N_2167,N_1908,N_396);
nand U2168 (N_2168,N_1972,N_327);
nand U2169 (N_2169,N_606,N_1956);
or U2170 (N_2170,N_1684,N_531);
nand U2171 (N_2171,N_1370,N_1503);
or U2172 (N_2172,N_1140,N_796);
nor U2173 (N_2173,N_1825,N_852);
nand U2174 (N_2174,N_1376,N_1349);
and U2175 (N_2175,N_1869,N_1860);
and U2176 (N_2176,N_955,N_1364);
nand U2177 (N_2177,N_1830,N_469);
nor U2178 (N_2178,N_1625,N_666);
nor U2179 (N_2179,N_1215,N_1800);
nor U2180 (N_2180,N_1585,N_1644);
or U2181 (N_2181,N_1729,N_1365);
or U2182 (N_2182,N_754,N_302);
nor U2183 (N_2183,N_966,N_1711);
or U2184 (N_2184,N_1921,N_736);
nor U2185 (N_2185,N_984,N_49);
or U2186 (N_2186,N_1749,N_1107);
nor U2187 (N_2187,N_506,N_1385);
and U2188 (N_2188,N_1978,N_1106);
or U2189 (N_2189,N_17,N_1328);
or U2190 (N_2190,N_876,N_1655);
and U2191 (N_2191,N_1621,N_1778);
nor U2192 (N_2192,N_1064,N_979);
nor U2193 (N_2193,N_441,N_362);
or U2194 (N_2194,N_1092,N_1117);
nor U2195 (N_2195,N_1192,N_1264);
nand U2196 (N_2196,N_459,N_243);
nand U2197 (N_2197,N_306,N_637);
nand U2198 (N_2198,N_1036,N_1639);
and U2199 (N_2199,N_141,N_389);
nand U2200 (N_2200,N_1133,N_368);
and U2201 (N_2201,N_759,N_1909);
and U2202 (N_2202,N_1102,N_1517);
or U2203 (N_2203,N_166,N_725);
nor U2204 (N_2204,N_1419,N_1787);
nor U2205 (N_2205,N_1029,N_1629);
and U2206 (N_2206,N_1314,N_215);
or U2207 (N_2207,N_312,N_915);
nand U2208 (N_2208,N_214,N_511);
and U2209 (N_2209,N_1991,N_484);
nand U2210 (N_2210,N_890,N_939);
nand U2211 (N_2211,N_938,N_655);
nand U2212 (N_2212,N_1281,N_1835);
nor U2213 (N_2213,N_1618,N_866);
xor U2214 (N_2214,N_613,N_1610);
or U2215 (N_2215,N_1131,N_348);
and U2216 (N_2216,N_1352,N_480);
and U2217 (N_2217,N_224,N_1212);
nor U2218 (N_2218,N_1809,N_328);
or U2219 (N_2219,N_1220,N_851);
nor U2220 (N_2220,N_602,N_240);
or U2221 (N_2221,N_1506,N_85);
nor U2222 (N_2222,N_1678,N_1261);
nor U2223 (N_2223,N_1084,N_1706);
nor U2224 (N_2224,N_1757,N_1487);
and U2225 (N_2225,N_1721,N_198);
and U2226 (N_2226,N_1145,N_1864);
nor U2227 (N_2227,N_1270,N_400);
and U2228 (N_2228,N_879,N_1578);
or U2229 (N_2229,N_882,N_342);
or U2230 (N_2230,N_6,N_1077);
nand U2231 (N_2231,N_130,N_126);
nand U2232 (N_2232,N_801,N_1200);
or U2233 (N_2233,N_933,N_61);
and U2234 (N_2234,N_834,N_405);
nor U2235 (N_2235,N_947,N_60);
and U2236 (N_2236,N_1132,N_626);
or U2237 (N_2237,N_838,N_275);
nand U2238 (N_2238,N_1663,N_496);
nand U2239 (N_2239,N_1626,N_435);
nand U2240 (N_2240,N_358,N_1460);
nor U2241 (N_2241,N_1899,N_317);
nor U2242 (N_2242,N_386,N_1671);
and U2243 (N_2243,N_1701,N_1358);
nand U2244 (N_2244,N_1732,N_1482);
or U2245 (N_2245,N_147,N_1408);
nand U2246 (N_2246,N_344,N_927);
or U2247 (N_2247,N_1485,N_523);
nor U2248 (N_2248,N_253,N_758);
nand U2249 (N_2249,N_311,N_960);
nand U2250 (N_2250,N_802,N_825);
and U2251 (N_2251,N_340,N_1054);
nor U2252 (N_2252,N_1166,N_1542);
or U2253 (N_2253,N_740,N_76);
or U2254 (N_2254,N_1967,N_1951);
or U2255 (N_2255,N_1556,N_1875);
or U2256 (N_2256,N_1417,N_1890);
and U2257 (N_2257,N_1263,N_832);
or U2258 (N_2258,N_1813,N_1406);
nand U2259 (N_2259,N_835,N_31);
nor U2260 (N_2260,N_1815,N_1535);
or U2261 (N_2261,N_1901,N_1836);
nand U2262 (N_2262,N_1905,N_950);
and U2263 (N_2263,N_1498,N_1891);
nand U2264 (N_2264,N_1319,N_1345);
and U2265 (N_2265,N_52,N_722);
and U2266 (N_2266,N_175,N_799);
and U2267 (N_2267,N_461,N_139);
or U2268 (N_2268,N_1730,N_167);
or U2269 (N_2269,N_483,N_83);
nand U2270 (N_2270,N_818,N_1619);
and U2271 (N_2271,N_528,N_514);
and U2272 (N_2272,N_1938,N_212);
nand U2273 (N_2273,N_1603,N_334);
nand U2274 (N_2274,N_1085,N_1634);
and U2275 (N_2275,N_360,N_809);
or U2276 (N_2276,N_1026,N_503);
nor U2277 (N_2277,N_1229,N_1747);
nor U2278 (N_2278,N_887,N_847);
and U2279 (N_2279,N_630,N_972);
and U2280 (N_2280,N_1313,N_378);
or U2281 (N_2281,N_1130,N_196);
and U2282 (N_2282,N_238,N_1718);
xor U2283 (N_2283,N_1686,N_478);
nor U2284 (N_2284,N_182,N_793);
nor U2285 (N_2285,N_1301,N_1447);
nor U2286 (N_2286,N_550,N_65);
nor U2287 (N_2287,N_447,N_1700);
or U2288 (N_2288,N_1737,N_1180);
xor U2289 (N_2289,N_1926,N_1083);
nand U2290 (N_2290,N_71,N_460);
or U2291 (N_2291,N_579,N_369);
or U2292 (N_2292,N_981,N_814);
or U2293 (N_2293,N_522,N_632);
nand U2294 (N_2294,N_720,N_1595);
and U2295 (N_2295,N_1812,N_433);
or U2296 (N_2296,N_1652,N_319);
and U2297 (N_2297,N_1395,N_1023);
nor U2298 (N_2298,N_1123,N_1753);
and U2299 (N_2299,N_956,N_1043);
and U2300 (N_2300,N_1653,N_268);
or U2301 (N_2301,N_22,N_227);
and U2302 (N_2302,N_495,N_1019);
nand U2303 (N_2303,N_418,N_928);
nor U2304 (N_2304,N_2,N_989);
or U2305 (N_2305,N_1524,N_677);
nand U2306 (N_2306,N_1690,N_190);
nor U2307 (N_2307,N_10,N_1296);
and U2308 (N_2308,N_246,N_210);
nor U2309 (N_2309,N_121,N_1260);
and U2310 (N_2310,N_335,N_1742);
nand U2311 (N_2311,N_774,N_1002);
and U2312 (N_2312,N_80,N_644);
and U2313 (N_2313,N_153,N_1845);
and U2314 (N_2314,N_1360,N_208);
nor U2315 (N_2315,N_990,N_505);
and U2316 (N_2316,N_865,N_1894);
or U2317 (N_2317,N_1068,N_1705);
or U2318 (N_2318,N_1526,N_787);
or U2319 (N_2319,N_1834,N_1147);
nand U2320 (N_2320,N_204,N_1509);
or U2321 (N_2321,N_341,N_231);
or U2322 (N_2322,N_1687,N_1602);
nand U2323 (N_2323,N_743,N_1615);
nor U2324 (N_2324,N_1251,N_1694);
xor U2325 (N_2325,N_780,N_128);
or U2326 (N_2326,N_1601,N_407);
nor U2327 (N_2327,N_1072,N_1295);
and U2328 (N_2328,N_1050,N_1943);
nand U2329 (N_2329,N_1548,N_487);
nor U2330 (N_2330,N_1470,N_1016);
or U2331 (N_2331,N_225,N_336);
and U2332 (N_2332,N_1824,N_1143);
or U2333 (N_2333,N_997,N_476);
nand U2334 (N_2334,N_1351,N_826);
or U2335 (N_2335,N_36,N_1493);
nand U2336 (N_2336,N_247,N_1481);
nand U2337 (N_2337,N_585,N_1129);
and U2338 (N_2338,N_14,N_1897);
and U2339 (N_2339,N_1197,N_1960);
nor U2340 (N_2340,N_479,N_1179);
or U2341 (N_2341,N_656,N_1623);
or U2342 (N_2342,N_1765,N_1555);
nand U2343 (N_2343,N_1088,N_1560);
and U2344 (N_2344,N_206,N_1309);
nor U2345 (N_2345,N_116,N_1288);
nand U2346 (N_2346,N_1381,N_1045);
or U2347 (N_2347,N_72,N_1124);
and U2348 (N_2348,N_267,N_1640);
nor U2349 (N_2349,N_1703,N_888);
nand U2350 (N_2350,N_1822,N_1386);
or U2351 (N_2351,N_1252,N_428);
or U2352 (N_2352,N_1681,N_1582);
and U2353 (N_2353,N_1713,N_1469);
and U2354 (N_2354,N_131,N_554);
or U2355 (N_2355,N_127,N_679);
and U2356 (N_2356,N_1564,N_604);
and U2357 (N_2357,N_1160,N_1505);
or U2358 (N_2358,N_1038,N_1680);
nor U2359 (N_2359,N_629,N_864);
nor U2360 (N_2360,N_1552,N_25);
nor U2361 (N_2361,N_1025,N_1674);
and U2362 (N_2362,N_1394,N_77);
or U2363 (N_2363,N_544,N_59);
nor U2364 (N_2364,N_412,N_397);
nand U2365 (N_2365,N_1677,N_1468);
or U2366 (N_2366,N_525,N_414);
and U2367 (N_2367,N_1923,N_1444);
and U2368 (N_2368,N_636,N_698);
nand U2369 (N_2369,N_1249,N_436);
and U2370 (N_2370,N_1420,N_1190);
xnor U2371 (N_2371,N_1633,N_1636);
and U2372 (N_2372,N_1048,N_1277);
and U2373 (N_2373,N_23,N_498);
nand U2374 (N_2374,N_1734,N_338);
nand U2375 (N_2375,N_1682,N_870);
nand U2376 (N_2376,N_949,N_194);
and U2377 (N_2377,N_1529,N_605);
nor U2378 (N_2378,N_1586,N_186);
xor U2379 (N_2379,N_1355,N_1372);
and U2380 (N_2380,N_1209,N_1488);
nor U2381 (N_2381,N_1356,N_1217);
or U2382 (N_2382,N_734,N_1719);
nor U2383 (N_2383,N_850,N_164);
or U2384 (N_2384,N_830,N_129);
or U2385 (N_2385,N_1780,N_1112);
nand U2386 (N_2386,N_1391,N_1187);
or U2387 (N_2387,N_970,N_1672);
and U2388 (N_2388,N_444,N_354);
nor U2389 (N_2389,N_538,N_1702);
nor U2390 (N_2390,N_491,N_1973);
nor U2391 (N_2391,N_1781,N_546);
nand U2392 (N_2392,N_1593,N_905);
and U2393 (N_2393,N_1475,N_583);
or U2394 (N_2394,N_508,N_1081);
or U2395 (N_2395,N_1243,N_1900);
nand U2396 (N_2396,N_1766,N_1887);
and U2397 (N_2397,N_1858,N_1942);
and U2398 (N_2398,N_1916,N_195);
nand U2399 (N_2399,N_289,N_1750);
and U2400 (N_2400,N_468,N_1008);
and U2401 (N_2401,N_1486,N_785);
nor U2402 (N_2402,N_1863,N_1874);
nor U2403 (N_2403,N_533,N_155);
or U2404 (N_2404,N_482,N_1463);
nor U2405 (N_2405,N_1992,N_1013);
or U2406 (N_2406,N_873,N_1594);
nand U2407 (N_2407,N_738,N_821);
nor U2408 (N_2408,N_1413,N_1318);
or U2409 (N_2409,N_107,N_1940);
or U2410 (N_2410,N_1389,N_1012);
and U2411 (N_2411,N_245,N_1530);
nor U2412 (N_2412,N_1483,N_615);
and U2413 (N_2413,N_1521,N_842);
nand U2414 (N_2414,N_1903,N_1794);
and U2415 (N_2415,N_466,N_363);
nor U2416 (N_2416,N_420,N_1040);
nand U2417 (N_2417,N_569,N_923);
nor U2418 (N_2418,N_1675,N_161);
and U2419 (N_2419,N_988,N_1138);
or U2420 (N_2420,N_1977,N_1095);
nor U2421 (N_2421,N_499,N_1218);
and U2422 (N_2422,N_1227,N_1359);
and U2423 (N_2423,N_207,N_472);
and U2424 (N_2424,N_34,N_1326);
and U2425 (N_2425,N_1067,N_761);
nor U2426 (N_2426,N_1993,N_1870);
nand U2427 (N_2427,N_1271,N_791);
nor U2428 (N_2428,N_1308,N_1259);
nor U2429 (N_2429,N_46,N_30);
and U2430 (N_2430,N_179,N_1518);
nand U2431 (N_2431,N_1738,N_1779);
or U2432 (N_2432,N_929,N_370);
and U2433 (N_2433,N_1811,N_1377);
and U2434 (N_2434,N_957,N_726);
nor U2435 (N_2435,N_764,N_1331);
or U2436 (N_2436,N_716,N_1871);
and U2437 (N_2437,N_1110,N_1557);
or U2438 (N_2438,N_507,N_470);
and U2439 (N_2439,N_900,N_1589);
or U2440 (N_2440,N_1802,N_410);
nor U2441 (N_2441,N_361,N_883);
and U2442 (N_2442,N_1312,N_114);
nor U2443 (N_2443,N_671,N_271);
nor U2444 (N_2444,N_1975,N_1466);
nand U2445 (N_2445,N_1071,N_1176);
and U2446 (N_2446,N_1775,N_730);
nor U2447 (N_2447,N_530,N_1248);
nor U2448 (N_2448,N_282,N_903);
or U2449 (N_2449,N_1559,N_1857);
and U2450 (N_2450,N_353,N_559);
or U2451 (N_2451,N_920,N_1425);
nand U2452 (N_2452,N_1646,N_1437);
nor U2453 (N_2453,N_1846,N_1816);
or U2454 (N_2454,N_385,N_1371);
nor U2455 (N_2455,N_678,N_1127);
nand U2456 (N_2456,N_1445,N_1832);
nor U2457 (N_2457,N_1158,N_1790);
and U2458 (N_2458,N_856,N_160);
nand U2459 (N_2459,N_1717,N_763);
and U2460 (N_2460,N_1722,N_324);
nor U2461 (N_2461,N_1688,N_1987);
and U2462 (N_2462,N_393,N_1404);
nor U2463 (N_2463,N_1744,N_1416);
nand U2464 (N_2464,N_1888,N_355);
nand U2465 (N_2465,N_1459,N_859);
or U2466 (N_2466,N_44,N_607);
and U2467 (N_2467,N_15,N_1104);
nand U2468 (N_2468,N_157,N_19);
or U2469 (N_2469,N_1808,N_1924);
and U2470 (N_2470,N_1329,N_628);
nand U2471 (N_2471,N_26,N_703);
and U2472 (N_2472,N_1171,N_1240);
or U2473 (N_2473,N_1198,N_1547);
and U2474 (N_2474,N_230,N_113);
or U2475 (N_2475,N_577,N_1635);
and U2476 (N_2476,N_1103,N_1069);
nand U2477 (N_2477,N_1597,N_1925);
nand U2478 (N_2478,N_610,N_226);
and U2479 (N_2479,N_1826,N_1527);
nand U2480 (N_2480,N_1429,N_169);
nor U2481 (N_2481,N_1402,N_1037);
or U2482 (N_2482,N_151,N_753);
nor U2483 (N_2483,N_485,N_20);
nor U2484 (N_2484,N_566,N_995);
and U2485 (N_2485,N_1930,N_570);
nor U2486 (N_2486,N_1910,N_712);
nand U2487 (N_2487,N_612,N_697);
nor U2488 (N_2488,N_1983,N_293);
or U2489 (N_2489,N_1289,N_1211);
nand U2490 (N_2490,N_964,N_564);
nand U2491 (N_2491,N_912,N_1245);
nand U2492 (N_2492,N_1431,N_901);
and U2493 (N_2493,N_1152,N_1819);
or U2494 (N_2494,N_1275,N_674);
nand U2495 (N_2495,N_251,N_156);
nand U2496 (N_2496,N_117,N_1771);
and U2497 (N_2497,N_1508,N_1380);
nand U2498 (N_2498,N_1763,N_1414);
or U2499 (N_2499,N_1950,N_1203);
and U2500 (N_2500,N_1494,N_134);
nor U2501 (N_2501,N_668,N_1994);
or U2502 (N_2502,N_213,N_539);
nand U2503 (N_2503,N_1174,N_1279);
and U2504 (N_2504,N_346,N_584);
nor U2505 (N_2505,N_931,N_1453);
nand U2506 (N_2506,N_1867,N_1434);
or U2507 (N_2507,N_176,N_1238);
and U2508 (N_2508,N_1390,N_54);
and U2509 (N_2509,N_270,N_880);
and U2510 (N_2510,N_608,N_689);
and U2511 (N_2511,N_1015,N_220);
and U2512 (N_2512,N_684,N_148);
nor U2513 (N_2513,N_1448,N_581);
or U2514 (N_2514,N_259,N_1810);
nand U2515 (N_2515,N_1528,N_1510);
and U2516 (N_2516,N_326,N_415);
and U2517 (N_2517,N_1267,N_1569);
or U2518 (N_2518,N_892,N_737);
and U2519 (N_2519,N_1163,N_279);
nand U2520 (N_2520,N_1662,N_3);
nor U2521 (N_2521,N_1630,N_1821);
nand U2522 (N_2522,N_653,N_1430);
nand U2523 (N_2523,N_1743,N_1499);
nor U2524 (N_2524,N_421,N_229);
nor U2525 (N_2525,N_1581,N_1605);
and U2526 (N_2526,N_776,N_1144);
and U2527 (N_2527,N_1611,N_371);
nor U2528 (N_2528,N_1424,N_926);
nand U2529 (N_2529,N_66,N_1196);
nand U2530 (N_2530,N_1051,N_352);
nand U2531 (N_2531,N_688,N_343);
or U2532 (N_2532,N_862,N_1886);
nand U2533 (N_2533,N_1161,N_1707);
nand U2534 (N_2534,N_649,N_1944);
xor U2535 (N_2535,N_1758,N_1561);
or U2536 (N_2536,N_1185,N_462);
nand U2537 (N_2537,N_1216,N_266);
or U2538 (N_2538,N_844,N_911);
nor U2539 (N_2539,N_846,N_886);
xor U2540 (N_2540,N_1149,N_1058);
or U2541 (N_2541,N_1206,N_244);
or U2542 (N_2542,N_1657,N_1156);
nor U2543 (N_2543,N_778,N_910);
or U2544 (N_2544,N_233,N_1100);
or U2545 (N_2545,N_1407,N_239);
or U2546 (N_2546,N_249,N_403);
nand U2547 (N_2547,N_74,N_1344);
and U2548 (N_2548,N_173,N_9);
or U2549 (N_2549,N_640,N_895);
and U2550 (N_2550,N_1188,N_1704);
or U2551 (N_2551,N_596,N_292);
or U2552 (N_2552,N_1935,N_1213);
nor U2553 (N_2553,N_893,N_1105);
and U2554 (N_2554,N_1612,N_1065);
nor U2555 (N_2555,N_202,N_1035);
and U2556 (N_2556,N_143,N_200);
nand U2557 (N_2557,N_38,N_769);
or U2558 (N_2558,N_1201,N_1965);
nor U2559 (N_2559,N_489,N_1645);
nand U2560 (N_2560,N_183,N_1803);
nor U2561 (N_2561,N_654,N_1540);
and U2562 (N_2562,N_1762,N_1337);
nand U2563 (N_2563,N_765,N_1293);
nor U2564 (N_2564,N_1917,N_1397);
nand U2565 (N_2565,N_1096,N_1307);
nand U2566 (N_2566,N_1872,N_376);
or U2567 (N_2567,N_1962,N_1665);
or U2568 (N_2568,N_616,N_394);
nand U2569 (N_2569,N_1541,N_1239);
and U2570 (N_2570,N_1330,N_236);
nand U2571 (N_2571,N_974,N_1480);
or U2572 (N_2572,N_1731,N_1667);
and U2573 (N_2573,N_1342,N_1141);
nand U2574 (N_2574,N_728,N_1773);
or U2575 (N_2575,N_1053,N_62);
nor U2576 (N_2576,N_1996,N_878);
nor U2577 (N_2577,N_1847,N_771);
or U2578 (N_2578,N_1668,N_1878);
nand U2579 (N_2579,N_1643,N_614);
nor U2580 (N_2580,N_449,N_1234);
nand U2581 (N_2581,N_543,N_481);
or U2582 (N_2582,N_1028,N_1063);
nand U2583 (N_2583,N_1449,N_1327);
nand U2584 (N_2584,N_806,N_1683);
nand U2585 (N_2585,N_283,N_1080);
nor U2586 (N_2586,N_680,N_1949);
nand U2587 (N_2587,N_1057,N_1348);
and U2588 (N_2588,N_250,N_609);
or U2589 (N_2589,N_81,N_124);
and U2590 (N_2590,N_667,N_1862);
nor U2591 (N_2591,N_330,N_681);
nor U2592 (N_2592,N_708,N_1184);
nor U2593 (N_2593,N_1739,N_1333);
nor U2594 (N_2594,N_103,N_1998);
nand U2595 (N_2595,N_913,N_1151);
nor U2596 (N_2596,N_1724,N_316);
and U2597 (N_2597,N_1907,N_1490);
and U2598 (N_2598,N_154,N_1186);
nand U2599 (N_2599,N_388,N_339);
nand U2600 (N_2600,N_1627,N_416);
or U2601 (N_2601,N_560,N_1850);
and U2602 (N_2602,N_1727,N_597);
nand U2603 (N_2603,N_1817,N_1136);
or U2604 (N_2604,N_187,N_696);
nor U2605 (N_2605,N_1840,N_917);
nand U2606 (N_2606,N_1367,N_909);
nand U2607 (N_2607,N_1849,N_756);
and U2608 (N_2608,N_1232,N_1982);
or U2609 (N_2609,N_170,N_545);
and U2610 (N_2610,N_1346,N_1060);
nand U2611 (N_2611,N_1580,N_1953);
nor U2612 (N_2612,N_706,N_1570);
nor U2613 (N_2613,N_1538,N_1266);
nand U2614 (N_2614,N_8,N_33);
nand U2615 (N_2615,N_463,N_714);
nor U2616 (N_2616,N_744,N_1423);
nand U2617 (N_2617,N_1958,N_375);
nor U2618 (N_2618,N_652,N_1021);
or U2619 (N_2619,N_94,N_216);
nor U2620 (N_2620,N_1047,N_1788);
nor U2621 (N_2621,N_1004,N_1446);
nand U2622 (N_2622,N_301,N_504);
nor U2623 (N_2623,N_805,N_492);
nor U2624 (N_2624,N_1091,N_1076);
nand U2625 (N_2625,N_1959,N_556);
nor U2626 (N_2626,N_1421,N_1379);
and U2627 (N_2627,N_1320,N_104);
or U2628 (N_2628,N_16,N_254);
or U2629 (N_2629,N_828,N_1856);
nand U2630 (N_2630,N_1411,N_234);
and U2631 (N_2631,N_635,N_519);
or U2632 (N_2632,N_1046,N_458);
or U2633 (N_2633,N_757,N_924);
and U2634 (N_2634,N_1725,N_70);
and U2635 (N_2635,N_1861,N_1491);
nand U2636 (N_2636,N_0,N_845);
nor U2637 (N_2637,N_1914,N_1403);
and U2638 (N_2638,N_582,N_137);
or U2639 (N_2639,N_817,N_717);
nor U2640 (N_2640,N_1041,N_100);
and U2641 (N_2641,N_820,N_1056);
and U2642 (N_2642,N_969,N_520);
and U2643 (N_2643,N_443,N_1575);
nor U2644 (N_2644,N_1604,N_1988);
nor U2645 (N_2645,N_1554,N_907);
nand U2646 (N_2646,N_450,N_265);
or U2647 (N_2647,N_633,N_1432);
or U2648 (N_2648,N_88,N_1929);
nor U2649 (N_2649,N_975,N_857);
and U2650 (N_2650,N_996,N_603);
or U2651 (N_2651,N_211,N_562);
nand U2652 (N_2652,N_808,N_1755);
nor U2653 (N_2653,N_588,N_639);
or U2654 (N_2654,N_1116,N_32);
nand U2655 (N_2655,N_1079,N_881);
nor U2656 (N_2656,N_1654,N_1534);
or U2657 (N_2657,N_1150,N_555);
nand U2658 (N_2658,N_1945,N_1985);
nor U2659 (N_2659,N_586,N_1317);
and U2660 (N_2660,N_1462,N_889);
or U2661 (N_2661,N_1033,N_1165);
xor U2662 (N_2662,N_434,N_417);
or U2663 (N_2663,N_406,N_1855);
nand U2664 (N_2664,N_1086,N_1512);
nor U2665 (N_2665,N_1388,N_1254);
nand U2666 (N_2666,N_1139,N_79);
or U2667 (N_2667,N_427,N_1484);
or U2668 (N_2668,N_1321,N_537);
and U2669 (N_2669,N_1795,N_307);
or U2670 (N_2670,N_624,N_978);
nand U2671 (N_2671,N_67,N_854);
nor U2672 (N_2672,N_1452,N_1439);
nor U2673 (N_2673,N_185,N_473);
nand U2674 (N_2674,N_779,N_1532);
or U2675 (N_2675,N_682,N_1697);
nand U2676 (N_2676,N_232,N_1474);
nand U2677 (N_2677,N_40,N_1954);
nand U2678 (N_2678,N_729,N_257);
or U2679 (N_2679,N_1338,N_1438);
or U2680 (N_2680,N_163,N_1455);
nand U2681 (N_2681,N_325,N_408);
nor U2682 (N_2682,N_971,N_295);
nand U2683 (N_2683,N_1400,N_1546);
nor U2684 (N_2684,N_665,N_518);
nor U2685 (N_2685,N_1155,N_1761);
nand U2686 (N_2686,N_1347,N_395);
nand U2687 (N_2687,N_1286,N_263);
and U2688 (N_2688,N_1062,N_976);
nor U2689 (N_2689,N_1927,N_592);
or U2690 (N_2690,N_1536,N_748);
xor U2691 (N_2691,N_58,N_1896);
or U2692 (N_2692,N_683,N_1189);
nor U2693 (N_2693,N_1115,N_713);
nor U2694 (N_2694,N_651,N_1128);
or U2695 (N_2695,N_1748,N_320);
nand U2696 (N_2696,N_831,N_529);
nand U2697 (N_2697,N_286,N_1093);
nor U2698 (N_2698,N_1691,N_123);
nor U2699 (N_2699,N_840,N_1368);
nor U2700 (N_2700,N_823,N_551);
nand U2701 (N_2701,N_357,N_475);
and U2702 (N_2702,N_1157,N_573);
and U2703 (N_2703,N_1656,N_310);
nor U2704 (N_2704,N_108,N_125);
nand U2705 (N_2705,N_782,N_1912);
or U2706 (N_2706,N_1375,N_1545);
and U2707 (N_2707,N_465,N_477);
or U2708 (N_2708,N_999,N_242);
or U2709 (N_2709,N_1968,N_1642);
and U2710 (N_2710,N_723,N_78);
nor U2711 (N_2711,N_1976,N_1168);
nor U2712 (N_2712,N_1514,N_1027);
nand U2713 (N_2713,N_35,N_1928);
nand U2714 (N_2714,N_221,N_1173);
xor U2715 (N_2715,N_37,N_1415);
nor U2716 (N_2716,N_1979,N_1571);
nand U2717 (N_2717,N_1241,N_1785);
nand U2718 (N_2718,N_1543,N_133);
nor U2719 (N_2719,N_1523,N_961);
or U2720 (N_2720,N_290,N_48);
and U2721 (N_2721,N_1820,N_1464);
nor U2722 (N_2722,N_1833,N_526);
nand U2723 (N_2723,N_1427,N_837);
nor U2724 (N_2724,N_1786,N_109);
nor U2725 (N_2725,N_1191,N_1292);
xnor U2726 (N_2726,N_453,N_724);
nand U2727 (N_2727,N_308,N_122);
and U2728 (N_2728,N_991,N_184);
or U2729 (N_2729,N_1114,N_457);
and U2730 (N_2730,N_294,N_953);
and U2731 (N_2731,N_687,N_1378);
or U2732 (N_2732,N_1649,N_1199);
and U2733 (N_2733,N_1039,N_1373);
and U2734 (N_2734,N_715,N_1387);
or U2735 (N_2735,N_350,N_359);
nor U2736 (N_2736,N_1770,N_1660);
nor U2737 (N_2737,N_853,N_784);
and U2738 (N_2738,N_135,N_285);
or U2739 (N_2739,N_535,N_241);
nor U2740 (N_2740,N_943,N_347);
and U2741 (N_2741,N_423,N_875);
nand U2742 (N_2742,N_948,N_1736);
nor U2743 (N_2743,N_1274,N_510);
nor U2744 (N_2744,N_1177,N_56);
and U2745 (N_2745,N_1244,N_99);
nand U2746 (N_2746,N_591,N_1262);
nand U2747 (N_2747,N_672,N_440);
nand U2748 (N_2748,N_1451,N_1250);
and U2749 (N_2749,N_1568,N_1366);
nand U2750 (N_2750,N_1515,N_1310);
and U2751 (N_2751,N_1007,N_399);
xnor U2752 (N_2752,N_455,N_643);
nand U2753 (N_2753,N_276,N_1183);
or U2754 (N_2754,N_1018,N_619);
or U2755 (N_2755,N_1119,N_1596);
or U2756 (N_2756,N_1752,N_1574);
nor U2757 (N_2757,N_552,N_381);
nand U2758 (N_2758,N_1458,N_1478);
nor U2759 (N_2759,N_1607,N_106);
nor U2760 (N_2760,N_1664,N_411);
and U2761 (N_2761,N_1997,N_351);
nand U2762 (N_2762,N_1963,N_1099);
nor U2763 (N_2763,N_965,N_790);
nor U2764 (N_2764,N_497,N_429);
nand U2765 (N_2765,N_897,N_490);
and U2766 (N_2766,N_1631,N_445);
nor U2767 (N_2767,N_1955,N_1952);
and U2768 (N_2768,N_1915,N_663);
nand U2769 (N_2769,N_1695,N_673);
and U2770 (N_2770,N_1767,N_217);
or U2771 (N_2771,N_860,N_1628);
nand U2772 (N_2772,N_1489,N_1492);
nor U2773 (N_2773,N_150,N_260);
or U2774 (N_2774,N_1606,N_833);
nand U2775 (N_2775,N_1693,N_1214);
nand U2776 (N_2776,N_1969,N_575);
and U2777 (N_2777,N_1911,N_788);
or U2778 (N_2778,N_189,N_1500);
and U2779 (N_2779,N_1465,N_209);
nand U2780 (N_2780,N_140,N_942);
nor U2781 (N_2781,N_812,N_807);
or U2782 (N_2782,N_527,N_1842);
nor U2783 (N_2783,N_675,N_1221);
and U2784 (N_2784,N_1409,N_919);
nand U2785 (N_2785,N_1471,N_1741);
or U2786 (N_2786,N_1577,N_836);
or U2787 (N_2787,N_1572,N_39);
and U2788 (N_2788,N_1827,N_1551);
and U2789 (N_2789,N_219,N_727);
or U2790 (N_2790,N_502,N_1782);
xor U2791 (N_2791,N_549,N_1880);
or U2792 (N_2792,N_41,N_1476);
nand U2793 (N_2793,N_1507,N_1181);
and U2794 (N_2794,N_1418,N_967);
and U2795 (N_2795,N_1708,N_1501);
or U2796 (N_2796,N_541,N_1172);
nor U2797 (N_2797,N_1410,N_872);
or U2798 (N_2798,N_437,N_898);
nand U2799 (N_2799,N_1030,N_1723);
nor U2800 (N_2800,N_1964,N_1531);
nand U2801 (N_2801,N_1576,N_620);
nand U2802 (N_2802,N_1225,N_1658);
nand U2803 (N_2803,N_542,N_322);
nand U2804 (N_2804,N_1539,N_398);
or U2805 (N_2805,N_1094,N_384);
or U2806 (N_2806,N_1620,N_431);
and U2807 (N_2807,N_1384,N_739);
or U2808 (N_2808,N_1696,N_1859);
or U2809 (N_2809,N_994,N_1728);
and U2810 (N_2810,N_1005,N_1247);
nor U2811 (N_2811,N_1357,N_1883);
or U2812 (N_2812,N_404,N_650);
nand U2813 (N_2813,N_424,N_747);
and U2814 (N_2814,N_1223,N_815);
nor U2815 (N_2815,N_1178,N_1941);
or U2816 (N_2816,N_908,N_1497);
and U2817 (N_2817,N_1669,N_1591);
nand U2818 (N_2818,N_264,N_1913);
nand U2819 (N_2819,N_1137,N_1269);
nor U2820 (N_2820,N_732,N_1922);
or U2821 (N_2821,N_733,N_426);
and U2822 (N_2822,N_980,N_983);
and U2823 (N_2823,N_1791,N_278);
nor U2824 (N_2824,N_1966,N_1268);
nand U2825 (N_2825,N_305,N_1258);
and U2826 (N_2826,N_97,N_902);
nand U2827 (N_2827,N_598,N_1278);
or U2828 (N_2828,N_115,N_1354);
or U2829 (N_2829,N_314,N_707);
or U2830 (N_2830,N_488,N_464);
nand U2831 (N_2831,N_1283,N_1974);
nand U2832 (N_2832,N_1257,N_1255);
nand U2833 (N_2833,N_1933,N_1881);
or U2834 (N_2834,N_1006,N_657);
nand U2835 (N_2835,N_1383,N_1562);
and U2836 (N_2836,N_391,N_1735);
nor U2837 (N_2837,N_709,N_1533);
or U2838 (N_2838,N_992,N_11);
and U2839 (N_2839,N_1971,N_567);
nor U2840 (N_2840,N_1920,N_171);
nor U2841 (N_2841,N_701,N_1590);
and U2842 (N_2842,N_1866,N_177);
and U2843 (N_2843,N_1287,N_1884);
or U2844 (N_2844,N_1563,N_1792);
and U2845 (N_2845,N_84,N_1298);
or U2846 (N_2846,N_287,N_746);
and U2847 (N_2847,N_1401,N_1709);
or U2848 (N_2848,N_638,N_1066);
and U2849 (N_2849,N_1479,N_1120);
nor U2850 (N_2850,N_1316,N_634);
and U2851 (N_2851,N_641,N_1022);
nor U2852 (N_2852,N_509,N_1324);
and U2853 (N_2853,N_1285,N_1726);
nand U2854 (N_2854,N_1237,N_617);
or U2855 (N_2855,N_1504,N_1622);
and U2856 (N_2856,N_1613,N_849);
or U2857 (N_2857,N_1838,N_1898);
or U2858 (N_2858,N_646,N_534);
or U2859 (N_2859,N_1055,N_1745);
or U2860 (N_2860,N_1396,N_548);
nand U2861 (N_2861,N_521,N_1600);
xor U2862 (N_2862,N_1990,N_1332);
and U2863 (N_2863,N_1831,N_690);
nand U2864 (N_2864,N_1566,N_1793);
nor U2865 (N_2865,N_1989,N_1273);
nor U2866 (N_2866,N_1801,N_789);
or U2867 (N_2867,N_1676,N_493);
nand U2868 (N_2868,N_804,N_313);
and U2869 (N_2869,N_1126,N_1456);
and U2870 (N_2870,N_188,N_1740);
nand U2871 (N_2871,N_572,N_858);
nor U2872 (N_2872,N_1336,N_1712);
nor U2873 (N_2873,N_1868,N_1522);
or U2874 (N_2874,N_1284,N_1720);
or U2875 (N_2875,N_1879,N_1246);
or U2876 (N_2876,N_1892,N_1253);
or U2877 (N_2877,N_985,N_1609);
nand U2878 (N_2878,N_590,N_1774);
and U2879 (N_2879,N_987,N_685);
nand U2880 (N_2880,N_43,N_1353);
or U2881 (N_2881,N_1797,N_517);
nor U2882 (N_2882,N_786,N_704);
or U2883 (N_2883,N_5,N_935);
nand U2884 (N_2884,N_304,N_711);
and U2885 (N_2885,N_1716,N_1011);
or U2886 (N_2886,N_364,N_500);
and U2887 (N_2887,N_1768,N_843);
nor U2888 (N_2888,N_547,N_486);
nor U2889 (N_2889,N_318,N_1435);
or U2890 (N_2890,N_810,N_145);
or U2891 (N_2891,N_540,N_1135);
and U2892 (N_2892,N_1599,N_419);
or U2893 (N_2893,N_803,N_1692);
and U2894 (N_2894,N_345,N_642);
nand U2895 (N_2895,N_1957,N_1304);
nor U2896 (N_2896,N_1995,N_373);
nor U2897 (N_2897,N_824,N_741);
nand U2898 (N_2898,N_1553,N_622);
nand U2899 (N_2899,N_1804,N_281);
and U2900 (N_2900,N_274,N_291);
nor U2901 (N_2901,N_92,N_918);
nand U2902 (N_2902,N_1614,N_1412);
or U2903 (N_2903,N_1841,N_1544);
and U2904 (N_2904,N_1322,N_45);
or U2905 (N_2905,N_1851,N_451);
or U2906 (N_2906,N_587,N_1937);
nand U2907 (N_2907,N_248,N_1343);
or U2908 (N_2908,N_1113,N_568);
nor U2909 (N_2909,N_152,N_28);
nand U2910 (N_2910,N_1689,N_1714);
nand U2911 (N_2911,N_1276,N_331);
or U2912 (N_2912,N_773,N_1759);
or U2913 (N_2913,N_1075,N_822);
nand U2914 (N_2914,N_1919,N_1059);
or U2915 (N_2915,N_1398,N_1764);
nand U2916 (N_2916,N_710,N_868);
or U2917 (N_2917,N_968,N_138);
nor U2918 (N_2918,N_467,N_203);
and U2919 (N_2919,N_752,N_1235);
nand U2920 (N_2920,N_1659,N_1224);
nor U2921 (N_2921,N_1598,N_1710);
and U2922 (N_2922,N_827,N_916);
and U2923 (N_2923,N_1641,N_237);
nand U2924 (N_2924,N_1020,N_1311);
nor U2925 (N_2925,N_1567,N_1073);
nor U2926 (N_2926,N_986,N_885);
nand U2927 (N_2927,N_848,N_934);
and U2928 (N_2928,N_795,N_1666);
or U2929 (N_2929,N_940,N_1784);
nand U2930 (N_2930,N_1877,N_174);
or U2931 (N_2931,N_1440,N_87);
nand U2932 (N_2932,N_1513,N_1848);
or U2933 (N_2933,N_660,N_1299);
nor U2934 (N_2934,N_1362,N_1422);
nand U2935 (N_2935,N_1024,N_563);
nor U2936 (N_2936,N_1472,N_1885);
or U2937 (N_2937,N_574,N_53);
nand U2938 (N_2938,N_1843,N_47);
nor U2939 (N_2939,N_298,N_1426);
nand U2940 (N_2940,N_21,N_686);
or U2941 (N_2941,N_670,N_800);
nand U2942 (N_2942,N_760,N_829);
or U2943 (N_2943,N_1679,N_277);
or U2944 (N_2944,N_557,N_1202);
or U2945 (N_2945,N_1118,N_337);
nand U2946 (N_2946,N_1579,N_1549);
nor U2947 (N_2947,N_55,N_1511);
or U2948 (N_2948,N_1014,N_662);
nand U2949 (N_2949,N_1789,N_695);
and U2950 (N_2950,N_1583,N_379);
nor U2951 (N_2951,N_1334,N_1584);
or U2952 (N_2952,N_1382,N_1461);
and U2953 (N_2953,N_162,N_261);
or U2954 (N_2954,N_1363,N_474);
and U2955 (N_2955,N_168,N_1272);
nand U2956 (N_2956,N_631,N_413);
and U2957 (N_2957,N_1661,N_442);
nor U2958 (N_2958,N_731,N_372);
and U2959 (N_2959,N_1699,N_781);
or U2960 (N_2960,N_946,N_1936);
nand U2961 (N_2961,N_861,N_63);
nand U2962 (N_2962,N_82,N_402);
or U2963 (N_2963,N_456,N_751);
nand U2964 (N_2964,N_1167,N_1294);
nor U2965 (N_2965,N_1034,N_178);
and U2966 (N_2966,N_839,N_111);
and U2967 (N_2967,N_1769,N_941);
or U2968 (N_2968,N_1906,N_158);
or U2969 (N_2969,N_1291,N_223);
and U2970 (N_2970,N_1009,N_1242);
nand U2971 (N_2971,N_513,N_269);
nor U2972 (N_2972,N_1170,N_1673);
or U2973 (N_2973,N_1796,N_255);
nand U2974 (N_2974,N_1441,N_914);
nand U2975 (N_2975,N_69,N_1101);
and U2976 (N_2976,N_515,N_811);
xnor U2977 (N_2977,N_578,N_1931);
nor U2978 (N_2978,N_645,N_993);
nand U2979 (N_2979,N_1089,N_1087);
and U2980 (N_2980,N_767,N_775);
nand U2981 (N_2981,N_894,N_222);
and U2982 (N_2982,N_512,N_813);
nand U2983 (N_2983,N_1496,N_1918);
and U2984 (N_2984,N_454,N_691);
or U2985 (N_2985,N_1823,N_1805);
or U2986 (N_2986,N_896,N_146);
xor U2987 (N_2987,N_1837,N_192);
and U2988 (N_2988,N_315,N_1853);
nor U2989 (N_2989,N_1208,N_877);
nor U2990 (N_2990,N_1893,N_1519);
and U2991 (N_2991,N_27,N_871);
nor U2992 (N_2992,N_1265,N_159);
nor U2993 (N_2993,N_977,N_1442);
nor U2994 (N_2994,N_13,N_1341);
or U2995 (N_2995,N_1169,N_1648);
nor U2996 (N_2996,N_922,N_676);
nand U2997 (N_2997,N_661,N_119);
or U2998 (N_2998,N_1946,N_1670);
and U2999 (N_2999,N_180,N_694);
or U3000 (N_3000,N_273,N_408);
nor U3001 (N_3001,N_366,N_1614);
or U3002 (N_3002,N_35,N_1669);
nor U3003 (N_3003,N_709,N_1653);
or U3004 (N_3004,N_1618,N_228);
and U3005 (N_3005,N_1633,N_1198);
or U3006 (N_3006,N_986,N_233);
and U3007 (N_3007,N_1037,N_1336);
nand U3008 (N_3008,N_819,N_623);
nor U3009 (N_3009,N_1433,N_662);
or U3010 (N_3010,N_1435,N_360);
nor U3011 (N_3011,N_1562,N_187);
or U3012 (N_3012,N_1487,N_552);
nand U3013 (N_3013,N_635,N_1699);
or U3014 (N_3014,N_350,N_85);
nor U3015 (N_3015,N_630,N_844);
and U3016 (N_3016,N_1640,N_1474);
and U3017 (N_3017,N_391,N_1985);
nand U3018 (N_3018,N_1956,N_1138);
nand U3019 (N_3019,N_1673,N_86);
and U3020 (N_3020,N_1584,N_1382);
nor U3021 (N_3021,N_1564,N_85);
or U3022 (N_3022,N_1557,N_1536);
xor U3023 (N_3023,N_19,N_424);
and U3024 (N_3024,N_573,N_376);
or U3025 (N_3025,N_1777,N_535);
nand U3026 (N_3026,N_616,N_1716);
nor U3027 (N_3027,N_968,N_1614);
and U3028 (N_3028,N_1047,N_378);
nand U3029 (N_3029,N_894,N_982);
and U3030 (N_3030,N_616,N_600);
and U3031 (N_3031,N_1427,N_1122);
and U3032 (N_3032,N_638,N_1073);
and U3033 (N_3033,N_668,N_197);
and U3034 (N_3034,N_848,N_1200);
nor U3035 (N_3035,N_1544,N_839);
and U3036 (N_3036,N_328,N_198);
or U3037 (N_3037,N_553,N_1358);
nand U3038 (N_3038,N_841,N_1796);
nand U3039 (N_3039,N_1716,N_886);
nand U3040 (N_3040,N_1265,N_437);
nor U3041 (N_3041,N_1411,N_729);
nand U3042 (N_3042,N_760,N_203);
nor U3043 (N_3043,N_884,N_1862);
and U3044 (N_3044,N_1843,N_153);
nor U3045 (N_3045,N_1871,N_881);
or U3046 (N_3046,N_407,N_1869);
nand U3047 (N_3047,N_289,N_1508);
or U3048 (N_3048,N_46,N_1684);
or U3049 (N_3049,N_441,N_1475);
and U3050 (N_3050,N_1090,N_663);
or U3051 (N_3051,N_586,N_348);
nor U3052 (N_3052,N_1128,N_951);
and U3053 (N_3053,N_1968,N_1289);
or U3054 (N_3054,N_233,N_108);
nand U3055 (N_3055,N_105,N_709);
or U3056 (N_3056,N_64,N_942);
or U3057 (N_3057,N_1792,N_836);
or U3058 (N_3058,N_794,N_519);
nor U3059 (N_3059,N_1965,N_962);
nor U3060 (N_3060,N_1546,N_1553);
nand U3061 (N_3061,N_1987,N_151);
and U3062 (N_3062,N_1954,N_526);
and U3063 (N_3063,N_550,N_250);
or U3064 (N_3064,N_1239,N_132);
or U3065 (N_3065,N_1849,N_1683);
nand U3066 (N_3066,N_310,N_1173);
or U3067 (N_3067,N_705,N_1982);
nand U3068 (N_3068,N_703,N_1508);
or U3069 (N_3069,N_691,N_1875);
or U3070 (N_3070,N_225,N_1459);
nor U3071 (N_3071,N_1366,N_580);
nor U3072 (N_3072,N_1580,N_1401);
nand U3073 (N_3073,N_1208,N_1628);
nor U3074 (N_3074,N_487,N_1300);
nand U3075 (N_3075,N_1872,N_738);
and U3076 (N_3076,N_1785,N_1210);
nand U3077 (N_3077,N_1013,N_825);
nand U3078 (N_3078,N_1242,N_345);
nor U3079 (N_3079,N_996,N_1417);
nand U3080 (N_3080,N_407,N_23);
nand U3081 (N_3081,N_1555,N_86);
and U3082 (N_3082,N_630,N_1620);
or U3083 (N_3083,N_175,N_1588);
nor U3084 (N_3084,N_1905,N_651);
or U3085 (N_3085,N_1067,N_722);
nand U3086 (N_3086,N_848,N_1390);
nand U3087 (N_3087,N_1412,N_1607);
nand U3088 (N_3088,N_729,N_1562);
or U3089 (N_3089,N_1929,N_689);
nor U3090 (N_3090,N_1220,N_978);
and U3091 (N_3091,N_1024,N_143);
nor U3092 (N_3092,N_1000,N_942);
nand U3093 (N_3093,N_1700,N_710);
and U3094 (N_3094,N_882,N_490);
nand U3095 (N_3095,N_171,N_316);
nor U3096 (N_3096,N_525,N_1228);
nand U3097 (N_3097,N_507,N_28);
and U3098 (N_3098,N_1134,N_178);
or U3099 (N_3099,N_323,N_951);
nand U3100 (N_3100,N_908,N_187);
nand U3101 (N_3101,N_1380,N_280);
or U3102 (N_3102,N_1173,N_1683);
or U3103 (N_3103,N_692,N_150);
nor U3104 (N_3104,N_1366,N_370);
nor U3105 (N_3105,N_634,N_1485);
and U3106 (N_3106,N_739,N_1326);
nand U3107 (N_3107,N_542,N_63);
nor U3108 (N_3108,N_1001,N_386);
nor U3109 (N_3109,N_1207,N_964);
nand U3110 (N_3110,N_1729,N_1337);
nor U3111 (N_3111,N_657,N_802);
or U3112 (N_3112,N_637,N_1606);
and U3113 (N_3113,N_418,N_1475);
nor U3114 (N_3114,N_691,N_1318);
nor U3115 (N_3115,N_1307,N_242);
and U3116 (N_3116,N_2,N_176);
nand U3117 (N_3117,N_579,N_1380);
nor U3118 (N_3118,N_1444,N_1856);
nand U3119 (N_3119,N_1844,N_478);
or U3120 (N_3120,N_1272,N_1717);
or U3121 (N_3121,N_835,N_1058);
nor U3122 (N_3122,N_258,N_1973);
and U3123 (N_3123,N_559,N_692);
and U3124 (N_3124,N_1247,N_276);
nor U3125 (N_3125,N_75,N_319);
nand U3126 (N_3126,N_942,N_1624);
nor U3127 (N_3127,N_1911,N_1671);
or U3128 (N_3128,N_223,N_946);
nor U3129 (N_3129,N_1615,N_1249);
nor U3130 (N_3130,N_257,N_549);
and U3131 (N_3131,N_812,N_770);
nor U3132 (N_3132,N_1678,N_1297);
or U3133 (N_3133,N_1704,N_569);
and U3134 (N_3134,N_220,N_756);
nand U3135 (N_3135,N_182,N_1395);
nand U3136 (N_3136,N_973,N_263);
nor U3137 (N_3137,N_1481,N_1336);
nor U3138 (N_3138,N_145,N_944);
and U3139 (N_3139,N_1253,N_243);
nor U3140 (N_3140,N_867,N_1025);
and U3141 (N_3141,N_432,N_937);
nor U3142 (N_3142,N_1660,N_1059);
or U3143 (N_3143,N_620,N_1131);
nand U3144 (N_3144,N_983,N_61);
or U3145 (N_3145,N_1533,N_886);
and U3146 (N_3146,N_46,N_315);
or U3147 (N_3147,N_1222,N_1731);
nor U3148 (N_3148,N_1419,N_233);
nand U3149 (N_3149,N_1402,N_677);
nor U3150 (N_3150,N_1358,N_1242);
nand U3151 (N_3151,N_1247,N_1524);
and U3152 (N_3152,N_1414,N_786);
and U3153 (N_3153,N_1680,N_1432);
or U3154 (N_3154,N_1679,N_1885);
nand U3155 (N_3155,N_1851,N_1837);
or U3156 (N_3156,N_1287,N_1810);
or U3157 (N_3157,N_1604,N_1000);
and U3158 (N_3158,N_1975,N_626);
and U3159 (N_3159,N_948,N_601);
nor U3160 (N_3160,N_1616,N_1167);
nor U3161 (N_3161,N_851,N_794);
or U3162 (N_3162,N_646,N_1152);
or U3163 (N_3163,N_345,N_533);
or U3164 (N_3164,N_1824,N_1015);
or U3165 (N_3165,N_51,N_1895);
and U3166 (N_3166,N_655,N_631);
nand U3167 (N_3167,N_1857,N_648);
and U3168 (N_3168,N_1022,N_134);
nor U3169 (N_3169,N_253,N_2);
or U3170 (N_3170,N_1535,N_615);
and U3171 (N_3171,N_50,N_1462);
or U3172 (N_3172,N_1838,N_1653);
or U3173 (N_3173,N_1276,N_1779);
or U3174 (N_3174,N_1331,N_818);
and U3175 (N_3175,N_1726,N_1674);
and U3176 (N_3176,N_259,N_1287);
nor U3177 (N_3177,N_1035,N_1615);
nand U3178 (N_3178,N_1118,N_799);
nor U3179 (N_3179,N_368,N_290);
nor U3180 (N_3180,N_1414,N_316);
and U3181 (N_3181,N_440,N_861);
nand U3182 (N_3182,N_324,N_975);
nand U3183 (N_3183,N_1245,N_1049);
nand U3184 (N_3184,N_47,N_593);
or U3185 (N_3185,N_1420,N_1492);
and U3186 (N_3186,N_435,N_35);
nor U3187 (N_3187,N_565,N_774);
nor U3188 (N_3188,N_1397,N_1840);
nor U3189 (N_3189,N_1993,N_1827);
and U3190 (N_3190,N_278,N_452);
nand U3191 (N_3191,N_1974,N_529);
nand U3192 (N_3192,N_35,N_1672);
and U3193 (N_3193,N_1671,N_1681);
nor U3194 (N_3194,N_1694,N_1645);
nand U3195 (N_3195,N_824,N_827);
nand U3196 (N_3196,N_1878,N_1658);
or U3197 (N_3197,N_1048,N_396);
xor U3198 (N_3198,N_313,N_1105);
nand U3199 (N_3199,N_369,N_1419);
and U3200 (N_3200,N_742,N_1560);
or U3201 (N_3201,N_430,N_1940);
nand U3202 (N_3202,N_498,N_483);
nor U3203 (N_3203,N_665,N_726);
and U3204 (N_3204,N_1894,N_775);
and U3205 (N_3205,N_1324,N_751);
nand U3206 (N_3206,N_676,N_551);
and U3207 (N_3207,N_1760,N_223);
nor U3208 (N_3208,N_619,N_42);
nand U3209 (N_3209,N_1992,N_394);
nor U3210 (N_3210,N_1610,N_402);
nor U3211 (N_3211,N_1019,N_1428);
or U3212 (N_3212,N_628,N_1911);
and U3213 (N_3213,N_853,N_153);
nor U3214 (N_3214,N_1011,N_375);
nor U3215 (N_3215,N_677,N_328);
nand U3216 (N_3216,N_1516,N_1793);
nand U3217 (N_3217,N_1520,N_1430);
nand U3218 (N_3218,N_1665,N_1813);
nand U3219 (N_3219,N_1824,N_141);
and U3220 (N_3220,N_1402,N_299);
nand U3221 (N_3221,N_412,N_1749);
nand U3222 (N_3222,N_1099,N_645);
nor U3223 (N_3223,N_1443,N_1330);
nor U3224 (N_3224,N_1720,N_684);
and U3225 (N_3225,N_1362,N_448);
or U3226 (N_3226,N_1947,N_1274);
nor U3227 (N_3227,N_114,N_1804);
nand U3228 (N_3228,N_1810,N_104);
or U3229 (N_3229,N_1707,N_1958);
nor U3230 (N_3230,N_1888,N_1407);
or U3231 (N_3231,N_230,N_1683);
and U3232 (N_3232,N_1504,N_730);
and U3233 (N_3233,N_1911,N_185);
nor U3234 (N_3234,N_1640,N_1329);
nand U3235 (N_3235,N_780,N_1549);
nand U3236 (N_3236,N_642,N_178);
nand U3237 (N_3237,N_1753,N_481);
and U3238 (N_3238,N_871,N_1351);
nor U3239 (N_3239,N_330,N_776);
nor U3240 (N_3240,N_927,N_713);
or U3241 (N_3241,N_113,N_968);
nand U3242 (N_3242,N_362,N_100);
or U3243 (N_3243,N_1813,N_1249);
or U3244 (N_3244,N_1546,N_1046);
or U3245 (N_3245,N_1493,N_268);
or U3246 (N_3246,N_1081,N_334);
nand U3247 (N_3247,N_1968,N_1508);
nand U3248 (N_3248,N_726,N_1370);
or U3249 (N_3249,N_1089,N_1500);
or U3250 (N_3250,N_1218,N_1313);
nor U3251 (N_3251,N_382,N_1595);
nand U3252 (N_3252,N_1773,N_1293);
or U3253 (N_3253,N_1677,N_1028);
nand U3254 (N_3254,N_1270,N_967);
nand U3255 (N_3255,N_154,N_1893);
or U3256 (N_3256,N_1841,N_1370);
nor U3257 (N_3257,N_627,N_561);
and U3258 (N_3258,N_811,N_855);
and U3259 (N_3259,N_361,N_248);
or U3260 (N_3260,N_136,N_95);
nor U3261 (N_3261,N_1958,N_1174);
nand U3262 (N_3262,N_60,N_1045);
or U3263 (N_3263,N_1440,N_1428);
or U3264 (N_3264,N_938,N_1270);
nand U3265 (N_3265,N_675,N_628);
nor U3266 (N_3266,N_1038,N_1327);
nor U3267 (N_3267,N_95,N_1761);
nand U3268 (N_3268,N_1168,N_1665);
and U3269 (N_3269,N_36,N_1555);
and U3270 (N_3270,N_324,N_1119);
and U3271 (N_3271,N_1613,N_1941);
nor U3272 (N_3272,N_924,N_1701);
or U3273 (N_3273,N_290,N_1281);
or U3274 (N_3274,N_1887,N_1144);
nand U3275 (N_3275,N_817,N_453);
nor U3276 (N_3276,N_1607,N_1814);
or U3277 (N_3277,N_981,N_984);
and U3278 (N_3278,N_384,N_721);
nor U3279 (N_3279,N_1759,N_895);
nor U3280 (N_3280,N_1126,N_574);
nor U3281 (N_3281,N_660,N_1938);
and U3282 (N_3282,N_67,N_461);
nand U3283 (N_3283,N_378,N_1411);
and U3284 (N_3284,N_1777,N_1514);
and U3285 (N_3285,N_1042,N_1493);
nor U3286 (N_3286,N_1458,N_34);
nor U3287 (N_3287,N_533,N_287);
xor U3288 (N_3288,N_1219,N_1919);
and U3289 (N_3289,N_12,N_1981);
nor U3290 (N_3290,N_1051,N_1661);
or U3291 (N_3291,N_424,N_1487);
nand U3292 (N_3292,N_814,N_31);
and U3293 (N_3293,N_1246,N_126);
nand U3294 (N_3294,N_762,N_682);
nor U3295 (N_3295,N_1792,N_1975);
nor U3296 (N_3296,N_1728,N_133);
nor U3297 (N_3297,N_579,N_1335);
nor U3298 (N_3298,N_213,N_1872);
nor U3299 (N_3299,N_1230,N_738);
or U3300 (N_3300,N_1856,N_459);
and U3301 (N_3301,N_43,N_1538);
or U3302 (N_3302,N_917,N_1671);
and U3303 (N_3303,N_619,N_835);
and U3304 (N_3304,N_282,N_1354);
nor U3305 (N_3305,N_944,N_1731);
xnor U3306 (N_3306,N_1471,N_1168);
nor U3307 (N_3307,N_55,N_1840);
or U3308 (N_3308,N_1651,N_1084);
and U3309 (N_3309,N_1448,N_356);
nand U3310 (N_3310,N_596,N_535);
or U3311 (N_3311,N_608,N_755);
nand U3312 (N_3312,N_1233,N_1537);
nor U3313 (N_3313,N_789,N_1061);
and U3314 (N_3314,N_146,N_1066);
nand U3315 (N_3315,N_204,N_629);
nor U3316 (N_3316,N_542,N_308);
and U3317 (N_3317,N_608,N_683);
nor U3318 (N_3318,N_1174,N_1138);
nand U3319 (N_3319,N_1807,N_378);
and U3320 (N_3320,N_1026,N_1774);
nand U3321 (N_3321,N_813,N_98);
or U3322 (N_3322,N_1752,N_754);
nand U3323 (N_3323,N_105,N_747);
nor U3324 (N_3324,N_936,N_1380);
nand U3325 (N_3325,N_110,N_45);
nand U3326 (N_3326,N_323,N_408);
and U3327 (N_3327,N_833,N_1149);
or U3328 (N_3328,N_1146,N_880);
nor U3329 (N_3329,N_1414,N_11);
or U3330 (N_3330,N_1680,N_395);
nand U3331 (N_3331,N_1042,N_707);
nand U3332 (N_3332,N_1963,N_524);
nand U3333 (N_3333,N_769,N_680);
nor U3334 (N_3334,N_1864,N_1877);
xnor U3335 (N_3335,N_1045,N_1070);
nand U3336 (N_3336,N_903,N_659);
or U3337 (N_3337,N_741,N_648);
nand U3338 (N_3338,N_1200,N_1210);
nor U3339 (N_3339,N_723,N_861);
or U3340 (N_3340,N_1868,N_1208);
or U3341 (N_3341,N_742,N_249);
nor U3342 (N_3342,N_292,N_1802);
nor U3343 (N_3343,N_396,N_390);
or U3344 (N_3344,N_83,N_1676);
and U3345 (N_3345,N_442,N_198);
and U3346 (N_3346,N_1919,N_1494);
nand U3347 (N_3347,N_840,N_32);
or U3348 (N_3348,N_1584,N_707);
nand U3349 (N_3349,N_872,N_1435);
or U3350 (N_3350,N_630,N_420);
nor U3351 (N_3351,N_120,N_199);
or U3352 (N_3352,N_563,N_1605);
or U3353 (N_3353,N_902,N_403);
nand U3354 (N_3354,N_89,N_1673);
or U3355 (N_3355,N_566,N_325);
nand U3356 (N_3356,N_1074,N_986);
or U3357 (N_3357,N_885,N_1703);
or U3358 (N_3358,N_1214,N_1665);
nor U3359 (N_3359,N_1130,N_997);
or U3360 (N_3360,N_1415,N_712);
nor U3361 (N_3361,N_895,N_1490);
xnor U3362 (N_3362,N_773,N_1322);
and U3363 (N_3363,N_1771,N_1308);
nand U3364 (N_3364,N_693,N_1267);
nand U3365 (N_3365,N_259,N_1153);
and U3366 (N_3366,N_669,N_793);
or U3367 (N_3367,N_45,N_1334);
nand U3368 (N_3368,N_1244,N_1347);
or U3369 (N_3369,N_400,N_24);
nor U3370 (N_3370,N_1678,N_370);
and U3371 (N_3371,N_404,N_329);
or U3372 (N_3372,N_659,N_1857);
and U3373 (N_3373,N_1575,N_1889);
nor U3374 (N_3374,N_1040,N_1492);
nand U3375 (N_3375,N_1672,N_1724);
xor U3376 (N_3376,N_675,N_1969);
and U3377 (N_3377,N_1086,N_1720);
or U3378 (N_3378,N_1257,N_804);
or U3379 (N_3379,N_1192,N_426);
nand U3380 (N_3380,N_32,N_292);
nand U3381 (N_3381,N_818,N_1527);
nor U3382 (N_3382,N_100,N_908);
and U3383 (N_3383,N_1804,N_1176);
nor U3384 (N_3384,N_1602,N_331);
nor U3385 (N_3385,N_1064,N_1964);
and U3386 (N_3386,N_802,N_946);
nand U3387 (N_3387,N_1969,N_1031);
nor U3388 (N_3388,N_775,N_407);
xor U3389 (N_3389,N_1932,N_131);
nor U3390 (N_3390,N_692,N_46);
xor U3391 (N_3391,N_1359,N_748);
nor U3392 (N_3392,N_981,N_1199);
nor U3393 (N_3393,N_504,N_969);
nand U3394 (N_3394,N_1189,N_1115);
nand U3395 (N_3395,N_811,N_259);
and U3396 (N_3396,N_1595,N_572);
nor U3397 (N_3397,N_595,N_715);
nand U3398 (N_3398,N_1361,N_400);
nand U3399 (N_3399,N_1810,N_646);
and U3400 (N_3400,N_1691,N_55);
nor U3401 (N_3401,N_1775,N_875);
nor U3402 (N_3402,N_1628,N_874);
or U3403 (N_3403,N_1216,N_1898);
or U3404 (N_3404,N_689,N_1436);
nor U3405 (N_3405,N_1671,N_392);
xor U3406 (N_3406,N_1443,N_1251);
and U3407 (N_3407,N_1270,N_1139);
nor U3408 (N_3408,N_1292,N_963);
nor U3409 (N_3409,N_1407,N_670);
and U3410 (N_3410,N_1548,N_1732);
nand U3411 (N_3411,N_262,N_242);
nor U3412 (N_3412,N_347,N_1641);
or U3413 (N_3413,N_109,N_9);
or U3414 (N_3414,N_40,N_610);
and U3415 (N_3415,N_1634,N_1942);
or U3416 (N_3416,N_1155,N_1628);
and U3417 (N_3417,N_897,N_408);
nand U3418 (N_3418,N_1038,N_780);
and U3419 (N_3419,N_747,N_550);
nand U3420 (N_3420,N_121,N_605);
or U3421 (N_3421,N_1509,N_1723);
nor U3422 (N_3422,N_885,N_1775);
nor U3423 (N_3423,N_184,N_1237);
nand U3424 (N_3424,N_1921,N_1320);
or U3425 (N_3425,N_545,N_1658);
or U3426 (N_3426,N_61,N_685);
and U3427 (N_3427,N_807,N_1710);
nand U3428 (N_3428,N_50,N_116);
and U3429 (N_3429,N_536,N_456);
nor U3430 (N_3430,N_1159,N_772);
or U3431 (N_3431,N_272,N_1068);
or U3432 (N_3432,N_1943,N_1247);
nor U3433 (N_3433,N_1810,N_509);
and U3434 (N_3434,N_1627,N_1750);
nand U3435 (N_3435,N_1413,N_1626);
and U3436 (N_3436,N_1796,N_1885);
nand U3437 (N_3437,N_1606,N_1543);
or U3438 (N_3438,N_1796,N_1805);
or U3439 (N_3439,N_117,N_159);
nor U3440 (N_3440,N_1192,N_1146);
and U3441 (N_3441,N_1321,N_1228);
nand U3442 (N_3442,N_1055,N_1952);
and U3443 (N_3443,N_503,N_1246);
and U3444 (N_3444,N_237,N_290);
nand U3445 (N_3445,N_379,N_735);
or U3446 (N_3446,N_86,N_1385);
nor U3447 (N_3447,N_694,N_1337);
and U3448 (N_3448,N_1958,N_288);
nand U3449 (N_3449,N_1190,N_1104);
or U3450 (N_3450,N_348,N_1379);
nor U3451 (N_3451,N_1775,N_13);
or U3452 (N_3452,N_612,N_665);
nand U3453 (N_3453,N_592,N_1611);
nand U3454 (N_3454,N_1323,N_292);
or U3455 (N_3455,N_1735,N_388);
and U3456 (N_3456,N_56,N_328);
and U3457 (N_3457,N_1334,N_548);
and U3458 (N_3458,N_1882,N_835);
and U3459 (N_3459,N_734,N_104);
and U3460 (N_3460,N_311,N_1101);
and U3461 (N_3461,N_644,N_208);
or U3462 (N_3462,N_830,N_1687);
and U3463 (N_3463,N_737,N_661);
nor U3464 (N_3464,N_675,N_609);
or U3465 (N_3465,N_851,N_244);
nand U3466 (N_3466,N_529,N_492);
or U3467 (N_3467,N_756,N_801);
or U3468 (N_3468,N_37,N_1828);
or U3469 (N_3469,N_160,N_1500);
nor U3470 (N_3470,N_994,N_493);
nand U3471 (N_3471,N_656,N_1100);
and U3472 (N_3472,N_1301,N_818);
nor U3473 (N_3473,N_1545,N_1685);
and U3474 (N_3474,N_1687,N_413);
and U3475 (N_3475,N_491,N_426);
nand U3476 (N_3476,N_1694,N_1527);
nor U3477 (N_3477,N_858,N_1027);
nand U3478 (N_3478,N_208,N_125);
nor U3479 (N_3479,N_1953,N_48);
and U3480 (N_3480,N_957,N_22);
nand U3481 (N_3481,N_1898,N_1245);
nand U3482 (N_3482,N_1512,N_1269);
nand U3483 (N_3483,N_401,N_1902);
and U3484 (N_3484,N_1261,N_1984);
or U3485 (N_3485,N_789,N_1062);
nor U3486 (N_3486,N_1156,N_1017);
or U3487 (N_3487,N_966,N_685);
nand U3488 (N_3488,N_1686,N_1265);
or U3489 (N_3489,N_1337,N_893);
or U3490 (N_3490,N_1991,N_1390);
and U3491 (N_3491,N_1799,N_1025);
nor U3492 (N_3492,N_122,N_1035);
nor U3493 (N_3493,N_1962,N_1585);
nor U3494 (N_3494,N_1165,N_1318);
nand U3495 (N_3495,N_1996,N_67);
nor U3496 (N_3496,N_735,N_394);
nand U3497 (N_3497,N_306,N_824);
and U3498 (N_3498,N_1721,N_74);
nor U3499 (N_3499,N_1592,N_439);
or U3500 (N_3500,N_320,N_1363);
nor U3501 (N_3501,N_937,N_362);
or U3502 (N_3502,N_1175,N_715);
and U3503 (N_3503,N_1208,N_1429);
and U3504 (N_3504,N_1098,N_207);
and U3505 (N_3505,N_1542,N_1399);
or U3506 (N_3506,N_215,N_417);
and U3507 (N_3507,N_820,N_743);
or U3508 (N_3508,N_1022,N_1570);
nor U3509 (N_3509,N_1391,N_1510);
nor U3510 (N_3510,N_244,N_802);
nand U3511 (N_3511,N_692,N_58);
nand U3512 (N_3512,N_1220,N_894);
nand U3513 (N_3513,N_774,N_1601);
or U3514 (N_3514,N_205,N_906);
or U3515 (N_3515,N_37,N_297);
and U3516 (N_3516,N_1261,N_634);
and U3517 (N_3517,N_527,N_1700);
nand U3518 (N_3518,N_327,N_905);
nor U3519 (N_3519,N_1574,N_1087);
and U3520 (N_3520,N_1199,N_877);
nand U3521 (N_3521,N_654,N_39);
nor U3522 (N_3522,N_1294,N_1795);
nor U3523 (N_3523,N_990,N_1577);
nor U3524 (N_3524,N_1370,N_212);
or U3525 (N_3525,N_895,N_1735);
or U3526 (N_3526,N_46,N_228);
nand U3527 (N_3527,N_722,N_1365);
or U3528 (N_3528,N_941,N_373);
nor U3529 (N_3529,N_707,N_758);
or U3530 (N_3530,N_492,N_1783);
nand U3531 (N_3531,N_78,N_1032);
and U3532 (N_3532,N_1626,N_1295);
nor U3533 (N_3533,N_190,N_1238);
or U3534 (N_3534,N_641,N_163);
nand U3535 (N_3535,N_104,N_796);
nor U3536 (N_3536,N_1331,N_561);
or U3537 (N_3537,N_1322,N_1421);
nor U3538 (N_3538,N_677,N_212);
and U3539 (N_3539,N_46,N_280);
and U3540 (N_3540,N_383,N_477);
or U3541 (N_3541,N_1108,N_429);
nor U3542 (N_3542,N_101,N_1645);
nor U3543 (N_3543,N_1859,N_1353);
nand U3544 (N_3544,N_562,N_1437);
nand U3545 (N_3545,N_1242,N_509);
or U3546 (N_3546,N_1811,N_374);
and U3547 (N_3547,N_1282,N_934);
nor U3548 (N_3548,N_1675,N_71);
or U3549 (N_3549,N_729,N_1229);
nor U3550 (N_3550,N_20,N_1783);
or U3551 (N_3551,N_808,N_190);
and U3552 (N_3552,N_1541,N_9);
or U3553 (N_3553,N_917,N_1344);
nand U3554 (N_3554,N_662,N_1087);
or U3555 (N_3555,N_753,N_1519);
or U3556 (N_3556,N_593,N_1125);
nor U3557 (N_3557,N_673,N_1241);
nor U3558 (N_3558,N_1728,N_1737);
nor U3559 (N_3559,N_1976,N_1091);
or U3560 (N_3560,N_674,N_121);
nand U3561 (N_3561,N_1022,N_634);
nand U3562 (N_3562,N_1729,N_981);
nand U3563 (N_3563,N_1505,N_1675);
and U3564 (N_3564,N_582,N_1122);
nand U3565 (N_3565,N_280,N_1012);
nand U3566 (N_3566,N_402,N_888);
and U3567 (N_3567,N_1143,N_1338);
nor U3568 (N_3568,N_999,N_1336);
nor U3569 (N_3569,N_168,N_597);
or U3570 (N_3570,N_1979,N_1674);
or U3571 (N_3571,N_82,N_1114);
nor U3572 (N_3572,N_356,N_277);
nand U3573 (N_3573,N_303,N_1042);
nand U3574 (N_3574,N_1261,N_1686);
nand U3575 (N_3575,N_1777,N_1508);
nand U3576 (N_3576,N_695,N_766);
nor U3577 (N_3577,N_1452,N_426);
nand U3578 (N_3578,N_1611,N_1027);
nand U3579 (N_3579,N_1781,N_62);
nor U3580 (N_3580,N_544,N_507);
and U3581 (N_3581,N_418,N_1795);
and U3582 (N_3582,N_1779,N_1543);
and U3583 (N_3583,N_385,N_752);
or U3584 (N_3584,N_851,N_1230);
and U3585 (N_3585,N_103,N_139);
or U3586 (N_3586,N_490,N_1180);
xor U3587 (N_3587,N_1168,N_632);
and U3588 (N_3588,N_1658,N_406);
and U3589 (N_3589,N_520,N_89);
nand U3590 (N_3590,N_610,N_1393);
nand U3591 (N_3591,N_1958,N_309);
or U3592 (N_3592,N_1009,N_1234);
nand U3593 (N_3593,N_1414,N_880);
or U3594 (N_3594,N_500,N_1759);
or U3595 (N_3595,N_126,N_1200);
or U3596 (N_3596,N_391,N_61);
nor U3597 (N_3597,N_777,N_6);
or U3598 (N_3598,N_1124,N_373);
and U3599 (N_3599,N_45,N_101);
nand U3600 (N_3600,N_1324,N_1769);
nand U3601 (N_3601,N_517,N_1186);
nor U3602 (N_3602,N_1104,N_1506);
or U3603 (N_3603,N_742,N_1970);
nor U3604 (N_3604,N_1973,N_162);
nor U3605 (N_3605,N_1938,N_321);
and U3606 (N_3606,N_1969,N_1782);
nand U3607 (N_3607,N_424,N_98);
nor U3608 (N_3608,N_1665,N_1438);
nand U3609 (N_3609,N_1307,N_1686);
nand U3610 (N_3610,N_1106,N_1623);
nor U3611 (N_3611,N_1586,N_479);
and U3612 (N_3612,N_1610,N_422);
and U3613 (N_3613,N_525,N_688);
or U3614 (N_3614,N_1169,N_1694);
nor U3615 (N_3615,N_729,N_573);
nor U3616 (N_3616,N_241,N_1469);
and U3617 (N_3617,N_1968,N_378);
nand U3618 (N_3618,N_950,N_157);
or U3619 (N_3619,N_880,N_489);
nor U3620 (N_3620,N_118,N_540);
or U3621 (N_3621,N_1772,N_1184);
nand U3622 (N_3622,N_147,N_167);
and U3623 (N_3623,N_1968,N_878);
or U3624 (N_3624,N_1461,N_1334);
or U3625 (N_3625,N_613,N_430);
nand U3626 (N_3626,N_327,N_959);
or U3627 (N_3627,N_845,N_827);
nor U3628 (N_3628,N_779,N_406);
nor U3629 (N_3629,N_1221,N_7);
or U3630 (N_3630,N_1813,N_1806);
nor U3631 (N_3631,N_457,N_1725);
nor U3632 (N_3632,N_1443,N_1884);
or U3633 (N_3633,N_793,N_1802);
and U3634 (N_3634,N_280,N_615);
nand U3635 (N_3635,N_1657,N_773);
or U3636 (N_3636,N_1054,N_1358);
nand U3637 (N_3637,N_1556,N_1763);
nand U3638 (N_3638,N_1673,N_1415);
or U3639 (N_3639,N_1402,N_1721);
and U3640 (N_3640,N_240,N_1926);
nand U3641 (N_3641,N_1265,N_1455);
nand U3642 (N_3642,N_47,N_1595);
and U3643 (N_3643,N_1027,N_533);
nand U3644 (N_3644,N_1365,N_129);
and U3645 (N_3645,N_500,N_41);
xor U3646 (N_3646,N_1526,N_1213);
or U3647 (N_3647,N_1644,N_350);
nand U3648 (N_3648,N_366,N_1835);
and U3649 (N_3649,N_1039,N_79);
nand U3650 (N_3650,N_942,N_932);
nand U3651 (N_3651,N_954,N_1237);
nor U3652 (N_3652,N_1457,N_1605);
or U3653 (N_3653,N_965,N_1111);
nand U3654 (N_3654,N_1773,N_1644);
nand U3655 (N_3655,N_939,N_1478);
and U3656 (N_3656,N_1012,N_1988);
or U3657 (N_3657,N_956,N_1966);
or U3658 (N_3658,N_378,N_1393);
nor U3659 (N_3659,N_1326,N_256);
and U3660 (N_3660,N_1093,N_1012);
or U3661 (N_3661,N_1603,N_1058);
nand U3662 (N_3662,N_233,N_378);
and U3663 (N_3663,N_1073,N_1912);
nand U3664 (N_3664,N_6,N_1903);
nand U3665 (N_3665,N_415,N_1637);
nor U3666 (N_3666,N_962,N_1553);
and U3667 (N_3667,N_384,N_1051);
nand U3668 (N_3668,N_264,N_819);
nand U3669 (N_3669,N_1167,N_269);
nand U3670 (N_3670,N_855,N_1413);
nand U3671 (N_3671,N_473,N_879);
nand U3672 (N_3672,N_237,N_1366);
and U3673 (N_3673,N_1435,N_333);
or U3674 (N_3674,N_91,N_227);
and U3675 (N_3675,N_445,N_1852);
and U3676 (N_3676,N_564,N_968);
nor U3677 (N_3677,N_1054,N_1284);
nand U3678 (N_3678,N_1828,N_1516);
and U3679 (N_3679,N_252,N_1590);
nor U3680 (N_3680,N_686,N_1949);
nand U3681 (N_3681,N_1784,N_1702);
or U3682 (N_3682,N_1987,N_578);
nor U3683 (N_3683,N_119,N_141);
and U3684 (N_3684,N_908,N_1624);
and U3685 (N_3685,N_487,N_748);
and U3686 (N_3686,N_1697,N_940);
or U3687 (N_3687,N_701,N_1062);
nor U3688 (N_3688,N_1228,N_1449);
and U3689 (N_3689,N_34,N_1296);
and U3690 (N_3690,N_1790,N_1231);
nand U3691 (N_3691,N_1981,N_615);
xor U3692 (N_3692,N_447,N_1088);
or U3693 (N_3693,N_477,N_1043);
xnor U3694 (N_3694,N_965,N_1347);
nor U3695 (N_3695,N_1512,N_185);
nand U3696 (N_3696,N_920,N_1398);
or U3697 (N_3697,N_326,N_587);
nand U3698 (N_3698,N_198,N_10);
nand U3699 (N_3699,N_536,N_482);
nand U3700 (N_3700,N_816,N_1651);
nand U3701 (N_3701,N_1837,N_1552);
or U3702 (N_3702,N_1285,N_342);
and U3703 (N_3703,N_40,N_906);
and U3704 (N_3704,N_54,N_495);
nand U3705 (N_3705,N_452,N_819);
and U3706 (N_3706,N_1679,N_514);
and U3707 (N_3707,N_1340,N_649);
or U3708 (N_3708,N_135,N_1733);
and U3709 (N_3709,N_1286,N_659);
nor U3710 (N_3710,N_888,N_740);
nand U3711 (N_3711,N_499,N_1879);
nor U3712 (N_3712,N_1746,N_1476);
or U3713 (N_3713,N_1217,N_999);
and U3714 (N_3714,N_1260,N_1544);
and U3715 (N_3715,N_1284,N_1681);
nand U3716 (N_3716,N_1167,N_860);
nand U3717 (N_3717,N_724,N_1590);
nor U3718 (N_3718,N_1844,N_744);
nor U3719 (N_3719,N_1851,N_170);
and U3720 (N_3720,N_1316,N_361);
or U3721 (N_3721,N_1799,N_1540);
and U3722 (N_3722,N_1809,N_384);
nor U3723 (N_3723,N_913,N_1430);
nand U3724 (N_3724,N_1669,N_1089);
nor U3725 (N_3725,N_921,N_278);
or U3726 (N_3726,N_1684,N_572);
or U3727 (N_3727,N_921,N_1393);
nor U3728 (N_3728,N_1423,N_213);
nor U3729 (N_3729,N_472,N_1258);
nor U3730 (N_3730,N_709,N_1212);
and U3731 (N_3731,N_1816,N_514);
or U3732 (N_3732,N_1259,N_1139);
nor U3733 (N_3733,N_1955,N_1140);
or U3734 (N_3734,N_1280,N_562);
or U3735 (N_3735,N_1227,N_700);
or U3736 (N_3736,N_988,N_98);
and U3737 (N_3737,N_750,N_843);
nand U3738 (N_3738,N_17,N_21);
xnor U3739 (N_3739,N_733,N_502);
or U3740 (N_3740,N_793,N_185);
nor U3741 (N_3741,N_66,N_173);
nor U3742 (N_3742,N_1775,N_262);
and U3743 (N_3743,N_1012,N_1480);
and U3744 (N_3744,N_824,N_1343);
nand U3745 (N_3745,N_1931,N_1168);
and U3746 (N_3746,N_330,N_1492);
or U3747 (N_3747,N_454,N_1836);
nor U3748 (N_3748,N_955,N_1774);
nand U3749 (N_3749,N_4,N_202);
and U3750 (N_3750,N_585,N_1538);
or U3751 (N_3751,N_1989,N_417);
or U3752 (N_3752,N_123,N_286);
and U3753 (N_3753,N_1523,N_1892);
and U3754 (N_3754,N_1541,N_1621);
nand U3755 (N_3755,N_1009,N_1541);
nor U3756 (N_3756,N_399,N_1898);
nand U3757 (N_3757,N_32,N_71);
nor U3758 (N_3758,N_1528,N_1975);
nor U3759 (N_3759,N_1783,N_624);
nand U3760 (N_3760,N_625,N_446);
nor U3761 (N_3761,N_275,N_42);
nand U3762 (N_3762,N_776,N_40);
and U3763 (N_3763,N_1424,N_741);
nor U3764 (N_3764,N_1781,N_187);
or U3765 (N_3765,N_1237,N_814);
nand U3766 (N_3766,N_151,N_1741);
nand U3767 (N_3767,N_1261,N_495);
nand U3768 (N_3768,N_1444,N_343);
or U3769 (N_3769,N_515,N_970);
nand U3770 (N_3770,N_1659,N_740);
and U3771 (N_3771,N_1244,N_1605);
and U3772 (N_3772,N_852,N_447);
nor U3773 (N_3773,N_1157,N_474);
nand U3774 (N_3774,N_1068,N_242);
or U3775 (N_3775,N_1216,N_1161);
and U3776 (N_3776,N_321,N_1067);
and U3777 (N_3777,N_372,N_993);
and U3778 (N_3778,N_1180,N_1472);
nor U3779 (N_3779,N_1511,N_231);
nor U3780 (N_3780,N_1943,N_1889);
nand U3781 (N_3781,N_1717,N_693);
nor U3782 (N_3782,N_640,N_1607);
and U3783 (N_3783,N_1820,N_412);
and U3784 (N_3784,N_881,N_786);
or U3785 (N_3785,N_1418,N_935);
nand U3786 (N_3786,N_1759,N_139);
or U3787 (N_3787,N_913,N_1077);
nand U3788 (N_3788,N_152,N_642);
nor U3789 (N_3789,N_546,N_416);
nand U3790 (N_3790,N_1197,N_293);
nor U3791 (N_3791,N_1476,N_176);
and U3792 (N_3792,N_142,N_193);
and U3793 (N_3793,N_1766,N_316);
and U3794 (N_3794,N_1703,N_179);
nand U3795 (N_3795,N_1849,N_1293);
or U3796 (N_3796,N_847,N_382);
and U3797 (N_3797,N_35,N_1644);
nand U3798 (N_3798,N_1979,N_1466);
nand U3799 (N_3799,N_120,N_554);
and U3800 (N_3800,N_1390,N_1245);
nor U3801 (N_3801,N_1070,N_451);
nor U3802 (N_3802,N_1698,N_319);
nor U3803 (N_3803,N_901,N_397);
and U3804 (N_3804,N_821,N_1570);
nand U3805 (N_3805,N_289,N_1813);
and U3806 (N_3806,N_1964,N_860);
or U3807 (N_3807,N_469,N_1708);
nand U3808 (N_3808,N_732,N_24);
nand U3809 (N_3809,N_1989,N_736);
and U3810 (N_3810,N_1907,N_157);
or U3811 (N_3811,N_1503,N_2);
nand U3812 (N_3812,N_730,N_943);
nand U3813 (N_3813,N_1898,N_1824);
or U3814 (N_3814,N_1831,N_1473);
nand U3815 (N_3815,N_1797,N_1882);
and U3816 (N_3816,N_1438,N_1320);
and U3817 (N_3817,N_1608,N_137);
or U3818 (N_3818,N_582,N_1419);
and U3819 (N_3819,N_1586,N_397);
nor U3820 (N_3820,N_352,N_244);
nor U3821 (N_3821,N_1995,N_1192);
nand U3822 (N_3822,N_1079,N_833);
nand U3823 (N_3823,N_1884,N_1618);
or U3824 (N_3824,N_1671,N_1369);
and U3825 (N_3825,N_249,N_549);
nand U3826 (N_3826,N_1435,N_1912);
and U3827 (N_3827,N_1795,N_1767);
nor U3828 (N_3828,N_944,N_1648);
and U3829 (N_3829,N_618,N_1881);
nor U3830 (N_3830,N_1451,N_1147);
xor U3831 (N_3831,N_531,N_76);
or U3832 (N_3832,N_1009,N_416);
nand U3833 (N_3833,N_811,N_685);
nand U3834 (N_3834,N_752,N_1688);
nor U3835 (N_3835,N_1526,N_638);
nor U3836 (N_3836,N_1839,N_580);
or U3837 (N_3837,N_643,N_873);
xnor U3838 (N_3838,N_826,N_1301);
and U3839 (N_3839,N_1451,N_287);
and U3840 (N_3840,N_1153,N_1626);
nor U3841 (N_3841,N_130,N_1943);
nor U3842 (N_3842,N_1060,N_1004);
or U3843 (N_3843,N_1438,N_128);
nand U3844 (N_3844,N_1767,N_895);
nand U3845 (N_3845,N_722,N_1559);
or U3846 (N_3846,N_863,N_1639);
or U3847 (N_3847,N_1258,N_1042);
and U3848 (N_3848,N_1767,N_1072);
nor U3849 (N_3849,N_784,N_1985);
and U3850 (N_3850,N_81,N_194);
nor U3851 (N_3851,N_1776,N_840);
and U3852 (N_3852,N_1057,N_1304);
or U3853 (N_3853,N_1541,N_858);
or U3854 (N_3854,N_1865,N_1380);
and U3855 (N_3855,N_1597,N_1425);
nand U3856 (N_3856,N_120,N_691);
nor U3857 (N_3857,N_453,N_292);
nor U3858 (N_3858,N_1491,N_1608);
nor U3859 (N_3859,N_1570,N_328);
or U3860 (N_3860,N_1407,N_65);
or U3861 (N_3861,N_515,N_29);
and U3862 (N_3862,N_1873,N_140);
nand U3863 (N_3863,N_1802,N_266);
or U3864 (N_3864,N_428,N_1074);
nand U3865 (N_3865,N_1833,N_352);
or U3866 (N_3866,N_247,N_504);
or U3867 (N_3867,N_1388,N_188);
nand U3868 (N_3868,N_1678,N_1601);
nor U3869 (N_3869,N_1918,N_341);
nand U3870 (N_3870,N_1014,N_1604);
nand U3871 (N_3871,N_1846,N_1859);
or U3872 (N_3872,N_1334,N_1708);
or U3873 (N_3873,N_35,N_985);
nand U3874 (N_3874,N_1326,N_757);
or U3875 (N_3875,N_964,N_100);
nand U3876 (N_3876,N_1574,N_728);
or U3877 (N_3877,N_1560,N_153);
nor U3878 (N_3878,N_1864,N_1437);
nor U3879 (N_3879,N_1667,N_944);
and U3880 (N_3880,N_718,N_1544);
or U3881 (N_3881,N_1758,N_356);
nor U3882 (N_3882,N_494,N_1435);
nor U3883 (N_3883,N_310,N_1350);
or U3884 (N_3884,N_356,N_445);
nor U3885 (N_3885,N_515,N_1133);
or U3886 (N_3886,N_1273,N_1759);
nor U3887 (N_3887,N_1053,N_974);
xnor U3888 (N_3888,N_1388,N_1478);
nor U3889 (N_3889,N_338,N_1926);
or U3890 (N_3890,N_1302,N_1367);
nor U3891 (N_3891,N_334,N_813);
and U3892 (N_3892,N_176,N_913);
and U3893 (N_3893,N_315,N_1344);
nand U3894 (N_3894,N_809,N_907);
and U3895 (N_3895,N_1709,N_943);
nand U3896 (N_3896,N_1660,N_1443);
and U3897 (N_3897,N_1880,N_1319);
nand U3898 (N_3898,N_532,N_1017);
nor U3899 (N_3899,N_923,N_1797);
or U3900 (N_3900,N_1803,N_278);
and U3901 (N_3901,N_1943,N_218);
and U3902 (N_3902,N_1576,N_163);
or U3903 (N_3903,N_865,N_1397);
nor U3904 (N_3904,N_748,N_1426);
or U3905 (N_3905,N_651,N_863);
nor U3906 (N_3906,N_1206,N_1978);
nand U3907 (N_3907,N_1566,N_1682);
nand U3908 (N_3908,N_1955,N_782);
nand U3909 (N_3909,N_190,N_419);
and U3910 (N_3910,N_1884,N_175);
xnor U3911 (N_3911,N_1529,N_1953);
nand U3912 (N_3912,N_1753,N_494);
or U3913 (N_3913,N_199,N_1785);
or U3914 (N_3914,N_638,N_402);
nand U3915 (N_3915,N_1298,N_1884);
and U3916 (N_3916,N_945,N_1193);
nand U3917 (N_3917,N_1145,N_463);
or U3918 (N_3918,N_1482,N_1225);
nand U3919 (N_3919,N_877,N_510);
or U3920 (N_3920,N_644,N_1830);
nor U3921 (N_3921,N_687,N_895);
nor U3922 (N_3922,N_155,N_652);
nand U3923 (N_3923,N_1616,N_850);
nor U3924 (N_3924,N_1088,N_1564);
nand U3925 (N_3925,N_41,N_101);
nand U3926 (N_3926,N_85,N_375);
or U3927 (N_3927,N_718,N_1239);
and U3928 (N_3928,N_1954,N_621);
nor U3929 (N_3929,N_431,N_1696);
nand U3930 (N_3930,N_1876,N_1763);
or U3931 (N_3931,N_525,N_1279);
and U3932 (N_3932,N_139,N_1320);
nor U3933 (N_3933,N_1149,N_1800);
nand U3934 (N_3934,N_537,N_1779);
nand U3935 (N_3935,N_65,N_1241);
and U3936 (N_3936,N_1833,N_641);
nand U3937 (N_3937,N_1765,N_1178);
nor U3938 (N_3938,N_606,N_1520);
or U3939 (N_3939,N_566,N_68);
nand U3940 (N_3940,N_787,N_1558);
or U3941 (N_3941,N_190,N_1354);
nand U3942 (N_3942,N_1261,N_1207);
and U3943 (N_3943,N_371,N_1348);
nand U3944 (N_3944,N_1364,N_420);
and U3945 (N_3945,N_441,N_290);
or U3946 (N_3946,N_388,N_1180);
and U3947 (N_3947,N_1388,N_835);
nor U3948 (N_3948,N_374,N_1571);
nand U3949 (N_3949,N_1421,N_1212);
or U3950 (N_3950,N_719,N_253);
or U3951 (N_3951,N_1920,N_68);
nor U3952 (N_3952,N_1710,N_1498);
or U3953 (N_3953,N_903,N_800);
or U3954 (N_3954,N_95,N_504);
nand U3955 (N_3955,N_1237,N_1573);
nor U3956 (N_3956,N_57,N_135);
and U3957 (N_3957,N_350,N_1762);
nor U3958 (N_3958,N_1269,N_1167);
nor U3959 (N_3959,N_814,N_688);
nor U3960 (N_3960,N_1185,N_732);
nor U3961 (N_3961,N_1544,N_433);
nand U3962 (N_3962,N_1668,N_538);
and U3963 (N_3963,N_132,N_907);
or U3964 (N_3964,N_1530,N_1274);
xnor U3965 (N_3965,N_1403,N_1834);
xnor U3966 (N_3966,N_649,N_1090);
nand U3967 (N_3967,N_636,N_1579);
nand U3968 (N_3968,N_1551,N_1133);
and U3969 (N_3969,N_588,N_1741);
or U3970 (N_3970,N_62,N_1615);
or U3971 (N_3971,N_1490,N_885);
and U3972 (N_3972,N_1630,N_1927);
and U3973 (N_3973,N_1522,N_1291);
nor U3974 (N_3974,N_756,N_1298);
or U3975 (N_3975,N_945,N_829);
nor U3976 (N_3976,N_995,N_904);
nor U3977 (N_3977,N_109,N_1295);
nor U3978 (N_3978,N_1533,N_800);
xor U3979 (N_3979,N_747,N_1930);
and U3980 (N_3980,N_14,N_271);
nor U3981 (N_3981,N_51,N_1788);
and U3982 (N_3982,N_332,N_261);
or U3983 (N_3983,N_1774,N_1425);
and U3984 (N_3984,N_454,N_1120);
and U3985 (N_3985,N_559,N_1503);
or U3986 (N_3986,N_1203,N_1463);
nand U3987 (N_3987,N_344,N_899);
and U3988 (N_3988,N_11,N_1722);
or U3989 (N_3989,N_941,N_680);
or U3990 (N_3990,N_1526,N_253);
nor U3991 (N_3991,N_1758,N_1165);
nor U3992 (N_3992,N_180,N_868);
nor U3993 (N_3993,N_195,N_1611);
and U3994 (N_3994,N_289,N_1489);
nor U3995 (N_3995,N_158,N_414);
nor U3996 (N_3996,N_606,N_1359);
nand U3997 (N_3997,N_710,N_185);
and U3998 (N_3998,N_1225,N_1815);
nor U3999 (N_3999,N_742,N_751);
nand U4000 (N_4000,N_2211,N_3188);
and U4001 (N_4001,N_3234,N_2087);
and U4002 (N_4002,N_2550,N_2778);
or U4003 (N_4003,N_3448,N_3468);
and U4004 (N_4004,N_3558,N_3183);
and U4005 (N_4005,N_2802,N_2517);
or U4006 (N_4006,N_3884,N_3075);
nand U4007 (N_4007,N_3756,N_3310);
and U4008 (N_4008,N_3910,N_3587);
or U4009 (N_4009,N_2122,N_3164);
nand U4010 (N_4010,N_3335,N_3019);
nor U4011 (N_4011,N_2410,N_2880);
or U4012 (N_4012,N_2805,N_3155);
or U4013 (N_4013,N_3676,N_3305);
and U4014 (N_4014,N_3187,N_2417);
or U4015 (N_4015,N_3857,N_3431);
nor U4016 (N_4016,N_3201,N_2876);
or U4017 (N_4017,N_2169,N_2006);
and U4018 (N_4018,N_2634,N_2729);
and U4019 (N_4019,N_3500,N_3023);
and U4020 (N_4020,N_2633,N_3648);
or U4021 (N_4021,N_2845,N_2906);
nor U4022 (N_4022,N_3511,N_3510);
or U4023 (N_4023,N_2535,N_2280);
nor U4024 (N_4024,N_3858,N_2598);
nor U4025 (N_4025,N_3024,N_3400);
or U4026 (N_4026,N_2508,N_2033);
nand U4027 (N_4027,N_3039,N_2583);
nor U4028 (N_4028,N_2571,N_2999);
nand U4029 (N_4029,N_2506,N_2698);
and U4030 (N_4030,N_2034,N_2407);
nand U4031 (N_4031,N_3514,N_2430);
nor U4032 (N_4032,N_2115,N_2705);
nand U4033 (N_4033,N_3955,N_3983);
or U4034 (N_4034,N_3411,N_2723);
nor U4035 (N_4035,N_2300,N_3258);
nand U4036 (N_4036,N_2370,N_2128);
nor U4037 (N_4037,N_2458,N_3956);
nand U4038 (N_4038,N_2798,N_2526);
or U4039 (N_4039,N_3906,N_2946);
nand U4040 (N_4040,N_3592,N_3841);
nor U4041 (N_4041,N_2055,N_2467);
or U4042 (N_4042,N_2872,N_3087);
or U4043 (N_4043,N_3395,N_2806);
and U4044 (N_4044,N_2655,N_3576);
nand U4045 (N_4045,N_2786,N_2229);
nor U4046 (N_4046,N_3808,N_2735);
nand U4047 (N_4047,N_2542,N_2247);
and U4048 (N_4048,N_2897,N_2649);
or U4049 (N_4049,N_3766,N_2235);
nor U4050 (N_4050,N_2696,N_3390);
and U4051 (N_4051,N_2185,N_2887);
and U4052 (N_4052,N_2674,N_2401);
or U4053 (N_4053,N_2125,N_2869);
or U4054 (N_4054,N_3050,N_2249);
or U4055 (N_4055,N_2551,N_3089);
or U4056 (N_4056,N_3486,N_2252);
nor U4057 (N_4057,N_2708,N_2240);
or U4058 (N_4058,N_3373,N_3191);
and U4059 (N_4059,N_2656,N_2920);
nor U4060 (N_4060,N_2192,N_2236);
nor U4061 (N_4061,N_3540,N_2835);
nor U4062 (N_4062,N_3489,N_2913);
nor U4063 (N_4063,N_2476,N_3623);
or U4064 (N_4064,N_2673,N_3124);
or U4065 (N_4065,N_3774,N_3717);
nor U4066 (N_4066,N_2619,N_2677);
or U4067 (N_4067,N_3664,N_2340);
nor U4068 (N_4068,N_3119,N_3454);
nand U4069 (N_4069,N_3503,N_3784);
nor U4070 (N_4070,N_2027,N_3112);
nand U4071 (N_4071,N_3353,N_2525);
xnor U4072 (N_4072,N_3182,N_3755);
nor U4073 (N_4073,N_2973,N_2302);
and U4074 (N_4074,N_2414,N_3782);
nand U4075 (N_4075,N_2616,N_3973);
and U4076 (N_4076,N_3938,N_3833);
and U4077 (N_4077,N_2760,N_3150);
nor U4078 (N_4078,N_2321,N_2864);
and U4079 (N_4079,N_2475,N_3851);
nor U4080 (N_4080,N_3306,N_2565);
and U4081 (N_4081,N_2182,N_2409);
and U4082 (N_4082,N_3442,N_2593);
nand U4083 (N_4083,N_2568,N_2815);
or U4084 (N_4084,N_2781,N_2189);
nor U4085 (N_4085,N_2577,N_3765);
and U4086 (N_4086,N_3773,N_2818);
and U4087 (N_4087,N_2768,N_2661);
and U4088 (N_4088,N_3746,N_2053);
and U4089 (N_4089,N_3527,N_2951);
nor U4090 (N_4090,N_3297,N_2178);
nand U4091 (N_4091,N_3946,N_2595);
nand U4092 (N_4092,N_2803,N_2270);
nand U4093 (N_4093,N_3881,N_2045);
xnor U4094 (N_4094,N_3056,N_3965);
or U4095 (N_4095,N_3475,N_2246);
nor U4096 (N_4096,N_2640,N_3689);
or U4097 (N_4097,N_2731,N_3239);
or U4098 (N_4098,N_2186,N_2369);
nand U4099 (N_4099,N_2047,N_3953);
and U4100 (N_4100,N_2755,N_2224);
or U4101 (N_4101,N_2162,N_2328);
and U4102 (N_4102,N_3810,N_2342);
or U4103 (N_4103,N_3579,N_3654);
and U4104 (N_4104,N_3314,N_3271);
and U4105 (N_4105,N_2352,N_3122);
nand U4106 (N_4106,N_3602,N_2611);
or U4107 (N_4107,N_3238,N_2645);
or U4108 (N_4108,N_3409,N_3550);
nand U4109 (N_4109,N_3275,N_2706);
nand U4110 (N_4110,N_3030,N_3852);
nor U4111 (N_4111,N_3086,N_2081);
and U4112 (N_4112,N_2636,N_2040);
nor U4113 (N_4113,N_3362,N_2438);
nand U4114 (N_4114,N_3894,N_3135);
nand U4115 (N_4115,N_3978,N_3343);
or U4116 (N_4116,N_3360,N_2159);
and U4117 (N_4117,N_2434,N_2011);
or U4118 (N_4118,N_3117,N_2016);
and U4119 (N_4119,N_2491,N_2914);
and U4120 (N_4120,N_3914,N_2727);
or U4121 (N_4121,N_2949,N_3688);
and U4122 (N_4122,N_2048,N_3830);
nand U4123 (N_4123,N_2987,N_3590);
nand U4124 (N_4124,N_2623,N_3645);
nor U4125 (N_4125,N_2184,N_3499);
and U4126 (N_4126,N_2563,N_2724);
and U4127 (N_4127,N_3235,N_2347);
and U4128 (N_4128,N_3349,N_2371);
and U4129 (N_4129,N_3507,N_3116);
nand U4130 (N_4130,N_2683,N_2303);
and U4131 (N_4131,N_3708,N_3470);
or U4132 (N_4132,N_2286,N_2676);
or U4133 (N_4133,N_3989,N_3364);
and U4134 (N_4134,N_3725,N_2250);
nand U4135 (N_4135,N_3371,N_3331);
or U4136 (N_4136,N_2085,N_2956);
nor U4137 (N_4137,N_2305,N_2251);
nor U4138 (N_4138,N_2174,N_2360);
or U4139 (N_4139,N_2689,N_2770);
and U4140 (N_4140,N_3350,N_2493);
nor U4141 (N_4141,N_2843,N_2455);
and U4142 (N_4142,N_3516,N_3332);
nand U4143 (N_4143,N_2293,N_3711);
nor U4144 (N_4144,N_3873,N_2232);
nand U4145 (N_4145,N_2998,N_2747);
nor U4146 (N_4146,N_2970,N_2552);
nand U4147 (N_4147,N_2459,N_2715);
or U4148 (N_4148,N_2380,N_3449);
nand U4149 (N_4149,N_3814,N_3134);
nand U4150 (N_4150,N_3302,N_2097);
nor U4151 (N_4151,N_2559,N_2181);
or U4152 (N_4152,N_2935,N_2516);
or U4153 (N_4153,N_2877,N_3151);
nor U4154 (N_4154,N_3723,N_3458);
and U4155 (N_4155,N_3369,N_2167);
or U4156 (N_4156,N_3829,N_2701);
nor U4157 (N_4157,N_2642,N_3560);
or U4158 (N_4158,N_2112,N_2313);
nor U4159 (N_4159,N_2127,N_2852);
and U4160 (N_4160,N_3600,N_2145);
or U4161 (N_4161,N_3170,N_3451);
nor U4162 (N_4162,N_2242,N_2323);
or U4163 (N_4163,N_3713,N_2402);
and U4164 (N_4164,N_2855,N_2398);
nor U4165 (N_4165,N_3764,N_2136);
nand U4166 (N_4166,N_2483,N_3801);
or U4167 (N_4167,N_3236,N_2894);
nor U4168 (N_4168,N_3897,N_3107);
nor U4169 (N_4169,N_3408,N_3812);
or U4170 (N_4170,N_2839,N_2991);
and U4171 (N_4171,N_2967,N_3130);
nand U4172 (N_4172,N_2426,N_3303);
nor U4173 (N_4173,N_2324,N_3129);
or U4174 (N_4174,N_3673,N_2317);
or U4175 (N_4175,N_2785,N_3568);
and U4176 (N_4176,N_3518,N_2141);
nand U4177 (N_4177,N_3605,N_2707);
and U4178 (N_4178,N_3308,N_2886);
and U4179 (N_4179,N_2140,N_2111);
nor U4180 (N_4180,N_2346,N_2166);
and U4181 (N_4181,N_2981,N_3625);
or U4182 (N_4182,N_2432,N_2231);
nor U4183 (N_4183,N_2183,N_2173);
nor U4184 (N_4184,N_2160,N_3021);
or U4185 (N_4185,N_2714,N_2210);
xor U4186 (N_4186,N_3406,N_2326);
or U4187 (N_4187,N_3904,N_3142);
nand U4188 (N_4188,N_3044,N_3304);
nor U4189 (N_4189,N_2253,N_2233);
and U4190 (N_4190,N_3935,N_3316);
and U4191 (N_4191,N_2950,N_3613);
and U4192 (N_4192,N_3779,N_2553);
and U4193 (N_4193,N_3334,N_2857);
or U4194 (N_4194,N_3929,N_3900);
nand U4195 (N_4195,N_3656,N_3192);
or U4196 (N_4196,N_2329,N_2039);
nand U4197 (N_4197,N_3995,N_3103);
or U4198 (N_4198,N_3637,N_2536);
nand U4199 (N_4199,N_3534,N_2732);
nand U4200 (N_4200,N_2936,N_2681);
and U4201 (N_4201,N_3687,N_3068);
nor U4202 (N_4202,N_2754,N_3326);
nor U4203 (N_4203,N_2237,N_2827);
or U4204 (N_4204,N_2966,N_2154);
or U4205 (N_4205,N_3700,N_3655);
and U4206 (N_4206,N_3616,N_3724);
nand U4207 (N_4207,N_2416,N_2197);
nand U4208 (N_4208,N_2068,N_2738);
nand U4209 (N_4209,N_2041,N_3356);
nor U4210 (N_4210,N_3374,N_2100);
nor U4211 (N_4211,N_2761,N_3805);
or U4212 (N_4212,N_2244,N_3079);
or U4213 (N_4213,N_2297,N_2461);
and U4214 (N_4214,N_2927,N_3083);
nor U4215 (N_4215,N_2773,N_3261);
nor U4216 (N_4216,N_2691,N_3295);
and U4217 (N_4217,N_2982,N_2264);
nor U4218 (N_4218,N_2031,N_2528);
nand U4219 (N_4219,N_3966,N_2227);
nand U4220 (N_4220,N_2507,N_2963);
nor U4221 (N_4221,N_3478,N_2974);
or U4222 (N_4222,N_3545,N_2971);
nor U4223 (N_4223,N_3099,N_2163);
nand U4224 (N_4224,N_3490,N_2378);
nor U4225 (N_4225,N_2433,N_3570);
nand U4226 (N_4226,N_2670,N_2899);
and U4227 (N_4227,N_3078,N_3791);
nor U4228 (N_4228,N_2118,N_2938);
nor U4229 (N_4229,N_2556,N_3770);
or U4230 (N_4230,N_2071,N_2168);
and U4231 (N_4231,N_3060,N_2879);
or U4232 (N_4232,N_2107,N_2243);
or U4233 (N_4233,N_2064,N_3957);
and U4234 (N_4234,N_2700,N_3416);
or U4235 (N_4235,N_3787,N_3809);
or U4236 (N_4236,N_2969,N_3743);
nor U4237 (N_4237,N_2005,N_3113);
nor U4238 (N_4238,N_2110,N_3544);
nor U4239 (N_4239,N_2846,N_2978);
nand U4240 (N_4240,N_2934,N_2822);
or U4241 (N_4241,N_3960,N_3203);
nand U4242 (N_4242,N_2073,N_3925);
and U4243 (N_4243,N_2756,N_3108);
and U4244 (N_4244,N_2423,N_2278);
nor U4245 (N_4245,N_2309,N_2488);
or U4246 (N_4246,N_2549,N_3822);
or U4247 (N_4247,N_3509,N_3895);
nand U4248 (N_4248,N_3312,N_2449);
and U4249 (N_4249,N_3074,N_3292);
or U4250 (N_4250,N_2500,N_2161);
nor U4251 (N_4251,N_3175,N_3320);
nor U4252 (N_4252,N_2441,N_3788);
or U4253 (N_4253,N_3339,N_2911);
and U4254 (N_4254,N_2405,N_2008);
and U4255 (N_4255,N_2043,N_2498);
nor U4256 (N_4256,N_3469,N_3378);
nor U4257 (N_4257,N_3123,N_3761);
or U4258 (N_4258,N_2883,N_3606);
or U4259 (N_4259,N_3248,N_3853);
and U4260 (N_4260,N_2819,N_2713);
nor U4261 (N_4261,N_2617,N_2804);
nor U4262 (N_4262,N_2885,N_2123);
and U4263 (N_4263,N_2363,N_3430);
nor U4264 (N_4264,N_3002,N_2025);
and U4265 (N_4265,N_2259,N_3462);
or U4266 (N_4266,N_3461,N_3650);
and U4267 (N_4267,N_3426,N_2435);
nor U4268 (N_4268,N_2961,N_2685);
and U4269 (N_4269,N_3504,N_2630);
nor U4270 (N_4270,N_2216,N_3051);
nand U4271 (N_4271,N_2444,N_2716);
and U4272 (N_4272,N_3663,N_3529);
nand U4273 (N_4273,N_3190,N_2924);
nor U4274 (N_4274,N_2574,N_2465);
nand U4275 (N_4275,N_2907,N_3473);
nor U4276 (N_4276,N_3629,N_2279);
or U4277 (N_4277,N_3635,N_2922);
nand U4278 (N_4278,N_2620,N_2939);
nor U4279 (N_4279,N_3922,N_3920);
nor U4280 (N_4280,N_3189,N_2797);
nor U4281 (N_4281,N_3243,N_3666);
nand U4282 (N_4282,N_3612,N_2412);
and U4283 (N_4283,N_3806,N_3968);
or U4284 (N_4284,N_2215,N_3927);
nor U4285 (N_4285,N_2943,N_3754);
nand U4286 (N_4286,N_2443,N_3432);
and U4287 (N_4287,N_3911,N_2453);
and U4288 (N_4288,N_3001,N_3684);
nand U4289 (N_4289,N_3678,N_2203);
nand U4290 (N_4290,N_3230,N_2354);
or U4291 (N_4291,N_3481,N_2587);
nor U4292 (N_4292,N_3317,N_2665);
nor U4293 (N_4293,N_2796,N_2332);
nand U4294 (N_4294,N_2146,N_2120);
and U4295 (N_4295,N_2396,N_2810);
or U4296 (N_4296,N_3280,N_3538);
nand U4297 (N_4297,N_3970,N_3041);
nand U4298 (N_4298,N_3961,N_3618);
nor U4299 (N_4299,N_2497,N_2930);
nand U4300 (N_4300,N_3147,N_3028);
nand U4301 (N_4301,N_3453,N_2537);
and U4302 (N_4302,N_3241,N_2648);
nand U4303 (N_4303,N_2289,N_3971);
nor U4304 (N_4304,N_3993,N_2471);
nor U4305 (N_4305,N_3244,N_3345);
nor U4306 (N_4306,N_2867,N_2509);
nand U4307 (N_4307,N_3885,N_3608);
nor U4308 (N_4308,N_2372,N_3818);
or U4309 (N_4309,N_2230,N_3287);
and U4310 (N_4310,N_3215,N_3849);
nor U4311 (N_4311,N_3105,N_2589);
and U4312 (N_4312,N_3013,N_2072);
and U4313 (N_4313,N_3035,N_3936);
nand U4314 (N_4314,N_3523,N_2274);
nand U4315 (N_4315,N_3318,N_3571);
nand U4316 (N_4316,N_3166,N_2101);
nand U4317 (N_4317,N_3136,N_2776);
nand U4318 (N_4318,N_2176,N_3734);
nand U4319 (N_4319,N_3476,N_3226);
or U4320 (N_4320,N_2860,N_3706);
or U4321 (N_4321,N_2105,N_3073);
and U4322 (N_4322,N_2295,N_3803);
nand U4323 (N_4323,N_3156,N_2226);
or U4324 (N_4324,N_2789,N_2917);
or U4325 (N_4325,N_2472,N_2000);
nand U4326 (N_4326,N_2393,N_3380);
or U4327 (N_4327,N_2386,N_3820);
nor U4328 (N_4328,N_2666,N_3862);
nor U4329 (N_4329,N_3484,N_2024);
nor U4330 (N_4330,N_3152,N_2003);
or U4331 (N_4331,N_3262,N_2499);
and U4332 (N_4332,N_3218,N_3128);
or U4333 (N_4333,N_3415,N_3278);
nor U4334 (N_4334,N_2271,N_3047);
nand U4335 (N_4335,N_3254,N_3393);
or U4336 (N_4336,N_3916,N_3143);
nand U4337 (N_4337,N_2406,N_3918);
or U4338 (N_4338,N_2223,N_2940);
nand U4339 (N_4339,N_2030,N_3662);
nor U4340 (N_4340,N_2816,N_3546);
or U4341 (N_4341,N_3205,N_3566);
or U4342 (N_4342,N_3890,N_3437);
nand U4343 (N_4343,N_3644,N_2736);
or U4344 (N_4344,N_3361,N_3944);
or U4345 (N_4345,N_3628,N_3465);
and U4346 (N_4346,N_2638,N_2772);
and U4347 (N_4347,N_2667,N_2196);
and U4348 (N_4348,N_2099,N_3162);
and U4349 (N_4349,N_3111,N_2379);
and U4350 (N_4350,N_2831,N_3680);
and U4351 (N_4351,N_2466,N_3090);
and U4352 (N_4352,N_3264,N_3071);
or U4353 (N_4353,N_2065,N_3100);
and U4354 (N_4354,N_2282,N_3718);
nor U4355 (N_4355,N_3905,N_2021);
and U4356 (N_4356,N_2157,N_2557);
nand U4357 (N_4357,N_2296,N_2272);
and U4358 (N_4358,N_3627,N_2165);
nand U4359 (N_4359,N_2180,N_2947);
or U4360 (N_4360,N_3324,N_3671);
nor U4361 (N_4361,N_3338,N_3005);
nand U4362 (N_4362,N_2361,N_2292);
nor U4363 (N_4363,N_2844,N_3363);
and U4364 (N_4364,N_3531,N_3138);
and U4365 (N_4365,N_3246,N_2348);
or U4366 (N_4366,N_2900,N_3158);
nand U4367 (N_4367,N_2658,N_2383);
nor U4368 (N_4368,N_2408,N_3977);
or U4369 (N_4369,N_3325,N_3999);
nor U4370 (N_4370,N_3959,N_2903);
and U4371 (N_4371,N_3127,N_3515);
nor U4372 (N_4372,N_2790,N_3095);
nand U4373 (N_4373,N_2555,N_3508);
and U4374 (N_4374,N_2004,N_3367);
or U4375 (N_4375,N_2149,N_3383);
nand U4376 (N_4376,N_3892,N_2200);
nor U4377 (N_4377,N_3947,N_2096);
or U4378 (N_4378,N_3031,N_3964);
or U4379 (N_4379,N_3064,N_3365);
or U4380 (N_4380,N_2734,N_3564);
nand U4381 (N_4381,N_2958,N_3410);
nor U4382 (N_4382,N_3375,N_3728);
nand U4383 (N_4383,N_2600,N_3125);
or U4384 (N_4384,N_2809,N_2891);
nand U4385 (N_4385,N_3495,N_3266);
nor U4386 (N_4386,N_2377,N_2121);
nor U4387 (N_4387,N_2777,N_2984);
and U4388 (N_4388,N_2859,N_2905);
nand U4389 (N_4389,N_3585,N_3085);
or U4390 (N_4390,N_3554,N_2436);
and U4391 (N_4391,N_3455,N_2902);
or U4392 (N_4392,N_3845,N_2017);
and U4393 (N_4393,N_3668,N_3990);
and U4394 (N_4394,N_3731,N_2190);
or U4395 (N_4395,N_3982,N_3020);
or U4396 (N_4396,N_2693,N_2643);
and U4397 (N_4397,N_2762,N_3172);
or U4398 (N_4398,N_2874,N_2671);
and U4399 (N_4399,N_3962,N_2632);
and U4400 (N_4400,N_2743,N_2256);
or U4401 (N_4401,N_2767,N_3011);
nor U4402 (N_4402,N_2364,N_3980);
and U4403 (N_4403,N_3674,N_2993);
nand U4404 (N_4404,N_2463,N_2007);
nand U4405 (N_4405,N_2403,N_3670);
nor U4406 (N_4406,N_2546,N_3211);
nor U4407 (N_4407,N_2353,N_2775);
or U4408 (N_4408,N_3659,N_2257);
nor U4409 (N_4409,N_2928,N_3776);
or U4410 (N_4410,N_3154,N_2652);
and U4411 (N_4411,N_2425,N_3493);
and U4412 (N_4412,N_2607,N_3512);
or U4413 (N_4413,N_2069,N_3033);
nand U4414 (N_4414,N_3790,N_3300);
nand U4415 (N_4415,N_2909,N_3265);
or U4416 (N_4416,N_2799,N_3778);
nor U4417 (N_4417,N_2692,N_3753);
and U4418 (N_4418,N_3599,N_3963);
xnor U4419 (N_4419,N_3088,N_2892);
or U4420 (N_4420,N_2783,N_2720);
or U4421 (N_4421,N_2997,N_2420);
and U4422 (N_4422,N_2284,N_3062);
or U4423 (N_4423,N_2375,N_2605);
nand U4424 (N_4424,N_2304,N_3553);
nand U4425 (N_4425,N_3009,N_2544);
or U4426 (N_4426,N_3401,N_3744);
and U4427 (N_4427,N_3006,N_2513);
or U4428 (N_4428,N_3048,N_2758);
nand U4429 (N_4429,N_3607,N_3926);
nand U4430 (N_4430,N_2651,N_2134);
and U4431 (N_4431,N_2704,N_3876);
and U4432 (N_4432,N_3494,N_3501);
nor U4433 (N_4433,N_3157,N_2207);
or U4434 (N_4434,N_2972,N_3010);
nor U4435 (N_4435,N_3467,N_3975);
nor U4436 (N_4436,N_2910,N_3561);
nor U4437 (N_4437,N_2904,N_2757);
nor U4438 (N_4438,N_2518,N_3533);
nor U4439 (N_4439,N_2840,N_2564);
and U4440 (N_4440,N_3667,N_3025);
and U4441 (N_4441,N_2365,N_3034);
nor U4442 (N_4442,N_2037,N_2669);
or U4443 (N_4443,N_2114,N_2109);
or U4444 (N_4444,N_3485,N_2036);
and U4445 (N_4445,N_3562,N_3496);
nand U4446 (N_4446,N_2520,N_3252);
and U4447 (N_4447,N_3081,N_2061);
and U4448 (N_4448,N_2710,N_3682);
nor U4449 (N_4449,N_3707,N_3309);
nand U4450 (N_4450,N_3588,N_3757);
nor U4451 (N_4451,N_3169,N_2612);
and U4452 (N_4452,N_3018,N_3445);
or U4453 (N_4453,N_2531,N_3017);
nand U4454 (N_4454,N_3565,N_3930);
nand U4455 (N_4455,N_3832,N_3866);
and U4456 (N_4456,N_3837,N_3054);
nand U4457 (N_4457,N_2351,N_3433);
or U4458 (N_4458,N_2601,N_3665);
nand U4459 (N_4459,N_2046,N_2560);
nor U4460 (N_4460,N_2338,N_3732);
xor U4461 (N_4461,N_3070,N_3206);
and U4462 (N_4462,N_3574,N_3917);
xor U4463 (N_4463,N_3329,N_3855);
and U4464 (N_4464,N_3691,N_2012);
nor U4465 (N_4465,N_2175,N_2349);
nand U4466 (N_4466,N_3583,N_2322);
or U4467 (N_4467,N_3242,N_2929);
and U4468 (N_4468,N_3315,N_3272);
nor U4469 (N_4469,N_3595,N_2299);
or U4470 (N_4470,N_2325,N_2026);
and U4471 (N_4471,N_3093,N_2394);
or U4472 (N_4472,N_3559,N_3472);
or U4473 (N_4473,N_2357,N_2418);
nand U4474 (N_4474,N_2889,N_2281);
nand U4475 (N_4475,N_2908,N_3014);
or U4476 (N_4476,N_3556,N_3716);
and U4477 (N_4477,N_2013,N_3386);
nand U4478 (N_4478,N_2541,N_3022);
or U4479 (N_4479,N_3180,N_2925);
xnor U4480 (N_4480,N_2102,N_3860);
nor U4481 (N_4481,N_3615,N_3898);
and U4482 (N_4482,N_2694,N_2591);
and U4483 (N_4483,N_3823,N_2066);
and U4484 (N_4484,N_3807,N_2044);
nand U4485 (N_4485,N_3943,N_3165);
or U4486 (N_4486,N_2875,N_3357);
or U4487 (N_4487,N_2266,N_3377);
and U4488 (N_4488,N_3661,N_3783);
nand U4489 (N_4489,N_2641,N_3000);
and U4490 (N_4490,N_3026,N_3223);
or U4491 (N_4491,N_2511,N_2213);
nand U4492 (N_4492,N_2854,N_3657);
nand U4493 (N_4493,N_2079,N_3893);
xnor U4494 (N_4494,N_2091,N_2582);
nand U4495 (N_4495,N_3299,N_3065);
nand U4496 (N_4496,N_3948,N_3638);
nor U4497 (N_4497,N_3526,N_3878);
or U4498 (N_4498,N_2273,N_3392);
nor U4499 (N_4499,N_3256,N_2258);
or U4500 (N_4500,N_3301,N_3865);
nor U4501 (N_4501,N_2604,N_3077);
nor U4502 (N_4502,N_3626,N_2440);
nor U4503 (N_4503,N_2316,N_2586);
or U4504 (N_4504,N_2268,N_2477);
and U4505 (N_4505,N_3831,N_2817);
nand U4506 (N_4506,N_3049,N_2614);
and U4507 (N_4507,N_3498,N_2626);
nor U4508 (N_4508,N_3417,N_3008);
or U4509 (N_4509,N_2986,N_2311);
or U4510 (N_4510,N_2469,N_2771);
nand U4511 (N_4511,N_2702,N_3843);
or U4512 (N_4512,N_2171,N_3981);
and U4513 (N_4513,N_2334,N_3786);
nor U4514 (N_4514,N_3212,N_2937);
nand U4515 (N_4515,N_2422,N_2218);
and U4516 (N_4516,N_3213,N_2241);
or U4517 (N_4517,N_3701,N_2994);
nand U4518 (N_4518,N_3173,N_2077);
or U4519 (N_4519,N_2020,N_3348);
nand U4520 (N_4520,N_2679,N_3016);
nand U4521 (N_4521,N_3421,N_3696);
nand U4522 (N_4522,N_3221,N_2454);
or U4523 (N_4523,N_3998,N_3413);
and U4524 (N_4524,N_2580,N_3679);
nor U4525 (N_4525,N_3441,N_3148);
nor U4526 (N_4526,N_3854,N_3291);
and U4527 (N_4527,N_3313,N_3407);
and U4528 (N_4528,N_2054,N_2049);
and U4529 (N_4529,N_2090,N_2504);
and U4530 (N_4530,N_3586,N_3480);
nor U4531 (N_4531,N_3184,N_3307);
or U4532 (N_4532,N_2445,N_3802);
nor U4533 (N_4533,N_3958,N_2155);
and U4534 (N_4534,N_2801,N_3672);
nor U4535 (N_4535,N_3422,N_2462);
and U4536 (N_4536,N_2955,N_2355);
nor U4537 (N_4537,N_2384,N_2791);
or U4538 (N_4538,N_3738,N_3328);
nor U4539 (N_4539,N_3777,N_2709);
or U4540 (N_4540,N_2056,N_2050);
or U4541 (N_4541,N_2288,N_3185);
and U4542 (N_4542,N_2428,N_2078);
xor U4543 (N_4543,N_3863,N_2863);
nor U4544 (N_4544,N_2382,N_2356);
or U4545 (N_4545,N_3651,N_3032);
or U4546 (N_4546,N_3735,N_2138);
and U4547 (N_4547,N_3076,N_2823);
and U4548 (N_4548,N_3834,N_2554);
nor U4549 (N_4549,N_2621,N_3749);
and U4550 (N_4550,N_2415,N_3572);
nand U4551 (N_4551,N_2878,N_3193);
nand U4552 (N_4552,N_3660,N_3528);
and U4553 (N_4553,N_2569,N_2592);
or U4554 (N_4554,N_2042,N_3624);
nand U4555 (N_4555,N_2494,N_3435);
nand U4556 (N_4556,N_3952,N_3647);
or U4557 (N_4557,N_2343,N_3539);
xor U4558 (N_4558,N_3438,N_2646);
nor U4559 (N_4559,N_3228,N_3029);
or U4560 (N_4560,N_3387,N_3524);
or U4561 (N_4561,N_2117,N_2737);
nand U4562 (N_4562,N_2602,N_2489);
and U4563 (N_4563,N_2562,N_3772);
nor U4564 (N_4564,N_2850,N_2800);
and U4565 (N_4565,N_3525,N_3547);
and U4566 (N_4566,N_2307,N_3631);
or U4567 (N_4567,N_3969,N_2606);
nand U4568 (N_4568,N_3699,N_2276);
and U4569 (N_4569,N_3354,N_3340);
and U4570 (N_4570,N_3536,N_3424);
and U4571 (N_4571,N_3007,N_2825);
or U4572 (N_4572,N_2076,N_2941);
or U4573 (N_4573,N_2830,N_2719);
nor U4574 (N_4574,N_2267,N_3931);
nor U4575 (N_4575,N_3798,N_3284);
nor U4576 (N_4576,N_3388,N_3698);
nand U4577 (N_4577,N_3063,N_3781);
and U4578 (N_4578,N_2319,N_3619);
nand U4579 (N_4579,N_3276,N_2238);
or U4580 (N_4580,N_2495,N_3194);
and U4581 (N_4581,N_2590,N_2995);
and U4582 (N_4582,N_2558,N_2618);
and U4583 (N_4583,N_2898,N_2780);
nand U4584 (N_4584,N_3985,N_3907);
nor U4585 (N_4585,N_2964,N_3121);
nand U4586 (N_4586,N_2448,N_2283);
or U4587 (N_4587,N_2515,N_2644);
nor U4588 (N_4588,N_2306,N_3161);
nand U4589 (N_4589,N_3563,N_3140);
nand U4590 (N_4590,N_2527,N_3748);
nand U4591 (N_4591,N_3038,N_3281);
or U4592 (N_4592,N_2287,N_3763);
and U4593 (N_4593,N_3622,N_3084);
nand U4594 (N_4594,N_2538,N_3658);
and U4595 (N_4595,N_2942,N_2217);
nand U4596 (N_4596,N_3237,N_2022);
or U4597 (N_4597,N_2896,N_3859);
and U4598 (N_4598,N_2083,N_3521);
or U4599 (N_4599,N_3934,N_2629);
or U4600 (N_4600,N_2093,N_2387);
nor U4601 (N_4601,N_2547,N_2487);
or U4602 (N_4602,N_2687,N_3797);
or U4603 (N_4603,N_2341,N_2437);
nor U4604 (N_4604,N_3737,N_2254);
nor U4605 (N_4605,N_2567,N_3986);
and U4606 (N_4606,N_2853,N_2752);
and U4607 (N_4607,N_3712,N_3997);
or U4608 (N_4608,N_3091,N_3552);
nand U4609 (N_4609,N_3762,N_3347);
nand U4610 (N_4610,N_3555,N_2842);
nor U4611 (N_4611,N_3745,N_3994);
or U4612 (N_4612,N_2534,N_2748);
nand U4613 (N_4613,N_3160,N_3816);
nor U4614 (N_4614,N_3474,N_2074);
and U4615 (N_4615,N_3279,N_2739);
nor U4616 (N_4616,N_3839,N_3497);
or U4617 (N_4617,N_2659,N_3871);
and U4618 (N_4618,N_2484,N_2820);
and U4619 (N_4619,N_3259,N_2657);
nand U4620 (N_4620,N_2988,N_3856);
nand U4621 (N_4621,N_2139,N_3915);
nand U4622 (N_4622,N_2933,N_3043);
nand U4623 (N_4623,N_3004,N_3423);
nand U4624 (N_4624,N_3219,N_3045);
or U4625 (N_4625,N_2594,N_2653);
nor U4626 (N_4626,N_3888,N_3836);
or U4627 (N_4627,N_3229,N_2764);
nand U4628 (N_4628,N_3532,N_2960);
nor U4629 (N_4629,N_2373,N_3593);
nand U4630 (N_4630,N_3167,N_2865);
nand U4631 (N_4631,N_2962,N_3846);
and U4632 (N_4632,N_3681,N_2888);
nand U4633 (N_4633,N_2833,N_2486);
nor U4634 (N_4634,N_3412,N_2198);
nand U4635 (N_4635,N_2015,N_2208);
nor U4636 (N_4636,N_2793,N_2524);
nor U4637 (N_4637,N_3263,N_3249);
nand U4638 (N_4638,N_3352,N_3436);
nand U4639 (N_4639,N_2821,N_3273);
or U4640 (N_4640,N_2918,N_2452);
and U4641 (N_4641,N_3178,N_2837);
nand U4642 (N_4642,N_3652,N_2018);
nor U4643 (N_4643,N_2108,N_2262);
nand U4644 (N_4644,N_3551,N_2023);
nand U4645 (N_4645,N_2124,N_2882);
or U4646 (N_4646,N_3604,N_2826);
nor U4647 (N_4647,N_2092,N_3813);
nor U4648 (N_4648,N_2765,N_2052);
nand U4649 (N_4649,N_2718,N_2388);
xnor U4650 (N_4650,N_3641,N_2057);
nand U4651 (N_4651,N_2662,N_2539);
or U4652 (N_4652,N_3385,N_3181);
nor U4653 (N_4653,N_2385,N_3883);
or U4654 (N_4654,N_3382,N_2116);
nand U4655 (N_4655,N_2275,N_3359);
nand U4656 (N_4656,N_2836,N_3092);
nand U4657 (N_4657,N_3891,N_3636);
nand U4658 (N_4658,N_3220,N_3792);
nand U4659 (N_4659,N_3692,N_2152);
nand U4660 (N_4660,N_2829,N_2468);
or U4661 (N_4661,N_2312,N_2344);
nand U4662 (N_4662,N_3950,N_2624);
nor U4663 (N_4663,N_2579,N_3037);
and U4664 (N_4664,N_3541,N_2427);
and U4665 (N_4665,N_2532,N_3198);
or U4666 (N_4666,N_3053,N_2856);
nor U4667 (N_4667,N_2411,N_3596);
or U4668 (N_4668,N_3446,N_2106);
nor U4669 (N_4669,N_2750,N_2631);
or U4670 (N_4670,N_2890,N_3460);
nor U4671 (N_4671,N_2996,N_3176);
nand U4672 (N_4672,N_2543,N_2686);
or U4673 (N_4673,N_2923,N_2451);
or U4674 (N_4674,N_3537,N_2032);
or U4675 (N_4675,N_2861,N_2147);
and U4676 (N_4676,N_3492,N_3225);
nor U4677 (N_4677,N_3685,N_2419);
nor U4678 (N_4678,N_3463,N_2808);
or U4679 (N_4679,N_3145,N_2195);
or U4680 (N_4680,N_3815,N_2570);
and U4681 (N_4681,N_3677,N_3102);
or U4682 (N_4682,N_2572,N_2482);
or U4683 (N_4683,N_2177,N_3972);
or U4684 (N_4684,N_2751,N_3821);
and U4685 (N_4685,N_3069,N_2622);
nand U4686 (N_4686,N_2191,N_2450);
nor U4687 (N_4687,N_3742,N_3875);
or U4688 (N_4688,N_2290,N_3695);
or U4689 (N_4689,N_2588,N_2688);
or U4690 (N_4690,N_3601,N_3217);
nand U4691 (N_4691,N_2464,N_2094);
nor U4692 (N_4692,N_2742,N_3052);
nor U4693 (N_4693,N_2759,N_2164);
nand U4694 (N_4694,N_2205,N_2792);
or U4695 (N_4695,N_3394,N_2862);
or U4696 (N_4696,N_3282,N_2672);
or U4697 (N_4697,N_2725,N_3577);
or U4698 (N_4698,N_3277,N_3058);
and U4699 (N_4699,N_3945,N_3882);
or U4700 (N_4700,N_3840,N_2613);
and U4701 (N_4701,N_3889,N_2285);
nand U4702 (N_4702,N_3609,N_2548);
nand U4703 (N_4703,N_3722,N_2726);
and U4704 (N_4704,N_3232,N_2609);
or U4705 (N_4705,N_3780,N_3703);
nand U4706 (N_4706,N_2479,N_2529);
and U4707 (N_4707,N_2333,N_2985);
nor U4708 (N_4708,N_2001,N_3133);
or U4709 (N_4709,N_3727,N_3267);
nor U4710 (N_4710,N_3872,N_3824);
and U4711 (N_4711,N_2478,N_2220);
nand U4712 (N_4712,N_2851,N_3414);
nor U4713 (N_4713,N_2787,N_2413);
and U4714 (N_4714,N_2795,N_3799);
xor U4715 (N_4715,N_3877,N_3603);
and U4716 (N_4716,N_3705,N_3199);
and U4717 (N_4717,N_2221,N_3979);
and U4718 (N_4718,N_2519,N_3611);
and U4719 (N_4719,N_2881,N_2959);
nor U4720 (N_4720,N_3771,N_2366);
or U4721 (N_4721,N_3804,N_3769);
and U4722 (N_4722,N_3614,N_3697);
and U4723 (N_4723,N_3775,N_2038);
or U4724 (N_4724,N_3358,N_3204);
or U4725 (N_4725,N_3939,N_2699);
nand U4726 (N_4726,N_3149,N_3868);
nand U4727 (N_4727,N_3653,N_2143);
and U4728 (N_4728,N_3913,N_2834);
nor U4729 (N_4729,N_3080,N_2337);
nor U4730 (N_4730,N_2245,N_2512);
nor U4731 (N_4731,N_3132,N_3505);
nand U4732 (N_4732,N_3396,N_3549);
or U4733 (N_4733,N_3222,N_2660);
nor U4734 (N_4734,N_3887,N_3715);
nor U4735 (N_4735,N_2533,N_2019);
or U4736 (N_4736,N_3418,N_2866);
nand U4737 (N_4737,N_3381,N_3342);
nor U4738 (N_4738,N_3730,N_2331);
nand U4739 (N_4739,N_2584,N_3323);
nor U4740 (N_4740,N_2447,N_2753);
or U4741 (N_4741,N_2144,N_2838);
nor U4742 (N_4742,N_2490,N_3137);
and U4743 (N_4743,N_2132,N_3903);
or U4744 (N_4744,N_3759,N_3240);
nor U4745 (N_4745,N_3321,N_3646);
nand U4746 (N_4746,N_2082,N_2070);
nand U4747 (N_4747,N_3584,N_2610);
nand U4748 (N_4748,N_3838,N_2067);
or U4749 (N_4749,N_3932,N_3835);
or U4750 (N_4750,N_3337,N_2367);
or U4751 (N_4751,N_3171,N_2150);
nand U4752 (N_4752,N_3471,N_2968);
and U4753 (N_4753,N_2522,N_2431);
nor U4754 (N_4754,N_2214,N_3015);
nand U4755 (N_4755,N_3825,N_3429);
and U4756 (N_4756,N_3483,N_2921);
nor U4757 (N_4757,N_2404,N_2103);
nor U4758 (N_4758,N_3255,N_3996);
and U4759 (N_4759,N_2953,N_3207);
nand U4760 (N_4760,N_2744,N_3630);
nor U4761 (N_4761,N_3040,N_3351);
nor U4762 (N_4762,N_3163,N_3283);
and U4763 (N_4763,N_3311,N_3669);
nor U4764 (N_4764,N_2721,N_3923);
or U4765 (N_4765,N_3106,N_3114);
or U4766 (N_4766,N_3542,N_3767);
and U4767 (N_4767,N_3967,N_3260);
nor U4768 (N_4768,N_2391,N_2014);
and U4769 (N_4769,N_3168,N_2269);
nand U4770 (N_4770,N_3543,N_2298);
nor U4771 (N_4771,N_2301,N_3251);
nor U4772 (N_4772,N_3146,N_2142);
nand U4773 (N_4773,N_3795,N_2397);
and U4774 (N_4774,N_3988,N_2957);
nand U4775 (N_4775,N_3794,N_3450);
nor U4776 (N_4776,N_3253,N_2080);
nor U4777 (N_4777,N_2153,N_3942);
nand U4778 (N_4778,N_2222,N_3640);
nor U4779 (N_4779,N_2690,N_3693);
nand U4780 (N_4780,N_2779,N_2811);
and U4781 (N_4781,N_2470,N_3057);
nand U4782 (N_4782,N_2199,N_3344);
nor U4783 (N_4783,N_2848,N_3061);
or U4784 (N_4784,N_2399,N_3072);
or U4785 (N_4785,N_2362,N_2392);
or U4786 (N_4786,N_3402,N_3610);
nand U4787 (N_4787,N_3440,N_2884);
nand U4788 (N_4788,N_3739,N_2603);
and U4789 (N_4789,N_2740,N_3733);
or U4790 (N_4790,N_3522,N_2849);
and U4791 (N_4791,N_3589,N_3819);
and U4792 (N_4792,N_3082,N_3909);
nand U4793 (N_4793,N_2919,N_3346);
nand U4794 (N_4794,N_3594,N_3027);
nand U4795 (N_4795,N_3992,N_3880);
and U4796 (N_4796,N_3144,N_3399);
nand U4797 (N_4797,N_2063,N_3210);
or U4798 (N_4798,N_3848,N_2234);
nor U4799 (N_4799,N_3719,N_3270);
nand U4800 (N_4800,N_2749,N_2926);
and U4801 (N_4801,N_3591,N_3987);
or U4802 (N_4802,N_2104,N_2540);
or U4803 (N_4803,N_3096,N_3247);
nor U4804 (N_4804,N_3487,N_3368);
nor U4805 (N_4805,N_2975,N_3874);
nor U4806 (N_4806,N_3793,N_2314);
nor U4807 (N_4807,N_3427,N_3214);
nor U4808 (N_4808,N_3582,N_2585);
nand U4809 (N_4809,N_3617,N_3974);
and U4810 (N_4810,N_2330,N_3902);
and U4811 (N_4811,N_3828,N_3330);
or U4812 (N_4812,N_2668,N_3110);
nor U4813 (N_4813,N_3195,N_2133);
or U4814 (N_4814,N_3186,N_3789);
nand U4815 (N_4815,N_3901,N_3597);
or U4816 (N_4816,N_3949,N_2794);
or U4817 (N_4817,N_3428,N_2158);
and U4818 (N_4818,N_3067,N_2976);
or U4819 (N_4819,N_3322,N_2945);
xnor U4820 (N_4820,N_2578,N_3879);
nand U4821 (N_4821,N_3491,N_3012);
nor U4822 (N_4822,N_3506,N_3580);
nand U4823 (N_4823,N_3126,N_3937);
or U4824 (N_4824,N_3740,N_3319);
and U4825 (N_4825,N_2597,N_3456);
nor U4826 (N_4826,N_2530,N_3598);
and U4827 (N_4827,N_3268,N_2832);
or U4828 (N_4828,N_3634,N_3404);
nor U4829 (N_4829,N_3398,N_3290);
or U4830 (N_4830,N_3197,N_2389);
or U4831 (N_4831,N_2663,N_3336);
nor U4832 (N_4832,N_2980,N_3066);
and U4833 (N_4833,N_2009,N_3296);
nand U4834 (N_4834,N_2062,N_3447);
or U4835 (N_4835,N_3179,N_3118);
nor U4836 (N_4836,N_3196,N_3954);
and U4837 (N_4837,N_3046,N_2774);
nor U4838 (N_4838,N_2858,N_3924);
and U4839 (N_4839,N_3298,N_2277);
and U4840 (N_4840,N_3289,N_2680);
and U4841 (N_4841,N_3633,N_3569);
nor U4842 (N_4842,N_2089,N_2573);
or U4843 (N_4843,N_3216,N_2932);
and U4844 (N_4844,N_2400,N_3800);
nand U4845 (N_4845,N_3908,N_3333);
nand U4846 (N_4846,N_2172,N_2261);
nand U4847 (N_4847,N_3153,N_2029);
or U4848 (N_4848,N_3690,N_2188);
nor U4849 (N_4849,N_3097,N_3384);
or U4850 (N_4850,N_2944,N_2429);
nand U4851 (N_4851,N_2457,N_3419);
or U4852 (N_4852,N_3519,N_3912);
or U4853 (N_4853,N_2576,N_2390);
or U4854 (N_4854,N_3464,N_2733);
xnor U4855 (N_4855,N_2358,N_2682);
and U4856 (N_4856,N_2265,N_3991);
or U4857 (N_4857,N_3517,N_2566);
or U4858 (N_4858,N_2315,N_2460);
nand U4859 (N_4859,N_2912,N_2473);
and U4860 (N_4860,N_2113,N_2769);
nand U4861 (N_4861,N_3389,N_3439);
or U4862 (N_4862,N_2989,N_2075);
or U4863 (N_4863,N_2931,N_3269);
or U4864 (N_4864,N_2763,N_2635);
nand U4865 (N_4865,N_3479,N_3811);
and U4866 (N_4866,N_3928,N_3200);
nand U4867 (N_4867,N_2954,N_2130);
nand U4868 (N_4868,N_3861,N_3224);
or U4869 (N_4869,N_3827,N_2170);
or U4870 (N_4870,N_3288,N_2209);
nor U4871 (N_4871,N_3581,N_3886);
nor U4872 (N_4872,N_2675,N_3639);
or U4873 (N_4873,N_2722,N_3768);
nand U4874 (N_4874,N_2871,N_2684);
or U4875 (N_4875,N_3720,N_3104);
and U4876 (N_4876,N_3867,N_2421);
and U4877 (N_4877,N_3817,N_3443);
nor U4878 (N_4878,N_3710,N_3209);
and U4879 (N_4879,N_3844,N_2639);
and U4880 (N_4880,N_2336,N_3202);
nand U4881 (N_4881,N_2841,N_3459);
and U4882 (N_4882,N_3575,N_3286);
nand U4883 (N_4883,N_3376,N_2456);
and U4884 (N_4884,N_2294,N_3466);
and U4885 (N_4885,N_2156,N_3233);
nor U4886 (N_4886,N_2051,N_3921);
or U4887 (N_4887,N_2745,N_2187);
xor U4888 (N_4888,N_3120,N_2194);
nor U4889 (N_4889,N_3683,N_3366);
and U4890 (N_4890,N_3632,N_2948);
and U4891 (N_4891,N_2474,N_3557);
or U4892 (N_4892,N_3530,N_2028);
or U4893 (N_4893,N_3721,N_2204);
nor U4894 (N_4894,N_2893,N_2625);
or U4895 (N_4895,N_2310,N_3513);
or U4896 (N_4896,N_3573,N_2446);
and U4897 (N_4897,N_2212,N_2291);
nor U4898 (N_4898,N_2992,N_2376);
or U4899 (N_4899,N_3649,N_2712);
and U4900 (N_4900,N_2255,N_2788);
or U4901 (N_4901,N_3098,N_2766);
nor U4902 (N_4902,N_3869,N_3686);
or U4903 (N_4903,N_2784,N_2697);
nand U4904 (N_4904,N_3403,N_2201);
and U4905 (N_4905,N_2915,N_2828);
nand U4906 (N_4906,N_3785,N_3379);
or U4907 (N_4907,N_3751,N_2664);
and U4908 (N_4908,N_3976,N_3420);
or U4909 (N_4909,N_3250,N_3736);
and U4910 (N_4910,N_2979,N_3208);
nor U4911 (N_4911,N_3870,N_2060);
and U4912 (N_4912,N_2350,N_2812);
and U4913 (N_4913,N_2206,N_3372);
and U4914 (N_4914,N_3257,N_2695);
nor U4915 (N_4915,N_2717,N_3933);
nor U4916 (N_4916,N_2179,N_3094);
nor U4917 (N_4917,N_3704,N_2086);
nor U4918 (N_4918,N_2193,N_2654);
and U4919 (N_4919,N_2503,N_2059);
or U4920 (N_4920,N_2381,N_2990);
and U4921 (N_4921,N_3488,N_2901);
or U4922 (N_4922,N_2126,N_3548);
nand U4923 (N_4923,N_3675,N_2502);
nand U4924 (N_4924,N_3726,N_3620);
nor U4925 (N_4925,N_2730,N_3003);
and U4926 (N_4926,N_3941,N_2359);
nor U4927 (N_4927,N_3714,N_3227);
and U4928 (N_4928,N_3293,N_3984);
nand U4929 (N_4929,N_2308,N_3864);
nor U4930 (N_4930,N_3174,N_3274);
and U4931 (N_4931,N_2628,N_2327);
and U4932 (N_4932,N_2058,N_3452);
nand U4933 (N_4933,N_3141,N_2637);
and U4934 (N_4934,N_3327,N_3919);
and U4935 (N_4935,N_2492,N_2746);
and U4936 (N_4936,N_2596,N_3899);
and U4937 (N_4937,N_3482,N_3177);
nor U4938 (N_4938,N_3477,N_3457);
nand U4939 (N_4939,N_2248,N_2225);
nand U4940 (N_4940,N_2084,N_2952);
and U4941 (N_4941,N_3940,N_2345);
nand U4942 (N_4942,N_3535,N_2131);
and U4943 (N_4943,N_3042,N_3341);
nor U4944 (N_4944,N_2510,N_2202);
or U4945 (N_4945,N_3370,N_3055);
and U4946 (N_4946,N_2868,N_3760);
and U4947 (N_4947,N_2711,N_3245);
nand U4948 (N_4948,N_2481,N_2129);
nor U4949 (N_4949,N_3159,N_3520);
nand U4950 (N_4950,N_2983,N_2095);
nor U4951 (N_4951,N_3294,N_2728);
nor U4952 (N_4952,N_3842,N_3758);
nor U4953 (N_4953,N_3109,N_2135);
nor U4954 (N_4954,N_2137,N_2485);
and U4955 (N_4955,N_2782,N_3355);
and U4956 (N_4956,N_2496,N_2561);
nand U4957 (N_4957,N_2374,N_2615);
and U4958 (N_4958,N_2010,N_2741);
and U4959 (N_4959,N_2581,N_3826);
or U4960 (N_4960,N_2608,N_2260);
and U4961 (N_4961,N_2627,N_3847);
nand U4962 (N_4962,N_2977,N_2870);
and U4963 (N_4963,N_2814,N_3444);
or U4964 (N_4964,N_3747,N_2439);
nor U4965 (N_4965,N_2148,N_3750);
nand U4966 (N_4966,N_3434,N_3643);
or U4967 (N_4967,N_2916,N_2678);
or U4968 (N_4968,N_2505,N_3621);
nand U4969 (N_4969,N_3752,N_3694);
or U4970 (N_4970,N_2813,N_2335);
nand U4971 (N_4971,N_2965,N_3709);
and U4972 (N_4972,N_2521,N_3796);
nor U4973 (N_4973,N_2599,N_3951);
nand U4974 (N_4974,N_3036,N_3131);
nand U4975 (N_4975,N_3502,N_3397);
nand U4976 (N_4976,N_2824,N_2035);
nor U4977 (N_4977,N_2575,N_3115);
or U4978 (N_4978,N_2873,N_2650);
or U4979 (N_4979,N_2895,N_3391);
and U4980 (N_4980,N_3729,N_2647);
nor U4981 (N_4981,N_3567,N_2847);
and U4982 (N_4982,N_2320,N_2219);
nand U4983 (N_4983,N_2424,N_2703);
and U4984 (N_4984,N_2501,N_2395);
and U4985 (N_4985,N_3059,N_2119);
nor U4986 (N_4986,N_2339,N_2239);
nand U4987 (N_4987,N_3642,N_2442);
nor U4988 (N_4988,N_2151,N_2368);
nor U4989 (N_4989,N_2098,N_3139);
nand U4990 (N_4990,N_3578,N_3741);
or U4991 (N_4991,N_2523,N_3285);
nor U4992 (N_4992,N_2318,N_3101);
nor U4993 (N_4993,N_2545,N_3896);
nand U4994 (N_4994,N_2480,N_2807);
nor U4995 (N_4995,N_2088,N_2514);
nor U4996 (N_4996,N_2263,N_3702);
or U4997 (N_4997,N_2002,N_3425);
or U4998 (N_4998,N_3850,N_3405);
and U4999 (N_4999,N_2228,N_3231);
nor U5000 (N_5000,N_2148,N_3982);
or U5001 (N_5001,N_3004,N_2694);
or U5002 (N_5002,N_2200,N_2900);
or U5003 (N_5003,N_3407,N_3639);
or U5004 (N_5004,N_3860,N_3869);
nor U5005 (N_5005,N_3673,N_3386);
or U5006 (N_5006,N_2355,N_2021);
and U5007 (N_5007,N_2026,N_3749);
and U5008 (N_5008,N_3986,N_2685);
nor U5009 (N_5009,N_2700,N_3965);
nor U5010 (N_5010,N_2399,N_3042);
nand U5011 (N_5011,N_2515,N_2189);
and U5012 (N_5012,N_3388,N_3131);
nor U5013 (N_5013,N_2630,N_3136);
or U5014 (N_5014,N_2814,N_3649);
and U5015 (N_5015,N_2132,N_2526);
nand U5016 (N_5016,N_2842,N_2168);
nor U5017 (N_5017,N_2707,N_3620);
nor U5018 (N_5018,N_2619,N_2359);
nand U5019 (N_5019,N_3321,N_3513);
nor U5020 (N_5020,N_3436,N_3082);
nor U5021 (N_5021,N_3141,N_2818);
nand U5022 (N_5022,N_3144,N_2059);
or U5023 (N_5023,N_3993,N_2999);
nand U5024 (N_5024,N_2230,N_2013);
and U5025 (N_5025,N_3524,N_3123);
nand U5026 (N_5026,N_2987,N_2588);
and U5027 (N_5027,N_3804,N_3354);
nor U5028 (N_5028,N_2475,N_2426);
and U5029 (N_5029,N_2690,N_2820);
and U5030 (N_5030,N_2110,N_3929);
nand U5031 (N_5031,N_2652,N_2369);
or U5032 (N_5032,N_2273,N_3631);
nor U5033 (N_5033,N_3584,N_3626);
or U5034 (N_5034,N_2947,N_2484);
or U5035 (N_5035,N_3729,N_2523);
nand U5036 (N_5036,N_3165,N_3345);
nor U5037 (N_5037,N_3602,N_3984);
and U5038 (N_5038,N_2891,N_2569);
or U5039 (N_5039,N_3480,N_2611);
nor U5040 (N_5040,N_2692,N_2285);
or U5041 (N_5041,N_2260,N_3493);
or U5042 (N_5042,N_3415,N_2814);
nor U5043 (N_5043,N_2699,N_3763);
or U5044 (N_5044,N_2788,N_3995);
and U5045 (N_5045,N_3326,N_3981);
or U5046 (N_5046,N_2224,N_2794);
and U5047 (N_5047,N_3708,N_2800);
and U5048 (N_5048,N_2739,N_2598);
nor U5049 (N_5049,N_3610,N_3705);
nand U5050 (N_5050,N_2326,N_3362);
and U5051 (N_5051,N_2736,N_3981);
and U5052 (N_5052,N_2517,N_3195);
nand U5053 (N_5053,N_3516,N_2778);
and U5054 (N_5054,N_3797,N_3564);
or U5055 (N_5055,N_3747,N_3642);
nor U5056 (N_5056,N_2976,N_2227);
nand U5057 (N_5057,N_3910,N_2882);
and U5058 (N_5058,N_3030,N_3583);
nor U5059 (N_5059,N_3624,N_2552);
and U5060 (N_5060,N_3862,N_2921);
xnor U5061 (N_5061,N_3764,N_2343);
and U5062 (N_5062,N_2673,N_2791);
or U5063 (N_5063,N_3227,N_2149);
nor U5064 (N_5064,N_2345,N_3982);
xnor U5065 (N_5065,N_2731,N_3761);
or U5066 (N_5066,N_2125,N_2665);
nor U5067 (N_5067,N_3739,N_2140);
or U5068 (N_5068,N_3847,N_3585);
and U5069 (N_5069,N_3235,N_3522);
nand U5070 (N_5070,N_3378,N_3698);
nor U5071 (N_5071,N_3200,N_2624);
or U5072 (N_5072,N_3776,N_3230);
or U5073 (N_5073,N_2597,N_3782);
and U5074 (N_5074,N_3023,N_2763);
or U5075 (N_5075,N_3677,N_3089);
nor U5076 (N_5076,N_2677,N_2993);
or U5077 (N_5077,N_3271,N_3579);
nor U5078 (N_5078,N_2939,N_3765);
nand U5079 (N_5079,N_3550,N_2130);
and U5080 (N_5080,N_3930,N_3714);
or U5081 (N_5081,N_2780,N_2788);
and U5082 (N_5082,N_3837,N_2848);
or U5083 (N_5083,N_3526,N_3826);
and U5084 (N_5084,N_3098,N_3303);
or U5085 (N_5085,N_3238,N_2636);
nand U5086 (N_5086,N_2881,N_3159);
nand U5087 (N_5087,N_3521,N_2997);
and U5088 (N_5088,N_3574,N_2509);
nor U5089 (N_5089,N_3998,N_3788);
and U5090 (N_5090,N_3663,N_2324);
or U5091 (N_5091,N_2489,N_2798);
nand U5092 (N_5092,N_3142,N_2713);
or U5093 (N_5093,N_2413,N_3123);
nor U5094 (N_5094,N_2484,N_3110);
and U5095 (N_5095,N_3714,N_3334);
and U5096 (N_5096,N_2478,N_2497);
nor U5097 (N_5097,N_3202,N_3325);
xnor U5098 (N_5098,N_2124,N_3546);
or U5099 (N_5099,N_3157,N_2176);
and U5100 (N_5100,N_3717,N_3286);
nand U5101 (N_5101,N_3959,N_3363);
or U5102 (N_5102,N_2186,N_2861);
and U5103 (N_5103,N_2342,N_2013);
and U5104 (N_5104,N_2786,N_3090);
nor U5105 (N_5105,N_3966,N_3994);
or U5106 (N_5106,N_3782,N_3671);
nor U5107 (N_5107,N_3093,N_2815);
nand U5108 (N_5108,N_3006,N_2816);
nand U5109 (N_5109,N_2081,N_2264);
nand U5110 (N_5110,N_2395,N_2737);
or U5111 (N_5111,N_2808,N_3717);
nor U5112 (N_5112,N_2749,N_2671);
and U5113 (N_5113,N_3877,N_3606);
nand U5114 (N_5114,N_3287,N_2065);
or U5115 (N_5115,N_3249,N_3831);
or U5116 (N_5116,N_3374,N_2968);
or U5117 (N_5117,N_3654,N_2651);
nand U5118 (N_5118,N_2766,N_3980);
and U5119 (N_5119,N_3551,N_3663);
nor U5120 (N_5120,N_2214,N_3961);
or U5121 (N_5121,N_2534,N_3606);
and U5122 (N_5122,N_2744,N_3267);
nor U5123 (N_5123,N_3513,N_3366);
nand U5124 (N_5124,N_3407,N_2396);
and U5125 (N_5125,N_3179,N_3161);
or U5126 (N_5126,N_3042,N_3030);
nor U5127 (N_5127,N_3217,N_2350);
nor U5128 (N_5128,N_3867,N_2202);
and U5129 (N_5129,N_2362,N_3516);
nor U5130 (N_5130,N_2587,N_3444);
nor U5131 (N_5131,N_3174,N_3969);
nand U5132 (N_5132,N_3721,N_3088);
nor U5133 (N_5133,N_3100,N_3922);
nand U5134 (N_5134,N_2109,N_3401);
nand U5135 (N_5135,N_2503,N_3769);
nor U5136 (N_5136,N_3442,N_3822);
and U5137 (N_5137,N_2006,N_3841);
and U5138 (N_5138,N_2432,N_3795);
or U5139 (N_5139,N_3425,N_2345);
or U5140 (N_5140,N_3439,N_3079);
or U5141 (N_5141,N_2533,N_3574);
and U5142 (N_5142,N_2101,N_2138);
or U5143 (N_5143,N_2559,N_2070);
and U5144 (N_5144,N_2419,N_3278);
nand U5145 (N_5145,N_3065,N_3898);
nor U5146 (N_5146,N_2502,N_2945);
and U5147 (N_5147,N_3883,N_3637);
nand U5148 (N_5148,N_2288,N_3472);
or U5149 (N_5149,N_2042,N_2732);
nor U5150 (N_5150,N_3382,N_3931);
or U5151 (N_5151,N_2575,N_2250);
or U5152 (N_5152,N_3453,N_2938);
and U5153 (N_5153,N_3727,N_2437);
and U5154 (N_5154,N_2268,N_2719);
or U5155 (N_5155,N_2031,N_2222);
or U5156 (N_5156,N_2883,N_2670);
and U5157 (N_5157,N_3413,N_2731);
nand U5158 (N_5158,N_3639,N_2787);
or U5159 (N_5159,N_2647,N_2719);
nor U5160 (N_5160,N_3508,N_3627);
nor U5161 (N_5161,N_2434,N_3345);
and U5162 (N_5162,N_2218,N_2728);
and U5163 (N_5163,N_3021,N_2425);
or U5164 (N_5164,N_3453,N_3508);
nor U5165 (N_5165,N_2210,N_3991);
nand U5166 (N_5166,N_3886,N_3497);
and U5167 (N_5167,N_3538,N_3934);
or U5168 (N_5168,N_2118,N_2440);
and U5169 (N_5169,N_2403,N_3565);
or U5170 (N_5170,N_2957,N_3165);
nand U5171 (N_5171,N_2453,N_2891);
nand U5172 (N_5172,N_2463,N_3842);
or U5173 (N_5173,N_3395,N_2465);
nor U5174 (N_5174,N_2483,N_3727);
and U5175 (N_5175,N_2425,N_3382);
or U5176 (N_5176,N_2106,N_2203);
and U5177 (N_5177,N_2201,N_2117);
nor U5178 (N_5178,N_3054,N_2901);
or U5179 (N_5179,N_3173,N_2868);
and U5180 (N_5180,N_2115,N_3029);
nor U5181 (N_5181,N_2428,N_2922);
and U5182 (N_5182,N_3488,N_3287);
and U5183 (N_5183,N_3249,N_3874);
and U5184 (N_5184,N_3978,N_2184);
nor U5185 (N_5185,N_2527,N_3323);
and U5186 (N_5186,N_3304,N_2985);
nand U5187 (N_5187,N_3351,N_2910);
nand U5188 (N_5188,N_2061,N_3335);
nor U5189 (N_5189,N_2591,N_2974);
and U5190 (N_5190,N_2172,N_3692);
nor U5191 (N_5191,N_2719,N_3119);
and U5192 (N_5192,N_3051,N_3232);
or U5193 (N_5193,N_2328,N_3336);
nor U5194 (N_5194,N_2902,N_2202);
nor U5195 (N_5195,N_2521,N_3371);
nand U5196 (N_5196,N_2995,N_2925);
nor U5197 (N_5197,N_2185,N_2221);
and U5198 (N_5198,N_3332,N_3881);
nor U5199 (N_5199,N_3511,N_3030);
nor U5200 (N_5200,N_3408,N_2266);
nor U5201 (N_5201,N_2292,N_3533);
nand U5202 (N_5202,N_3850,N_3536);
nor U5203 (N_5203,N_3174,N_2518);
or U5204 (N_5204,N_3488,N_3057);
nor U5205 (N_5205,N_2348,N_2942);
nand U5206 (N_5206,N_2976,N_3783);
nand U5207 (N_5207,N_3654,N_3338);
and U5208 (N_5208,N_3771,N_2847);
or U5209 (N_5209,N_2757,N_2026);
or U5210 (N_5210,N_2714,N_3998);
xnor U5211 (N_5211,N_2874,N_3535);
nand U5212 (N_5212,N_3514,N_3460);
nor U5213 (N_5213,N_3870,N_3469);
or U5214 (N_5214,N_2266,N_2790);
or U5215 (N_5215,N_3337,N_3737);
nor U5216 (N_5216,N_3684,N_3182);
nand U5217 (N_5217,N_2145,N_2412);
or U5218 (N_5218,N_2272,N_3815);
and U5219 (N_5219,N_2543,N_3327);
and U5220 (N_5220,N_2099,N_3779);
nor U5221 (N_5221,N_2764,N_2831);
nand U5222 (N_5222,N_2689,N_2296);
nand U5223 (N_5223,N_3312,N_3492);
nand U5224 (N_5224,N_2923,N_3895);
nand U5225 (N_5225,N_2973,N_2134);
and U5226 (N_5226,N_3982,N_2087);
nand U5227 (N_5227,N_2133,N_2718);
nor U5228 (N_5228,N_3745,N_3452);
nor U5229 (N_5229,N_2759,N_2074);
nor U5230 (N_5230,N_2140,N_2332);
and U5231 (N_5231,N_3632,N_2203);
or U5232 (N_5232,N_3792,N_3952);
nand U5233 (N_5233,N_2823,N_2410);
and U5234 (N_5234,N_3381,N_3719);
and U5235 (N_5235,N_3736,N_2307);
nand U5236 (N_5236,N_3112,N_2787);
or U5237 (N_5237,N_3239,N_2152);
or U5238 (N_5238,N_3805,N_3328);
xnor U5239 (N_5239,N_3812,N_2385);
or U5240 (N_5240,N_2845,N_3284);
nor U5241 (N_5241,N_3713,N_2211);
nand U5242 (N_5242,N_2525,N_2794);
nand U5243 (N_5243,N_3191,N_3305);
nand U5244 (N_5244,N_3282,N_3138);
nor U5245 (N_5245,N_3337,N_3373);
nand U5246 (N_5246,N_2785,N_2318);
and U5247 (N_5247,N_3146,N_2868);
nor U5248 (N_5248,N_2241,N_3707);
and U5249 (N_5249,N_2937,N_2819);
and U5250 (N_5250,N_2329,N_3141);
nor U5251 (N_5251,N_2619,N_3982);
and U5252 (N_5252,N_2212,N_3560);
nor U5253 (N_5253,N_3084,N_3085);
and U5254 (N_5254,N_3621,N_3834);
nor U5255 (N_5255,N_3088,N_2192);
and U5256 (N_5256,N_2420,N_2429);
nand U5257 (N_5257,N_3817,N_2299);
nand U5258 (N_5258,N_3534,N_3715);
nor U5259 (N_5259,N_2889,N_2482);
nor U5260 (N_5260,N_2875,N_3210);
nor U5261 (N_5261,N_3563,N_2333);
or U5262 (N_5262,N_2699,N_3429);
or U5263 (N_5263,N_2969,N_3623);
or U5264 (N_5264,N_3541,N_2038);
nor U5265 (N_5265,N_2932,N_2393);
and U5266 (N_5266,N_2395,N_3508);
and U5267 (N_5267,N_2375,N_2463);
nand U5268 (N_5268,N_2794,N_3460);
and U5269 (N_5269,N_3252,N_2675);
or U5270 (N_5270,N_2185,N_3192);
nor U5271 (N_5271,N_3915,N_3555);
or U5272 (N_5272,N_3081,N_2969);
and U5273 (N_5273,N_2504,N_2654);
and U5274 (N_5274,N_3788,N_3025);
or U5275 (N_5275,N_3894,N_3573);
nor U5276 (N_5276,N_3484,N_3497);
nor U5277 (N_5277,N_3088,N_3753);
nor U5278 (N_5278,N_3200,N_3703);
or U5279 (N_5279,N_2715,N_3775);
xnor U5280 (N_5280,N_2283,N_3096);
nand U5281 (N_5281,N_2740,N_2148);
nand U5282 (N_5282,N_3564,N_3289);
nor U5283 (N_5283,N_2088,N_3413);
nor U5284 (N_5284,N_3050,N_2898);
nor U5285 (N_5285,N_3830,N_2038);
and U5286 (N_5286,N_2631,N_2545);
nor U5287 (N_5287,N_3219,N_3483);
nor U5288 (N_5288,N_3404,N_3949);
nand U5289 (N_5289,N_3520,N_3366);
nor U5290 (N_5290,N_3512,N_3754);
nand U5291 (N_5291,N_3881,N_2800);
and U5292 (N_5292,N_3236,N_3173);
nor U5293 (N_5293,N_2674,N_3028);
nor U5294 (N_5294,N_2901,N_2836);
nor U5295 (N_5295,N_2081,N_3423);
and U5296 (N_5296,N_2179,N_2428);
nor U5297 (N_5297,N_2587,N_2465);
or U5298 (N_5298,N_3023,N_3977);
nor U5299 (N_5299,N_2881,N_2297);
nor U5300 (N_5300,N_3917,N_2199);
or U5301 (N_5301,N_3370,N_2360);
and U5302 (N_5302,N_3156,N_3285);
or U5303 (N_5303,N_2089,N_3533);
nor U5304 (N_5304,N_3324,N_3800);
or U5305 (N_5305,N_2892,N_2298);
or U5306 (N_5306,N_2835,N_2586);
and U5307 (N_5307,N_2376,N_2256);
nand U5308 (N_5308,N_2372,N_3717);
nor U5309 (N_5309,N_3732,N_3611);
nand U5310 (N_5310,N_2033,N_3733);
or U5311 (N_5311,N_3216,N_3682);
and U5312 (N_5312,N_2956,N_3482);
and U5313 (N_5313,N_2462,N_3652);
nand U5314 (N_5314,N_2737,N_2591);
nand U5315 (N_5315,N_3577,N_3035);
nand U5316 (N_5316,N_2992,N_2965);
nand U5317 (N_5317,N_2256,N_2251);
nor U5318 (N_5318,N_2541,N_2940);
nor U5319 (N_5319,N_3791,N_3380);
nand U5320 (N_5320,N_3188,N_2121);
nor U5321 (N_5321,N_2243,N_2706);
nor U5322 (N_5322,N_3387,N_3217);
nor U5323 (N_5323,N_2812,N_2540);
or U5324 (N_5324,N_2601,N_3869);
and U5325 (N_5325,N_3814,N_3826);
nand U5326 (N_5326,N_2974,N_2262);
and U5327 (N_5327,N_2803,N_2911);
and U5328 (N_5328,N_2520,N_3963);
or U5329 (N_5329,N_3055,N_3867);
and U5330 (N_5330,N_3745,N_2902);
or U5331 (N_5331,N_2501,N_3787);
nor U5332 (N_5332,N_2592,N_2806);
or U5333 (N_5333,N_3311,N_2891);
or U5334 (N_5334,N_3373,N_2624);
nor U5335 (N_5335,N_2386,N_3900);
or U5336 (N_5336,N_2271,N_2429);
or U5337 (N_5337,N_2391,N_2287);
nor U5338 (N_5338,N_2860,N_2518);
nand U5339 (N_5339,N_2555,N_2587);
and U5340 (N_5340,N_2414,N_3319);
or U5341 (N_5341,N_3607,N_3744);
or U5342 (N_5342,N_2756,N_2312);
nand U5343 (N_5343,N_2437,N_2066);
nand U5344 (N_5344,N_3123,N_3889);
nand U5345 (N_5345,N_3381,N_3081);
nand U5346 (N_5346,N_3721,N_3015);
nor U5347 (N_5347,N_3568,N_2716);
and U5348 (N_5348,N_3821,N_2130);
and U5349 (N_5349,N_3435,N_2080);
and U5350 (N_5350,N_2917,N_2077);
nand U5351 (N_5351,N_3574,N_2501);
and U5352 (N_5352,N_3485,N_3946);
and U5353 (N_5353,N_2900,N_3330);
and U5354 (N_5354,N_2065,N_3292);
xor U5355 (N_5355,N_3191,N_3748);
nor U5356 (N_5356,N_2126,N_2929);
nor U5357 (N_5357,N_2334,N_2313);
and U5358 (N_5358,N_2992,N_2536);
and U5359 (N_5359,N_3403,N_2318);
nor U5360 (N_5360,N_3198,N_3102);
nor U5361 (N_5361,N_3217,N_2982);
or U5362 (N_5362,N_2342,N_2483);
nor U5363 (N_5363,N_3395,N_2301);
nand U5364 (N_5364,N_3440,N_3072);
or U5365 (N_5365,N_3895,N_2399);
nor U5366 (N_5366,N_2154,N_2210);
and U5367 (N_5367,N_3574,N_2070);
nor U5368 (N_5368,N_3684,N_3915);
and U5369 (N_5369,N_3458,N_2092);
or U5370 (N_5370,N_2962,N_3412);
nor U5371 (N_5371,N_2915,N_3066);
or U5372 (N_5372,N_3654,N_2539);
or U5373 (N_5373,N_2432,N_3307);
and U5374 (N_5374,N_2316,N_2198);
nand U5375 (N_5375,N_3327,N_2638);
nand U5376 (N_5376,N_2305,N_3165);
nor U5377 (N_5377,N_2543,N_2002);
nand U5378 (N_5378,N_2821,N_3635);
or U5379 (N_5379,N_3789,N_2389);
or U5380 (N_5380,N_3649,N_2420);
nor U5381 (N_5381,N_3292,N_3991);
and U5382 (N_5382,N_2212,N_3358);
nor U5383 (N_5383,N_2175,N_2067);
nand U5384 (N_5384,N_2060,N_2644);
nand U5385 (N_5385,N_2124,N_3629);
or U5386 (N_5386,N_2314,N_2293);
or U5387 (N_5387,N_2229,N_2766);
nand U5388 (N_5388,N_3824,N_2031);
nor U5389 (N_5389,N_2676,N_2129);
nand U5390 (N_5390,N_3634,N_2751);
nor U5391 (N_5391,N_2473,N_3358);
and U5392 (N_5392,N_3254,N_3638);
or U5393 (N_5393,N_2886,N_3180);
nand U5394 (N_5394,N_2351,N_2867);
nor U5395 (N_5395,N_3936,N_2656);
nor U5396 (N_5396,N_3509,N_2402);
nor U5397 (N_5397,N_2629,N_3445);
or U5398 (N_5398,N_2131,N_2555);
nand U5399 (N_5399,N_3635,N_2522);
or U5400 (N_5400,N_3474,N_2929);
nor U5401 (N_5401,N_3855,N_2428);
nand U5402 (N_5402,N_2696,N_3588);
or U5403 (N_5403,N_3560,N_2052);
nor U5404 (N_5404,N_2423,N_3529);
nor U5405 (N_5405,N_3138,N_3789);
nand U5406 (N_5406,N_2341,N_3558);
nand U5407 (N_5407,N_2529,N_3821);
or U5408 (N_5408,N_2614,N_2209);
and U5409 (N_5409,N_2231,N_2206);
and U5410 (N_5410,N_3293,N_3523);
nor U5411 (N_5411,N_2075,N_3687);
and U5412 (N_5412,N_3629,N_2025);
or U5413 (N_5413,N_3906,N_2551);
and U5414 (N_5414,N_3429,N_2372);
nand U5415 (N_5415,N_3436,N_2108);
and U5416 (N_5416,N_3220,N_2998);
nand U5417 (N_5417,N_2793,N_2124);
nand U5418 (N_5418,N_2023,N_3636);
nand U5419 (N_5419,N_2915,N_2728);
nor U5420 (N_5420,N_2431,N_2892);
nor U5421 (N_5421,N_3927,N_3133);
nand U5422 (N_5422,N_3505,N_3455);
or U5423 (N_5423,N_3644,N_3228);
or U5424 (N_5424,N_2220,N_3978);
or U5425 (N_5425,N_2528,N_3349);
nand U5426 (N_5426,N_3887,N_3332);
nand U5427 (N_5427,N_2587,N_2521);
nand U5428 (N_5428,N_3280,N_2661);
and U5429 (N_5429,N_3166,N_3340);
nor U5430 (N_5430,N_3708,N_2935);
and U5431 (N_5431,N_3228,N_2841);
nand U5432 (N_5432,N_3217,N_3612);
nand U5433 (N_5433,N_3776,N_3468);
and U5434 (N_5434,N_3317,N_2129);
or U5435 (N_5435,N_3882,N_2297);
nor U5436 (N_5436,N_3234,N_2001);
nand U5437 (N_5437,N_2848,N_2310);
and U5438 (N_5438,N_3273,N_3720);
or U5439 (N_5439,N_3293,N_3886);
nor U5440 (N_5440,N_3858,N_3849);
nand U5441 (N_5441,N_2897,N_2331);
and U5442 (N_5442,N_3326,N_2498);
nor U5443 (N_5443,N_2425,N_3085);
nor U5444 (N_5444,N_3491,N_2737);
and U5445 (N_5445,N_3295,N_3151);
or U5446 (N_5446,N_3812,N_3267);
nand U5447 (N_5447,N_3212,N_2121);
nor U5448 (N_5448,N_3389,N_3052);
and U5449 (N_5449,N_3446,N_3476);
or U5450 (N_5450,N_3759,N_2064);
and U5451 (N_5451,N_2804,N_3310);
and U5452 (N_5452,N_3993,N_2718);
nand U5453 (N_5453,N_2778,N_2158);
or U5454 (N_5454,N_2271,N_2242);
and U5455 (N_5455,N_3593,N_3541);
nor U5456 (N_5456,N_3422,N_3610);
nand U5457 (N_5457,N_2366,N_3050);
nor U5458 (N_5458,N_2585,N_2637);
or U5459 (N_5459,N_3978,N_3833);
xor U5460 (N_5460,N_2840,N_3664);
nor U5461 (N_5461,N_3422,N_2004);
nor U5462 (N_5462,N_2080,N_2453);
or U5463 (N_5463,N_3496,N_2740);
and U5464 (N_5464,N_3469,N_3185);
and U5465 (N_5465,N_3015,N_2151);
and U5466 (N_5466,N_2354,N_2616);
nand U5467 (N_5467,N_3341,N_2422);
and U5468 (N_5468,N_2268,N_2100);
nand U5469 (N_5469,N_2053,N_3526);
nor U5470 (N_5470,N_3901,N_2835);
or U5471 (N_5471,N_2305,N_3572);
nand U5472 (N_5472,N_3305,N_2948);
nor U5473 (N_5473,N_2914,N_2551);
or U5474 (N_5474,N_3396,N_3217);
or U5475 (N_5475,N_2134,N_2959);
nor U5476 (N_5476,N_3678,N_3853);
xnor U5477 (N_5477,N_2511,N_3028);
or U5478 (N_5478,N_2762,N_2266);
nand U5479 (N_5479,N_3774,N_2400);
nor U5480 (N_5480,N_2799,N_2504);
or U5481 (N_5481,N_2725,N_2105);
or U5482 (N_5482,N_2929,N_3148);
nor U5483 (N_5483,N_3614,N_2614);
nor U5484 (N_5484,N_3905,N_3466);
nand U5485 (N_5485,N_2146,N_3516);
and U5486 (N_5486,N_2686,N_3573);
and U5487 (N_5487,N_3151,N_3483);
nor U5488 (N_5488,N_3720,N_3477);
and U5489 (N_5489,N_3872,N_3070);
nand U5490 (N_5490,N_2938,N_2269);
nand U5491 (N_5491,N_3888,N_3536);
nor U5492 (N_5492,N_3621,N_3314);
or U5493 (N_5493,N_3337,N_3785);
nand U5494 (N_5494,N_3819,N_3668);
nor U5495 (N_5495,N_3754,N_3603);
and U5496 (N_5496,N_2825,N_3557);
xor U5497 (N_5497,N_3869,N_2276);
or U5498 (N_5498,N_3990,N_3421);
and U5499 (N_5499,N_2240,N_2636);
nand U5500 (N_5500,N_3383,N_2488);
nand U5501 (N_5501,N_2350,N_2335);
nor U5502 (N_5502,N_2983,N_3071);
nor U5503 (N_5503,N_2140,N_2325);
or U5504 (N_5504,N_3173,N_3053);
nand U5505 (N_5505,N_2104,N_2079);
and U5506 (N_5506,N_3811,N_2203);
nand U5507 (N_5507,N_2891,N_3904);
nor U5508 (N_5508,N_3217,N_2125);
nand U5509 (N_5509,N_2829,N_2709);
or U5510 (N_5510,N_2804,N_3409);
or U5511 (N_5511,N_2438,N_3345);
nor U5512 (N_5512,N_2382,N_3641);
nor U5513 (N_5513,N_3018,N_3972);
xnor U5514 (N_5514,N_3221,N_2671);
nand U5515 (N_5515,N_3997,N_2795);
or U5516 (N_5516,N_3361,N_3173);
and U5517 (N_5517,N_3292,N_3024);
nor U5518 (N_5518,N_3747,N_2778);
nor U5519 (N_5519,N_3598,N_2925);
nor U5520 (N_5520,N_2521,N_2472);
nand U5521 (N_5521,N_2402,N_3247);
nand U5522 (N_5522,N_2971,N_2149);
and U5523 (N_5523,N_2813,N_3389);
nor U5524 (N_5524,N_3854,N_2468);
and U5525 (N_5525,N_3446,N_3519);
nand U5526 (N_5526,N_2971,N_2688);
or U5527 (N_5527,N_3199,N_3628);
or U5528 (N_5528,N_3585,N_3825);
xor U5529 (N_5529,N_2103,N_3927);
or U5530 (N_5530,N_2961,N_2528);
nor U5531 (N_5531,N_2687,N_3064);
nand U5532 (N_5532,N_3999,N_3954);
or U5533 (N_5533,N_2418,N_2827);
or U5534 (N_5534,N_3042,N_2519);
nand U5535 (N_5535,N_3284,N_2960);
nor U5536 (N_5536,N_3508,N_3476);
and U5537 (N_5537,N_2063,N_3233);
nand U5538 (N_5538,N_3067,N_3333);
and U5539 (N_5539,N_3649,N_2386);
or U5540 (N_5540,N_3104,N_3797);
nand U5541 (N_5541,N_2311,N_3853);
or U5542 (N_5542,N_2757,N_3969);
and U5543 (N_5543,N_3824,N_3455);
nor U5544 (N_5544,N_2964,N_2214);
or U5545 (N_5545,N_2208,N_2767);
or U5546 (N_5546,N_3626,N_3759);
and U5547 (N_5547,N_2758,N_3574);
nor U5548 (N_5548,N_3804,N_2515);
or U5549 (N_5549,N_2478,N_3810);
and U5550 (N_5550,N_3663,N_3260);
xor U5551 (N_5551,N_2115,N_3862);
nor U5552 (N_5552,N_2147,N_3112);
nand U5553 (N_5553,N_2746,N_3359);
or U5554 (N_5554,N_3753,N_2429);
nand U5555 (N_5555,N_3942,N_2599);
nor U5556 (N_5556,N_3181,N_3534);
nand U5557 (N_5557,N_3197,N_2978);
nor U5558 (N_5558,N_3500,N_2721);
nor U5559 (N_5559,N_3318,N_3013);
nand U5560 (N_5560,N_3097,N_3186);
and U5561 (N_5561,N_2870,N_2558);
nor U5562 (N_5562,N_3928,N_3085);
or U5563 (N_5563,N_3401,N_3929);
and U5564 (N_5564,N_3282,N_3187);
nand U5565 (N_5565,N_3891,N_2647);
nand U5566 (N_5566,N_2406,N_2439);
and U5567 (N_5567,N_3379,N_3366);
nand U5568 (N_5568,N_3403,N_3022);
or U5569 (N_5569,N_3755,N_3315);
or U5570 (N_5570,N_2744,N_3508);
nor U5571 (N_5571,N_3305,N_3395);
xor U5572 (N_5572,N_2969,N_2550);
and U5573 (N_5573,N_2650,N_2579);
and U5574 (N_5574,N_3990,N_2391);
and U5575 (N_5575,N_2563,N_3871);
or U5576 (N_5576,N_2011,N_2388);
nor U5577 (N_5577,N_2530,N_2382);
nand U5578 (N_5578,N_3331,N_2098);
nand U5579 (N_5579,N_2509,N_3385);
nor U5580 (N_5580,N_3603,N_3972);
nor U5581 (N_5581,N_3466,N_3003);
and U5582 (N_5582,N_3989,N_2360);
and U5583 (N_5583,N_2224,N_3436);
nor U5584 (N_5584,N_3566,N_2617);
and U5585 (N_5585,N_3505,N_2591);
xnor U5586 (N_5586,N_2158,N_2505);
or U5587 (N_5587,N_2967,N_3342);
and U5588 (N_5588,N_2770,N_2488);
and U5589 (N_5589,N_2885,N_3611);
nor U5590 (N_5590,N_2275,N_2731);
and U5591 (N_5591,N_2703,N_2176);
nor U5592 (N_5592,N_3466,N_3055);
and U5593 (N_5593,N_2381,N_3862);
nand U5594 (N_5594,N_3274,N_3470);
nand U5595 (N_5595,N_3788,N_2035);
nand U5596 (N_5596,N_2529,N_2066);
xor U5597 (N_5597,N_3350,N_3119);
nand U5598 (N_5598,N_3928,N_3192);
and U5599 (N_5599,N_2909,N_2512);
nor U5600 (N_5600,N_2680,N_2622);
nand U5601 (N_5601,N_2432,N_3132);
or U5602 (N_5602,N_2666,N_3711);
nor U5603 (N_5603,N_2856,N_2202);
nand U5604 (N_5604,N_2630,N_3808);
nand U5605 (N_5605,N_2985,N_3831);
and U5606 (N_5606,N_3382,N_2499);
or U5607 (N_5607,N_3105,N_3233);
and U5608 (N_5608,N_2545,N_2364);
or U5609 (N_5609,N_3625,N_2726);
and U5610 (N_5610,N_2068,N_2264);
or U5611 (N_5611,N_2622,N_2147);
nand U5612 (N_5612,N_3553,N_2184);
and U5613 (N_5613,N_2016,N_3547);
and U5614 (N_5614,N_2280,N_2954);
nand U5615 (N_5615,N_2458,N_2298);
or U5616 (N_5616,N_2052,N_3911);
nand U5617 (N_5617,N_2407,N_3961);
nand U5618 (N_5618,N_3172,N_3407);
and U5619 (N_5619,N_2197,N_3240);
or U5620 (N_5620,N_2174,N_3392);
nor U5621 (N_5621,N_2676,N_2798);
or U5622 (N_5622,N_2628,N_2466);
nor U5623 (N_5623,N_2691,N_3513);
nor U5624 (N_5624,N_3105,N_2415);
or U5625 (N_5625,N_2014,N_2613);
nor U5626 (N_5626,N_3372,N_3056);
nor U5627 (N_5627,N_3530,N_3451);
nand U5628 (N_5628,N_3186,N_3963);
and U5629 (N_5629,N_2568,N_3291);
nor U5630 (N_5630,N_3175,N_2482);
nand U5631 (N_5631,N_3120,N_3614);
nand U5632 (N_5632,N_3388,N_2188);
nand U5633 (N_5633,N_3071,N_3921);
and U5634 (N_5634,N_2985,N_2935);
and U5635 (N_5635,N_3471,N_3023);
and U5636 (N_5636,N_3840,N_3092);
nor U5637 (N_5637,N_3127,N_3685);
nand U5638 (N_5638,N_2863,N_3381);
nor U5639 (N_5639,N_3697,N_2526);
or U5640 (N_5640,N_2494,N_3183);
or U5641 (N_5641,N_3615,N_3476);
nand U5642 (N_5642,N_2167,N_2047);
nand U5643 (N_5643,N_3945,N_2228);
and U5644 (N_5644,N_2237,N_3053);
nor U5645 (N_5645,N_3784,N_3346);
nor U5646 (N_5646,N_2508,N_2125);
and U5647 (N_5647,N_2209,N_2412);
nor U5648 (N_5648,N_3188,N_3763);
and U5649 (N_5649,N_2452,N_2225);
or U5650 (N_5650,N_3143,N_3601);
or U5651 (N_5651,N_2008,N_3305);
nand U5652 (N_5652,N_2744,N_3613);
and U5653 (N_5653,N_2222,N_2811);
nand U5654 (N_5654,N_2880,N_3050);
or U5655 (N_5655,N_2868,N_2518);
or U5656 (N_5656,N_2102,N_2157);
or U5657 (N_5657,N_2275,N_3972);
nor U5658 (N_5658,N_3069,N_3113);
nand U5659 (N_5659,N_2001,N_3991);
and U5660 (N_5660,N_2584,N_2085);
nor U5661 (N_5661,N_2653,N_2806);
or U5662 (N_5662,N_3004,N_2776);
or U5663 (N_5663,N_2978,N_2061);
nor U5664 (N_5664,N_3119,N_3096);
or U5665 (N_5665,N_2936,N_3299);
and U5666 (N_5666,N_3994,N_3231);
or U5667 (N_5667,N_2223,N_3228);
and U5668 (N_5668,N_3219,N_3661);
nand U5669 (N_5669,N_2190,N_2695);
nand U5670 (N_5670,N_3680,N_2568);
or U5671 (N_5671,N_2645,N_2574);
and U5672 (N_5672,N_2796,N_2427);
and U5673 (N_5673,N_2630,N_2872);
nand U5674 (N_5674,N_3888,N_2625);
and U5675 (N_5675,N_2666,N_3229);
and U5676 (N_5676,N_2650,N_3272);
or U5677 (N_5677,N_2152,N_3413);
or U5678 (N_5678,N_3565,N_3170);
and U5679 (N_5679,N_2550,N_3167);
or U5680 (N_5680,N_3363,N_3464);
nor U5681 (N_5681,N_3053,N_3208);
nor U5682 (N_5682,N_2957,N_2232);
and U5683 (N_5683,N_3236,N_3625);
and U5684 (N_5684,N_2972,N_3632);
and U5685 (N_5685,N_3330,N_2654);
and U5686 (N_5686,N_2866,N_3262);
nor U5687 (N_5687,N_3296,N_2919);
or U5688 (N_5688,N_3334,N_2527);
nand U5689 (N_5689,N_2717,N_3268);
or U5690 (N_5690,N_2807,N_3539);
nand U5691 (N_5691,N_3751,N_3201);
and U5692 (N_5692,N_3526,N_3187);
nor U5693 (N_5693,N_2508,N_3276);
xnor U5694 (N_5694,N_2873,N_3534);
nor U5695 (N_5695,N_2565,N_3137);
and U5696 (N_5696,N_2471,N_3717);
nor U5697 (N_5697,N_2284,N_3612);
or U5698 (N_5698,N_2663,N_2549);
nand U5699 (N_5699,N_3421,N_3296);
and U5700 (N_5700,N_2770,N_2048);
and U5701 (N_5701,N_3056,N_2006);
nor U5702 (N_5702,N_3099,N_2365);
nand U5703 (N_5703,N_2057,N_3613);
and U5704 (N_5704,N_2457,N_3831);
nor U5705 (N_5705,N_3512,N_3113);
xor U5706 (N_5706,N_3689,N_2437);
nor U5707 (N_5707,N_3516,N_2930);
nor U5708 (N_5708,N_2106,N_3691);
and U5709 (N_5709,N_3543,N_3479);
nor U5710 (N_5710,N_2236,N_2815);
nor U5711 (N_5711,N_2863,N_3012);
nor U5712 (N_5712,N_2297,N_3658);
or U5713 (N_5713,N_3252,N_3362);
and U5714 (N_5714,N_2956,N_3034);
or U5715 (N_5715,N_2727,N_2092);
nor U5716 (N_5716,N_2075,N_2451);
nand U5717 (N_5717,N_2052,N_3506);
nor U5718 (N_5718,N_3570,N_3555);
and U5719 (N_5719,N_3846,N_3305);
or U5720 (N_5720,N_2621,N_3614);
or U5721 (N_5721,N_3834,N_2652);
or U5722 (N_5722,N_3247,N_2701);
or U5723 (N_5723,N_3378,N_3849);
nor U5724 (N_5724,N_2309,N_2595);
nand U5725 (N_5725,N_3811,N_2724);
nor U5726 (N_5726,N_2188,N_3304);
or U5727 (N_5727,N_2652,N_3769);
or U5728 (N_5728,N_2019,N_3248);
or U5729 (N_5729,N_3090,N_3201);
or U5730 (N_5730,N_2562,N_2565);
nand U5731 (N_5731,N_3390,N_3717);
nor U5732 (N_5732,N_2002,N_3929);
nand U5733 (N_5733,N_3155,N_2935);
and U5734 (N_5734,N_3487,N_3066);
nand U5735 (N_5735,N_3012,N_3418);
nor U5736 (N_5736,N_3170,N_2400);
nand U5737 (N_5737,N_2528,N_2320);
nand U5738 (N_5738,N_2078,N_3023);
nor U5739 (N_5739,N_3516,N_2854);
and U5740 (N_5740,N_3866,N_3313);
or U5741 (N_5741,N_2651,N_3777);
nand U5742 (N_5742,N_3556,N_3300);
nand U5743 (N_5743,N_3374,N_2556);
nor U5744 (N_5744,N_3360,N_2591);
nor U5745 (N_5745,N_3712,N_3409);
nor U5746 (N_5746,N_2324,N_3297);
nand U5747 (N_5747,N_2148,N_3679);
and U5748 (N_5748,N_3010,N_2004);
nor U5749 (N_5749,N_2546,N_3698);
nand U5750 (N_5750,N_3925,N_2955);
or U5751 (N_5751,N_2126,N_3218);
nor U5752 (N_5752,N_3471,N_2439);
or U5753 (N_5753,N_2357,N_2283);
nand U5754 (N_5754,N_2373,N_3160);
or U5755 (N_5755,N_2213,N_2496);
nand U5756 (N_5756,N_3662,N_2852);
nand U5757 (N_5757,N_3589,N_2622);
nor U5758 (N_5758,N_3910,N_3651);
and U5759 (N_5759,N_2281,N_2292);
or U5760 (N_5760,N_3158,N_3157);
or U5761 (N_5761,N_3902,N_3815);
nor U5762 (N_5762,N_2529,N_2234);
nor U5763 (N_5763,N_2625,N_2188);
nand U5764 (N_5764,N_3284,N_2855);
nor U5765 (N_5765,N_3684,N_3423);
or U5766 (N_5766,N_3194,N_2680);
and U5767 (N_5767,N_2052,N_3949);
and U5768 (N_5768,N_3768,N_3242);
nor U5769 (N_5769,N_2423,N_2021);
nor U5770 (N_5770,N_2424,N_2737);
nor U5771 (N_5771,N_3492,N_2865);
nor U5772 (N_5772,N_2046,N_3829);
or U5773 (N_5773,N_2879,N_3432);
or U5774 (N_5774,N_2487,N_3661);
and U5775 (N_5775,N_2049,N_2555);
or U5776 (N_5776,N_3735,N_3165);
and U5777 (N_5777,N_3765,N_2567);
nand U5778 (N_5778,N_3492,N_3944);
and U5779 (N_5779,N_3230,N_2063);
nor U5780 (N_5780,N_3030,N_2665);
and U5781 (N_5781,N_3141,N_3923);
nor U5782 (N_5782,N_3321,N_3314);
and U5783 (N_5783,N_3812,N_3495);
nor U5784 (N_5784,N_2286,N_2032);
nand U5785 (N_5785,N_2768,N_2304);
or U5786 (N_5786,N_3982,N_2112);
and U5787 (N_5787,N_2314,N_2308);
or U5788 (N_5788,N_3084,N_3158);
nor U5789 (N_5789,N_3750,N_2761);
nand U5790 (N_5790,N_3042,N_2746);
or U5791 (N_5791,N_2112,N_2100);
nand U5792 (N_5792,N_2486,N_3770);
xor U5793 (N_5793,N_3314,N_2841);
and U5794 (N_5794,N_3241,N_2383);
nor U5795 (N_5795,N_3432,N_2547);
nor U5796 (N_5796,N_3028,N_2927);
and U5797 (N_5797,N_3119,N_2456);
nor U5798 (N_5798,N_3809,N_2936);
or U5799 (N_5799,N_3615,N_3366);
and U5800 (N_5800,N_3614,N_3503);
or U5801 (N_5801,N_3944,N_2935);
nor U5802 (N_5802,N_2303,N_2726);
or U5803 (N_5803,N_2531,N_3496);
and U5804 (N_5804,N_3187,N_3574);
nand U5805 (N_5805,N_2480,N_2848);
and U5806 (N_5806,N_3285,N_2902);
or U5807 (N_5807,N_2083,N_2217);
or U5808 (N_5808,N_2371,N_2679);
nor U5809 (N_5809,N_2766,N_2403);
or U5810 (N_5810,N_3191,N_2126);
or U5811 (N_5811,N_3543,N_2770);
nand U5812 (N_5812,N_3988,N_3613);
nand U5813 (N_5813,N_2103,N_3196);
and U5814 (N_5814,N_2070,N_2153);
nand U5815 (N_5815,N_3019,N_3475);
and U5816 (N_5816,N_2888,N_3613);
nand U5817 (N_5817,N_2006,N_2615);
nand U5818 (N_5818,N_2865,N_3485);
or U5819 (N_5819,N_2695,N_3843);
nand U5820 (N_5820,N_3126,N_3166);
nor U5821 (N_5821,N_2486,N_3431);
and U5822 (N_5822,N_3126,N_2655);
nand U5823 (N_5823,N_2923,N_3072);
and U5824 (N_5824,N_3376,N_2753);
and U5825 (N_5825,N_3760,N_3745);
and U5826 (N_5826,N_2602,N_3167);
or U5827 (N_5827,N_3194,N_2982);
or U5828 (N_5828,N_2974,N_3970);
and U5829 (N_5829,N_2890,N_2255);
nand U5830 (N_5830,N_3786,N_2869);
and U5831 (N_5831,N_2220,N_3027);
nor U5832 (N_5832,N_2181,N_3614);
nand U5833 (N_5833,N_2960,N_2308);
nor U5834 (N_5834,N_2124,N_3222);
and U5835 (N_5835,N_3758,N_3387);
or U5836 (N_5836,N_3900,N_3256);
nor U5837 (N_5837,N_2305,N_2276);
or U5838 (N_5838,N_2972,N_2207);
and U5839 (N_5839,N_3110,N_2893);
or U5840 (N_5840,N_2659,N_3296);
nor U5841 (N_5841,N_2708,N_3477);
nand U5842 (N_5842,N_3880,N_2114);
nor U5843 (N_5843,N_2160,N_3766);
and U5844 (N_5844,N_2466,N_2279);
or U5845 (N_5845,N_2812,N_3790);
or U5846 (N_5846,N_3568,N_3604);
nand U5847 (N_5847,N_2562,N_2427);
nand U5848 (N_5848,N_3147,N_2315);
and U5849 (N_5849,N_3342,N_2432);
and U5850 (N_5850,N_2580,N_3773);
nand U5851 (N_5851,N_2502,N_3063);
nand U5852 (N_5852,N_2973,N_3842);
nor U5853 (N_5853,N_2710,N_3105);
nor U5854 (N_5854,N_3750,N_2397);
nand U5855 (N_5855,N_3577,N_2129);
nor U5856 (N_5856,N_2788,N_2572);
nor U5857 (N_5857,N_3142,N_2944);
or U5858 (N_5858,N_2172,N_2847);
nor U5859 (N_5859,N_2906,N_2555);
and U5860 (N_5860,N_3534,N_2795);
nor U5861 (N_5861,N_3880,N_3943);
nand U5862 (N_5862,N_3895,N_3198);
or U5863 (N_5863,N_3740,N_2145);
nand U5864 (N_5864,N_2015,N_2010);
nor U5865 (N_5865,N_2551,N_2089);
nor U5866 (N_5866,N_3637,N_2860);
or U5867 (N_5867,N_3397,N_2478);
or U5868 (N_5868,N_3643,N_2991);
nor U5869 (N_5869,N_3400,N_2920);
xnor U5870 (N_5870,N_3450,N_2832);
or U5871 (N_5871,N_3791,N_3650);
and U5872 (N_5872,N_3584,N_3761);
nor U5873 (N_5873,N_3319,N_3100);
nor U5874 (N_5874,N_2615,N_2201);
nand U5875 (N_5875,N_3960,N_3934);
nand U5876 (N_5876,N_2942,N_2444);
nand U5877 (N_5877,N_3961,N_2151);
and U5878 (N_5878,N_3419,N_2395);
or U5879 (N_5879,N_2485,N_3496);
nor U5880 (N_5880,N_2312,N_3604);
nor U5881 (N_5881,N_2308,N_3776);
and U5882 (N_5882,N_2709,N_2953);
or U5883 (N_5883,N_3148,N_3275);
or U5884 (N_5884,N_2410,N_3442);
nand U5885 (N_5885,N_2718,N_2972);
nand U5886 (N_5886,N_2699,N_3673);
nor U5887 (N_5887,N_2348,N_3400);
nand U5888 (N_5888,N_3958,N_3525);
or U5889 (N_5889,N_3128,N_2419);
and U5890 (N_5890,N_3393,N_2934);
and U5891 (N_5891,N_2837,N_3691);
or U5892 (N_5892,N_3573,N_3925);
nand U5893 (N_5893,N_3650,N_2598);
nand U5894 (N_5894,N_2076,N_3295);
nor U5895 (N_5895,N_2606,N_2116);
nor U5896 (N_5896,N_2561,N_3257);
and U5897 (N_5897,N_2775,N_2405);
or U5898 (N_5898,N_3191,N_3102);
nand U5899 (N_5899,N_3542,N_3895);
and U5900 (N_5900,N_2511,N_2379);
and U5901 (N_5901,N_2628,N_2562);
and U5902 (N_5902,N_2766,N_2823);
and U5903 (N_5903,N_2625,N_3303);
nor U5904 (N_5904,N_2623,N_2326);
or U5905 (N_5905,N_3591,N_3906);
nor U5906 (N_5906,N_2957,N_2836);
and U5907 (N_5907,N_3393,N_2608);
and U5908 (N_5908,N_2453,N_2022);
nor U5909 (N_5909,N_3858,N_2332);
nor U5910 (N_5910,N_3119,N_3709);
and U5911 (N_5911,N_2781,N_3626);
and U5912 (N_5912,N_2199,N_3873);
nand U5913 (N_5913,N_3826,N_2926);
and U5914 (N_5914,N_3510,N_2449);
nor U5915 (N_5915,N_2565,N_3157);
nor U5916 (N_5916,N_3085,N_2642);
and U5917 (N_5917,N_3700,N_3146);
or U5918 (N_5918,N_2167,N_2865);
or U5919 (N_5919,N_2954,N_2988);
or U5920 (N_5920,N_2797,N_3740);
nor U5921 (N_5921,N_2893,N_2783);
nand U5922 (N_5922,N_2586,N_3877);
and U5923 (N_5923,N_2480,N_2528);
or U5924 (N_5924,N_2635,N_3950);
and U5925 (N_5925,N_2613,N_2345);
nand U5926 (N_5926,N_3999,N_3778);
nor U5927 (N_5927,N_3714,N_3797);
nand U5928 (N_5928,N_2069,N_2851);
nand U5929 (N_5929,N_2194,N_2509);
or U5930 (N_5930,N_2487,N_2630);
and U5931 (N_5931,N_2372,N_3125);
or U5932 (N_5932,N_3008,N_2075);
and U5933 (N_5933,N_2287,N_2224);
and U5934 (N_5934,N_2822,N_3615);
nor U5935 (N_5935,N_3069,N_2218);
or U5936 (N_5936,N_3011,N_3776);
and U5937 (N_5937,N_3307,N_3811);
or U5938 (N_5938,N_3039,N_2679);
and U5939 (N_5939,N_3443,N_3917);
or U5940 (N_5940,N_3581,N_2719);
nand U5941 (N_5941,N_3966,N_2470);
and U5942 (N_5942,N_2959,N_3972);
nor U5943 (N_5943,N_3196,N_3962);
nor U5944 (N_5944,N_2257,N_2778);
or U5945 (N_5945,N_2537,N_3501);
or U5946 (N_5946,N_3003,N_2724);
nand U5947 (N_5947,N_2418,N_2234);
or U5948 (N_5948,N_3501,N_2092);
or U5949 (N_5949,N_2911,N_3338);
nor U5950 (N_5950,N_2431,N_2895);
or U5951 (N_5951,N_3656,N_3073);
nand U5952 (N_5952,N_3458,N_3782);
or U5953 (N_5953,N_3662,N_2188);
or U5954 (N_5954,N_3636,N_2861);
nand U5955 (N_5955,N_2514,N_3909);
nor U5956 (N_5956,N_2258,N_2726);
nand U5957 (N_5957,N_3148,N_3437);
nor U5958 (N_5958,N_2798,N_2510);
or U5959 (N_5959,N_3021,N_2165);
or U5960 (N_5960,N_2611,N_3748);
or U5961 (N_5961,N_2830,N_3303);
or U5962 (N_5962,N_2174,N_3529);
nor U5963 (N_5963,N_2949,N_2537);
nand U5964 (N_5964,N_2615,N_3592);
and U5965 (N_5965,N_2631,N_2038);
nand U5966 (N_5966,N_2267,N_2232);
and U5967 (N_5967,N_3258,N_3577);
and U5968 (N_5968,N_3505,N_3220);
nand U5969 (N_5969,N_3196,N_2747);
nor U5970 (N_5970,N_2378,N_2714);
or U5971 (N_5971,N_3475,N_2769);
nor U5972 (N_5972,N_2417,N_2474);
nand U5973 (N_5973,N_3762,N_3349);
nor U5974 (N_5974,N_2748,N_2526);
nand U5975 (N_5975,N_2545,N_2336);
nor U5976 (N_5976,N_2887,N_3614);
or U5977 (N_5977,N_3163,N_2797);
nor U5978 (N_5978,N_2600,N_2620);
nor U5979 (N_5979,N_2560,N_3068);
nand U5980 (N_5980,N_2477,N_2713);
nor U5981 (N_5981,N_2990,N_3566);
nand U5982 (N_5982,N_3822,N_2372);
nand U5983 (N_5983,N_3310,N_3944);
nor U5984 (N_5984,N_2747,N_3015);
or U5985 (N_5985,N_3538,N_3272);
and U5986 (N_5986,N_3137,N_3657);
and U5987 (N_5987,N_2840,N_2580);
nor U5988 (N_5988,N_3069,N_3660);
nor U5989 (N_5989,N_2252,N_2980);
or U5990 (N_5990,N_3868,N_3699);
nand U5991 (N_5991,N_2112,N_3160);
and U5992 (N_5992,N_2217,N_3599);
or U5993 (N_5993,N_2497,N_2378);
nor U5994 (N_5994,N_2122,N_3763);
and U5995 (N_5995,N_3023,N_3143);
nor U5996 (N_5996,N_2067,N_2571);
or U5997 (N_5997,N_3161,N_2926);
nand U5998 (N_5998,N_3747,N_2973);
nand U5999 (N_5999,N_3905,N_2248);
and U6000 (N_6000,N_4075,N_5634);
and U6001 (N_6001,N_4809,N_4685);
nand U6002 (N_6002,N_5685,N_4625);
or U6003 (N_6003,N_5477,N_4042);
or U6004 (N_6004,N_5647,N_5441);
and U6005 (N_6005,N_5842,N_4238);
nor U6006 (N_6006,N_4921,N_4356);
or U6007 (N_6007,N_4343,N_4613);
nand U6008 (N_6008,N_5101,N_5870);
and U6009 (N_6009,N_5872,N_4846);
nand U6010 (N_6010,N_4569,N_5233);
nand U6011 (N_6011,N_4676,N_4265);
and U6012 (N_6012,N_4035,N_5817);
or U6013 (N_6013,N_4241,N_4568);
and U6014 (N_6014,N_4318,N_5253);
and U6015 (N_6015,N_5025,N_4611);
and U6016 (N_6016,N_5498,N_5232);
nor U6017 (N_6017,N_5262,N_5071);
nand U6018 (N_6018,N_4380,N_5329);
or U6019 (N_6019,N_5367,N_4235);
nand U6020 (N_6020,N_4192,N_5493);
and U6021 (N_6021,N_5650,N_4558);
nand U6022 (N_6022,N_5887,N_4375);
or U6023 (N_6023,N_4572,N_4877);
and U6024 (N_6024,N_5421,N_4421);
and U6025 (N_6025,N_5463,N_4755);
nor U6026 (N_6026,N_4324,N_5768);
or U6027 (N_6027,N_4830,N_5107);
or U6028 (N_6028,N_4453,N_5403);
nor U6029 (N_6029,N_5045,N_5763);
nor U6030 (N_6030,N_4562,N_4945);
nor U6031 (N_6031,N_5955,N_5093);
nor U6032 (N_6032,N_5428,N_5147);
and U6033 (N_6033,N_5626,N_5427);
nand U6034 (N_6034,N_4418,N_5109);
or U6035 (N_6035,N_5316,N_4423);
and U6036 (N_6036,N_5694,N_5234);
and U6037 (N_6037,N_4458,N_4696);
and U6038 (N_6038,N_5519,N_4160);
nand U6039 (N_6039,N_5119,N_5240);
or U6040 (N_6040,N_4591,N_5724);
nor U6041 (N_6041,N_4072,N_4826);
or U6042 (N_6042,N_4068,N_4483);
nand U6043 (N_6043,N_5116,N_5079);
nor U6044 (N_6044,N_5016,N_4783);
nor U6045 (N_6045,N_5348,N_5118);
and U6046 (N_6046,N_4105,N_5690);
nor U6047 (N_6047,N_5141,N_4911);
nor U6048 (N_6048,N_4659,N_4110);
nand U6049 (N_6049,N_5143,N_5127);
or U6050 (N_6050,N_5556,N_4994);
and U6051 (N_6051,N_4024,N_5569);
and U6052 (N_6052,N_5576,N_4440);
or U6053 (N_6053,N_4976,N_4387);
nor U6054 (N_6054,N_5604,N_4504);
nand U6055 (N_6055,N_4530,N_5973);
nor U6056 (N_6056,N_4066,N_5005);
nand U6057 (N_6057,N_5711,N_4347);
and U6058 (N_6058,N_5136,N_5571);
nor U6059 (N_6059,N_5040,N_4478);
nor U6060 (N_6060,N_5757,N_4654);
nor U6061 (N_6061,N_5582,N_5713);
nor U6062 (N_6062,N_5976,N_5611);
nor U6063 (N_6063,N_4801,N_5165);
nor U6064 (N_6064,N_5824,N_5283);
or U6065 (N_6065,N_4379,N_5264);
nand U6066 (N_6066,N_4284,N_5776);
and U6067 (N_6067,N_4632,N_4106);
and U6068 (N_6068,N_4782,N_4793);
nand U6069 (N_6069,N_4836,N_5935);
and U6070 (N_6070,N_4847,N_5511);
nor U6071 (N_6071,N_4660,N_4109);
nor U6072 (N_6072,N_4372,N_4353);
or U6073 (N_6073,N_5873,N_5307);
or U6074 (N_6074,N_4884,N_5178);
or U6075 (N_6075,N_4381,N_5564);
nand U6076 (N_6076,N_4193,N_4986);
nand U6077 (N_6077,N_5875,N_5432);
nor U6078 (N_6078,N_4533,N_4792);
and U6079 (N_6079,N_4052,N_4463);
nand U6080 (N_6080,N_5628,N_4887);
nand U6081 (N_6081,N_4842,N_4780);
nand U6082 (N_6082,N_4998,N_4816);
nor U6083 (N_6083,N_5522,N_4184);
nand U6084 (N_6084,N_5619,N_5394);
and U6085 (N_6085,N_5720,N_4722);
and U6086 (N_6086,N_4490,N_4694);
nand U6087 (N_6087,N_4438,N_5054);
nand U6088 (N_6088,N_4889,N_5066);
nor U6089 (N_6089,N_4634,N_5204);
and U6090 (N_6090,N_5485,N_5134);
or U6091 (N_6091,N_4690,N_5954);
or U6092 (N_6092,N_5814,N_4876);
nand U6093 (N_6093,N_4899,N_4173);
or U6094 (N_6094,N_5645,N_4371);
and U6095 (N_6095,N_4195,N_5219);
and U6096 (N_6096,N_5524,N_5745);
and U6097 (N_6097,N_4506,N_5530);
nor U6098 (N_6098,N_4981,N_4328);
and U6099 (N_6099,N_4408,N_4701);
nor U6100 (N_6100,N_5704,N_5220);
nand U6101 (N_6101,N_5506,N_5431);
and U6102 (N_6102,N_5466,N_5339);
nor U6103 (N_6103,N_4599,N_4181);
nand U6104 (N_6104,N_4788,N_5507);
or U6105 (N_6105,N_4773,N_5950);
nand U6106 (N_6106,N_5004,N_4271);
nand U6107 (N_6107,N_5526,N_5105);
and U6108 (N_6108,N_4187,N_5275);
nand U6109 (N_6109,N_5797,N_5122);
and U6110 (N_6110,N_4206,N_5207);
and U6111 (N_6111,N_5010,N_4635);
nor U6112 (N_6112,N_5154,N_4255);
and U6113 (N_6113,N_4957,N_4010);
and U6114 (N_6114,N_4096,N_4363);
nor U6115 (N_6115,N_4071,N_4406);
nor U6116 (N_6116,N_5562,N_5175);
nand U6117 (N_6117,N_5000,N_5881);
nor U6118 (N_6118,N_5717,N_5335);
and U6119 (N_6119,N_4711,N_5691);
nand U6120 (N_6120,N_5110,N_5245);
or U6121 (N_6121,N_4224,N_5050);
nand U6122 (N_6122,N_5958,N_4014);
or U6123 (N_6123,N_5680,N_5971);
nor U6124 (N_6124,N_4620,N_5282);
nor U6125 (N_6125,N_4333,N_5419);
and U6126 (N_6126,N_4201,N_5953);
and U6127 (N_6127,N_5087,N_4200);
and U6128 (N_6128,N_4564,N_5822);
nand U6129 (N_6129,N_5589,N_5674);
nand U6130 (N_6130,N_4776,N_5867);
or U6131 (N_6131,N_4751,N_5877);
or U6132 (N_6132,N_4939,N_5957);
nor U6133 (N_6133,N_4172,N_4213);
and U6134 (N_6134,N_4189,N_4481);
or U6135 (N_6135,N_5227,N_5221);
nor U6136 (N_6136,N_4435,N_5649);
nor U6137 (N_6137,N_5820,N_4983);
nand U6138 (N_6138,N_4529,N_4401);
and U6139 (N_6139,N_5601,N_4606);
nand U6140 (N_6140,N_4285,N_5012);
nand U6141 (N_6141,N_4474,N_4411);
and U6142 (N_6142,N_5360,N_4516);
or U6143 (N_6143,N_5613,N_4320);
nor U6144 (N_6144,N_5492,N_4051);
and U6145 (N_6145,N_5575,N_5076);
nand U6146 (N_6146,N_5144,N_5780);
or U6147 (N_6147,N_4405,N_4101);
and U6148 (N_6148,N_4441,N_4044);
nor U6149 (N_6149,N_4592,N_5978);
nor U6150 (N_6150,N_5860,N_5151);
nand U6151 (N_6151,N_4825,N_4774);
nor U6152 (N_6152,N_5969,N_5859);
and U6153 (N_6153,N_4342,N_4236);
nand U6154 (N_6154,N_5377,N_4869);
or U6155 (N_6155,N_5807,N_5944);
nor U6156 (N_6156,N_5901,N_4671);
and U6157 (N_6157,N_4571,N_5566);
and U6158 (N_6158,N_5907,N_4159);
xor U6159 (N_6159,N_5987,N_5533);
nand U6160 (N_6160,N_5451,N_4389);
and U6161 (N_6161,N_5783,N_5523);
nor U6162 (N_6162,N_4539,N_5250);
and U6163 (N_6163,N_5811,N_5315);
nor U6164 (N_6164,N_4429,N_5084);
nor U6165 (N_6165,N_4289,N_5060);
and U6166 (N_6166,N_5515,N_4849);
and U6167 (N_6167,N_4698,N_4305);
nor U6168 (N_6168,N_5149,N_4581);
nand U6169 (N_6169,N_5750,N_4848);
and U6170 (N_6170,N_5454,N_4057);
nand U6171 (N_6171,N_4146,N_4731);
or U6172 (N_6172,N_5209,N_5413);
and U6173 (N_6173,N_4442,N_5180);
and U6174 (N_6174,N_5903,N_5673);
nor U6175 (N_6175,N_4856,N_5073);
nor U6176 (N_6176,N_5146,N_4756);
or U6177 (N_6177,N_5892,N_5248);
or U6178 (N_6178,N_4009,N_5319);
and U6179 (N_6179,N_4242,N_5839);
nor U6180 (N_6180,N_5011,N_5679);
or U6181 (N_6181,N_4695,N_4872);
nand U6182 (N_6182,N_4777,N_4416);
or U6183 (N_6183,N_4894,N_5462);
or U6184 (N_6184,N_4575,N_4230);
nand U6185 (N_6185,N_5979,N_4934);
nand U6186 (N_6186,N_4732,N_5900);
or U6187 (N_6187,N_4963,N_5682);
or U6188 (N_6188,N_4439,N_5085);
and U6189 (N_6189,N_5023,N_4153);
nor U6190 (N_6190,N_5921,N_5376);
and U6191 (N_6191,N_4706,N_5932);
and U6192 (N_6192,N_5026,N_4541);
and U6193 (N_6193,N_5627,N_4639);
or U6194 (N_6194,N_4133,N_4913);
nor U6195 (N_6195,N_4393,N_5622);
xor U6196 (N_6196,N_5125,N_4013);
nand U6197 (N_6197,N_4352,N_5959);
or U6198 (N_6198,N_5746,N_5672);
nand U6199 (N_6199,N_4480,N_4145);
or U6200 (N_6200,N_4107,N_4080);
or U6201 (N_6201,N_5764,N_5265);
or U6202 (N_6202,N_5064,N_4443);
nor U6203 (N_6203,N_4031,N_5847);
nor U6204 (N_6204,N_4345,N_4287);
nor U6205 (N_6205,N_4740,N_4518);
nor U6206 (N_6206,N_5001,N_4707);
nor U6207 (N_6207,N_4337,N_4741);
nor U6208 (N_6208,N_4126,N_5553);
nand U6209 (N_6209,N_5112,N_4309);
nor U6210 (N_6210,N_4736,N_4355);
or U6211 (N_6211,N_4155,N_4244);
nand U6212 (N_6212,N_4798,N_5631);
or U6213 (N_6213,N_4467,N_5276);
nand U6214 (N_6214,N_5198,N_4447);
nor U6215 (N_6215,N_4007,N_4972);
nand U6216 (N_6216,N_5467,N_5997);
or U6217 (N_6217,N_5366,N_5405);
nor U6218 (N_6218,N_4662,N_5081);
and U6219 (N_6219,N_5237,N_4770);
and U6220 (N_6220,N_4665,N_5555);
nor U6221 (N_6221,N_4188,N_4391);
and U6222 (N_6222,N_5755,N_5879);
or U6223 (N_6223,N_5929,N_4338);
nor U6224 (N_6224,N_4114,N_5810);
or U6225 (N_6225,N_4283,N_4938);
xnor U6226 (N_6226,N_4603,N_4962);
nand U6227 (N_6227,N_5398,N_5430);
nor U6228 (N_6228,N_5261,N_5215);
nand U6229 (N_6229,N_4484,N_5057);
nand U6230 (N_6230,N_5835,N_4807);
nor U6231 (N_6231,N_5106,N_4502);
or U6232 (N_6232,N_5707,N_5718);
nand U6233 (N_6233,N_5470,N_5925);
nor U6234 (N_6234,N_5365,N_4473);
nor U6235 (N_6235,N_5429,N_4931);
nor U6236 (N_6236,N_5472,N_5490);
nor U6237 (N_6237,N_5597,N_4609);
nor U6238 (N_6238,N_4087,N_5020);
nand U6239 (N_6239,N_5699,N_5323);
nor U6240 (N_6240,N_5346,N_5998);
or U6241 (N_6241,N_5074,N_5314);
or U6242 (N_6242,N_5374,N_5696);
or U6243 (N_6243,N_4871,N_5423);
nand U6244 (N_6244,N_4813,N_5471);
and U6245 (N_6245,N_4012,N_4944);
or U6246 (N_6246,N_5934,N_4745);
or U6247 (N_6247,N_4070,N_5868);
nand U6248 (N_6248,N_5637,N_4692);
nand U6249 (N_6249,N_4078,N_5591);
nor U6250 (N_6250,N_4651,N_4705);
nand U6251 (N_6251,N_5623,N_5244);
nand U6252 (N_6252,N_4055,N_4177);
and U6253 (N_6253,N_5804,N_4319);
nor U6254 (N_6254,N_4488,N_5318);
and U6255 (N_6255,N_5858,N_4648);
nand U6256 (N_6256,N_5225,N_5167);
or U6257 (N_6257,N_4434,N_4163);
nand U6258 (N_6258,N_5529,N_4302);
nand U6259 (N_6259,N_5362,N_5547);
and U6260 (N_6260,N_4689,N_4403);
nand U6261 (N_6261,N_5563,N_5205);
and U6262 (N_6262,N_4536,N_4626);
nand U6263 (N_6263,N_4002,N_5516);
and U6264 (N_6264,N_5743,N_5864);
and U6265 (N_6265,N_4143,N_5038);
and U6266 (N_6266,N_4112,N_5211);
and U6267 (N_6267,N_4041,N_5422);
or U6268 (N_6268,N_4935,N_5482);
and U6269 (N_6269,N_5538,N_4566);
nand U6270 (N_6270,N_5551,N_4225);
or U6271 (N_6271,N_4125,N_4322);
nor U6272 (N_6272,N_4821,N_5917);
nor U6273 (N_6273,N_5322,N_5852);
nor U6274 (N_6274,N_4532,N_4420);
nor U6275 (N_6275,N_4679,N_5310);
nor U6276 (N_6276,N_4446,N_5036);
nand U6277 (N_6277,N_5407,N_4641);
nor U6278 (N_6278,N_4321,N_5171);
nor U6279 (N_6279,N_5606,N_4062);
nand U6280 (N_6280,N_5665,N_4968);
and U6281 (N_6281,N_4053,N_5426);
and U6282 (N_6282,N_5210,N_4489);
or U6283 (N_6283,N_4185,N_4384);
nor U6284 (N_6284,N_5689,N_4924);
nor U6285 (N_6285,N_4191,N_4797);
and U6286 (N_6286,N_5657,N_4227);
nand U6287 (N_6287,N_5368,N_5799);
nor U6288 (N_6288,N_5381,N_4901);
and U6289 (N_6289,N_5208,N_4396);
or U6290 (N_6290,N_5196,N_4307);
nor U6291 (N_6291,N_4892,N_4282);
nand U6292 (N_6292,N_5200,N_4266);
and U6293 (N_6293,N_4514,N_5988);
or U6294 (N_6294,N_5187,N_4079);
nor U6295 (N_6295,N_4221,N_4469);
nor U6296 (N_6296,N_4708,N_4958);
nand U6297 (N_6297,N_4388,N_5939);
nor U6298 (N_6298,N_4428,N_4147);
or U6299 (N_6299,N_5919,N_5782);
and U6300 (N_6300,N_4169,N_4234);
nand U6301 (N_6301,N_5061,N_5383);
and U6302 (N_6302,N_4590,N_5840);
nand U6303 (N_6303,N_4269,N_5653);
and U6304 (N_6304,N_4702,N_5252);
or U6305 (N_6305,N_4883,N_5385);
nor U6306 (N_6306,N_5294,N_4315);
nand U6307 (N_6307,N_4157,N_5108);
nand U6308 (N_6308,N_4025,N_5642);
nand U6309 (N_6309,N_4373,N_4930);
nand U6310 (N_6310,N_5734,N_5308);
nand U6311 (N_6311,N_4312,N_5838);
or U6312 (N_6312,N_5951,N_4989);
or U6313 (N_6313,N_5813,N_4802);
nand U6314 (N_6314,N_5758,N_5766);
nand U6315 (N_6315,N_4865,N_5521);
and U6316 (N_6316,N_4805,N_4205);
nor U6317 (N_6317,N_5296,N_5725);
nand U6318 (N_6318,N_5334,N_5386);
or U6319 (N_6319,N_4559,N_5594);
nand U6320 (N_6320,N_4997,N_4210);
or U6321 (N_6321,N_5042,N_5798);
and U6322 (N_6322,N_4404,N_5818);
xnor U6323 (N_6323,N_5800,N_5793);
or U6324 (N_6324,N_4982,N_4531);
or U6325 (N_6325,N_5371,N_4067);
nand U6326 (N_6326,N_5188,N_5819);
nor U6327 (N_6327,N_5305,N_4601);
and U6328 (N_6328,N_5358,N_5448);
nand U6329 (N_6329,N_5595,N_5588);
or U6330 (N_6330,N_4619,N_4605);
nor U6331 (N_6331,N_4602,N_4941);
and U6332 (N_6332,N_5052,N_4642);
nor U6333 (N_6333,N_5779,N_5787);
or U6334 (N_6334,N_5640,N_4973);
nor U6335 (N_6335,N_5695,N_4064);
and U6336 (N_6336,N_5982,N_5920);
nor U6337 (N_6337,N_5655,N_5177);
and U6338 (N_6338,N_4710,N_5285);
nor U6339 (N_6339,N_4135,N_4553);
or U6340 (N_6340,N_4425,N_4882);
nor U6341 (N_6341,N_5910,N_5028);
nor U6342 (N_6342,N_4525,N_4008);
and U6343 (N_6343,N_4392,N_5573);
and U6344 (N_6344,N_5128,N_5222);
nand U6345 (N_6345,N_5508,N_5436);
nor U6346 (N_6346,N_4546,N_4190);
or U6347 (N_6347,N_4340,N_4419);
and U6348 (N_6348,N_5461,N_4256);
or U6349 (N_6349,N_5558,N_4699);
or U6350 (N_6350,N_4127,N_5351);
nand U6351 (N_6351,N_5384,N_5948);
nor U6352 (N_6352,N_4000,N_5053);
and U6353 (N_6353,N_5051,N_4231);
and U6354 (N_6354,N_4618,N_5778);
nor U6355 (N_6355,N_4296,N_5224);
nand U6356 (N_6356,N_4890,N_4688);
or U6357 (N_6357,N_4011,N_4682);
and U6358 (N_6358,N_5754,N_4917);
nor U6359 (N_6359,N_5644,N_5828);
or U6360 (N_6360,N_5639,N_4974);
and U6361 (N_6361,N_4175,N_5473);
or U6362 (N_6362,N_4542,N_4327);
and U6363 (N_6363,N_5259,N_5476);
or U6364 (N_6364,N_5671,N_5534);
nand U6365 (N_6365,N_5048,N_5115);
and U6366 (N_6366,N_4663,N_5455);
or U6367 (N_6367,N_5829,N_5843);
nor U6368 (N_6368,N_4902,N_4034);
or U6369 (N_6369,N_5702,N_4017);
nand U6370 (N_6370,N_5017,N_4757);
and U6371 (N_6371,N_4383,N_4593);
or U6372 (N_6372,N_5034,N_5130);
nand U6373 (N_6373,N_5239,N_4527);
nor U6374 (N_6374,N_5014,N_4158);
or U6375 (N_6375,N_5412,N_5044);
nand U6376 (N_6376,N_4300,N_5340);
or U6377 (N_6377,N_4713,N_5914);
nand U6378 (N_6378,N_4932,N_5229);
and U6379 (N_6379,N_4223,N_5388);
nor U6380 (N_6380,N_5796,N_4850);
nand U6381 (N_6381,N_5856,N_4295);
and U6382 (N_6382,N_5369,N_4775);
or U6383 (N_6383,N_5625,N_5520);
nand U6384 (N_6384,N_5343,N_4717);
nor U6385 (N_6385,N_4259,N_5893);
or U6386 (N_6386,N_4376,N_4402);
and U6387 (N_6387,N_5181,N_5037);
or U6388 (N_6388,N_5401,N_5667);
nand U6389 (N_6389,N_4116,N_4927);
or U6390 (N_6390,N_5578,N_5077);
nand U6391 (N_6391,N_5603,N_4839);
or U6392 (N_6392,N_5321,N_5945);
nand U6393 (N_6393,N_5111,N_5503);
nor U6394 (N_6394,N_4073,N_5007);
nand U6395 (N_6395,N_4113,N_5280);
and U6396 (N_6396,N_5882,N_4170);
nor U6397 (N_6397,N_4728,N_4604);
or U6398 (N_6398,N_5697,N_5458);
nand U6399 (N_6399,N_4407,N_5936);
nor U6400 (N_6400,N_5056,N_4270);
nand U6401 (N_6401,N_5156,N_4645);
and U6402 (N_6402,N_5687,N_4646);
nor U6403 (N_6403,N_5035,N_4712);
nor U6404 (N_6404,N_5311,N_5668);
or U6405 (N_6405,N_5616,N_5480);
or U6406 (N_6406,N_5841,N_4834);
nor U6407 (N_6407,N_4936,N_5654);
nand U6408 (N_6408,N_5542,N_5816);
and U6409 (N_6409,N_4900,N_4655);
nand U6410 (N_6410,N_4908,N_5583);
or U6411 (N_6411,N_5646,N_4048);
and U6412 (N_6412,N_4033,N_5356);
or U6413 (N_6413,N_5131,N_5536);
and U6414 (N_6414,N_4432,N_5297);
and U6415 (N_6415,N_5703,N_4140);
nand U6416 (N_6416,N_5347,N_5943);
nor U6417 (N_6417,N_4864,N_5228);
nand U6418 (N_6418,N_5303,N_5173);
nand U6419 (N_6419,N_4971,N_4537);
nor U6420 (N_6420,N_5324,N_5692);
nand U6421 (N_6421,N_4505,N_4137);
and U6422 (N_6422,N_4669,N_4043);
or U6423 (N_6423,N_4716,N_4683);
or U6424 (N_6424,N_5565,N_5965);
and U6425 (N_6425,N_5541,N_5008);
nor U6426 (N_6426,N_5152,N_4584);
or U6427 (N_6427,N_4812,N_5747);
and U6428 (N_6428,N_5592,N_4246);
and U6429 (N_6429,N_5981,N_5281);
and U6430 (N_6430,N_5391,N_5357);
and U6431 (N_6431,N_4059,N_5527);
or U6432 (N_6432,N_5518,N_5584);
or U6433 (N_6433,N_5086,N_4228);
nand U6434 (N_6434,N_5486,N_5930);
nor U6435 (N_6435,N_5664,N_4720);
and U6436 (N_6436,N_5602,N_5065);
nand U6437 (N_6437,N_4909,N_4560);
or U6438 (N_6438,N_4885,N_4739);
or U6439 (N_6439,N_4250,N_4186);
nand U6440 (N_6440,N_5306,N_4528);
nand U6441 (N_6441,N_5532,N_5390);
nand U6442 (N_6442,N_4721,N_5719);
nor U6443 (N_6443,N_4583,N_5202);
and U6444 (N_6444,N_4766,N_4464);
nand U6445 (N_6445,N_5009,N_5496);
nor U6446 (N_6446,N_4161,N_5710);
and U6447 (N_6447,N_4975,N_5621);
nor U6448 (N_6448,N_4207,N_4422);
and U6449 (N_6449,N_5815,N_5777);
and U6450 (N_6450,N_4999,N_4022);
nand U6451 (N_6451,N_4629,N_4152);
nor U6452 (N_6452,N_5162,N_4964);
nor U6453 (N_6453,N_5505,N_5886);
or U6454 (N_6454,N_5600,N_4395);
or U6455 (N_6455,N_4519,N_4748);
or U6456 (N_6456,N_5803,N_5918);
nor U6457 (N_6457,N_5442,N_4273);
nor U6458 (N_6458,N_4354,N_5133);
or U6459 (N_6459,N_4961,N_5206);
and U6460 (N_6460,N_4517,N_5773);
nand U6461 (N_6461,N_4074,N_5715);
nand U6462 (N_6462,N_5022,N_4500);
or U6463 (N_6463,N_5299,N_5142);
nor U6464 (N_6464,N_4491,N_5537);
nor U6465 (N_6465,N_4677,N_4299);
nand U6466 (N_6466,N_4578,N_5185);
and U6467 (N_6467,N_4959,N_4183);
nor U6468 (N_6468,N_5608,N_4102);
nor U6469 (N_6469,N_4510,N_4507);
nand U6470 (N_6470,N_4681,N_5420);
nor U6471 (N_6471,N_5577,N_4746);
nand U6472 (N_6472,N_5795,N_5434);
or U6473 (N_6473,N_5402,N_4955);
nor U6474 (N_6474,N_5666,N_5182);
and U6475 (N_6475,N_4279,N_4753);
and U6476 (N_6476,N_4637,N_4522);
nand U6477 (N_6477,N_5304,N_4151);
nand U6478 (N_6478,N_4752,N_4866);
nor U6479 (N_6479,N_5909,N_4245);
and U6480 (N_6480,N_4647,N_4498);
nor U6481 (N_6481,N_5585,N_5406);
or U6482 (N_6482,N_4579,N_5145);
nand U6483 (N_6483,N_4946,N_4278);
or U6484 (N_6484,N_4167,N_5610);
and U6485 (N_6485,N_5433,N_5861);
and U6486 (N_6486,N_5096,N_5191);
or U6487 (N_6487,N_5094,N_5906);
and U6488 (N_6488,N_5579,N_4311);
nor U6489 (N_6489,N_5922,N_4949);
nand U6490 (N_6490,N_4288,N_4627);
nand U6491 (N_6491,N_5453,N_4535);
nand U6492 (N_6492,N_4859,N_4208);
and U6493 (N_6493,N_5693,N_5236);
or U6494 (N_6494,N_5298,N_5629);
nand U6495 (N_6495,N_5067,N_5410);
nor U6496 (N_6496,N_4803,N_4215);
or U6497 (N_6497,N_4680,N_5716);
and U6498 (N_6498,N_5956,N_4703);
and U6499 (N_6499,N_5139,N_5006);
nand U6500 (N_6500,N_5288,N_5761);
nand U6501 (N_6501,N_5823,N_5212);
nand U6502 (N_6502,N_4118,N_4764);
nand U6503 (N_6503,N_5509,N_4824);
xor U6504 (N_6504,N_4082,N_4589);
xnor U6505 (N_6505,N_4557,N_4880);
and U6506 (N_6506,N_4436,N_4386);
or U6507 (N_6507,N_4100,N_5003);
nor U6508 (N_6508,N_4240,N_5338);
nand U6509 (N_6509,N_4750,N_4670);
nor U6510 (N_6510,N_5418,N_4367);
xnor U6511 (N_6511,N_4838,N_5947);
and U6512 (N_6512,N_4050,N_5784);
nand U6513 (N_6513,N_4622,N_4948);
or U6514 (N_6514,N_5726,N_5554);
and U6515 (N_6515,N_4493,N_4444);
and U6516 (N_6516,N_5337,N_4487);
nor U6517 (N_6517,N_4769,N_5735);
and U6518 (N_6518,N_4687,N_5242);
or U6519 (N_6519,N_4268,N_5706);
nand U6520 (N_6520,N_5382,N_5850);
and U6521 (N_6521,N_5652,N_4840);
nor U6522 (N_6522,N_4744,N_4896);
or U6523 (N_6523,N_4099,N_5605);
or U6524 (N_6524,N_5379,N_5489);
or U6525 (N_6525,N_4657,N_4897);
and U6526 (N_6526,N_5733,N_4226);
and U6527 (N_6527,N_5157,N_5063);
and U6528 (N_6528,N_4357,N_5874);
and U6529 (N_6529,N_4538,N_5812);
nor U6530 (N_6530,N_5174,N_5435);
nor U6531 (N_6531,N_5465,N_4123);
and U6532 (N_6532,N_4212,N_4551);
or U6533 (N_6533,N_5082,N_5928);
nand U6534 (N_6534,N_4217,N_4729);
nand U6535 (N_6535,N_4374,N_4003);
and U6536 (N_6536,N_5251,N_5124);
or U6537 (N_6537,N_4704,N_4115);
and U6538 (N_6538,N_4454,N_4323);
nor U6539 (N_6539,N_4977,N_4233);
nor U6540 (N_6540,N_5883,N_5373);
or U6541 (N_6541,N_5705,N_4329);
nand U6542 (N_6542,N_4179,N_4359);
nand U6543 (N_6543,N_5479,N_4313);
nand U6544 (N_6544,N_5751,N_4810);
nand U6545 (N_6545,N_5968,N_4800);
nand U6546 (N_6546,N_4451,N_4984);
and U6547 (N_6547,N_5395,N_5326);
xnor U6548 (N_6548,N_4719,N_4026);
nor U6549 (N_6549,N_4365,N_5164);
nand U6550 (N_6550,N_4199,N_4351);
nand U6551 (N_6551,N_5150,N_4806);
nor U6552 (N_6552,N_5794,N_5730);
nor U6553 (N_6553,N_4565,N_4979);
and U6554 (N_6554,N_4263,N_5552);
nor U6555 (N_6555,N_4122,N_4804);
nor U6556 (N_6556,N_4501,N_4653);
and U6557 (N_6557,N_4445,N_4308);
xor U6558 (N_6558,N_4317,N_5996);
nor U6559 (N_6559,N_5273,N_4926);
and U6560 (N_6560,N_5443,N_5638);
nor U6561 (N_6561,N_5805,N_4743);
nor U6562 (N_6562,N_5927,N_5549);
and U6563 (N_6563,N_5752,N_5895);
nand U6564 (N_6564,N_4820,N_5539);
nor U6565 (N_6565,N_4738,N_4861);
nand U6566 (N_6566,N_5739,N_4814);
and U6567 (N_6567,N_4249,N_5574);
and U6568 (N_6568,N_4397,N_4808);
and U6569 (N_6569,N_4142,N_4316);
nand U6570 (N_6570,N_4771,N_5825);
nand U6571 (N_6571,N_5938,N_5972);
nor U6572 (N_6572,N_4652,N_5027);
and U6573 (N_6573,N_4928,N_5059);
nand U6574 (N_6574,N_4960,N_5137);
nand U6575 (N_6575,N_5762,N_5409);
nor U6576 (N_6576,N_4216,N_5030);
nand U6577 (N_6577,N_4426,N_5771);
and U6578 (N_6578,N_4130,N_4919);
or U6579 (N_6579,N_4991,N_5159);
nor U6580 (N_6580,N_5809,N_5456);
and U6581 (N_6581,N_5658,N_4497);
nand U6582 (N_6582,N_5727,N_4253);
nand U6583 (N_6583,N_5355,N_5214);
or U6584 (N_6584,N_4947,N_5514);
and U6585 (N_6585,N_4929,N_5216);
nand U6586 (N_6586,N_5363,N_5651);
and U6587 (N_6587,N_4638,N_5912);
nor U6588 (N_6588,N_4156,N_4725);
nand U6589 (N_6589,N_4254,N_5681);
and U6590 (N_6590,N_5400,N_5975);
or U6591 (N_6591,N_4992,N_5031);
or U6592 (N_6592,N_4427,N_4297);
nand U6593 (N_6593,N_4595,N_5223);
nor U6594 (N_6594,N_5287,N_4084);
and U6595 (N_6595,N_5531,N_4086);
and U6596 (N_6596,N_4503,N_5126);
and U6597 (N_6597,N_4475,N_4141);
and U6598 (N_6598,N_4906,N_5290);
and U6599 (N_6599,N_4893,N_4950);
and U6600 (N_6600,N_4633,N_5104);
or U6601 (N_6601,N_5510,N_4985);
nor U6602 (N_6602,N_5612,N_4916);
nand U6603 (N_6603,N_5714,N_4449);
and U6604 (N_6604,N_5190,N_4724);
nor U6605 (N_6605,N_4277,N_4197);
or U6606 (N_6606,N_4171,N_4366);
and U6607 (N_6607,N_4796,N_4433);
nor U6608 (N_6608,N_4164,N_4841);
nand U6609 (N_6609,N_4512,N_5169);
nand U6610 (N_6610,N_4092,N_4413);
nor U6611 (N_6611,N_4093,N_5459);
nor U6612 (N_6612,N_5424,N_5439);
or U6613 (N_6613,N_5163,N_4586);
and U6614 (N_6614,N_4831,N_4953);
or U6615 (N_6615,N_5738,N_5700);
nor U6616 (N_6616,N_4144,N_4784);
nor U6617 (N_6617,N_5317,N_4730);
nor U6618 (N_6618,N_4239,N_4219);
and U6619 (N_6619,N_4237,N_5989);
nor U6620 (N_6620,N_5046,N_5924);
nor U6621 (N_6621,N_5849,N_5494);
nor U6622 (N_6622,N_4540,N_4749);
nor U6623 (N_6623,N_4049,N_4377);
and U6624 (N_6624,N_5946,N_5272);
or U6625 (N_6625,N_4495,N_5559);
nand U6626 (N_6626,N_5291,N_4854);
or U6627 (N_6627,N_5176,N_5279);
and U6628 (N_6628,N_5183,N_5408);
nor U6629 (N_6629,N_5641,N_4430);
nor U6630 (N_6630,N_5179,N_5772);
or U6631 (N_6631,N_5662,N_4686);
nand U6632 (N_6632,N_4585,N_4369);
and U6633 (N_6633,N_4176,N_4661);
nand U6634 (N_6634,N_5160,N_5263);
or U6635 (N_6635,N_4058,N_5940);
or U6636 (N_6636,N_4361,N_5117);
nand U6637 (N_6637,N_5884,N_5095);
and U6638 (N_6638,N_5129,N_4040);
nand U6639 (N_6639,N_5256,N_5121);
nor U6640 (N_6640,N_4570,N_5380);
or U6641 (N_6641,N_4513,N_4996);
nand U6642 (N_6642,N_4649,N_4845);
nand U6643 (N_6643,N_4039,N_5888);
nor U6644 (N_6644,N_5425,N_5019);
and U6645 (N_6645,N_5744,N_5457);
or U6646 (N_6646,N_4594,N_4910);
or U6647 (N_6647,N_5354,N_4001);
or U6648 (N_6648,N_4465,N_4857);
and U6649 (N_6649,N_5732,N_5438);
nor U6650 (N_6650,N_4499,N_4543);
nand U6651 (N_6651,N_5502,N_4523);
or U6652 (N_6652,N_4600,N_5543);
nor U6653 (N_6653,N_5964,N_4995);
or U6654 (N_6654,N_5683,N_4886);
or U6655 (N_6655,N_5790,N_5481);
or U6656 (N_6656,N_4063,N_4667);
nor U6657 (N_6657,N_4378,N_4247);
or U6658 (N_6658,N_4214,N_5960);
and U6659 (N_6659,N_5896,N_4768);
or U6660 (N_6660,N_4956,N_4567);
nor U6661 (N_6661,N_4612,N_4090);
nand U6662 (N_6662,N_4823,N_4988);
nor U6663 (N_6663,N_5284,N_5361);
or U6664 (N_6664,N_5013,N_5931);
or U6665 (N_6665,N_4534,N_4668);
nor U6666 (N_6666,N_5015,N_4550);
nor U6667 (N_6667,N_4789,N_5899);
nor U6668 (N_6668,N_5869,N_5092);
nand U6669 (N_6669,N_5995,N_5721);
nand U6670 (N_6670,N_4344,N_4742);
nor U6671 (N_6671,N_4149,N_5484);
or U6672 (N_6672,N_5099,N_5123);
nand U6673 (N_6673,N_4524,N_4350);
xor U6674 (N_6674,N_5986,N_5213);
nor U6675 (N_6675,N_5741,N_5833);
xor U6676 (N_6676,N_4098,N_4644);
or U6677 (N_6677,N_4760,N_5327);
nor U6678 (N_6678,N_4117,N_5723);
or U6679 (N_6679,N_4471,N_4656);
or U6680 (N_6680,N_4095,N_5548);
nor U6681 (N_6681,N_5670,N_4829);
nand U6682 (N_6682,N_5500,N_5857);
nand U6683 (N_6683,N_4485,N_5257);
nand U6684 (N_6684,N_4616,N_5344);
nor U6685 (N_6685,N_4873,N_4276);
and U6686 (N_6686,N_4410,N_4672);
or U6687 (N_6687,N_4089,N_4111);
nand U6688 (N_6688,N_4545,N_5632);
nand U6689 (N_6689,N_4614,N_5648);
nand U6690 (N_6690,N_4723,N_4905);
and U6691 (N_6691,N_4879,N_4486);
and U6692 (N_6692,N_5517,N_5238);
nand U6693 (N_6693,N_5753,N_4735);
nor U6694 (N_6694,N_5199,N_5246);
nand U6695 (N_6695,N_4414,N_4267);
or U6696 (N_6696,N_4417,N_5659);
nor U6697 (N_6697,N_5630,N_4954);
and U6698 (N_6698,N_4274,N_4832);
nor U6699 (N_6699,N_4103,N_5661);
nand U6700 (N_6700,N_5942,N_5089);
or U6701 (N_6701,N_5330,N_4980);
nand U6702 (N_6702,N_4952,N_5274);
and U6703 (N_6703,N_4650,N_4178);
and U6704 (N_6704,N_4509,N_4370);
nand U6705 (N_6705,N_4335,N_5148);
nand U6706 (N_6706,N_4220,N_4462);
nand U6707 (N_6707,N_4174,N_5189);
and U6708 (N_6708,N_5767,N_5468);
nor U6709 (N_6709,N_5587,N_4673);
xnor U6710 (N_6710,N_5913,N_4623);
nor U6711 (N_6711,N_5267,N_5078);
nand U6712 (N_6712,N_4196,N_4032);
and U6713 (N_6713,N_5446,N_4511);
or U6714 (N_6714,N_5984,N_5487);
nor U6715 (N_6715,N_5786,N_5488);
or U6716 (N_6716,N_5991,N_5615);
and U6717 (N_6717,N_4697,N_4325);
or U6718 (N_6718,N_4257,N_5618);
and U6719 (N_6719,N_5161,N_5293);
nor U6720 (N_6720,N_5512,N_5962);
or U6721 (N_6721,N_5155,N_4085);
or U6722 (N_6722,N_4211,N_4920);
nor U6723 (N_6723,N_4693,N_4904);
or U6724 (N_6724,N_4833,N_4097);
and U6725 (N_6725,N_5834,N_4054);
nand U6726 (N_6726,N_5742,N_4636);
and U6727 (N_6727,N_5226,N_4264);
and U6728 (N_6728,N_4811,N_4431);
or U6729 (N_6729,N_4588,N_4631);
or U6730 (N_6730,N_5194,N_5770);
or U6731 (N_6731,N_5643,N_5871);
nand U6732 (N_6732,N_5075,N_5072);
and U6733 (N_6733,N_5332,N_4914);
nor U6734 (N_6734,N_5342,N_5581);
and U6735 (N_6735,N_5974,N_4166);
or U6736 (N_6736,N_4094,N_4358);
nor U6737 (N_6737,N_4330,N_4852);
and U6738 (N_6738,N_4132,N_5449);
or U6739 (N_6739,N_5450,N_5460);
or U6740 (N_6740,N_5268,N_4021);
and U6741 (N_6741,N_4482,N_4791);
and U6742 (N_6742,N_5620,N_4124);
or U6743 (N_6743,N_5908,N_4943);
or U6744 (N_6744,N_4004,N_4582);
nor U6745 (N_6745,N_5271,N_4867);
nand U6746 (N_6746,N_5499,N_4348);
nor U6747 (N_6747,N_4772,N_4596);
and U6748 (N_6748,N_4903,N_5320);
xnor U6749 (N_6749,N_4734,N_4978);
or U6750 (N_6750,N_4580,N_4455);
nand U6751 (N_6751,N_4468,N_5635);
and U6752 (N_6752,N_5897,N_5058);
and U6753 (N_6753,N_4202,N_4339);
nand U6754 (N_6754,N_5230,N_4346);
nor U6755 (N_6755,N_4822,N_5218);
xor U6756 (N_6756,N_5417,N_5756);
or U6757 (N_6757,N_4281,N_4933);
or U6758 (N_6758,N_5193,N_4382);
or U6759 (N_6759,N_4298,N_5688);
and U6760 (N_6760,N_5474,N_4028);
and U6761 (N_6761,N_5392,N_4286);
nor U6762 (N_6762,N_5677,N_5158);
nand U6763 (N_6763,N_4563,N_4548);
nor U6764 (N_6764,N_5983,N_4969);
and U6765 (N_6765,N_4967,N_5801);
and U6766 (N_6766,N_5100,N_5266);
nand U6767 (N_6767,N_5802,N_4452);
nand U6768 (N_6768,N_5832,N_5774);
or U6769 (N_6769,N_4060,N_5617);
nand U6770 (N_6770,N_5295,N_5249);
or U6771 (N_6771,N_5201,N_5080);
and U6772 (N_6772,N_5999,N_4617);
or U6773 (N_6773,N_5260,N_5243);
nand U6774 (N_6774,N_4180,N_5378);
nor U6775 (N_6775,N_4326,N_4334);
and U6776 (N_6776,N_4229,N_5540);
or U6777 (N_6777,N_4630,N_5269);
or U6778 (N_6778,N_4765,N_4678);
nand U6779 (N_6779,N_4045,N_4232);
nor U6780 (N_6780,N_5331,N_5926);
or U6781 (N_6781,N_5195,N_4088);
nor U6782 (N_6782,N_4301,N_5941);
or U6783 (N_6783,N_4029,N_4272);
nor U6784 (N_6784,N_5255,N_5197);
nand U6785 (N_6785,N_5475,N_5967);
nor U6786 (N_6786,N_4942,N_4194);
nor U6787 (N_6787,N_4912,N_4615);
or U6788 (N_6788,N_5663,N_5890);
nand U6789 (N_6789,N_5043,N_5286);
nand U6790 (N_6790,N_5041,N_5029);
and U6791 (N_6791,N_4077,N_5977);
or U6792 (N_6792,N_4222,N_4252);
nor U6793 (N_6793,N_4336,N_4203);
and U6794 (N_6794,N_4907,N_4747);
and U6795 (N_6795,N_5088,N_5836);
and U6796 (N_6796,N_5372,N_5985);
nand U6797 (N_6797,N_4767,N_5483);
nor U6798 (N_6798,N_5341,N_5049);
and U6799 (N_6799,N_4762,N_4385);
and U6800 (N_6800,N_4477,N_4990);
nor U6801 (N_6801,N_4508,N_5876);
and U6802 (N_6802,N_4065,N_5916);
nand U6803 (N_6803,N_4293,N_4023);
or U6804 (N_6804,N_4556,N_5091);
or U6805 (N_6805,N_4754,N_4409);
nand U6806 (N_6806,N_5312,N_4733);
or U6807 (N_6807,N_4666,N_5596);
or U6808 (N_6808,N_5166,N_5399);
nor U6809 (N_6809,N_5328,N_5846);
nor U6810 (N_6810,N_4691,N_4863);
nand U6811 (N_6811,N_4362,N_5349);
nand U6812 (N_6812,N_5102,N_4855);
nor U6813 (N_6813,N_5712,N_5277);
nand U6814 (N_6814,N_5364,N_5325);
xnor U6815 (N_6815,N_5586,N_4598);
or U6816 (N_6816,N_4450,N_4494);
and U6817 (N_6817,N_5570,N_4785);
nand U6818 (N_6818,N_5168,N_4815);
and U6819 (N_6819,N_5103,N_5607);
nand U6820 (N_6820,N_4310,N_4056);
nor U6821 (N_6821,N_4868,N_5359);
and U6822 (N_6822,N_4168,N_5083);
nand U6823 (N_6823,N_5336,N_5731);
nand U6824 (N_6824,N_5546,N_5848);
nor U6825 (N_6825,N_4006,N_5333);
nor U6826 (N_6826,N_5863,N_5055);
and U6827 (N_6827,N_4260,N_4019);
or U6828 (N_6828,N_4400,N_4314);
nor U6829 (N_6829,N_5827,N_4574);
and U6830 (N_6830,N_4709,N_4794);
and U6831 (N_6831,N_4292,N_5153);
nand U6832 (N_6832,N_4875,N_4965);
nor U6833 (N_6833,N_4552,N_4870);
or U6834 (N_6834,N_4069,N_4758);
nand U6835 (N_6835,N_5270,N_5002);
or U6836 (N_6836,N_4104,N_5120);
nand U6837 (N_6837,N_5808,N_4844);
and U6838 (N_6838,N_4818,N_5292);
or U6839 (N_6839,N_4294,N_4038);
nand U6840 (N_6840,N_5495,N_5135);
nand U6841 (N_6841,N_4456,N_4332);
nor U6842 (N_6842,N_5980,N_4878);
nor U6843 (N_6843,N_4304,N_5478);
and U6844 (N_6844,N_5590,N_5593);
nor U6845 (N_6845,N_5113,N_5609);
or U6846 (N_6846,N_5992,N_4479);
and U6847 (N_6847,N_5387,N_5785);
nor U6848 (N_6848,N_4737,N_4076);
or U6849 (N_6849,N_4521,N_5831);
nand U6850 (N_6850,N_5047,N_5669);
and U6851 (N_6851,N_4951,N_4218);
nor U6852 (N_6852,N_5729,N_5097);
nand U6853 (N_6853,N_4922,N_4470);
or U6854 (N_6854,N_5865,N_4862);
nor U6855 (N_6855,N_4827,N_4526);
and U6856 (N_6856,N_4364,N_4966);
nor U6857 (N_6857,N_4555,N_5963);
or U6858 (N_6858,N_5070,N_4781);
and U6859 (N_6859,N_5415,N_4915);
nor U6860 (N_6860,N_4837,N_4587);
xnor U6861 (N_6861,N_5032,N_5375);
or U6862 (N_6862,N_5132,N_5994);
nor U6863 (N_6863,N_4675,N_4851);
nand U6864 (N_6864,N_5203,N_4674);
and U6865 (N_6865,N_4496,N_5024);
nor U6866 (N_6866,N_4843,N_4628);
and U6867 (N_6867,N_5447,N_4121);
and U6868 (N_6868,N_5862,N_4061);
nor U6869 (N_6869,N_4016,N_4290);
or U6870 (N_6870,N_4291,N_5891);
nand U6871 (N_6871,N_5923,N_4036);
nor U6872 (N_6872,N_4554,N_5961);
or U6873 (N_6873,N_5904,N_5018);
or U6874 (N_6874,N_5830,N_4120);
nand U6875 (N_6875,N_4597,N_5172);
and U6876 (N_6876,N_5970,N_5885);
and U6877 (N_6877,N_4037,N_4787);
nand U6878 (N_6878,N_5821,N_5021);
nand U6879 (N_6879,N_4005,N_4828);
nand U6880 (N_6880,N_5090,N_4331);
and U6881 (N_6881,N_5633,N_4027);
and U6882 (N_6882,N_4204,N_5254);
nor U6883 (N_6883,N_4993,N_4727);
xor U6884 (N_6884,N_4608,N_5788);
nand U6885 (N_6885,N_4162,N_4261);
nand U6886 (N_6886,N_4020,N_5736);
nand U6887 (N_6887,N_5497,N_4561);
nor U6888 (N_6888,N_5186,N_5765);
nand U6889 (N_6889,N_4790,N_4925);
or U6890 (N_6890,N_5792,N_4763);
and U6891 (N_6891,N_4853,N_4799);
and U6892 (N_6892,N_4251,N_4714);
nor U6893 (N_6893,N_4891,N_5370);
xor U6894 (N_6894,N_4547,N_5915);
or U6895 (N_6895,N_5235,N_5313);
or U6896 (N_6896,N_4786,N_5684);
nor U6897 (N_6897,N_5837,N_4303);
nand U6898 (N_6898,N_5708,N_5911);
nand U6899 (N_6899,N_5678,N_5309);
nand U6900 (N_6900,N_5599,N_4415);
nor U6901 (N_6901,N_5614,N_4544);
nor U6902 (N_6902,N_4390,N_5550);
nor U6903 (N_6903,N_5300,N_4128);
and U6904 (N_6904,N_4874,N_5140);
or U6905 (N_6905,N_5568,N_4198);
or U6906 (N_6906,N_4437,N_4154);
and U6907 (N_6907,N_5937,N_5278);
or U6908 (N_6908,N_5404,N_5760);
nand U6909 (N_6909,N_4715,N_5769);
nor U6910 (N_6910,N_5728,N_4761);
or U6911 (N_6911,N_4119,N_4209);
nor U6912 (N_6912,N_5397,N_5709);
and U6913 (N_6913,N_4136,N_5389);
and U6914 (N_6914,N_5560,N_5844);
or U6915 (N_6915,N_4515,N_4083);
nand U6916 (N_6916,N_4576,N_5039);
or U6917 (N_6917,N_5855,N_5170);
or U6918 (N_6918,N_5464,N_5525);
nor U6919 (N_6919,N_5789,N_4476);
nand U6920 (N_6920,N_5759,N_4275);
nor U6921 (N_6921,N_4778,N_5301);
or U6922 (N_6922,N_4817,N_4881);
nor U6923 (N_6923,N_4461,N_4937);
nand U6924 (N_6924,N_4394,N_4349);
nor U6925 (N_6925,N_4607,N_4460);
nor U6926 (N_6926,N_5686,N_5504);
or U6927 (N_6927,N_4987,N_5894);
nor U6928 (N_6928,N_5952,N_4148);
nand U6929 (N_6929,N_4970,N_5350);
and U6930 (N_6930,N_5393,N_4658);
nand U6931 (N_6931,N_4015,N_4046);
nor U6932 (N_6932,N_4424,N_5247);
and U6933 (N_6933,N_5491,N_5880);
nor U6934 (N_6934,N_5289,N_5069);
and U6935 (N_6935,N_5749,N_5933);
and U6936 (N_6936,N_5878,N_5545);
nor U6937 (N_6937,N_5258,N_4165);
nand U6938 (N_6938,N_4718,N_4726);
or U6939 (N_6939,N_5748,N_4018);
or U6940 (N_6940,N_5675,N_4306);
or U6941 (N_6941,N_4448,N_5445);
nor U6942 (N_6942,N_4399,N_5949);
or U6943 (N_6943,N_5806,N_5737);
nand U6944 (N_6944,N_4858,N_4182);
or U6945 (N_6945,N_5452,N_4923);
nand U6946 (N_6946,N_4610,N_5469);
nor U6947 (N_6947,N_4459,N_5184);
or U6948 (N_6948,N_5352,N_4108);
nor U6949 (N_6949,N_5993,N_5701);
nand U6950 (N_6950,N_5561,N_5902);
xnor U6951 (N_6951,N_4457,N_4472);
nor U6952 (N_6952,N_4129,N_5396);
or U6953 (N_6953,N_5345,N_5353);
nor U6954 (N_6954,N_5656,N_5217);
nor U6955 (N_6955,N_5033,N_4398);
nand U6956 (N_6956,N_5698,N_5437);
and U6957 (N_6957,N_4835,N_4341);
or U6958 (N_6958,N_5624,N_4091);
or U6959 (N_6959,N_5501,N_4898);
nand U6960 (N_6960,N_5854,N_5302);
nor U6961 (N_6961,N_4643,N_5557);
xor U6962 (N_6962,N_4030,N_5567);
or U6963 (N_6963,N_4492,N_4573);
or U6964 (N_6964,N_5853,N_4412);
nor U6965 (N_6965,N_4640,N_4918);
or U6966 (N_6966,N_4700,N_4819);
and U6967 (N_6967,N_4150,N_5990);
nor U6968 (N_6968,N_5513,N_4860);
nor U6969 (N_6969,N_5966,N_4243);
or U6970 (N_6970,N_4248,N_5740);
nor U6971 (N_6971,N_5572,N_5138);
nor U6972 (N_6972,N_5722,N_5866);
or U6973 (N_6973,N_5544,N_5231);
or U6974 (N_6974,N_5416,N_4759);
and U6975 (N_6975,N_5580,N_5781);
and U6976 (N_6976,N_5241,N_4888);
or U6977 (N_6977,N_5775,N_4134);
nor U6978 (N_6978,N_5845,N_4795);
and U6979 (N_6979,N_5528,N_5440);
and U6980 (N_6980,N_5851,N_4895);
nor U6981 (N_6981,N_5889,N_4258);
nor U6982 (N_6982,N_5098,N_5411);
nand U6983 (N_6983,N_5636,N_4466);
nor U6984 (N_6984,N_4549,N_4139);
nor U6985 (N_6985,N_4081,N_4047);
nor U6986 (N_6986,N_4779,N_4664);
nor U6987 (N_6987,N_4624,N_5114);
nand U6988 (N_6988,N_5535,N_4280);
or U6989 (N_6989,N_5898,N_4684);
nand U6990 (N_6990,N_5444,N_5068);
nor U6991 (N_6991,N_5660,N_4577);
nand U6992 (N_6992,N_4138,N_4621);
or U6993 (N_6993,N_4368,N_4262);
and U6994 (N_6994,N_5676,N_5905);
nor U6995 (N_6995,N_5062,N_4940);
and U6996 (N_6996,N_5791,N_4520);
and U6997 (N_6997,N_5192,N_4360);
nor U6998 (N_6998,N_5826,N_4131);
nand U6999 (N_6999,N_5598,N_5414);
nor U7000 (N_7000,N_5965,N_4847);
nand U7001 (N_7001,N_5192,N_4854);
and U7002 (N_7002,N_4598,N_4733);
nor U7003 (N_7003,N_4165,N_5261);
and U7004 (N_7004,N_4901,N_4189);
and U7005 (N_7005,N_5904,N_5106);
nor U7006 (N_7006,N_4518,N_5589);
nand U7007 (N_7007,N_5705,N_4706);
nor U7008 (N_7008,N_4156,N_4988);
or U7009 (N_7009,N_5680,N_4942);
and U7010 (N_7010,N_5255,N_4254);
and U7011 (N_7011,N_5022,N_5077);
nand U7012 (N_7012,N_5353,N_4028);
and U7013 (N_7013,N_4861,N_5190);
nor U7014 (N_7014,N_4798,N_5917);
xnor U7015 (N_7015,N_5173,N_5479);
nand U7016 (N_7016,N_5903,N_4507);
nor U7017 (N_7017,N_5530,N_4903);
or U7018 (N_7018,N_5915,N_5518);
nand U7019 (N_7019,N_4911,N_4039);
and U7020 (N_7020,N_5937,N_4909);
or U7021 (N_7021,N_5526,N_4055);
nor U7022 (N_7022,N_4921,N_5952);
nand U7023 (N_7023,N_4785,N_5593);
nand U7024 (N_7024,N_5671,N_4487);
or U7025 (N_7025,N_5304,N_4690);
or U7026 (N_7026,N_5383,N_4988);
or U7027 (N_7027,N_4843,N_4523);
nor U7028 (N_7028,N_5266,N_4183);
and U7029 (N_7029,N_5280,N_4472);
and U7030 (N_7030,N_4878,N_4869);
nand U7031 (N_7031,N_5991,N_4703);
xnor U7032 (N_7032,N_5448,N_4300);
nor U7033 (N_7033,N_5700,N_4367);
nand U7034 (N_7034,N_5365,N_4246);
nor U7035 (N_7035,N_5794,N_5430);
nor U7036 (N_7036,N_5540,N_5327);
nor U7037 (N_7037,N_5602,N_5739);
and U7038 (N_7038,N_4147,N_5025);
nand U7039 (N_7039,N_4657,N_4568);
nand U7040 (N_7040,N_5091,N_5206);
and U7041 (N_7041,N_5688,N_5859);
and U7042 (N_7042,N_4706,N_5733);
or U7043 (N_7043,N_4876,N_5384);
and U7044 (N_7044,N_5824,N_5890);
nand U7045 (N_7045,N_5238,N_4146);
nor U7046 (N_7046,N_5477,N_5582);
and U7047 (N_7047,N_4282,N_4927);
or U7048 (N_7048,N_5329,N_5013);
and U7049 (N_7049,N_5175,N_4055);
nand U7050 (N_7050,N_4833,N_4447);
xor U7051 (N_7051,N_5659,N_5364);
nor U7052 (N_7052,N_5454,N_4217);
nand U7053 (N_7053,N_4124,N_5689);
nand U7054 (N_7054,N_4450,N_4365);
nand U7055 (N_7055,N_5454,N_4845);
nor U7056 (N_7056,N_5910,N_5525);
and U7057 (N_7057,N_4663,N_5648);
nor U7058 (N_7058,N_4248,N_5189);
or U7059 (N_7059,N_5960,N_5560);
and U7060 (N_7060,N_4093,N_4744);
and U7061 (N_7061,N_5122,N_4910);
nand U7062 (N_7062,N_5342,N_5647);
and U7063 (N_7063,N_4139,N_5580);
nand U7064 (N_7064,N_5427,N_5269);
or U7065 (N_7065,N_4386,N_4209);
nor U7066 (N_7066,N_5329,N_5045);
nand U7067 (N_7067,N_4593,N_4034);
or U7068 (N_7068,N_5655,N_4857);
or U7069 (N_7069,N_4165,N_5920);
nor U7070 (N_7070,N_5656,N_5969);
nand U7071 (N_7071,N_5053,N_5835);
nand U7072 (N_7072,N_5803,N_4924);
nor U7073 (N_7073,N_5371,N_4987);
and U7074 (N_7074,N_5337,N_5466);
or U7075 (N_7075,N_4425,N_4317);
nor U7076 (N_7076,N_5764,N_4727);
and U7077 (N_7077,N_5578,N_4647);
nor U7078 (N_7078,N_5997,N_4334);
and U7079 (N_7079,N_4837,N_4369);
nand U7080 (N_7080,N_5913,N_4514);
nand U7081 (N_7081,N_5031,N_5883);
nand U7082 (N_7082,N_4480,N_5513);
and U7083 (N_7083,N_4967,N_4073);
nand U7084 (N_7084,N_5267,N_5278);
nor U7085 (N_7085,N_5868,N_5980);
nor U7086 (N_7086,N_5127,N_5377);
or U7087 (N_7087,N_4132,N_5373);
or U7088 (N_7088,N_5681,N_5130);
or U7089 (N_7089,N_5150,N_4525);
and U7090 (N_7090,N_4670,N_4841);
nand U7091 (N_7091,N_4800,N_4623);
nand U7092 (N_7092,N_4829,N_5993);
nor U7093 (N_7093,N_5827,N_5663);
nor U7094 (N_7094,N_5409,N_4715);
nand U7095 (N_7095,N_5493,N_5637);
nor U7096 (N_7096,N_5477,N_5622);
nand U7097 (N_7097,N_4959,N_5184);
and U7098 (N_7098,N_5696,N_4397);
or U7099 (N_7099,N_4085,N_5426);
nor U7100 (N_7100,N_4907,N_4374);
and U7101 (N_7101,N_5028,N_5054);
nand U7102 (N_7102,N_5066,N_5146);
nor U7103 (N_7103,N_4544,N_5926);
and U7104 (N_7104,N_4788,N_5874);
or U7105 (N_7105,N_4914,N_4459);
nor U7106 (N_7106,N_4124,N_5414);
nor U7107 (N_7107,N_4292,N_5026);
or U7108 (N_7108,N_5834,N_5659);
or U7109 (N_7109,N_4607,N_4132);
nand U7110 (N_7110,N_4243,N_5147);
nor U7111 (N_7111,N_5091,N_5100);
or U7112 (N_7112,N_5287,N_5707);
nand U7113 (N_7113,N_5994,N_5895);
or U7114 (N_7114,N_5435,N_4883);
or U7115 (N_7115,N_5585,N_5142);
nand U7116 (N_7116,N_4519,N_5061);
or U7117 (N_7117,N_5544,N_5954);
or U7118 (N_7118,N_5452,N_5391);
and U7119 (N_7119,N_4797,N_5892);
nor U7120 (N_7120,N_5921,N_5546);
nor U7121 (N_7121,N_5231,N_4868);
nor U7122 (N_7122,N_5510,N_5338);
nand U7123 (N_7123,N_4014,N_4575);
nand U7124 (N_7124,N_4045,N_5488);
and U7125 (N_7125,N_4187,N_4598);
nor U7126 (N_7126,N_5953,N_4376);
and U7127 (N_7127,N_4327,N_5409);
or U7128 (N_7128,N_4426,N_4550);
or U7129 (N_7129,N_4513,N_4814);
nor U7130 (N_7130,N_4100,N_4919);
and U7131 (N_7131,N_5358,N_4438);
nand U7132 (N_7132,N_5063,N_4653);
nand U7133 (N_7133,N_4356,N_5493);
nand U7134 (N_7134,N_5289,N_4258);
and U7135 (N_7135,N_5353,N_5569);
nor U7136 (N_7136,N_4327,N_5128);
and U7137 (N_7137,N_4531,N_5400);
nor U7138 (N_7138,N_4846,N_5803);
and U7139 (N_7139,N_5225,N_5137);
nor U7140 (N_7140,N_4199,N_4403);
or U7141 (N_7141,N_4132,N_4713);
or U7142 (N_7142,N_4890,N_5997);
and U7143 (N_7143,N_4794,N_4030);
or U7144 (N_7144,N_4333,N_4278);
and U7145 (N_7145,N_4506,N_5223);
nor U7146 (N_7146,N_4371,N_5695);
or U7147 (N_7147,N_5541,N_5075);
nor U7148 (N_7148,N_5049,N_5350);
or U7149 (N_7149,N_5532,N_5336);
or U7150 (N_7150,N_4400,N_5109);
nand U7151 (N_7151,N_5234,N_5628);
nand U7152 (N_7152,N_5260,N_4522);
and U7153 (N_7153,N_4434,N_5852);
or U7154 (N_7154,N_5337,N_5522);
nor U7155 (N_7155,N_5102,N_5561);
nor U7156 (N_7156,N_4933,N_5538);
nand U7157 (N_7157,N_5770,N_5289);
nor U7158 (N_7158,N_5525,N_4276);
and U7159 (N_7159,N_5109,N_4584);
nor U7160 (N_7160,N_5638,N_4602);
nor U7161 (N_7161,N_5242,N_4578);
and U7162 (N_7162,N_5464,N_5381);
or U7163 (N_7163,N_5967,N_4420);
or U7164 (N_7164,N_5305,N_5172);
and U7165 (N_7165,N_5434,N_5085);
nand U7166 (N_7166,N_4024,N_4331);
nand U7167 (N_7167,N_4001,N_5399);
nand U7168 (N_7168,N_5915,N_5800);
and U7169 (N_7169,N_5626,N_4828);
or U7170 (N_7170,N_4134,N_4863);
and U7171 (N_7171,N_5553,N_4097);
or U7172 (N_7172,N_4352,N_5106);
or U7173 (N_7173,N_4446,N_4025);
or U7174 (N_7174,N_4952,N_4857);
nor U7175 (N_7175,N_4180,N_5136);
nor U7176 (N_7176,N_5426,N_5120);
or U7177 (N_7177,N_4863,N_5376);
or U7178 (N_7178,N_4013,N_4764);
and U7179 (N_7179,N_4308,N_5581);
or U7180 (N_7180,N_4160,N_4633);
and U7181 (N_7181,N_4341,N_5707);
or U7182 (N_7182,N_4222,N_5747);
nand U7183 (N_7183,N_4447,N_4731);
or U7184 (N_7184,N_4051,N_5359);
and U7185 (N_7185,N_5736,N_5649);
or U7186 (N_7186,N_5413,N_5995);
and U7187 (N_7187,N_4255,N_5411);
and U7188 (N_7188,N_4659,N_4242);
or U7189 (N_7189,N_4327,N_4896);
xnor U7190 (N_7190,N_5764,N_4410);
nand U7191 (N_7191,N_5532,N_5414);
nor U7192 (N_7192,N_5506,N_4312);
xor U7193 (N_7193,N_4418,N_4750);
nand U7194 (N_7194,N_4352,N_5397);
nand U7195 (N_7195,N_5795,N_4738);
or U7196 (N_7196,N_4849,N_5160);
nor U7197 (N_7197,N_5698,N_4924);
nor U7198 (N_7198,N_4392,N_4023);
nand U7199 (N_7199,N_4970,N_5692);
nor U7200 (N_7200,N_5490,N_5110);
nor U7201 (N_7201,N_4348,N_4961);
or U7202 (N_7202,N_4879,N_5682);
nor U7203 (N_7203,N_4300,N_5176);
xnor U7204 (N_7204,N_4279,N_5893);
nand U7205 (N_7205,N_5553,N_5038);
and U7206 (N_7206,N_5402,N_4079);
or U7207 (N_7207,N_5955,N_4308);
nor U7208 (N_7208,N_5360,N_5680);
nor U7209 (N_7209,N_4087,N_5000);
or U7210 (N_7210,N_5364,N_5959);
nand U7211 (N_7211,N_5377,N_5393);
nor U7212 (N_7212,N_4539,N_5217);
and U7213 (N_7213,N_4076,N_4345);
nor U7214 (N_7214,N_5131,N_4538);
nor U7215 (N_7215,N_5103,N_5135);
and U7216 (N_7216,N_5053,N_4434);
or U7217 (N_7217,N_5761,N_4550);
nand U7218 (N_7218,N_4711,N_5208);
nand U7219 (N_7219,N_4088,N_4724);
or U7220 (N_7220,N_5840,N_5678);
nand U7221 (N_7221,N_5850,N_5101);
nand U7222 (N_7222,N_4044,N_4013);
and U7223 (N_7223,N_5615,N_4260);
and U7224 (N_7224,N_4021,N_5404);
and U7225 (N_7225,N_4329,N_4940);
nor U7226 (N_7226,N_4320,N_4333);
nand U7227 (N_7227,N_5492,N_5349);
nor U7228 (N_7228,N_4080,N_4413);
and U7229 (N_7229,N_4402,N_4940);
or U7230 (N_7230,N_4586,N_4084);
nor U7231 (N_7231,N_5395,N_5501);
nor U7232 (N_7232,N_5912,N_4205);
and U7233 (N_7233,N_4948,N_5224);
nand U7234 (N_7234,N_4386,N_5526);
or U7235 (N_7235,N_4987,N_5593);
and U7236 (N_7236,N_5572,N_4605);
nor U7237 (N_7237,N_4639,N_4194);
or U7238 (N_7238,N_4242,N_4980);
nand U7239 (N_7239,N_5609,N_5863);
and U7240 (N_7240,N_4636,N_4945);
nor U7241 (N_7241,N_4188,N_4655);
and U7242 (N_7242,N_5253,N_4234);
nand U7243 (N_7243,N_4920,N_4784);
nand U7244 (N_7244,N_5034,N_5719);
nor U7245 (N_7245,N_4130,N_5547);
nand U7246 (N_7246,N_5594,N_4626);
and U7247 (N_7247,N_5296,N_4749);
or U7248 (N_7248,N_5480,N_5690);
or U7249 (N_7249,N_5604,N_5041);
or U7250 (N_7250,N_4904,N_5001);
nand U7251 (N_7251,N_4935,N_4162);
and U7252 (N_7252,N_4566,N_5699);
nand U7253 (N_7253,N_5221,N_5141);
nor U7254 (N_7254,N_4347,N_5268);
nand U7255 (N_7255,N_5681,N_5470);
nand U7256 (N_7256,N_4760,N_5464);
and U7257 (N_7257,N_4382,N_5665);
or U7258 (N_7258,N_4013,N_5355);
or U7259 (N_7259,N_4786,N_5229);
and U7260 (N_7260,N_4439,N_4603);
nor U7261 (N_7261,N_4999,N_5453);
nor U7262 (N_7262,N_5621,N_4406);
nor U7263 (N_7263,N_5676,N_5766);
nand U7264 (N_7264,N_5835,N_5396);
nor U7265 (N_7265,N_5108,N_5959);
or U7266 (N_7266,N_4507,N_4310);
nor U7267 (N_7267,N_5619,N_5470);
nor U7268 (N_7268,N_5164,N_5803);
nand U7269 (N_7269,N_4189,N_4367);
nor U7270 (N_7270,N_4785,N_4626);
or U7271 (N_7271,N_4044,N_5614);
nor U7272 (N_7272,N_5652,N_4362);
and U7273 (N_7273,N_5701,N_5409);
and U7274 (N_7274,N_4475,N_4915);
nor U7275 (N_7275,N_4722,N_4785);
and U7276 (N_7276,N_4997,N_4312);
and U7277 (N_7277,N_5631,N_4701);
nand U7278 (N_7278,N_5955,N_4762);
nor U7279 (N_7279,N_4693,N_4605);
nor U7280 (N_7280,N_4036,N_5324);
nand U7281 (N_7281,N_5816,N_4613);
nand U7282 (N_7282,N_5848,N_5235);
nor U7283 (N_7283,N_4366,N_5697);
nor U7284 (N_7284,N_4380,N_5496);
nand U7285 (N_7285,N_4848,N_4555);
and U7286 (N_7286,N_4755,N_4930);
or U7287 (N_7287,N_4380,N_5571);
and U7288 (N_7288,N_5301,N_5692);
or U7289 (N_7289,N_4643,N_4258);
xnor U7290 (N_7290,N_5218,N_5002);
nand U7291 (N_7291,N_4687,N_5854);
or U7292 (N_7292,N_5219,N_5103);
nand U7293 (N_7293,N_4343,N_4515);
nand U7294 (N_7294,N_4799,N_5635);
nand U7295 (N_7295,N_5810,N_4426);
nand U7296 (N_7296,N_4178,N_4321);
nor U7297 (N_7297,N_4667,N_4928);
or U7298 (N_7298,N_5376,N_5621);
nand U7299 (N_7299,N_4709,N_5451);
nand U7300 (N_7300,N_4591,N_4434);
and U7301 (N_7301,N_5668,N_4793);
nor U7302 (N_7302,N_5160,N_4048);
and U7303 (N_7303,N_5945,N_4061);
nor U7304 (N_7304,N_4054,N_5560);
or U7305 (N_7305,N_5663,N_5035);
or U7306 (N_7306,N_5034,N_4119);
nand U7307 (N_7307,N_4122,N_4165);
and U7308 (N_7308,N_4351,N_4506);
and U7309 (N_7309,N_5650,N_4004);
and U7310 (N_7310,N_4819,N_4739);
nand U7311 (N_7311,N_5171,N_4503);
nand U7312 (N_7312,N_5740,N_4170);
nand U7313 (N_7313,N_4471,N_4341);
and U7314 (N_7314,N_4925,N_4726);
nand U7315 (N_7315,N_5390,N_4375);
or U7316 (N_7316,N_4868,N_5681);
nand U7317 (N_7317,N_5074,N_5353);
or U7318 (N_7318,N_4792,N_5437);
and U7319 (N_7319,N_5423,N_5830);
nand U7320 (N_7320,N_4108,N_5872);
nand U7321 (N_7321,N_4167,N_4239);
nor U7322 (N_7322,N_5136,N_5851);
and U7323 (N_7323,N_4283,N_5372);
and U7324 (N_7324,N_5636,N_4993);
nand U7325 (N_7325,N_5256,N_5566);
nor U7326 (N_7326,N_4167,N_4260);
and U7327 (N_7327,N_4407,N_4871);
xnor U7328 (N_7328,N_5393,N_4214);
and U7329 (N_7329,N_5042,N_5689);
nor U7330 (N_7330,N_5367,N_4104);
or U7331 (N_7331,N_4419,N_4696);
nand U7332 (N_7332,N_4666,N_4482);
nor U7333 (N_7333,N_4607,N_5204);
nand U7334 (N_7334,N_5365,N_5680);
and U7335 (N_7335,N_5803,N_4893);
nor U7336 (N_7336,N_4138,N_4460);
nor U7337 (N_7337,N_4512,N_5500);
and U7338 (N_7338,N_5745,N_4244);
or U7339 (N_7339,N_4792,N_5583);
or U7340 (N_7340,N_4158,N_5930);
or U7341 (N_7341,N_5590,N_5699);
or U7342 (N_7342,N_5146,N_4145);
and U7343 (N_7343,N_5156,N_4144);
nor U7344 (N_7344,N_4009,N_4115);
and U7345 (N_7345,N_5568,N_5466);
or U7346 (N_7346,N_4203,N_5182);
or U7347 (N_7347,N_5466,N_5443);
nand U7348 (N_7348,N_4726,N_4221);
or U7349 (N_7349,N_5920,N_5828);
nand U7350 (N_7350,N_4509,N_4954);
or U7351 (N_7351,N_5442,N_5176);
or U7352 (N_7352,N_4095,N_4188);
or U7353 (N_7353,N_4670,N_5530);
or U7354 (N_7354,N_5138,N_5379);
or U7355 (N_7355,N_4987,N_4113);
nand U7356 (N_7356,N_5249,N_4423);
nand U7357 (N_7357,N_4690,N_5777);
nand U7358 (N_7358,N_5868,N_5607);
nor U7359 (N_7359,N_5146,N_4153);
and U7360 (N_7360,N_4029,N_4712);
nand U7361 (N_7361,N_4357,N_5120);
and U7362 (N_7362,N_4948,N_4320);
and U7363 (N_7363,N_4845,N_4736);
or U7364 (N_7364,N_4047,N_5437);
or U7365 (N_7365,N_4604,N_4548);
or U7366 (N_7366,N_4301,N_5504);
and U7367 (N_7367,N_4789,N_5360);
and U7368 (N_7368,N_5540,N_5083);
nand U7369 (N_7369,N_4486,N_4270);
and U7370 (N_7370,N_5089,N_5074);
or U7371 (N_7371,N_5662,N_5611);
and U7372 (N_7372,N_4112,N_5565);
or U7373 (N_7373,N_5306,N_5432);
or U7374 (N_7374,N_5647,N_5112);
nor U7375 (N_7375,N_5217,N_5602);
and U7376 (N_7376,N_5096,N_5259);
and U7377 (N_7377,N_5712,N_4686);
nand U7378 (N_7378,N_5010,N_5939);
nand U7379 (N_7379,N_4969,N_4362);
nor U7380 (N_7380,N_4352,N_4761);
nor U7381 (N_7381,N_4215,N_4683);
and U7382 (N_7382,N_4139,N_4261);
or U7383 (N_7383,N_4920,N_4189);
nand U7384 (N_7384,N_4217,N_4417);
and U7385 (N_7385,N_4421,N_4832);
nor U7386 (N_7386,N_4033,N_4516);
and U7387 (N_7387,N_4751,N_5774);
and U7388 (N_7388,N_4691,N_4529);
and U7389 (N_7389,N_4688,N_5300);
or U7390 (N_7390,N_5784,N_5806);
nand U7391 (N_7391,N_5669,N_4241);
or U7392 (N_7392,N_4077,N_4589);
nand U7393 (N_7393,N_5911,N_4876);
or U7394 (N_7394,N_4843,N_5160);
nand U7395 (N_7395,N_4722,N_4168);
or U7396 (N_7396,N_5046,N_4249);
and U7397 (N_7397,N_5426,N_4197);
and U7398 (N_7398,N_5939,N_5869);
nand U7399 (N_7399,N_4700,N_4318);
and U7400 (N_7400,N_5416,N_4075);
nand U7401 (N_7401,N_5890,N_4469);
nand U7402 (N_7402,N_4000,N_5323);
nand U7403 (N_7403,N_4797,N_5049);
nor U7404 (N_7404,N_4514,N_4215);
nor U7405 (N_7405,N_4659,N_5917);
or U7406 (N_7406,N_4949,N_4431);
nor U7407 (N_7407,N_4638,N_5979);
and U7408 (N_7408,N_5113,N_5829);
nor U7409 (N_7409,N_4432,N_4536);
and U7410 (N_7410,N_4574,N_4850);
and U7411 (N_7411,N_5202,N_5737);
nand U7412 (N_7412,N_4792,N_5401);
or U7413 (N_7413,N_5470,N_4681);
nand U7414 (N_7414,N_4300,N_4498);
nand U7415 (N_7415,N_5269,N_4739);
nor U7416 (N_7416,N_4423,N_4914);
nor U7417 (N_7417,N_5137,N_5247);
and U7418 (N_7418,N_5625,N_4881);
and U7419 (N_7419,N_4555,N_4063);
and U7420 (N_7420,N_4337,N_4884);
nand U7421 (N_7421,N_5131,N_4058);
nor U7422 (N_7422,N_5713,N_5611);
nor U7423 (N_7423,N_5786,N_4393);
nor U7424 (N_7424,N_4747,N_5538);
or U7425 (N_7425,N_5124,N_5840);
and U7426 (N_7426,N_5045,N_5307);
or U7427 (N_7427,N_4876,N_5025);
nand U7428 (N_7428,N_5559,N_4328);
and U7429 (N_7429,N_5514,N_4890);
or U7430 (N_7430,N_5124,N_4551);
nand U7431 (N_7431,N_4407,N_5918);
and U7432 (N_7432,N_4848,N_5485);
or U7433 (N_7433,N_5309,N_4102);
or U7434 (N_7434,N_5171,N_4496);
and U7435 (N_7435,N_5113,N_4322);
and U7436 (N_7436,N_5551,N_4744);
or U7437 (N_7437,N_5555,N_4850);
and U7438 (N_7438,N_5110,N_4430);
or U7439 (N_7439,N_4793,N_4352);
or U7440 (N_7440,N_4062,N_4814);
nor U7441 (N_7441,N_5030,N_4291);
nand U7442 (N_7442,N_4938,N_5058);
and U7443 (N_7443,N_5240,N_5756);
or U7444 (N_7444,N_5914,N_4371);
or U7445 (N_7445,N_5019,N_5011);
nand U7446 (N_7446,N_5664,N_5172);
nor U7447 (N_7447,N_5193,N_5668);
nor U7448 (N_7448,N_4730,N_4514);
or U7449 (N_7449,N_5167,N_5685);
and U7450 (N_7450,N_4663,N_4063);
nand U7451 (N_7451,N_4088,N_4639);
nand U7452 (N_7452,N_4885,N_4954);
or U7453 (N_7453,N_4887,N_5745);
or U7454 (N_7454,N_5144,N_4418);
nand U7455 (N_7455,N_5513,N_5536);
nand U7456 (N_7456,N_5729,N_5100);
or U7457 (N_7457,N_4758,N_4507);
nor U7458 (N_7458,N_4378,N_4586);
nor U7459 (N_7459,N_5595,N_4966);
nand U7460 (N_7460,N_4478,N_4373);
nor U7461 (N_7461,N_5134,N_5300);
and U7462 (N_7462,N_4408,N_5239);
nor U7463 (N_7463,N_4362,N_5649);
and U7464 (N_7464,N_5202,N_5392);
nand U7465 (N_7465,N_5099,N_4937);
nor U7466 (N_7466,N_5465,N_5908);
or U7467 (N_7467,N_4301,N_4091);
and U7468 (N_7468,N_4801,N_4880);
nand U7469 (N_7469,N_5912,N_4544);
nand U7470 (N_7470,N_5904,N_5563);
or U7471 (N_7471,N_5634,N_5365);
nor U7472 (N_7472,N_5038,N_5026);
nor U7473 (N_7473,N_4339,N_5541);
and U7474 (N_7474,N_5304,N_4829);
and U7475 (N_7475,N_4448,N_4701);
nand U7476 (N_7476,N_4981,N_4699);
or U7477 (N_7477,N_5989,N_4558);
nand U7478 (N_7478,N_5203,N_4731);
and U7479 (N_7479,N_4906,N_4998);
or U7480 (N_7480,N_4134,N_4661);
nand U7481 (N_7481,N_5270,N_5925);
nor U7482 (N_7482,N_5209,N_5927);
nor U7483 (N_7483,N_4484,N_4426);
nand U7484 (N_7484,N_5354,N_5980);
and U7485 (N_7485,N_5654,N_4536);
nand U7486 (N_7486,N_4898,N_5725);
or U7487 (N_7487,N_4949,N_5177);
and U7488 (N_7488,N_4545,N_5609);
nor U7489 (N_7489,N_4898,N_4816);
and U7490 (N_7490,N_5976,N_4238);
nand U7491 (N_7491,N_5624,N_5146);
or U7492 (N_7492,N_4551,N_4880);
nor U7493 (N_7493,N_4648,N_4609);
or U7494 (N_7494,N_4595,N_4629);
or U7495 (N_7495,N_4618,N_5738);
nor U7496 (N_7496,N_5509,N_4939);
and U7497 (N_7497,N_5774,N_4371);
nor U7498 (N_7498,N_4647,N_4365);
nor U7499 (N_7499,N_4302,N_4873);
nor U7500 (N_7500,N_5251,N_4140);
and U7501 (N_7501,N_5871,N_4650);
nor U7502 (N_7502,N_5882,N_5255);
or U7503 (N_7503,N_5937,N_4794);
nor U7504 (N_7504,N_5041,N_4791);
or U7505 (N_7505,N_5284,N_5213);
nor U7506 (N_7506,N_5180,N_5030);
and U7507 (N_7507,N_4889,N_4738);
or U7508 (N_7508,N_4535,N_5817);
nor U7509 (N_7509,N_4281,N_5647);
or U7510 (N_7510,N_4181,N_4014);
or U7511 (N_7511,N_5078,N_5473);
nor U7512 (N_7512,N_5686,N_5405);
or U7513 (N_7513,N_5278,N_4329);
and U7514 (N_7514,N_5656,N_5899);
nor U7515 (N_7515,N_4875,N_4712);
nand U7516 (N_7516,N_4876,N_5127);
nand U7517 (N_7517,N_4928,N_5875);
nor U7518 (N_7518,N_5878,N_5298);
nand U7519 (N_7519,N_5169,N_5524);
or U7520 (N_7520,N_4032,N_4929);
and U7521 (N_7521,N_5544,N_4893);
or U7522 (N_7522,N_5538,N_5849);
and U7523 (N_7523,N_4354,N_4292);
and U7524 (N_7524,N_4340,N_4053);
and U7525 (N_7525,N_4199,N_5354);
and U7526 (N_7526,N_4662,N_4495);
nand U7527 (N_7527,N_4816,N_5525);
and U7528 (N_7528,N_4288,N_4803);
nand U7529 (N_7529,N_5772,N_4856);
nor U7530 (N_7530,N_4876,N_4734);
nand U7531 (N_7531,N_5157,N_5946);
nand U7532 (N_7532,N_4338,N_4471);
nor U7533 (N_7533,N_5452,N_5161);
nand U7534 (N_7534,N_4074,N_4829);
and U7535 (N_7535,N_5344,N_5737);
and U7536 (N_7536,N_5263,N_4383);
or U7537 (N_7537,N_5726,N_5139);
nand U7538 (N_7538,N_4013,N_5293);
or U7539 (N_7539,N_5471,N_4182);
nand U7540 (N_7540,N_5942,N_4596);
or U7541 (N_7541,N_4876,N_5322);
nand U7542 (N_7542,N_5326,N_4895);
nand U7543 (N_7543,N_4916,N_4677);
nor U7544 (N_7544,N_5658,N_4297);
and U7545 (N_7545,N_4269,N_5165);
or U7546 (N_7546,N_5695,N_4927);
nor U7547 (N_7547,N_4867,N_5182);
nand U7548 (N_7548,N_4948,N_4147);
nand U7549 (N_7549,N_4198,N_4332);
nor U7550 (N_7550,N_5296,N_4837);
and U7551 (N_7551,N_5842,N_4745);
nand U7552 (N_7552,N_5995,N_4607);
nor U7553 (N_7553,N_5511,N_4846);
nand U7554 (N_7554,N_5601,N_4049);
nand U7555 (N_7555,N_4633,N_4709);
nor U7556 (N_7556,N_5590,N_5382);
nor U7557 (N_7557,N_4211,N_5157);
nand U7558 (N_7558,N_5703,N_4288);
and U7559 (N_7559,N_4324,N_4233);
or U7560 (N_7560,N_4784,N_5951);
nor U7561 (N_7561,N_5493,N_4348);
or U7562 (N_7562,N_5437,N_4756);
and U7563 (N_7563,N_4676,N_4348);
nor U7564 (N_7564,N_5079,N_4863);
or U7565 (N_7565,N_4368,N_5381);
nand U7566 (N_7566,N_4969,N_5327);
or U7567 (N_7567,N_4249,N_5880);
nand U7568 (N_7568,N_4334,N_4275);
and U7569 (N_7569,N_5934,N_5516);
nor U7570 (N_7570,N_4141,N_4513);
and U7571 (N_7571,N_4012,N_4602);
or U7572 (N_7572,N_5069,N_4299);
and U7573 (N_7573,N_5131,N_4945);
nand U7574 (N_7574,N_4369,N_4758);
nand U7575 (N_7575,N_5903,N_4979);
and U7576 (N_7576,N_4806,N_5573);
nor U7577 (N_7577,N_5795,N_4950);
and U7578 (N_7578,N_4717,N_5291);
nand U7579 (N_7579,N_5728,N_4830);
and U7580 (N_7580,N_5686,N_5481);
or U7581 (N_7581,N_5273,N_4133);
or U7582 (N_7582,N_5725,N_4667);
nand U7583 (N_7583,N_4349,N_4982);
and U7584 (N_7584,N_5407,N_5150);
or U7585 (N_7585,N_5750,N_4401);
nand U7586 (N_7586,N_5381,N_5829);
or U7587 (N_7587,N_4778,N_4081);
or U7588 (N_7588,N_4059,N_4330);
nand U7589 (N_7589,N_4540,N_4829);
and U7590 (N_7590,N_5664,N_5403);
and U7591 (N_7591,N_5808,N_5368);
nand U7592 (N_7592,N_4486,N_5077);
nand U7593 (N_7593,N_4800,N_4945);
and U7594 (N_7594,N_5741,N_5853);
nor U7595 (N_7595,N_4384,N_4350);
and U7596 (N_7596,N_5026,N_5018);
and U7597 (N_7597,N_5860,N_4367);
xnor U7598 (N_7598,N_4479,N_5793);
or U7599 (N_7599,N_4061,N_5338);
nand U7600 (N_7600,N_5140,N_5299);
nor U7601 (N_7601,N_4182,N_5167);
and U7602 (N_7602,N_4131,N_4867);
and U7603 (N_7603,N_4776,N_4768);
nor U7604 (N_7604,N_4328,N_4935);
or U7605 (N_7605,N_4130,N_5934);
and U7606 (N_7606,N_5076,N_5816);
nor U7607 (N_7607,N_5393,N_5722);
nor U7608 (N_7608,N_5305,N_4653);
nor U7609 (N_7609,N_5181,N_5595);
nor U7610 (N_7610,N_4865,N_4599);
and U7611 (N_7611,N_5364,N_4794);
nand U7612 (N_7612,N_5650,N_4486);
nand U7613 (N_7613,N_5510,N_4225);
or U7614 (N_7614,N_4025,N_5346);
nor U7615 (N_7615,N_4460,N_5009);
nor U7616 (N_7616,N_4120,N_4094);
nor U7617 (N_7617,N_4917,N_4076);
nand U7618 (N_7618,N_5398,N_4574);
nand U7619 (N_7619,N_5800,N_4445);
nand U7620 (N_7620,N_5237,N_4333);
and U7621 (N_7621,N_5078,N_5310);
nand U7622 (N_7622,N_5739,N_5095);
or U7623 (N_7623,N_4942,N_5512);
nor U7624 (N_7624,N_4498,N_5887);
nor U7625 (N_7625,N_5518,N_4230);
and U7626 (N_7626,N_4613,N_4760);
or U7627 (N_7627,N_5815,N_5613);
nor U7628 (N_7628,N_4772,N_5387);
or U7629 (N_7629,N_4147,N_5177);
nor U7630 (N_7630,N_4546,N_5822);
and U7631 (N_7631,N_5273,N_4365);
nor U7632 (N_7632,N_5594,N_4437);
and U7633 (N_7633,N_4756,N_4842);
nand U7634 (N_7634,N_4134,N_5902);
and U7635 (N_7635,N_5968,N_4625);
nand U7636 (N_7636,N_4343,N_5700);
nand U7637 (N_7637,N_5017,N_4503);
or U7638 (N_7638,N_4266,N_5694);
and U7639 (N_7639,N_4417,N_5000);
nand U7640 (N_7640,N_5490,N_5396);
and U7641 (N_7641,N_4374,N_4353);
or U7642 (N_7642,N_4462,N_4104);
or U7643 (N_7643,N_5310,N_5646);
nand U7644 (N_7644,N_4551,N_4496);
or U7645 (N_7645,N_5688,N_5077);
nand U7646 (N_7646,N_5387,N_4874);
nor U7647 (N_7647,N_4817,N_5721);
and U7648 (N_7648,N_4200,N_4421);
or U7649 (N_7649,N_4458,N_5119);
nor U7650 (N_7650,N_4437,N_4570);
and U7651 (N_7651,N_4464,N_4952);
and U7652 (N_7652,N_5363,N_4455);
or U7653 (N_7653,N_4226,N_4690);
nor U7654 (N_7654,N_4847,N_4940);
nor U7655 (N_7655,N_4422,N_5192);
nor U7656 (N_7656,N_5801,N_4938);
nand U7657 (N_7657,N_4912,N_4821);
nor U7658 (N_7658,N_5941,N_5095);
nand U7659 (N_7659,N_5795,N_5622);
nor U7660 (N_7660,N_4769,N_5342);
nand U7661 (N_7661,N_5243,N_4479);
nor U7662 (N_7662,N_5465,N_5039);
and U7663 (N_7663,N_5432,N_5198);
nor U7664 (N_7664,N_4950,N_5473);
nand U7665 (N_7665,N_5477,N_4080);
nor U7666 (N_7666,N_5195,N_4908);
or U7667 (N_7667,N_5826,N_4083);
and U7668 (N_7668,N_4272,N_5475);
nand U7669 (N_7669,N_5105,N_5070);
nor U7670 (N_7670,N_5291,N_4780);
or U7671 (N_7671,N_5440,N_4505);
and U7672 (N_7672,N_4203,N_5267);
and U7673 (N_7673,N_5621,N_4899);
xor U7674 (N_7674,N_5606,N_4453);
nand U7675 (N_7675,N_5590,N_5989);
nand U7676 (N_7676,N_5318,N_4889);
nor U7677 (N_7677,N_4064,N_5512);
or U7678 (N_7678,N_5932,N_5077);
nand U7679 (N_7679,N_5462,N_5542);
nand U7680 (N_7680,N_4343,N_4757);
or U7681 (N_7681,N_5147,N_4448);
and U7682 (N_7682,N_5997,N_4578);
nor U7683 (N_7683,N_4928,N_4205);
or U7684 (N_7684,N_4940,N_5042);
nand U7685 (N_7685,N_5988,N_5034);
nand U7686 (N_7686,N_4383,N_4885);
nor U7687 (N_7687,N_5607,N_4236);
or U7688 (N_7688,N_4376,N_5902);
or U7689 (N_7689,N_5216,N_5295);
xnor U7690 (N_7690,N_4237,N_4997);
nand U7691 (N_7691,N_5855,N_4802);
and U7692 (N_7692,N_5808,N_5476);
and U7693 (N_7693,N_4868,N_4794);
and U7694 (N_7694,N_5116,N_5781);
or U7695 (N_7695,N_5530,N_4494);
nand U7696 (N_7696,N_4333,N_4565);
nor U7697 (N_7697,N_4848,N_5736);
nand U7698 (N_7698,N_4548,N_5207);
nor U7699 (N_7699,N_4683,N_4862);
nand U7700 (N_7700,N_5107,N_5689);
nand U7701 (N_7701,N_4290,N_5899);
or U7702 (N_7702,N_4867,N_4234);
and U7703 (N_7703,N_4402,N_4863);
or U7704 (N_7704,N_4864,N_5401);
nand U7705 (N_7705,N_5167,N_5489);
nand U7706 (N_7706,N_5551,N_5706);
or U7707 (N_7707,N_4970,N_5263);
and U7708 (N_7708,N_5246,N_5610);
nand U7709 (N_7709,N_4527,N_4719);
nand U7710 (N_7710,N_5917,N_5820);
nand U7711 (N_7711,N_4681,N_4890);
nor U7712 (N_7712,N_4114,N_5496);
nor U7713 (N_7713,N_4697,N_4490);
and U7714 (N_7714,N_5741,N_4711);
nand U7715 (N_7715,N_5618,N_5268);
or U7716 (N_7716,N_5035,N_5522);
nand U7717 (N_7717,N_5449,N_4509);
nand U7718 (N_7718,N_5705,N_5302);
nand U7719 (N_7719,N_5514,N_5988);
and U7720 (N_7720,N_5806,N_4502);
and U7721 (N_7721,N_5818,N_5861);
and U7722 (N_7722,N_5046,N_4744);
nor U7723 (N_7723,N_4628,N_5905);
nand U7724 (N_7724,N_5885,N_5903);
and U7725 (N_7725,N_5230,N_5630);
nor U7726 (N_7726,N_5687,N_5480);
nand U7727 (N_7727,N_4696,N_4871);
xnor U7728 (N_7728,N_4854,N_4678);
and U7729 (N_7729,N_4547,N_4055);
nor U7730 (N_7730,N_5999,N_5534);
nor U7731 (N_7731,N_4173,N_5023);
nand U7732 (N_7732,N_5518,N_5300);
nand U7733 (N_7733,N_5559,N_4303);
or U7734 (N_7734,N_5369,N_5947);
or U7735 (N_7735,N_4235,N_5735);
nand U7736 (N_7736,N_5090,N_4495);
or U7737 (N_7737,N_4447,N_4118);
nor U7738 (N_7738,N_4610,N_5793);
nor U7739 (N_7739,N_5469,N_5338);
nand U7740 (N_7740,N_5286,N_5433);
and U7741 (N_7741,N_5060,N_5554);
and U7742 (N_7742,N_5958,N_5488);
nor U7743 (N_7743,N_5808,N_5129);
and U7744 (N_7744,N_4605,N_5404);
nor U7745 (N_7745,N_4546,N_5151);
and U7746 (N_7746,N_4668,N_5337);
nor U7747 (N_7747,N_5702,N_4628);
nand U7748 (N_7748,N_4925,N_5379);
and U7749 (N_7749,N_4866,N_4706);
nor U7750 (N_7750,N_4785,N_4045);
or U7751 (N_7751,N_5094,N_4572);
nand U7752 (N_7752,N_4134,N_4430);
nor U7753 (N_7753,N_4844,N_4933);
nand U7754 (N_7754,N_4325,N_4973);
nand U7755 (N_7755,N_5900,N_4587);
and U7756 (N_7756,N_4289,N_4292);
nand U7757 (N_7757,N_4185,N_4651);
and U7758 (N_7758,N_4869,N_4526);
nor U7759 (N_7759,N_4198,N_5985);
nor U7760 (N_7760,N_5711,N_4988);
nand U7761 (N_7761,N_5718,N_4254);
or U7762 (N_7762,N_5708,N_4895);
and U7763 (N_7763,N_4890,N_5665);
or U7764 (N_7764,N_5919,N_5203);
nand U7765 (N_7765,N_4935,N_4652);
nor U7766 (N_7766,N_4701,N_4539);
or U7767 (N_7767,N_4014,N_4112);
and U7768 (N_7768,N_5920,N_4982);
nor U7769 (N_7769,N_5939,N_5903);
or U7770 (N_7770,N_4734,N_4811);
nor U7771 (N_7771,N_4759,N_4587);
or U7772 (N_7772,N_4077,N_4755);
and U7773 (N_7773,N_4709,N_5060);
or U7774 (N_7774,N_4512,N_5450);
nand U7775 (N_7775,N_4665,N_4152);
and U7776 (N_7776,N_5525,N_4845);
or U7777 (N_7777,N_5903,N_4015);
or U7778 (N_7778,N_5879,N_5198);
nand U7779 (N_7779,N_5913,N_5191);
nand U7780 (N_7780,N_4637,N_4712);
or U7781 (N_7781,N_4562,N_4666);
and U7782 (N_7782,N_4859,N_5805);
and U7783 (N_7783,N_5189,N_5395);
nand U7784 (N_7784,N_4096,N_4308);
nand U7785 (N_7785,N_5661,N_5555);
nand U7786 (N_7786,N_4845,N_5459);
and U7787 (N_7787,N_5949,N_4788);
and U7788 (N_7788,N_5253,N_4900);
nor U7789 (N_7789,N_4566,N_4326);
and U7790 (N_7790,N_5648,N_5949);
and U7791 (N_7791,N_4451,N_4823);
and U7792 (N_7792,N_4763,N_4908);
and U7793 (N_7793,N_5814,N_5471);
or U7794 (N_7794,N_4210,N_4686);
nand U7795 (N_7795,N_4243,N_5727);
or U7796 (N_7796,N_4429,N_4228);
nor U7797 (N_7797,N_5316,N_4756);
nor U7798 (N_7798,N_5241,N_5308);
nand U7799 (N_7799,N_5828,N_4184);
nor U7800 (N_7800,N_5295,N_5604);
xnor U7801 (N_7801,N_4165,N_5268);
or U7802 (N_7802,N_4889,N_5866);
nand U7803 (N_7803,N_5506,N_5437);
and U7804 (N_7804,N_5785,N_5163);
and U7805 (N_7805,N_4405,N_4582);
nor U7806 (N_7806,N_4800,N_4490);
nor U7807 (N_7807,N_4338,N_5560);
or U7808 (N_7808,N_5892,N_4969);
nand U7809 (N_7809,N_4231,N_4247);
nor U7810 (N_7810,N_4409,N_5669);
nand U7811 (N_7811,N_4472,N_5146);
nand U7812 (N_7812,N_4723,N_5515);
or U7813 (N_7813,N_4597,N_5914);
nand U7814 (N_7814,N_5071,N_5850);
nor U7815 (N_7815,N_5265,N_4842);
nand U7816 (N_7816,N_5630,N_4587);
or U7817 (N_7817,N_5214,N_5170);
nand U7818 (N_7818,N_5561,N_5690);
or U7819 (N_7819,N_5267,N_4999);
and U7820 (N_7820,N_4279,N_4507);
nand U7821 (N_7821,N_4722,N_4422);
or U7822 (N_7822,N_5718,N_4099);
and U7823 (N_7823,N_4889,N_5352);
nand U7824 (N_7824,N_5897,N_4654);
nand U7825 (N_7825,N_5303,N_5625);
nand U7826 (N_7826,N_4971,N_5656);
or U7827 (N_7827,N_4317,N_4369);
nand U7828 (N_7828,N_5513,N_4473);
xor U7829 (N_7829,N_5012,N_4221);
nor U7830 (N_7830,N_5152,N_4421);
nor U7831 (N_7831,N_5371,N_5164);
nand U7832 (N_7832,N_4062,N_5077);
or U7833 (N_7833,N_5327,N_5355);
nand U7834 (N_7834,N_5459,N_4862);
or U7835 (N_7835,N_5471,N_4394);
nor U7836 (N_7836,N_5038,N_4616);
nor U7837 (N_7837,N_4845,N_5711);
and U7838 (N_7838,N_4853,N_5138);
nor U7839 (N_7839,N_4689,N_5879);
nand U7840 (N_7840,N_5678,N_4585);
nand U7841 (N_7841,N_5925,N_4390);
nand U7842 (N_7842,N_5779,N_4349);
and U7843 (N_7843,N_5354,N_4243);
nor U7844 (N_7844,N_4628,N_5238);
and U7845 (N_7845,N_4075,N_4759);
and U7846 (N_7846,N_4769,N_4210);
or U7847 (N_7847,N_4442,N_5109);
nor U7848 (N_7848,N_4209,N_4079);
nand U7849 (N_7849,N_4586,N_4312);
and U7850 (N_7850,N_5588,N_4211);
or U7851 (N_7851,N_5241,N_4669);
nor U7852 (N_7852,N_4368,N_4881);
and U7853 (N_7853,N_4681,N_4290);
and U7854 (N_7854,N_4672,N_5650);
nand U7855 (N_7855,N_5613,N_4694);
nand U7856 (N_7856,N_5187,N_5848);
or U7857 (N_7857,N_5635,N_4387);
nor U7858 (N_7858,N_5338,N_4466);
nor U7859 (N_7859,N_5346,N_4716);
nand U7860 (N_7860,N_5849,N_4339);
and U7861 (N_7861,N_5418,N_5283);
nor U7862 (N_7862,N_4534,N_4011);
and U7863 (N_7863,N_4102,N_5903);
nand U7864 (N_7864,N_5019,N_4076);
nand U7865 (N_7865,N_5079,N_5430);
or U7866 (N_7866,N_4152,N_4485);
or U7867 (N_7867,N_5241,N_4692);
nor U7868 (N_7868,N_5872,N_4662);
or U7869 (N_7869,N_4917,N_4252);
or U7870 (N_7870,N_5156,N_4235);
and U7871 (N_7871,N_5675,N_5100);
nor U7872 (N_7872,N_4910,N_4147);
nor U7873 (N_7873,N_4549,N_5248);
and U7874 (N_7874,N_5038,N_5781);
and U7875 (N_7875,N_4787,N_5229);
nor U7876 (N_7876,N_5188,N_5583);
nor U7877 (N_7877,N_4487,N_5851);
nand U7878 (N_7878,N_4728,N_5737);
nor U7879 (N_7879,N_5789,N_5844);
nand U7880 (N_7880,N_4711,N_5023);
nand U7881 (N_7881,N_5783,N_5674);
nand U7882 (N_7882,N_5343,N_4442);
nor U7883 (N_7883,N_4089,N_4153);
or U7884 (N_7884,N_5201,N_5913);
nand U7885 (N_7885,N_4519,N_4329);
nand U7886 (N_7886,N_4518,N_5374);
nand U7887 (N_7887,N_4503,N_4518);
nand U7888 (N_7888,N_5740,N_5749);
or U7889 (N_7889,N_5029,N_4665);
nor U7890 (N_7890,N_4431,N_5314);
and U7891 (N_7891,N_5992,N_4666);
nand U7892 (N_7892,N_5750,N_5073);
nor U7893 (N_7893,N_4963,N_4533);
or U7894 (N_7894,N_4616,N_5365);
or U7895 (N_7895,N_4746,N_5680);
and U7896 (N_7896,N_5463,N_4238);
nor U7897 (N_7897,N_5827,N_4572);
and U7898 (N_7898,N_4881,N_5391);
and U7899 (N_7899,N_5930,N_4745);
nor U7900 (N_7900,N_4460,N_5151);
nand U7901 (N_7901,N_5506,N_5079);
and U7902 (N_7902,N_5944,N_5282);
nor U7903 (N_7903,N_5274,N_4762);
nor U7904 (N_7904,N_4277,N_5920);
and U7905 (N_7905,N_5418,N_4221);
nand U7906 (N_7906,N_4622,N_4081);
nand U7907 (N_7907,N_5658,N_5897);
and U7908 (N_7908,N_5571,N_5458);
nor U7909 (N_7909,N_4831,N_4047);
nand U7910 (N_7910,N_4694,N_4024);
xor U7911 (N_7911,N_4962,N_4122);
nor U7912 (N_7912,N_4713,N_4256);
nor U7913 (N_7913,N_4689,N_5123);
and U7914 (N_7914,N_5526,N_5679);
or U7915 (N_7915,N_4108,N_5518);
or U7916 (N_7916,N_4682,N_5423);
nand U7917 (N_7917,N_5934,N_5094);
nor U7918 (N_7918,N_5177,N_4365);
nand U7919 (N_7919,N_4305,N_5257);
nor U7920 (N_7920,N_5747,N_4750);
or U7921 (N_7921,N_4512,N_5242);
or U7922 (N_7922,N_4957,N_4368);
nor U7923 (N_7923,N_5002,N_4433);
and U7924 (N_7924,N_4372,N_4135);
or U7925 (N_7925,N_4163,N_4283);
nand U7926 (N_7926,N_4423,N_4446);
or U7927 (N_7927,N_4729,N_5058);
nand U7928 (N_7928,N_4331,N_5308);
and U7929 (N_7929,N_5747,N_4678);
nand U7930 (N_7930,N_5286,N_4742);
nand U7931 (N_7931,N_5416,N_4128);
nand U7932 (N_7932,N_5776,N_4533);
nand U7933 (N_7933,N_4698,N_4349);
nor U7934 (N_7934,N_4289,N_4324);
and U7935 (N_7935,N_5777,N_5649);
and U7936 (N_7936,N_5101,N_4815);
and U7937 (N_7937,N_4137,N_4737);
nor U7938 (N_7938,N_5929,N_5912);
nor U7939 (N_7939,N_4172,N_5837);
and U7940 (N_7940,N_5569,N_5107);
nor U7941 (N_7941,N_5950,N_5730);
and U7942 (N_7942,N_4059,N_5189);
nand U7943 (N_7943,N_5719,N_5121);
and U7944 (N_7944,N_5176,N_5209);
xnor U7945 (N_7945,N_4387,N_5761);
nor U7946 (N_7946,N_5751,N_5242);
nor U7947 (N_7947,N_5506,N_4474);
nand U7948 (N_7948,N_5436,N_5980);
or U7949 (N_7949,N_4528,N_4757);
xor U7950 (N_7950,N_5057,N_5186);
and U7951 (N_7951,N_4866,N_5267);
nand U7952 (N_7952,N_5701,N_4501);
or U7953 (N_7953,N_5832,N_5841);
nor U7954 (N_7954,N_4771,N_5653);
nand U7955 (N_7955,N_4734,N_5381);
and U7956 (N_7956,N_4922,N_5673);
and U7957 (N_7957,N_4397,N_5181);
nand U7958 (N_7958,N_4810,N_4470);
and U7959 (N_7959,N_4084,N_4842);
or U7960 (N_7960,N_4424,N_5932);
and U7961 (N_7961,N_4200,N_5183);
nor U7962 (N_7962,N_4795,N_4248);
or U7963 (N_7963,N_4974,N_4787);
and U7964 (N_7964,N_4516,N_5928);
or U7965 (N_7965,N_5863,N_4372);
nand U7966 (N_7966,N_4022,N_5038);
and U7967 (N_7967,N_4609,N_4573);
nand U7968 (N_7968,N_4966,N_4089);
or U7969 (N_7969,N_4984,N_4954);
nor U7970 (N_7970,N_4756,N_5897);
nor U7971 (N_7971,N_4057,N_5514);
and U7972 (N_7972,N_5216,N_5643);
nand U7973 (N_7973,N_5115,N_5728);
nor U7974 (N_7974,N_5721,N_4344);
nand U7975 (N_7975,N_5474,N_5330);
and U7976 (N_7976,N_4736,N_5601);
or U7977 (N_7977,N_5070,N_4658);
or U7978 (N_7978,N_5110,N_4606);
nand U7979 (N_7979,N_5132,N_5694);
nor U7980 (N_7980,N_4258,N_4740);
nand U7981 (N_7981,N_4336,N_5481);
nor U7982 (N_7982,N_5884,N_5669);
nor U7983 (N_7983,N_5902,N_5168);
or U7984 (N_7984,N_5311,N_5301);
or U7985 (N_7985,N_5029,N_5886);
and U7986 (N_7986,N_5979,N_4074);
and U7987 (N_7987,N_4086,N_5285);
nor U7988 (N_7988,N_4113,N_4712);
nand U7989 (N_7989,N_5708,N_5424);
nand U7990 (N_7990,N_5671,N_4615);
and U7991 (N_7991,N_5785,N_5043);
and U7992 (N_7992,N_5193,N_4747);
nand U7993 (N_7993,N_4904,N_5488);
and U7994 (N_7994,N_5644,N_4034);
nor U7995 (N_7995,N_5725,N_4006);
nor U7996 (N_7996,N_5982,N_5111);
or U7997 (N_7997,N_4587,N_4296);
nand U7998 (N_7998,N_5045,N_5552);
nor U7999 (N_7999,N_5142,N_5503);
or U8000 (N_8000,N_6851,N_7021);
nor U8001 (N_8001,N_6932,N_6833);
and U8002 (N_8002,N_7098,N_6868);
or U8003 (N_8003,N_6338,N_6030);
and U8004 (N_8004,N_7140,N_7097);
and U8005 (N_8005,N_7378,N_6057);
or U8006 (N_8006,N_6545,N_6707);
nor U8007 (N_8007,N_6308,N_6233);
or U8008 (N_8008,N_7786,N_7458);
and U8009 (N_8009,N_7347,N_6579);
nand U8010 (N_8010,N_6509,N_6417);
or U8011 (N_8011,N_6746,N_6780);
or U8012 (N_8012,N_6538,N_7778);
nand U8013 (N_8013,N_6229,N_7246);
or U8014 (N_8014,N_7586,N_7269);
nand U8015 (N_8015,N_7732,N_7627);
nor U8016 (N_8016,N_7951,N_6255);
nand U8017 (N_8017,N_7884,N_7689);
nand U8018 (N_8018,N_6155,N_6343);
and U8019 (N_8019,N_6477,N_7820);
or U8020 (N_8020,N_7675,N_6305);
nand U8021 (N_8021,N_6906,N_7795);
or U8022 (N_8022,N_6345,N_6694);
or U8023 (N_8023,N_6239,N_7183);
or U8024 (N_8024,N_6668,N_6626);
or U8025 (N_8025,N_7741,N_6216);
xor U8026 (N_8026,N_7197,N_7060);
nand U8027 (N_8027,N_6635,N_6652);
nand U8028 (N_8028,N_6681,N_7574);
and U8029 (N_8029,N_7931,N_6376);
or U8030 (N_8030,N_6195,N_6601);
or U8031 (N_8031,N_7075,N_7946);
nor U8032 (N_8032,N_7356,N_6574);
nand U8033 (N_8033,N_7108,N_7463);
nor U8034 (N_8034,N_6299,N_7350);
nor U8035 (N_8035,N_6341,N_7735);
nand U8036 (N_8036,N_6528,N_7855);
or U8037 (N_8037,N_7189,N_6661);
nor U8038 (N_8038,N_7917,N_6420);
nor U8039 (N_8039,N_7312,N_7056);
nor U8040 (N_8040,N_7083,N_6535);
or U8041 (N_8041,N_7986,N_7292);
or U8042 (N_8042,N_6953,N_7699);
nand U8043 (N_8043,N_6859,N_6739);
nand U8044 (N_8044,N_7006,N_6867);
or U8045 (N_8045,N_7327,N_7670);
nand U8046 (N_8046,N_6440,N_6560);
and U8047 (N_8047,N_6736,N_6543);
and U8048 (N_8048,N_7115,N_6261);
nand U8049 (N_8049,N_7760,N_7817);
and U8050 (N_8050,N_6294,N_6823);
nand U8051 (N_8051,N_6516,N_6609);
or U8052 (N_8052,N_7811,N_7828);
or U8053 (N_8053,N_7572,N_6174);
and U8054 (N_8054,N_6905,N_6331);
nor U8055 (N_8055,N_7095,N_7185);
nor U8056 (N_8056,N_6835,N_7927);
and U8057 (N_8057,N_6593,N_7859);
nor U8058 (N_8058,N_6242,N_6200);
or U8059 (N_8059,N_6252,N_6850);
and U8060 (N_8060,N_6900,N_7219);
nor U8061 (N_8061,N_7159,N_7646);
nor U8062 (N_8062,N_7093,N_6041);
nor U8063 (N_8063,N_7211,N_7285);
nor U8064 (N_8064,N_6045,N_7110);
nand U8065 (N_8065,N_7294,N_6813);
nand U8066 (N_8066,N_7141,N_6575);
nor U8067 (N_8067,N_6125,N_7215);
nand U8068 (N_8068,N_6256,N_7370);
nand U8069 (N_8069,N_7477,N_7125);
nor U8070 (N_8070,N_7540,N_7372);
or U8071 (N_8071,N_7615,N_6323);
nor U8072 (N_8072,N_7612,N_7174);
and U8073 (N_8073,N_7799,N_6191);
and U8074 (N_8074,N_6260,N_6066);
or U8075 (N_8075,N_6334,N_6017);
nand U8076 (N_8076,N_7429,N_7309);
or U8077 (N_8077,N_6327,N_6786);
nor U8078 (N_8078,N_7013,N_7548);
or U8079 (N_8079,N_6837,N_7385);
nor U8080 (N_8080,N_7239,N_6364);
nand U8081 (N_8081,N_6686,N_6268);
and U8082 (N_8082,N_7445,N_6840);
and U8083 (N_8083,N_6978,N_7713);
xor U8084 (N_8084,N_7149,N_7263);
nor U8085 (N_8085,N_7768,N_6358);
nor U8086 (N_8086,N_6482,N_7284);
and U8087 (N_8087,N_7777,N_7161);
and U8088 (N_8088,N_7256,N_7692);
nor U8089 (N_8089,N_6505,N_6107);
and U8090 (N_8090,N_7121,N_7867);
nand U8091 (N_8091,N_7084,N_7305);
nor U8092 (N_8092,N_7621,N_6199);
nand U8093 (N_8093,N_6075,N_6036);
and U8094 (N_8094,N_7836,N_6640);
and U8095 (N_8095,N_7672,N_7575);
nor U8096 (N_8096,N_7600,N_6103);
nand U8097 (N_8097,N_7418,N_6437);
or U8098 (N_8098,N_6092,N_7900);
nand U8099 (N_8099,N_6207,N_7489);
or U8100 (N_8100,N_6211,N_6181);
nor U8101 (N_8101,N_6682,N_6457);
and U8102 (N_8102,N_6597,N_7532);
and U8103 (N_8103,N_7396,N_7935);
nor U8104 (N_8104,N_6144,N_6785);
nand U8105 (N_8105,N_6462,N_7224);
and U8106 (N_8106,N_7776,N_7187);
nor U8107 (N_8107,N_7415,N_7259);
or U8108 (N_8108,N_6806,N_7071);
or U8109 (N_8109,N_7346,N_7381);
or U8110 (N_8110,N_7339,N_6287);
and U8111 (N_8111,N_7580,N_6012);
or U8112 (N_8112,N_7065,N_7365);
and U8113 (N_8113,N_6800,N_6855);
nand U8114 (N_8114,N_6361,N_7780);
nand U8115 (N_8115,N_7980,N_7503);
nor U8116 (N_8116,N_7452,N_6767);
and U8117 (N_8117,N_6168,N_6866);
nand U8118 (N_8118,N_6600,N_7920);
or U8119 (N_8119,N_6546,N_7020);
nand U8120 (N_8120,N_7593,N_6554);
or U8121 (N_8121,N_7897,N_7667);
or U8122 (N_8122,N_7969,N_7684);
nand U8123 (N_8123,N_6756,N_7922);
and U8124 (N_8124,N_6071,N_7230);
nor U8125 (N_8125,N_6020,N_6858);
or U8126 (N_8126,N_7974,N_6830);
and U8127 (N_8127,N_6647,N_6754);
and U8128 (N_8128,N_7911,N_6100);
or U8129 (N_8129,N_6377,N_7085);
and U8130 (N_8130,N_7873,N_6826);
or U8131 (N_8131,N_6770,N_7077);
nand U8132 (N_8132,N_6413,N_6108);
nor U8133 (N_8133,N_6824,N_7886);
nand U8134 (N_8134,N_6118,N_6908);
or U8135 (N_8135,N_6102,N_7982);
and U8136 (N_8136,N_7734,N_6023);
and U8137 (N_8137,N_6086,N_7634);
nand U8138 (N_8138,N_7529,N_6662);
or U8139 (N_8139,N_7571,N_7526);
or U8140 (N_8140,N_6585,N_6675);
nor U8141 (N_8141,N_7119,N_6316);
nand U8142 (N_8142,N_6992,N_6499);
or U8143 (N_8143,N_6390,N_7374);
and U8144 (N_8144,N_7271,N_7521);
nor U8145 (N_8145,N_6997,N_6192);
and U8146 (N_8146,N_6180,N_6067);
nand U8147 (N_8147,N_7552,N_7959);
or U8148 (N_8148,N_6497,N_6881);
nand U8149 (N_8149,N_7547,N_7644);
nand U8150 (N_8150,N_7724,N_6958);
or U8151 (N_8151,N_7983,N_7858);
or U8152 (N_8152,N_7072,N_7279);
nor U8153 (N_8153,N_7422,N_7751);
nand U8154 (N_8154,N_7376,N_7943);
or U8155 (N_8155,N_7104,N_6741);
nand U8156 (N_8156,N_7938,N_6816);
nand U8157 (N_8157,N_6183,N_6533);
nand U8158 (N_8158,N_6949,N_6653);
nand U8159 (N_8159,N_6524,N_6379);
and U8160 (N_8160,N_7049,N_7382);
or U8161 (N_8161,N_7486,N_6044);
nor U8162 (N_8162,N_7516,N_7332);
and U8163 (N_8163,N_7304,N_7543);
nand U8164 (N_8164,N_7490,N_7815);
nor U8165 (N_8165,N_6368,N_6553);
and U8166 (N_8166,N_6649,N_6454);
or U8167 (N_8167,N_6265,N_6356);
or U8168 (N_8168,N_7460,N_7630);
or U8169 (N_8169,N_7390,N_6937);
nand U8170 (N_8170,N_7447,N_6219);
or U8171 (N_8171,N_7813,N_7905);
or U8172 (N_8172,N_7524,N_6853);
nor U8173 (N_8173,N_6808,N_7923);
and U8174 (N_8174,N_6088,N_7725);
nand U8175 (N_8175,N_7267,N_6400);
nor U8176 (N_8176,N_7078,N_7875);
and U8177 (N_8177,N_6349,N_6981);
xnor U8178 (N_8178,N_7178,N_7403);
and U8179 (N_8179,N_6470,N_7832);
and U8180 (N_8180,N_6369,N_7235);
and U8181 (N_8181,N_6373,N_6724);
nand U8182 (N_8182,N_7970,N_6685);
nand U8183 (N_8183,N_7156,N_6383);
nor U8184 (N_8184,N_7377,N_7879);
xnor U8185 (N_8185,N_6014,N_6002);
and U8186 (N_8186,N_7054,N_6494);
nor U8187 (N_8187,N_7479,N_6674);
and U8188 (N_8188,N_6312,N_7352);
nand U8189 (N_8189,N_7788,N_7413);
nor U8190 (N_8190,N_6515,N_6719);
nand U8191 (N_8191,N_6438,N_7299);
or U8192 (N_8192,N_6781,N_6970);
and U8193 (N_8193,N_6371,N_7744);
and U8194 (N_8194,N_7929,N_7889);
nand U8195 (N_8195,N_7947,N_6104);
nand U8196 (N_8196,N_6692,N_7694);
nand U8197 (N_8197,N_6946,N_6650);
nand U8198 (N_8198,N_6033,N_6884);
or U8199 (N_8199,N_6160,N_6606);
nor U8200 (N_8200,N_7220,N_7375);
and U8201 (N_8201,N_6988,N_7202);
and U8202 (N_8202,N_7433,N_6836);
or U8203 (N_8203,N_7248,N_7782);
or U8204 (N_8204,N_6977,N_6424);
nor U8205 (N_8205,N_6995,N_7633);
or U8206 (N_8206,N_6306,N_7669);
nor U8207 (N_8207,N_6895,N_6274);
or U8208 (N_8208,N_6520,N_6202);
nor U8209 (N_8209,N_6101,N_6415);
nand U8210 (N_8210,N_7565,N_6936);
and U8211 (N_8211,N_7283,N_7919);
nand U8212 (N_8212,N_6121,N_6656);
and U8213 (N_8213,N_7373,N_7293);
nor U8214 (N_8214,N_7229,N_6493);
or U8215 (N_8215,N_7993,N_6339);
or U8216 (N_8216,N_7026,N_7467);
nand U8217 (N_8217,N_6196,N_7620);
or U8218 (N_8218,N_7209,N_6514);
and U8219 (N_8219,N_6963,N_7231);
or U8220 (N_8220,N_7175,N_7846);
and U8221 (N_8221,N_6009,N_6464);
and U8222 (N_8222,N_6580,N_6564);
or U8223 (N_8223,N_7155,N_7142);
nand U8224 (N_8224,N_7310,N_7136);
nor U8225 (N_8225,N_6070,N_7144);
nor U8226 (N_8226,N_6698,N_7029);
or U8227 (N_8227,N_6729,N_7818);
and U8228 (N_8228,N_7740,N_7924);
nor U8229 (N_8229,N_7994,N_7590);
or U8230 (N_8230,N_7150,N_7186);
or U8231 (N_8231,N_7932,N_7465);
and U8232 (N_8232,N_7344,N_7319);
or U8233 (N_8233,N_7316,N_7254);
nor U8234 (N_8234,N_6603,N_6592);
nor U8235 (N_8235,N_6938,N_7213);
and U8236 (N_8236,N_7567,N_7647);
nor U8237 (N_8237,N_7916,N_6904);
and U8238 (N_8238,N_6034,N_7910);
nor U8239 (N_8239,N_7861,N_7443);
nor U8240 (N_8240,N_7693,N_7325);
or U8241 (N_8241,N_6458,N_6056);
nor U8242 (N_8242,N_7308,N_6311);
nor U8243 (N_8243,N_6720,N_7088);
nand U8244 (N_8244,N_6511,N_6631);
and U8245 (N_8245,N_6394,N_6414);
nor U8246 (N_8246,N_6248,N_6847);
and U8247 (N_8247,N_6666,N_6975);
nand U8248 (N_8248,N_6636,N_6087);
nand U8249 (N_8249,N_7090,N_7160);
and U8250 (N_8250,N_7587,N_7723);
or U8251 (N_8251,N_6179,N_7157);
nand U8252 (N_8252,N_7240,N_6042);
nand U8253 (N_8253,N_6857,N_6445);
nor U8254 (N_8254,N_6779,N_6957);
nand U8255 (N_8255,N_6024,N_7329);
and U8256 (N_8256,N_6003,N_6139);
nand U8257 (N_8257,N_7466,N_6864);
and U8258 (N_8258,N_7247,N_6004);
and U8259 (N_8259,N_7518,N_7424);
and U8260 (N_8260,N_6271,N_6874);
and U8261 (N_8261,N_6777,N_6621);
and U8262 (N_8262,N_7148,N_7225);
and U8263 (N_8263,N_7000,N_7893);
nor U8264 (N_8264,N_7653,N_6915);
or U8265 (N_8265,N_6796,N_7027);
nand U8266 (N_8266,N_7041,N_6986);
nand U8267 (N_8267,N_7686,N_6098);
nor U8268 (N_8268,N_7985,N_6352);
or U8269 (N_8269,N_6419,N_7704);
or U8270 (N_8270,N_6269,N_6584);
nand U8271 (N_8271,N_6841,N_7454);
nor U8272 (N_8272,N_6022,N_7793);
nor U8273 (N_8273,N_6266,N_7515);
nand U8274 (N_8274,N_7639,N_6049);
nor U8275 (N_8275,N_7996,N_6328);
and U8276 (N_8276,N_7772,N_6644);
nand U8277 (N_8277,N_6116,N_6917);
or U8278 (N_8278,N_6537,N_7362);
and U8279 (N_8279,N_6998,N_6620);
or U8280 (N_8280,N_6093,N_7096);
nor U8281 (N_8281,N_6871,N_7210);
nand U8282 (N_8282,N_6643,N_6709);
xnor U8283 (N_8283,N_7173,N_7908);
nor U8284 (N_8284,N_6130,N_7208);
and U8285 (N_8285,N_6576,N_7816);
nand U8286 (N_8286,N_7641,N_6184);
nor U8287 (N_8287,N_6106,N_6141);
and U8288 (N_8288,N_7555,N_7481);
nor U8289 (N_8289,N_7198,N_6298);
or U8290 (N_8290,N_6629,N_7371);
nand U8291 (N_8291,N_7367,N_7756);
and U8292 (N_8292,N_7257,N_7336);
and U8293 (N_8293,N_6446,N_6406);
nand U8294 (N_8294,N_7031,N_7718);
and U8295 (N_8295,N_6945,N_6138);
and U8296 (N_8296,N_6326,N_7829);
nand U8297 (N_8297,N_6799,N_7169);
nand U8298 (N_8298,N_7509,N_6570);
nand U8299 (N_8299,N_7448,N_7080);
and U8300 (N_8300,N_6916,N_7823);
and U8301 (N_8301,N_6539,N_6562);
nor U8302 (N_8302,N_6190,N_7773);
and U8303 (N_8303,N_7449,N_7895);
or U8304 (N_8304,N_7296,N_6398);
nand U8305 (N_8305,N_7640,N_6865);
or U8306 (N_8306,N_6611,N_7322);
nor U8307 (N_8307,N_6348,N_6828);
nand U8308 (N_8308,N_6987,N_6498);
or U8309 (N_8309,N_7009,N_6583);
and U8310 (N_8310,N_7264,N_7966);
nand U8311 (N_8311,N_6894,N_7888);
nor U8312 (N_8312,N_6966,N_6476);
or U8313 (N_8313,N_6461,N_7514);
or U8314 (N_8314,N_7874,N_6572);
and U8315 (N_8315,N_7674,N_7369);
nor U8316 (N_8316,N_6544,N_7955);
or U8317 (N_8317,N_6877,N_6433);
nor U8318 (N_8318,N_6443,N_7517);
nand U8319 (N_8319,N_6676,N_7255);
and U8320 (N_8320,N_7745,N_7934);
nor U8321 (N_8321,N_7488,N_7082);
and U8322 (N_8322,N_6083,N_6818);
nor U8323 (N_8323,N_7949,N_6503);
or U8324 (N_8324,N_6532,N_6386);
or U8325 (N_8325,N_7392,N_6639);
and U8326 (N_8326,N_6010,N_7722);
nand U8327 (N_8327,N_7482,N_7249);
and U8328 (N_8328,N_6911,N_7663);
or U8329 (N_8329,N_6028,N_7758);
nand U8330 (N_8330,N_7607,N_6885);
or U8331 (N_8331,N_7203,N_6210);
or U8332 (N_8332,N_6689,N_7991);
and U8333 (N_8333,N_7495,N_6693);
and U8334 (N_8334,N_6319,N_6309);
nor U8335 (N_8335,N_6965,N_7005);
nor U8336 (N_8336,N_7783,N_7589);
nand U8337 (N_8337,N_6472,N_7904);
nor U8338 (N_8338,N_6473,N_7266);
or U8339 (N_8339,N_7583,N_6436);
nor U8340 (N_8340,N_7856,N_6401);
and U8341 (N_8341,N_6891,N_7216);
or U8342 (N_8342,N_6185,N_7559);
nand U8343 (N_8343,N_6096,N_7290);
or U8344 (N_8344,N_7854,N_7643);
or U8345 (N_8345,N_7987,N_6717);
nor U8346 (N_8346,N_7914,N_6764);
nor U8347 (N_8347,N_7560,N_6578);
nor U8348 (N_8348,N_7550,N_6220);
or U8349 (N_8349,N_7536,N_7303);
nor U8350 (N_8350,N_7480,N_7671);
or U8351 (N_8351,N_7340,N_6923);
and U8352 (N_8352,N_6161,N_6820);
or U8353 (N_8353,N_7909,N_6145);
and U8354 (N_8354,N_7930,N_6872);
nor U8355 (N_8355,N_7800,N_6730);
or U8356 (N_8356,N_7742,N_6931);
and U8357 (N_8357,N_6007,N_7801);
and U8358 (N_8358,N_7541,N_6079);
or U8359 (N_8359,N_6205,N_6586);
and U8360 (N_8360,N_6731,N_6588);
nand U8361 (N_8361,N_6052,N_7790);
and U8362 (N_8362,N_6602,N_7595);
nand U8363 (N_8363,N_7493,N_6984);
nand U8364 (N_8364,N_7055,N_7839);
and U8365 (N_8365,N_7469,N_7796);
nor U8366 (N_8366,N_7826,N_6934);
nand U8367 (N_8367,N_6423,N_6618);
or U8368 (N_8368,N_6297,N_6127);
nand U8369 (N_8369,N_7569,N_6976);
and U8370 (N_8370,N_6752,N_6076);
nand U8371 (N_8371,N_7218,N_6705);
nand U8372 (N_8372,N_6566,N_7348);
nor U8373 (N_8373,N_7926,N_6819);
and U8374 (N_8374,N_7270,N_6659);
or U8375 (N_8375,N_7331,N_7170);
nor U8376 (N_8376,N_6702,N_6114);
nand U8377 (N_8377,N_6362,N_7494);
and U8378 (N_8378,N_7401,N_6000);
nand U8379 (N_8379,N_6124,N_6166);
nor U8380 (N_8380,N_7101,N_6301);
nor U8381 (N_8381,N_6637,N_6375);
or U8382 (N_8382,N_7767,N_7945);
nor U8383 (N_8383,N_7045,N_7333);
nor U8384 (N_8384,N_7400,N_6622);
or U8385 (N_8385,N_7852,N_7131);
or U8386 (N_8386,N_6531,N_6448);
nor U8387 (N_8387,N_7957,N_7973);
nand U8388 (N_8388,N_7116,N_6721);
or U8389 (N_8389,N_6809,N_7512);
nor U8390 (N_8390,N_7601,N_7566);
nor U8391 (N_8391,N_7033,N_6292);
or U8392 (N_8392,N_6225,N_6869);
nor U8393 (N_8393,N_6072,N_6815);
nand U8394 (N_8394,N_6534,N_6598);
or U8395 (N_8395,N_7002,N_6723);
nand U8396 (N_8396,N_6149,N_6791);
nand U8397 (N_8397,N_6842,N_7990);
nor U8398 (N_8398,N_6090,N_6188);
nor U8399 (N_8399,N_7207,N_7729);
nand U8400 (N_8400,N_6541,N_7898);
or U8401 (N_8401,N_6757,N_7577);
nor U8402 (N_8402,N_7570,N_6839);
nand U8403 (N_8403,N_6447,N_7631);
nor U8404 (N_8404,N_6948,N_6590);
or U8405 (N_8405,N_6927,N_6870);
nor U8406 (N_8406,N_6393,N_7289);
nor U8407 (N_8407,N_7534,N_6950);
nor U8408 (N_8408,N_6018,N_7242);
or U8409 (N_8409,N_6834,N_6336);
and U8410 (N_8410,N_7007,N_6412);
and U8411 (N_8411,N_6614,N_7791);
or U8412 (N_8412,N_6712,N_6568);
nor U8413 (N_8413,N_6706,N_6441);
or U8414 (N_8414,N_7139,N_6113);
nand U8415 (N_8415,N_7166,N_6700);
nand U8416 (N_8416,N_7062,N_7081);
nand U8417 (N_8417,N_7492,N_7564);
or U8418 (N_8418,N_6737,N_6158);
or U8419 (N_8419,N_7195,N_6983);
or U8420 (N_8420,N_7129,N_7695);
and U8421 (N_8421,N_6755,N_7585);
and U8422 (N_8422,N_6536,N_6912);
or U8423 (N_8423,N_7107,N_7696);
and U8424 (N_8424,N_7921,N_6811);
and U8425 (N_8425,N_7720,N_7624);
and U8426 (N_8426,N_7635,N_6463);
and U8427 (N_8427,N_7747,N_6381);
nand U8428 (N_8428,N_7214,N_7181);
or U8429 (N_8429,N_6318,N_6696);
and U8430 (N_8430,N_7794,N_6787);
or U8431 (N_8431,N_7086,N_7655);
or U8432 (N_8432,N_6425,N_6317);
nor U8433 (N_8433,N_6234,N_6996);
nand U8434 (N_8434,N_7673,N_6843);
and U8435 (N_8435,N_6774,N_7349);
and U8436 (N_8436,N_7451,N_6725);
nor U8437 (N_8437,N_7753,N_6043);
nor U8438 (N_8438,N_7700,N_6432);
and U8439 (N_8439,N_7167,N_7953);
and U8440 (N_8440,N_6670,N_7395);
or U8441 (N_8441,N_7386,N_6907);
nor U8442 (N_8442,N_6047,N_6684);
nor U8443 (N_8443,N_6466,N_7483);
nand U8444 (N_8444,N_6549,N_7298);
nor U8445 (N_8445,N_7530,N_6314);
and U8446 (N_8446,N_6411,N_7952);
nor U8447 (N_8447,N_6893,N_7277);
nor U8448 (N_8448,N_6587,N_7971);
nor U8449 (N_8449,N_7581,N_6395);
or U8450 (N_8450,N_6861,N_7533);
nor U8451 (N_8451,N_6197,N_7960);
and U8452 (N_8452,N_7619,N_7406);
or U8453 (N_8453,N_6021,N_7302);
and U8454 (N_8454,N_6484,N_6758);
or U8455 (N_8455,N_7180,N_6055);
nor U8456 (N_8456,N_6247,N_6344);
and U8457 (N_8457,N_7387,N_7188);
or U8458 (N_8458,N_6634,N_6175);
or U8459 (N_8459,N_7992,N_6716);
and U8460 (N_8460,N_6667,N_6887);
and U8461 (N_8461,N_6335,N_7608);
and U8462 (N_8462,N_7297,N_6596);
nor U8463 (N_8463,N_6387,N_6749);
nand U8464 (N_8464,N_6745,N_7501);
and U8465 (N_8465,N_6801,N_6360);
nor U8466 (N_8466,N_6935,N_7831);
nor U8467 (N_8467,N_7925,N_6273);
nand U8468 (N_8468,N_7940,N_6396);
and U8469 (N_8469,N_7074,N_7659);
nor U8470 (N_8470,N_6152,N_6782);
or U8471 (N_8471,N_7427,N_7535);
nor U8472 (N_8472,N_6886,N_7276);
or U8473 (N_8473,N_7775,N_6888);
nor U8474 (N_8474,N_7066,N_6264);
and U8475 (N_8475,N_6176,N_6198);
and U8476 (N_8476,N_7411,N_6228);
nor U8477 (N_8477,N_6065,N_7473);
or U8478 (N_8478,N_7845,N_7453);
nand U8479 (N_8479,N_6506,N_7044);
nand U8480 (N_8480,N_7833,N_6284);
nand U8481 (N_8481,N_6734,N_7779);
and U8482 (N_8482,N_7105,N_6170);
or U8483 (N_8483,N_6272,N_6980);
or U8484 (N_8484,N_7666,N_6735);
nand U8485 (N_8485,N_6409,N_6077);
nor U8486 (N_8486,N_7809,N_7414);
nand U8487 (N_8487,N_7222,N_6985);
nor U8488 (N_8488,N_7407,N_7891);
or U8489 (N_8489,N_7683,N_7423);
or U8490 (N_8490,N_6496,N_6763);
nand U8491 (N_8491,N_7527,N_6140);
and U8492 (N_8492,N_7282,N_7227);
and U8493 (N_8493,N_7301,N_6365);
nor U8494 (N_8494,N_6929,N_7053);
or U8495 (N_8495,N_7802,N_6404);
nand U8496 (N_8496,N_6177,N_7334);
and U8497 (N_8497,N_6910,N_7668);
nor U8498 (N_8498,N_6060,N_7330);
nor U8499 (N_8499,N_7948,N_6821);
nor U8500 (N_8500,N_7151,N_6703);
nor U8501 (N_8501,N_7665,N_6027);
nor U8502 (N_8502,N_7113,N_6969);
nor U8503 (N_8503,N_7883,N_7645);
or U8504 (N_8504,N_7103,N_7439);
nor U8505 (N_8505,N_6483,N_7730);
nor U8506 (N_8506,N_7037,N_7748);
or U8507 (N_8507,N_7604,N_6468);
nor U8508 (N_8508,N_6627,N_7597);
or U8509 (N_8509,N_6822,N_6542);
nand U8510 (N_8510,N_6825,N_6812);
nand U8511 (N_8511,N_7496,N_6926);
and U8512 (N_8512,N_7877,N_6664);
nand U8513 (N_8513,N_7573,N_7358);
or U8514 (N_8514,N_6844,N_6402);
xnor U8515 (N_8515,N_7656,N_7164);
or U8516 (N_8516,N_7317,N_6508);
nand U8517 (N_8517,N_7885,N_7238);
xnor U8518 (N_8518,N_7591,N_7193);
nand U8519 (N_8519,N_7359,N_7967);
and U8520 (N_8520,N_7004,N_6035);
nand U8521 (N_8521,N_7632,N_7754);
or U8522 (N_8522,N_6961,N_6982);
nand U8523 (N_8523,N_6920,N_6651);
nor U8524 (N_8524,N_6204,N_6955);
or U8525 (N_8525,N_6921,N_7746);
or U8526 (N_8526,N_7409,N_7528);
nor U8527 (N_8527,N_6960,N_7068);
nor U8528 (N_8528,N_6903,N_7456);
nand U8529 (N_8529,N_6701,N_6153);
or U8530 (N_8530,N_6302,N_6909);
nor U8531 (N_8531,N_7623,N_6240);
or U8532 (N_8532,N_7288,N_6074);
nand U8533 (N_8533,N_6633,N_7497);
or U8534 (N_8534,N_6530,N_6378);
nand U8535 (N_8535,N_7939,N_7710);
xor U8536 (N_8536,N_6550,N_6434);
or U8537 (N_8537,N_6206,N_6453);
or U8538 (N_8538,N_6439,N_6263);
or U8539 (N_8539,N_6189,N_6491);
nand U8540 (N_8540,N_6994,N_6350);
or U8541 (N_8541,N_7638,N_6346);
nor U8542 (N_8542,N_7907,N_7011);
nor U8543 (N_8543,N_7506,N_6474);
nand U8544 (N_8544,N_6146,N_6159);
nand U8545 (N_8545,N_7281,N_6979);
and U8546 (N_8546,N_7658,N_7976);
nand U8547 (N_8547,N_6053,N_6789);
nand U8548 (N_8548,N_7416,N_6805);
nand U8549 (N_8549,N_7024,N_6250);
nand U8550 (N_8550,N_7245,N_6944);
nor U8551 (N_8551,N_7426,N_6407);
nand U8552 (N_8552,N_6342,N_6226);
and U8553 (N_8553,N_7513,N_7063);
nor U8554 (N_8554,N_6137,N_7706);
nor U8555 (N_8555,N_6069,N_7774);
nor U8556 (N_8556,N_6253,N_6320);
nor U8557 (N_8557,N_6591,N_7275);
nor U8558 (N_8558,N_6129,N_6525);
nand U8559 (N_8559,N_7977,N_7163);
or U8560 (N_8560,N_6186,N_7172);
nor U8561 (N_8561,N_7337,N_6275);
nand U8562 (N_8562,N_7810,N_7765);
nand U8563 (N_8563,N_7520,N_6321);
nor U8564 (N_8564,N_7067,N_6262);
xnor U8565 (N_8565,N_6006,N_7784);
or U8566 (N_8566,N_6663,N_6026);
nand U8567 (N_8567,N_6467,N_7705);
nand U8568 (N_8568,N_7662,N_6971);
nand U8569 (N_8569,N_7507,N_7300);
or U8570 (N_8570,N_7648,N_6638);
or U8571 (N_8571,N_6829,N_6630);
nand U8572 (N_8572,N_6479,N_6001);
or U8573 (N_8573,N_7539,N_6648);
and U8574 (N_8574,N_7162,N_7708);
nor U8575 (N_8575,N_7199,N_7944);
nor U8576 (N_8576,N_6325,N_7610);
nand U8577 (N_8577,N_6300,N_7759);
nor U8578 (N_8578,N_7500,N_7179);
nor U8579 (N_8579,N_7383,N_6178);
and U8580 (N_8580,N_7200,N_6288);
or U8581 (N_8581,N_6039,N_6050);
nand U8582 (N_8582,N_6019,N_6577);
or U8583 (N_8583,N_7380,N_7019);
nand U8584 (N_8584,N_6235,N_6135);
nand U8585 (N_8585,N_7519,N_7763);
or U8586 (N_8586,N_7862,N_7402);
nor U8587 (N_8587,N_7318,N_7474);
and U8588 (N_8588,N_6005,N_7251);
nand U8589 (N_8589,N_7637,N_6224);
nand U8590 (N_8590,N_6792,N_7425);
nand U8591 (N_8591,N_6171,N_7614);
nand U8592 (N_8592,N_6392,N_7023);
and U8593 (N_8593,N_6860,N_7609);
or U8594 (N_8594,N_6245,N_6061);
nand U8595 (N_8595,N_7736,N_7738);
nor U8596 (N_8596,N_6282,N_6182);
nor U8597 (N_8597,N_6416,N_7324);
nand U8598 (N_8598,N_7089,N_6973);
nor U8599 (N_8599,N_7733,N_7070);
nand U8600 (N_8600,N_7903,N_7135);
nand U8601 (N_8601,N_6089,N_6848);
and U8602 (N_8602,N_7950,N_7870);
nand U8603 (N_8603,N_6278,N_7069);
nand U8604 (N_8604,N_6492,N_7691);
and U8605 (N_8605,N_7578,N_6128);
nor U8606 (N_8606,N_7998,N_6157);
nor U8607 (N_8607,N_6513,N_7205);
nand U8608 (N_8608,N_7558,N_6552);
nand U8609 (N_8609,N_7430,N_6254);
and U8610 (N_8610,N_7761,N_7126);
nor U8611 (N_8611,N_7568,N_7702);
nand U8612 (N_8612,N_6919,N_6744);
nand U8613 (N_8613,N_6429,N_7092);
and U8614 (N_8614,N_6660,N_6459);
nor U8615 (N_8615,N_7118,N_6501);
nand U8616 (N_8616,N_6212,N_6507);
nor U8617 (N_8617,N_6340,N_7192);
nor U8618 (N_8618,N_6296,N_6991);
nor U8619 (N_8619,N_7177,N_6040);
and U8620 (N_8620,N_7311,N_6347);
nor U8621 (N_8621,N_6222,N_7864);
nor U8622 (N_8622,N_7968,N_6115);
nand U8623 (N_8623,N_7504,N_7408);
nand U8624 (N_8624,N_7769,N_7052);
or U8625 (N_8625,N_6671,N_6751);
and U8626 (N_8626,N_6029,N_7476);
nand U8627 (N_8627,N_6523,N_6873);
or U8628 (N_8628,N_7871,N_7345);
nand U8629 (N_8629,N_7261,N_6571);
nand U8630 (N_8630,N_6431,N_6704);
or U8631 (N_8631,N_6876,N_7484);
or U8632 (N_8632,N_6046,N_7576);
or U8633 (N_8633,N_6449,N_7545);
or U8634 (N_8634,N_6594,N_7217);
and U8635 (N_8635,N_7388,N_6283);
nand U8636 (N_8636,N_6422,N_6722);
and U8637 (N_8637,N_7419,N_6418);
or U8638 (N_8638,N_7335,N_7690);
nor U8639 (N_8639,N_6993,N_6173);
nand U8640 (N_8640,N_7236,N_6038);
nor U8641 (N_8641,N_6558,N_6095);
nand U8642 (N_8642,N_7123,N_7860);
nor U8643 (N_8643,N_7954,N_7602);
or U8644 (N_8644,N_6489,N_6581);
nor U8645 (N_8645,N_7355,N_6713);
or U8646 (N_8646,N_7654,N_6285);
and U8647 (N_8647,N_6013,N_7434);
nor U8648 (N_8648,N_6604,N_7844);
and U8649 (N_8649,N_6478,N_7933);
or U8650 (N_8650,N_7307,N_6354);
nor U8651 (N_8651,N_6697,N_7721);
nor U8652 (N_8652,N_6708,N_7204);
or U8653 (N_8653,N_7420,N_7711);
and U8654 (N_8654,N_7306,N_6832);
or U8655 (N_8655,N_7843,N_6625);
and U8656 (N_8656,N_7857,N_6561);
nor U8657 (N_8657,N_7030,N_6526);
nor U8658 (N_8658,N_6519,N_7226);
and U8659 (N_8659,N_7397,N_7100);
or U8660 (N_8660,N_6154,N_6658);
and U8661 (N_8661,N_7538,N_7379);
nor U8662 (N_8662,N_6391,N_6372);
or U8663 (N_8663,N_6452,N_7094);
and U8664 (N_8664,N_7357,N_6642);
xnor U8665 (N_8665,N_7028,N_6270);
or U8666 (N_8666,N_6281,N_6203);
and U8667 (N_8667,N_7853,N_6132);
or U8668 (N_8668,N_6068,N_7531);
and U8669 (N_8669,N_7824,N_6277);
nor U8670 (N_8670,N_6430,N_7896);
and U8671 (N_8671,N_6728,N_7471);
and U8672 (N_8672,N_7232,N_6964);
or U8673 (N_8673,N_6522,N_7064);
nor U8674 (N_8674,N_6258,N_7739);
nand U8675 (N_8675,N_6512,N_6223);
and U8676 (N_8676,N_6097,N_6122);
or U8677 (N_8677,N_7995,N_6357);
and U8678 (N_8678,N_6942,N_6619);
nor U8679 (N_8679,N_6783,N_6827);
or U8680 (N_8680,N_6126,N_6972);
nand U8681 (N_8681,N_6862,N_7132);
nand U8682 (N_8682,N_6748,N_6119);
nor U8683 (N_8683,N_6954,N_7880);
or U8684 (N_8684,N_7727,N_7618);
or U8685 (N_8685,N_7039,N_6892);
and U8686 (N_8686,N_7341,N_7685);
and U8687 (N_8687,N_6112,N_7678);
nand U8688 (N_8688,N_6110,N_7561);
nand U8689 (N_8689,N_7182,N_6081);
nor U8690 (N_8690,N_6286,N_6925);
or U8691 (N_8691,N_7596,N_7364);
nor U8692 (N_8692,N_7726,N_6645);
and U8693 (N_8693,N_7657,N_6772);
and U8694 (N_8694,N_7629,N_7314);
nor U8695 (N_8695,N_7363,N_7018);
nand U8696 (N_8696,N_6810,N_6952);
nand U8697 (N_8697,N_7137,N_7017);
or U8698 (N_8698,N_6902,N_7394);
nor U8699 (N_8699,N_7553,N_6941);
or U8700 (N_8700,N_7268,N_6773);
nand U8701 (N_8701,N_6502,N_6761);
or U8702 (N_8702,N_6846,N_7837);
and U8703 (N_8703,N_6733,N_6804);
or U8704 (N_8704,N_7703,N_7731);
nand U8705 (N_8705,N_7048,N_6615);
nor U8706 (N_8706,N_6616,N_7153);
nor U8707 (N_8707,N_6363,N_6896);
nor U8708 (N_8708,N_6267,N_6169);
and U8709 (N_8709,N_6257,N_7438);
nor U8710 (N_8710,N_6718,N_6172);
nor U8711 (N_8711,N_6147,N_7894);
nand U8712 (N_8712,N_6117,N_7827);
and U8713 (N_8713,N_7650,N_7059);
nor U8714 (N_8714,N_6099,N_7291);
or U8715 (N_8715,N_6798,N_6091);
or U8716 (N_8716,N_7417,N_7114);
or U8717 (N_8717,N_6548,N_6293);
or U8718 (N_8718,N_7450,N_6759);
nor U8719 (N_8719,N_7076,N_7253);
nand U8720 (N_8720,N_7244,N_6589);
nand U8721 (N_8721,N_6607,N_7981);
nand U8722 (N_8722,N_7636,N_7676);
nand U8723 (N_8723,N_7680,N_6276);
nand U8724 (N_8724,N_7015,N_7360);
and U8725 (N_8725,N_6504,N_6599);
xor U8726 (N_8726,N_7792,N_6054);
nor U8727 (N_8727,N_7962,N_7384);
and U8728 (N_8728,N_7866,N_6563);
nor U8729 (N_8729,N_7755,N_7848);
and U8730 (N_8730,N_6085,N_6487);
or U8731 (N_8731,N_7250,N_7191);
nor U8732 (N_8732,N_7036,N_6797);
xor U8733 (N_8733,N_6131,N_6959);
or U8734 (N_8734,N_7579,N_6460);
or U8735 (N_8735,N_6939,N_6726);
nand U8736 (N_8736,N_6672,N_7804);
nor U8737 (N_8737,N_6517,N_6241);
and U8738 (N_8738,N_6403,N_7260);
nand U8739 (N_8739,N_6251,N_6230);
and U8740 (N_8740,N_7764,N_6665);
nand U8741 (N_8741,N_6882,N_7546);
and U8742 (N_8742,N_6683,N_7988);
nand U8743 (N_8743,N_6974,N_6148);
and U8744 (N_8744,N_7913,N_7628);
and U8745 (N_8745,N_7825,N_7805);
nand U8746 (N_8746,N_7234,N_6442);
nor U8747 (N_8747,N_7942,N_6307);
and U8748 (N_8748,N_7989,N_7032);
or U8749 (N_8749,N_6678,N_6064);
or U8750 (N_8750,N_7410,N_7798);
and U8751 (N_8751,N_6333,N_7603);
or U8752 (N_8752,N_6680,N_7878);
or U8753 (N_8753,N_7881,N_7313);
and U8754 (N_8754,N_6901,N_6209);
or U8755 (N_8755,N_7399,N_6315);
nor U8756 (N_8756,N_6760,N_7461);
or U8757 (N_8757,N_7681,N_6359);
nor U8758 (N_8758,N_7431,N_7797);
nand U8759 (N_8759,N_6769,N_6740);
and U8760 (N_8760,N_6408,N_7508);
and U8761 (N_8761,N_6465,N_6495);
nor U8762 (N_8762,N_6628,N_7679);
or U8763 (N_8763,N_6924,N_7715);
nor U8764 (N_8764,N_6111,N_6329);
nand U8765 (N_8765,N_7280,N_7034);
or U8766 (N_8766,N_7351,N_6727);
nor U8767 (N_8767,N_7393,N_7444);
nand U8768 (N_8768,N_6208,N_7470);
or U8769 (N_8769,N_6244,N_7701);
and U8770 (N_8770,N_7404,N_7812);
nand U8771 (N_8771,N_6610,N_6303);
and U8772 (N_8772,N_6456,N_6807);
and U8773 (N_8773,N_6753,N_7171);
nor U8774 (N_8774,N_7743,N_7842);
xnor U8775 (N_8775,N_6142,N_6897);
nor U8776 (N_8776,N_7965,N_6710);
nand U8777 (N_8777,N_7485,N_6351);
and U8778 (N_8778,N_6898,N_6569);
and U8779 (N_8779,N_6573,N_6062);
nand U8780 (N_8780,N_6374,N_7087);
or U8781 (N_8781,N_6032,N_7040);
nor U8782 (N_8782,N_7542,N_7464);
or U8783 (N_8783,N_6747,N_7323);
or U8784 (N_8784,N_6073,N_6555);
nand U8785 (N_8785,N_7117,N_7446);
nand U8786 (N_8786,N_6510,N_7556);
nand U8787 (N_8787,N_6094,N_6031);
or U8788 (N_8788,N_7326,N_6218);
nand U8789 (N_8789,N_7562,N_7979);
nor U8790 (N_8790,N_6366,N_7221);
and U8791 (N_8791,N_6217,N_7851);
nor U8792 (N_8792,N_7057,N_7468);
or U8793 (N_8793,N_7432,N_6854);
or U8794 (N_8794,N_6488,N_7505);
nand U8795 (N_8795,N_7252,N_6084);
and U8796 (N_8796,N_7127,N_7714);
or U8797 (N_8797,N_7785,N_6291);
nand U8798 (N_8798,N_6427,N_7958);
or U8799 (N_8799,N_7719,N_7502);
nand U8800 (N_8800,N_6565,N_7134);
and U8801 (N_8801,N_6990,N_7237);
and U8802 (N_8802,N_7343,N_6444);
nor U8803 (N_8803,N_6899,N_7523);
nor U8804 (N_8804,N_6641,N_7158);
and U8805 (N_8805,N_7598,N_7262);
or U8806 (N_8806,N_6943,N_7544);
and U8807 (N_8807,N_7956,N_6451);
or U8808 (N_8808,N_6933,N_7014);
nor U8809 (N_8809,N_6058,N_6687);
nand U8810 (N_8810,N_6133,N_6455);
nor U8811 (N_8811,N_6310,N_6059);
and U8812 (N_8812,N_7421,N_7652);
nand U8813 (N_8813,N_7102,N_6435);
nand U8814 (N_8814,N_6521,N_6405);
or U8815 (N_8815,N_7841,N_7295);
nor U8816 (N_8816,N_7687,N_7664);
or U8817 (N_8817,N_6016,N_6187);
and U8818 (N_8818,N_6715,N_6863);
and U8819 (N_8819,N_6711,N_6889);
xnor U8820 (N_8820,N_7152,N_7130);
or U8821 (N_8821,N_7272,N_7757);
or U8822 (N_8822,N_6237,N_6623);
nand U8823 (N_8823,N_7320,N_7752);
nor U8824 (N_8824,N_6669,N_6123);
or U8825 (N_8825,N_6605,N_7582);
nand U8826 (N_8826,N_7243,N_7168);
nand U8827 (N_8827,N_7599,N_6164);
nand U8828 (N_8828,N_7834,N_7398);
and U8829 (N_8829,N_6654,N_7912);
nor U8830 (N_8830,N_6471,N_7022);
nand U8831 (N_8831,N_7212,N_6280);
nor U8832 (N_8832,N_6913,N_6426);
nand U8833 (N_8833,N_7850,N_7819);
and U8834 (N_8834,N_6290,N_7876);
and U8835 (N_8835,N_6011,N_7814);
and U8836 (N_8836,N_6008,N_6120);
nor U8837 (N_8837,N_7626,N_7972);
or U8838 (N_8838,N_6410,N_7928);
nand U8839 (N_8839,N_6940,N_7830);
nor U8840 (N_8840,N_6790,N_6612);
or U8841 (N_8841,N_7287,N_6613);
and U8842 (N_8842,N_6690,N_6962);
or U8843 (N_8843,N_6330,N_6322);
nor U8844 (N_8844,N_6397,N_7770);
and U8845 (N_8845,N_6165,N_7808);
nand U8846 (N_8846,N_7265,N_7058);
and U8847 (N_8847,N_7892,N_6475);
nand U8848 (N_8848,N_6657,N_6421);
nor U8849 (N_8849,N_6236,N_6367);
nor U8850 (N_8850,N_7128,N_7258);
or U8851 (N_8851,N_6214,N_7428);
and U8852 (N_8852,N_7551,N_7457);
nand U8853 (N_8853,N_6567,N_7025);
nor U8854 (N_8854,N_7233,N_7697);
and U8855 (N_8855,N_6213,N_7525);
nor U8856 (N_8856,N_6388,N_6080);
nor U8857 (N_8857,N_7887,N_6078);
or U8858 (N_8858,N_7997,N_6469);
and U8859 (N_8859,N_7441,N_7865);
or U8860 (N_8860,N_7737,N_6922);
nand U8861 (N_8861,N_7455,N_7677);
and U8862 (N_8862,N_6399,N_6485);
and U8863 (N_8863,N_7592,N_6556);
or U8864 (N_8864,N_7906,N_6691);
and U8865 (N_8865,N_6450,N_6246);
or U8866 (N_8866,N_7712,N_6243);
nand U8867 (N_8867,N_6193,N_6765);
or U8868 (N_8868,N_7717,N_6389);
and U8869 (N_8869,N_6540,N_6875);
or U8870 (N_8870,N_6150,N_7051);
nor U8871 (N_8871,N_7557,N_6778);
and U8872 (N_8872,N_6879,N_6037);
nand U8873 (N_8873,N_6486,N_6817);
or U8874 (N_8874,N_7849,N_7522);
or U8875 (N_8875,N_6852,N_7042);
xnor U8876 (N_8876,N_7642,N_7984);
or U8877 (N_8877,N_6743,N_7391);
and U8878 (N_8878,N_6109,N_6582);
nor U8879 (N_8879,N_7594,N_6784);
nor U8880 (N_8880,N_7046,N_7016);
nand U8881 (N_8881,N_6802,N_7196);
nand U8882 (N_8882,N_7918,N_7613);
and U8883 (N_8883,N_7124,N_6849);
nor U8884 (N_8884,N_7975,N_7709);
or U8885 (N_8885,N_6878,N_6151);
nand U8886 (N_8886,N_7050,N_6370);
and U8887 (N_8887,N_7442,N_6632);
nor U8888 (N_8888,N_6231,N_6688);
or U8889 (N_8889,N_7194,N_7616);
nand U8890 (N_8890,N_7043,N_7472);
nor U8891 (N_8891,N_7437,N_7286);
nand U8892 (N_8892,N_6355,N_6136);
nand U8893 (N_8893,N_6793,N_7537);
nand U8894 (N_8894,N_6156,N_7688);
nor U8895 (N_8895,N_6856,N_7120);
nand U8896 (N_8896,N_7368,N_6238);
nor U8897 (N_8897,N_7902,N_7807);
nor U8898 (N_8898,N_6428,N_6551);
nand U8899 (N_8899,N_6788,N_7003);
nand U8900 (N_8900,N_7147,N_7223);
and U8901 (N_8901,N_7915,N_7554);
and U8902 (N_8902,N_6732,N_7112);
and U8903 (N_8903,N_6714,N_7278);
nor U8904 (N_8904,N_6063,N_7273);
and U8905 (N_8905,N_7588,N_6167);
or U8906 (N_8906,N_7605,N_6143);
nor U8907 (N_8907,N_7475,N_7361);
nand U8908 (N_8908,N_6015,N_7122);
nor U8909 (N_8909,N_7682,N_7840);
nor U8910 (N_8910,N_7617,N_7999);
nand U8911 (N_8911,N_7510,N_6313);
nand U8912 (N_8912,N_7133,N_6776);
or U8913 (N_8913,N_7106,N_7651);
nand U8914 (N_8914,N_7806,N_6385);
nand U8915 (N_8915,N_6617,N_6051);
or U8916 (N_8916,N_7803,N_6646);
nand U8917 (N_8917,N_6914,N_7964);
nor U8918 (N_8918,N_7863,N_7206);
or U8919 (N_8919,N_6775,N_7771);
nor U8920 (N_8920,N_7963,N_7079);
nand U8921 (N_8921,N_7176,N_6547);
and U8922 (N_8922,N_6795,N_7061);
nor U8923 (N_8923,N_6738,N_6232);
and U8924 (N_8924,N_6766,N_6227);
and U8925 (N_8925,N_6201,N_6480);
nor U8926 (N_8926,N_7008,N_7491);
nor U8927 (N_8927,N_6918,N_6332);
nor U8928 (N_8928,N_6967,N_6771);
nand U8929 (N_8929,N_7868,N_6337);
nand U8930 (N_8930,N_7498,N_6518);
or U8931 (N_8931,N_6883,N_7145);
or U8932 (N_8932,N_7099,N_7487);
nand U8933 (N_8933,N_7462,N_7901);
or U8934 (N_8934,N_7781,N_6134);
nand U8935 (N_8935,N_6221,N_7869);
nor U8936 (N_8936,N_6215,N_6279);
nor U8937 (N_8937,N_6490,N_6803);
or U8938 (N_8938,N_7012,N_7412);
and U8939 (N_8939,N_6595,N_6289);
nand U8940 (N_8940,N_6750,N_7459);
nor U8941 (N_8941,N_7822,N_6082);
nand U8942 (N_8942,N_7190,N_7838);
and U8943 (N_8943,N_6500,N_6794);
or U8944 (N_8944,N_6930,N_6890);
and U8945 (N_8945,N_6928,N_7789);
nand U8946 (N_8946,N_6353,N_7511);
and U8947 (N_8947,N_7478,N_6527);
nor U8948 (N_8948,N_7625,N_7750);
and U8949 (N_8949,N_7111,N_7661);
nand U8950 (N_8950,N_6989,N_6845);
and U8951 (N_8951,N_6557,N_6673);
xor U8952 (N_8952,N_7549,N_7342);
or U8953 (N_8953,N_7649,N_7978);
nor U8954 (N_8954,N_6838,N_7766);
or U8955 (N_8955,N_7154,N_7047);
or U8956 (N_8956,N_6968,N_7366);
nor U8957 (N_8957,N_6624,N_6742);
nand U8958 (N_8958,N_6699,N_7606);
nand U8959 (N_8959,N_7835,N_7882);
nand U8960 (N_8960,N_7184,N_6768);
and U8961 (N_8961,N_6194,N_7698);
nand U8962 (N_8962,N_7937,N_7611);
and U8963 (N_8963,N_7435,N_6249);
nand U8964 (N_8964,N_7146,N_7201);
nand U8965 (N_8965,N_6814,N_7961);
or U8966 (N_8966,N_6384,N_7787);
and U8967 (N_8967,N_7001,N_6956);
and U8968 (N_8968,N_7274,N_6559);
and U8969 (N_8969,N_7941,N_7440);
nor U8970 (N_8970,N_6380,N_7091);
nor U8971 (N_8971,N_7707,N_6324);
or U8972 (N_8972,N_6162,N_7499);
nand U8973 (N_8973,N_6999,N_7315);
nor U8974 (N_8974,N_7109,N_7010);
and U8975 (N_8975,N_7353,N_6259);
nand U8976 (N_8976,N_7228,N_6304);
and U8977 (N_8977,N_7584,N_6105);
and U8978 (N_8978,N_7890,N_7936);
and U8979 (N_8979,N_7073,N_7038);
nor U8980 (N_8980,N_6295,N_6529);
nor U8981 (N_8981,N_6608,N_7035);
nor U8982 (N_8982,N_6677,N_7749);
or U8983 (N_8983,N_7762,N_7354);
nor U8984 (N_8984,N_7389,N_6947);
and U8985 (N_8985,N_7563,N_7241);
or U8986 (N_8986,N_6695,N_7436);
nor U8987 (N_8987,N_7728,N_7328);
nand U8988 (N_8988,N_7660,N_7847);
or U8989 (N_8989,N_6679,N_7899);
nand U8990 (N_8990,N_7321,N_6951);
nand U8991 (N_8991,N_7405,N_6880);
or U8992 (N_8992,N_7165,N_6762);
nand U8993 (N_8993,N_7716,N_7338);
and U8994 (N_8994,N_7872,N_6655);
nor U8995 (N_8995,N_7143,N_6481);
and U8996 (N_8996,N_7821,N_6163);
or U8997 (N_8997,N_6382,N_7138);
or U8998 (N_8998,N_6025,N_6048);
and U8999 (N_8999,N_7622,N_6831);
or U9000 (N_9000,N_7866,N_7746);
nand U9001 (N_9001,N_6636,N_6053);
nand U9002 (N_9002,N_7614,N_7348);
nand U9003 (N_9003,N_6057,N_7740);
and U9004 (N_9004,N_6516,N_6212);
or U9005 (N_9005,N_6480,N_6767);
nand U9006 (N_9006,N_6480,N_7889);
and U9007 (N_9007,N_7267,N_6291);
and U9008 (N_9008,N_7024,N_7101);
nand U9009 (N_9009,N_7971,N_7756);
nand U9010 (N_9010,N_6364,N_7398);
and U9011 (N_9011,N_6521,N_6310);
nand U9012 (N_9012,N_7938,N_7909);
and U9013 (N_9013,N_6181,N_6169);
xor U9014 (N_9014,N_6521,N_6020);
nand U9015 (N_9015,N_7580,N_6813);
and U9016 (N_9016,N_6611,N_6860);
nand U9017 (N_9017,N_6173,N_7974);
nand U9018 (N_9018,N_6819,N_7619);
nand U9019 (N_9019,N_7446,N_6338);
and U9020 (N_9020,N_6643,N_6154);
or U9021 (N_9021,N_6656,N_6484);
nor U9022 (N_9022,N_6408,N_6881);
or U9023 (N_9023,N_6164,N_6529);
or U9024 (N_9024,N_6080,N_7203);
nor U9025 (N_9025,N_7430,N_6264);
nor U9026 (N_9026,N_7558,N_7521);
nand U9027 (N_9027,N_6959,N_7440);
or U9028 (N_9028,N_6451,N_6712);
nor U9029 (N_9029,N_6803,N_7835);
and U9030 (N_9030,N_7966,N_6955);
or U9031 (N_9031,N_6704,N_7420);
nand U9032 (N_9032,N_7544,N_6578);
nand U9033 (N_9033,N_6828,N_6837);
nor U9034 (N_9034,N_7368,N_7291);
or U9035 (N_9035,N_7924,N_6061);
or U9036 (N_9036,N_6468,N_6407);
and U9037 (N_9037,N_6959,N_7085);
nor U9038 (N_9038,N_7238,N_7791);
nand U9039 (N_9039,N_7932,N_6234);
nand U9040 (N_9040,N_7797,N_6165);
or U9041 (N_9041,N_6326,N_6537);
or U9042 (N_9042,N_6474,N_6698);
nand U9043 (N_9043,N_6746,N_7320);
or U9044 (N_9044,N_6326,N_6105);
or U9045 (N_9045,N_6321,N_7701);
and U9046 (N_9046,N_6513,N_6263);
nand U9047 (N_9047,N_7070,N_6304);
or U9048 (N_9048,N_7914,N_6842);
nor U9049 (N_9049,N_6688,N_6483);
xnor U9050 (N_9050,N_6326,N_6644);
and U9051 (N_9051,N_6864,N_6647);
or U9052 (N_9052,N_7569,N_6167);
nor U9053 (N_9053,N_6505,N_7468);
and U9054 (N_9054,N_7940,N_7767);
or U9055 (N_9055,N_6647,N_6107);
or U9056 (N_9056,N_6165,N_6563);
nand U9057 (N_9057,N_7954,N_7256);
nand U9058 (N_9058,N_6316,N_7760);
or U9059 (N_9059,N_7988,N_6048);
xnor U9060 (N_9060,N_6060,N_7382);
nor U9061 (N_9061,N_7871,N_7454);
or U9062 (N_9062,N_7687,N_6044);
xor U9063 (N_9063,N_6427,N_7988);
nand U9064 (N_9064,N_6858,N_7332);
nand U9065 (N_9065,N_6745,N_7184);
nor U9066 (N_9066,N_6736,N_6589);
nor U9067 (N_9067,N_7086,N_6227);
or U9068 (N_9068,N_7148,N_7064);
or U9069 (N_9069,N_7161,N_7863);
or U9070 (N_9070,N_7221,N_6153);
and U9071 (N_9071,N_7089,N_7706);
or U9072 (N_9072,N_7436,N_7637);
nor U9073 (N_9073,N_7175,N_7425);
nor U9074 (N_9074,N_7897,N_6545);
nor U9075 (N_9075,N_7106,N_6685);
nor U9076 (N_9076,N_7915,N_6995);
or U9077 (N_9077,N_7509,N_6140);
and U9078 (N_9078,N_6990,N_7629);
nand U9079 (N_9079,N_7861,N_7909);
nand U9080 (N_9080,N_7380,N_7391);
nand U9081 (N_9081,N_7955,N_6475);
nor U9082 (N_9082,N_6283,N_7755);
nand U9083 (N_9083,N_6066,N_7884);
or U9084 (N_9084,N_7471,N_6146);
nor U9085 (N_9085,N_7463,N_7512);
nor U9086 (N_9086,N_7892,N_6470);
nand U9087 (N_9087,N_7047,N_7452);
and U9088 (N_9088,N_7890,N_6838);
nand U9089 (N_9089,N_7476,N_6446);
and U9090 (N_9090,N_7700,N_6805);
nor U9091 (N_9091,N_7503,N_7752);
nand U9092 (N_9092,N_7697,N_6835);
and U9093 (N_9093,N_6821,N_6760);
nand U9094 (N_9094,N_7064,N_7038);
nor U9095 (N_9095,N_6420,N_7488);
and U9096 (N_9096,N_7903,N_7278);
nand U9097 (N_9097,N_6818,N_6564);
nor U9098 (N_9098,N_6035,N_7062);
and U9099 (N_9099,N_7591,N_6478);
or U9100 (N_9100,N_7087,N_6429);
nand U9101 (N_9101,N_6565,N_6307);
and U9102 (N_9102,N_7844,N_6194);
and U9103 (N_9103,N_6728,N_7729);
nand U9104 (N_9104,N_7512,N_7844);
nand U9105 (N_9105,N_6821,N_6265);
nand U9106 (N_9106,N_6986,N_6836);
and U9107 (N_9107,N_6603,N_6465);
nor U9108 (N_9108,N_6541,N_7868);
or U9109 (N_9109,N_7160,N_6331);
nor U9110 (N_9110,N_6476,N_6154);
or U9111 (N_9111,N_7797,N_6057);
or U9112 (N_9112,N_7066,N_6667);
xor U9113 (N_9113,N_6507,N_7839);
or U9114 (N_9114,N_7821,N_7461);
or U9115 (N_9115,N_6164,N_7569);
nand U9116 (N_9116,N_6536,N_6579);
nand U9117 (N_9117,N_7699,N_7805);
xnor U9118 (N_9118,N_7523,N_7584);
and U9119 (N_9119,N_7136,N_6772);
and U9120 (N_9120,N_6367,N_7933);
nand U9121 (N_9121,N_6695,N_6748);
and U9122 (N_9122,N_7375,N_6804);
nor U9123 (N_9123,N_7543,N_7945);
and U9124 (N_9124,N_6914,N_6185);
nand U9125 (N_9125,N_7814,N_7872);
or U9126 (N_9126,N_6412,N_7475);
nand U9127 (N_9127,N_6187,N_6024);
or U9128 (N_9128,N_6441,N_7568);
and U9129 (N_9129,N_7676,N_7236);
xnor U9130 (N_9130,N_6614,N_7744);
or U9131 (N_9131,N_6000,N_6895);
or U9132 (N_9132,N_6732,N_6487);
nor U9133 (N_9133,N_6864,N_7189);
and U9134 (N_9134,N_6511,N_7923);
and U9135 (N_9135,N_6363,N_7947);
nand U9136 (N_9136,N_7983,N_7464);
or U9137 (N_9137,N_6392,N_6894);
and U9138 (N_9138,N_6488,N_7295);
or U9139 (N_9139,N_6694,N_6272);
nand U9140 (N_9140,N_7234,N_7774);
and U9141 (N_9141,N_6831,N_7058);
and U9142 (N_9142,N_7514,N_6148);
and U9143 (N_9143,N_7136,N_6918);
nand U9144 (N_9144,N_7048,N_7522);
nand U9145 (N_9145,N_7121,N_6590);
nand U9146 (N_9146,N_7845,N_7373);
nand U9147 (N_9147,N_6312,N_7905);
and U9148 (N_9148,N_7011,N_7230);
nor U9149 (N_9149,N_7635,N_7813);
nand U9150 (N_9150,N_6437,N_6802);
nand U9151 (N_9151,N_7719,N_7528);
nand U9152 (N_9152,N_6469,N_7472);
and U9153 (N_9153,N_7495,N_7561);
and U9154 (N_9154,N_7682,N_7390);
nand U9155 (N_9155,N_6908,N_6108);
or U9156 (N_9156,N_7271,N_7842);
or U9157 (N_9157,N_7438,N_6125);
and U9158 (N_9158,N_6813,N_6194);
nand U9159 (N_9159,N_7613,N_7824);
nand U9160 (N_9160,N_7123,N_7549);
nor U9161 (N_9161,N_7530,N_6649);
nor U9162 (N_9162,N_6374,N_6768);
nand U9163 (N_9163,N_6972,N_6913);
and U9164 (N_9164,N_6540,N_7558);
and U9165 (N_9165,N_6010,N_7011);
and U9166 (N_9166,N_7235,N_6770);
and U9167 (N_9167,N_7058,N_6813);
nand U9168 (N_9168,N_7317,N_7090);
and U9169 (N_9169,N_6978,N_7041);
or U9170 (N_9170,N_7657,N_7495);
and U9171 (N_9171,N_6564,N_7482);
and U9172 (N_9172,N_7492,N_7599);
and U9173 (N_9173,N_6922,N_6561);
or U9174 (N_9174,N_7838,N_7242);
and U9175 (N_9175,N_7543,N_6593);
or U9176 (N_9176,N_6650,N_6532);
nand U9177 (N_9177,N_7202,N_7035);
or U9178 (N_9178,N_6928,N_7524);
nor U9179 (N_9179,N_6488,N_6558);
and U9180 (N_9180,N_6572,N_7854);
and U9181 (N_9181,N_6316,N_6947);
or U9182 (N_9182,N_6722,N_7345);
and U9183 (N_9183,N_6838,N_7255);
nor U9184 (N_9184,N_7769,N_6011);
nor U9185 (N_9185,N_7260,N_6772);
or U9186 (N_9186,N_7924,N_6055);
nand U9187 (N_9187,N_6971,N_6095);
nand U9188 (N_9188,N_7169,N_7320);
nand U9189 (N_9189,N_6195,N_7619);
and U9190 (N_9190,N_7281,N_7202);
or U9191 (N_9191,N_6962,N_6695);
and U9192 (N_9192,N_7959,N_7030);
nor U9193 (N_9193,N_6883,N_6745);
nand U9194 (N_9194,N_7024,N_7532);
and U9195 (N_9195,N_7084,N_7075);
nand U9196 (N_9196,N_7568,N_6933);
xor U9197 (N_9197,N_7997,N_6355);
nor U9198 (N_9198,N_7949,N_7180);
nor U9199 (N_9199,N_7688,N_6894);
and U9200 (N_9200,N_7241,N_7292);
and U9201 (N_9201,N_6739,N_6363);
or U9202 (N_9202,N_6355,N_6421);
nand U9203 (N_9203,N_7722,N_6950);
or U9204 (N_9204,N_6897,N_6571);
nor U9205 (N_9205,N_6080,N_6387);
and U9206 (N_9206,N_7370,N_7083);
nor U9207 (N_9207,N_7098,N_6538);
nor U9208 (N_9208,N_6182,N_7507);
nor U9209 (N_9209,N_6576,N_7370);
or U9210 (N_9210,N_7974,N_7748);
and U9211 (N_9211,N_7477,N_6210);
nand U9212 (N_9212,N_6476,N_7654);
or U9213 (N_9213,N_7780,N_6955);
and U9214 (N_9214,N_6404,N_6052);
and U9215 (N_9215,N_6569,N_7664);
and U9216 (N_9216,N_6372,N_7551);
nor U9217 (N_9217,N_7604,N_7897);
nor U9218 (N_9218,N_6594,N_7952);
or U9219 (N_9219,N_6195,N_7048);
nor U9220 (N_9220,N_6678,N_6256);
and U9221 (N_9221,N_6583,N_7613);
or U9222 (N_9222,N_7563,N_6881);
nor U9223 (N_9223,N_7592,N_6091);
nor U9224 (N_9224,N_6283,N_6480);
nand U9225 (N_9225,N_7375,N_6786);
nand U9226 (N_9226,N_7690,N_7433);
nand U9227 (N_9227,N_6197,N_6229);
nor U9228 (N_9228,N_7039,N_6121);
nor U9229 (N_9229,N_7844,N_6134);
nand U9230 (N_9230,N_7380,N_6552);
nor U9231 (N_9231,N_6732,N_7420);
and U9232 (N_9232,N_7923,N_6764);
nand U9233 (N_9233,N_7454,N_7702);
nor U9234 (N_9234,N_6331,N_7202);
nand U9235 (N_9235,N_6594,N_7247);
and U9236 (N_9236,N_6867,N_6671);
and U9237 (N_9237,N_7097,N_7820);
nor U9238 (N_9238,N_6084,N_7510);
or U9239 (N_9239,N_7202,N_7883);
or U9240 (N_9240,N_6642,N_6325);
and U9241 (N_9241,N_6035,N_7284);
nand U9242 (N_9242,N_6900,N_7598);
or U9243 (N_9243,N_7170,N_7127);
or U9244 (N_9244,N_6178,N_7997);
nor U9245 (N_9245,N_6850,N_6332);
nand U9246 (N_9246,N_7094,N_7866);
nand U9247 (N_9247,N_6295,N_6651);
and U9248 (N_9248,N_6870,N_7171);
nand U9249 (N_9249,N_6343,N_6510);
and U9250 (N_9250,N_6105,N_6759);
or U9251 (N_9251,N_7204,N_7920);
or U9252 (N_9252,N_7681,N_7541);
or U9253 (N_9253,N_6784,N_7363);
nor U9254 (N_9254,N_7760,N_7776);
nor U9255 (N_9255,N_7877,N_7202);
nor U9256 (N_9256,N_7082,N_7466);
and U9257 (N_9257,N_7349,N_6442);
nor U9258 (N_9258,N_7334,N_6866);
or U9259 (N_9259,N_7879,N_6423);
nor U9260 (N_9260,N_7200,N_7527);
nor U9261 (N_9261,N_6309,N_6695);
nor U9262 (N_9262,N_7558,N_7876);
and U9263 (N_9263,N_6486,N_7339);
and U9264 (N_9264,N_6301,N_6805);
and U9265 (N_9265,N_7209,N_6775);
or U9266 (N_9266,N_7419,N_7052);
nor U9267 (N_9267,N_7317,N_7842);
nor U9268 (N_9268,N_6810,N_6745);
or U9269 (N_9269,N_6311,N_6810);
nand U9270 (N_9270,N_6399,N_7721);
and U9271 (N_9271,N_6214,N_7936);
nand U9272 (N_9272,N_7046,N_7456);
nor U9273 (N_9273,N_7013,N_7838);
and U9274 (N_9274,N_6173,N_7892);
nor U9275 (N_9275,N_7106,N_6631);
nor U9276 (N_9276,N_7802,N_7065);
and U9277 (N_9277,N_7703,N_6957);
and U9278 (N_9278,N_7762,N_6829);
and U9279 (N_9279,N_6677,N_7314);
or U9280 (N_9280,N_7848,N_7074);
and U9281 (N_9281,N_6747,N_6263);
nor U9282 (N_9282,N_6659,N_7912);
nor U9283 (N_9283,N_6692,N_6279);
or U9284 (N_9284,N_7671,N_6629);
and U9285 (N_9285,N_7647,N_7946);
nor U9286 (N_9286,N_7711,N_6130);
and U9287 (N_9287,N_6893,N_6789);
nand U9288 (N_9288,N_6525,N_7712);
nand U9289 (N_9289,N_6260,N_7425);
or U9290 (N_9290,N_6401,N_7799);
and U9291 (N_9291,N_7681,N_6235);
nor U9292 (N_9292,N_7975,N_6763);
and U9293 (N_9293,N_7873,N_7065);
or U9294 (N_9294,N_6661,N_7028);
nor U9295 (N_9295,N_7960,N_7170);
or U9296 (N_9296,N_7135,N_6186);
and U9297 (N_9297,N_7502,N_7760);
nand U9298 (N_9298,N_7539,N_6209);
nand U9299 (N_9299,N_6040,N_6369);
or U9300 (N_9300,N_7104,N_6123);
and U9301 (N_9301,N_7666,N_7524);
nand U9302 (N_9302,N_7491,N_7584);
nor U9303 (N_9303,N_7174,N_7656);
nand U9304 (N_9304,N_6209,N_6399);
and U9305 (N_9305,N_6978,N_6773);
nor U9306 (N_9306,N_6064,N_7738);
nand U9307 (N_9307,N_7681,N_7112);
and U9308 (N_9308,N_7331,N_6815);
or U9309 (N_9309,N_6032,N_7661);
and U9310 (N_9310,N_7145,N_6574);
nand U9311 (N_9311,N_7759,N_6186);
nor U9312 (N_9312,N_7414,N_6024);
and U9313 (N_9313,N_7120,N_7122);
nor U9314 (N_9314,N_7924,N_7460);
or U9315 (N_9315,N_7430,N_6322);
nor U9316 (N_9316,N_7119,N_6093);
nor U9317 (N_9317,N_7480,N_7455);
nor U9318 (N_9318,N_7418,N_6212);
nor U9319 (N_9319,N_7473,N_6333);
nor U9320 (N_9320,N_7314,N_7108);
nand U9321 (N_9321,N_6653,N_7335);
or U9322 (N_9322,N_6388,N_7132);
and U9323 (N_9323,N_7928,N_6816);
nand U9324 (N_9324,N_7098,N_6524);
nor U9325 (N_9325,N_7112,N_6353);
nand U9326 (N_9326,N_7568,N_6960);
nor U9327 (N_9327,N_6788,N_6011);
xnor U9328 (N_9328,N_6235,N_7685);
nor U9329 (N_9329,N_6710,N_6706);
nand U9330 (N_9330,N_6253,N_7368);
nor U9331 (N_9331,N_6123,N_6524);
nor U9332 (N_9332,N_7911,N_6492);
nor U9333 (N_9333,N_6737,N_7823);
and U9334 (N_9334,N_6228,N_6489);
nor U9335 (N_9335,N_7806,N_7673);
nand U9336 (N_9336,N_6448,N_6954);
or U9337 (N_9337,N_6509,N_6350);
nor U9338 (N_9338,N_6816,N_6872);
nor U9339 (N_9339,N_6478,N_6690);
nand U9340 (N_9340,N_6679,N_6367);
and U9341 (N_9341,N_7120,N_7209);
nor U9342 (N_9342,N_6399,N_7621);
and U9343 (N_9343,N_7376,N_7930);
nand U9344 (N_9344,N_7798,N_7095);
or U9345 (N_9345,N_7084,N_7581);
nand U9346 (N_9346,N_7565,N_7829);
nor U9347 (N_9347,N_6832,N_6260);
nand U9348 (N_9348,N_6688,N_7703);
or U9349 (N_9349,N_7287,N_6832);
nor U9350 (N_9350,N_7527,N_6432);
and U9351 (N_9351,N_7129,N_7970);
nand U9352 (N_9352,N_7633,N_6050);
nand U9353 (N_9353,N_6311,N_6425);
nand U9354 (N_9354,N_7421,N_6275);
nand U9355 (N_9355,N_7589,N_6888);
nand U9356 (N_9356,N_7389,N_7183);
nor U9357 (N_9357,N_6553,N_7970);
or U9358 (N_9358,N_6990,N_7027);
and U9359 (N_9359,N_6801,N_6690);
nand U9360 (N_9360,N_7174,N_7712);
nor U9361 (N_9361,N_6332,N_6974);
or U9362 (N_9362,N_6404,N_7860);
or U9363 (N_9363,N_7117,N_6377);
or U9364 (N_9364,N_6271,N_6320);
nor U9365 (N_9365,N_7686,N_6249);
nor U9366 (N_9366,N_7829,N_7138);
nor U9367 (N_9367,N_6102,N_6843);
nor U9368 (N_9368,N_7974,N_7785);
nand U9369 (N_9369,N_6484,N_7757);
nor U9370 (N_9370,N_7092,N_6736);
nand U9371 (N_9371,N_7558,N_6614);
and U9372 (N_9372,N_7897,N_6601);
and U9373 (N_9373,N_7350,N_7242);
or U9374 (N_9374,N_7567,N_7931);
nand U9375 (N_9375,N_7057,N_6777);
nand U9376 (N_9376,N_7965,N_7364);
nand U9377 (N_9377,N_7408,N_6324);
nor U9378 (N_9378,N_6948,N_6833);
or U9379 (N_9379,N_6691,N_7023);
or U9380 (N_9380,N_7409,N_7229);
nor U9381 (N_9381,N_7410,N_7510);
nor U9382 (N_9382,N_7119,N_6899);
nor U9383 (N_9383,N_7415,N_7354);
nor U9384 (N_9384,N_7040,N_6090);
and U9385 (N_9385,N_7184,N_7817);
nand U9386 (N_9386,N_7331,N_6996);
and U9387 (N_9387,N_6413,N_7010);
and U9388 (N_9388,N_7522,N_7055);
and U9389 (N_9389,N_6724,N_6706);
nand U9390 (N_9390,N_7666,N_7920);
or U9391 (N_9391,N_6217,N_6144);
nand U9392 (N_9392,N_7100,N_7228);
or U9393 (N_9393,N_7589,N_7140);
nor U9394 (N_9394,N_7033,N_7437);
and U9395 (N_9395,N_6643,N_7638);
or U9396 (N_9396,N_7257,N_7833);
nand U9397 (N_9397,N_7803,N_6131);
nand U9398 (N_9398,N_6811,N_6411);
nor U9399 (N_9399,N_7135,N_7842);
nor U9400 (N_9400,N_7099,N_6941);
nor U9401 (N_9401,N_7765,N_7303);
nand U9402 (N_9402,N_7881,N_6848);
and U9403 (N_9403,N_7918,N_7665);
and U9404 (N_9404,N_7639,N_6159);
nor U9405 (N_9405,N_6068,N_7905);
nor U9406 (N_9406,N_6843,N_6829);
nor U9407 (N_9407,N_6138,N_7504);
nor U9408 (N_9408,N_6714,N_6659);
nor U9409 (N_9409,N_6421,N_6907);
or U9410 (N_9410,N_7802,N_6709);
or U9411 (N_9411,N_7238,N_6847);
or U9412 (N_9412,N_7570,N_6569);
nand U9413 (N_9413,N_7052,N_7075);
and U9414 (N_9414,N_6736,N_7730);
xor U9415 (N_9415,N_6597,N_7334);
and U9416 (N_9416,N_6033,N_6979);
nand U9417 (N_9417,N_7346,N_6811);
nand U9418 (N_9418,N_7971,N_7138);
nand U9419 (N_9419,N_7259,N_7427);
or U9420 (N_9420,N_6013,N_6331);
nor U9421 (N_9421,N_6169,N_7562);
nand U9422 (N_9422,N_7952,N_7362);
nand U9423 (N_9423,N_7938,N_6798);
nand U9424 (N_9424,N_6490,N_7501);
and U9425 (N_9425,N_6227,N_6320);
or U9426 (N_9426,N_7411,N_7880);
or U9427 (N_9427,N_6955,N_6396);
and U9428 (N_9428,N_7313,N_6098);
nand U9429 (N_9429,N_7397,N_7846);
and U9430 (N_9430,N_7735,N_7924);
and U9431 (N_9431,N_6262,N_6637);
or U9432 (N_9432,N_7930,N_6631);
nor U9433 (N_9433,N_7126,N_6475);
nor U9434 (N_9434,N_7408,N_6654);
and U9435 (N_9435,N_7300,N_7332);
and U9436 (N_9436,N_7726,N_6357);
or U9437 (N_9437,N_6944,N_6992);
nand U9438 (N_9438,N_6782,N_6085);
nand U9439 (N_9439,N_7770,N_7027);
nor U9440 (N_9440,N_6282,N_7950);
nor U9441 (N_9441,N_7599,N_7109);
nor U9442 (N_9442,N_6979,N_7701);
or U9443 (N_9443,N_7292,N_6578);
and U9444 (N_9444,N_6963,N_7250);
nand U9445 (N_9445,N_7065,N_7894);
and U9446 (N_9446,N_7420,N_6114);
or U9447 (N_9447,N_6166,N_7735);
and U9448 (N_9448,N_7021,N_6883);
or U9449 (N_9449,N_6452,N_7526);
nor U9450 (N_9450,N_7525,N_6249);
and U9451 (N_9451,N_7411,N_6599);
nor U9452 (N_9452,N_6462,N_7176);
and U9453 (N_9453,N_7842,N_6379);
nand U9454 (N_9454,N_6282,N_7859);
or U9455 (N_9455,N_6870,N_6550);
nor U9456 (N_9456,N_7533,N_7027);
nor U9457 (N_9457,N_6472,N_7105);
or U9458 (N_9458,N_7946,N_6073);
and U9459 (N_9459,N_6037,N_6642);
nand U9460 (N_9460,N_6842,N_6346);
nor U9461 (N_9461,N_6734,N_6335);
and U9462 (N_9462,N_7897,N_6851);
nor U9463 (N_9463,N_6517,N_6632);
nand U9464 (N_9464,N_6477,N_6616);
nor U9465 (N_9465,N_6882,N_7343);
nand U9466 (N_9466,N_6082,N_6124);
and U9467 (N_9467,N_7266,N_7640);
nor U9468 (N_9468,N_6826,N_6422);
nand U9469 (N_9469,N_7668,N_7977);
and U9470 (N_9470,N_7448,N_6212);
xor U9471 (N_9471,N_7268,N_7732);
xnor U9472 (N_9472,N_6254,N_6260);
or U9473 (N_9473,N_7268,N_7129);
or U9474 (N_9474,N_6716,N_7192);
and U9475 (N_9475,N_7687,N_7748);
or U9476 (N_9476,N_7657,N_7349);
nand U9477 (N_9477,N_7848,N_6546);
nand U9478 (N_9478,N_6886,N_6914);
or U9479 (N_9479,N_6971,N_7929);
and U9480 (N_9480,N_7160,N_6159);
nor U9481 (N_9481,N_7922,N_7611);
nor U9482 (N_9482,N_7602,N_6875);
nand U9483 (N_9483,N_7614,N_6293);
and U9484 (N_9484,N_6028,N_6690);
and U9485 (N_9485,N_6713,N_6808);
nor U9486 (N_9486,N_6007,N_7659);
and U9487 (N_9487,N_6211,N_7484);
and U9488 (N_9488,N_6410,N_6000);
or U9489 (N_9489,N_6332,N_6431);
or U9490 (N_9490,N_6606,N_7967);
nand U9491 (N_9491,N_7084,N_6725);
nand U9492 (N_9492,N_6586,N_7732);
or U9493 (N_9493,N_6688,N_7268);
nor U9494 (N_9494,N_7082,N_6010);
nand U9495 (N_9495,N_6278,N_6352);
or U9496 (N_9496,N_6556,N_6004);
nor U9497 (N_9497,N_7418,N_7696);
nand U9498 (N_9498,N_7343,N_6201);
nand U9499 (N_9499,N_7382,N_7275);
and U9500 (N_9500,N_6858,N_6037);
and U9501 (N_9501,N_7592,N_7403);
or U9502 (N_9502,N_7692,N_6211);
nor U9503 (N_9503,N_6244,N_7777);
nor U9504 (N_9504,N_6068,N_7453);
or U9505 (N_9505,N_7751,N_6556);
nand U9506 (N_9506,N_7514,N_6784);
and U9507 (N_9507,N_7079,N_6841);
and U9508 (N_9508,N_7942,N_7488);
nor U9509 (N_9509,N_7714,N_6918);
nor U9510 (N_9510,N_7314,N_6543);
nand U9511 (N_9511,N_7215,N_7867);
and U9512 (N_9512,N_7952,N_6653);
nand U9513 (N_9513,N_7077,N_6058);
nand U9514 (N_9514,N_7520,N_7755);
nand U9515 (N_9515,N_7373,N_6286);
or U9516 (N_9516,N_6105,N_6180);
and U9517 (N_9517,N_7927,N_7699);
or U9518 (N_9518,N_7185,N_7925);
or U9519 (N_9519,N_6205,N_7278);
nor U9520 (N_9520,N_6989,N_7320);
nor U9521 (N_9521,N_6024,N_7082);
or U9522 (N_9522,N_6105,N_6508);
or U9523 (N_9523,N_7095,N_7601);
or U9524 (N_9524,N_7221,N_6248);
and U9525 (N_9525,N_6148,N_6718);
or U9526 (N_9526,N_6088,N_6782);
nor U9527 (N_9527,N_7530,N_7418);
or U9528 (N_9528,N_6416,N_7819);
nand U9529 (N_9529,N_7327,N_6759);
nand U9530 (N_9530,N_7386,N_6908);
or U9531 (N_9531,N_7951,N_6137);
and U9532 (N_9532,N_7676,N_6434);
nor U9533 (N_9533,N_7419,N_7071);
or U9534 (N_9534,N_6788,N_6149);
nand U9535 (N_9535,N_6168,N_6615);
or U9536 (N_9536,N_6437,N_6509);
or U9537 (N_9537,N_6686,N_6975);
nor U9538 (N_9538,N_7656,N_7592);
nor U9539 (N_9539,N_6419,N_7844);
nor U9540 (N_9540,N_6229,N_6127);
nand U9541 (N_9541,N_7166,N_7346);
nor U9542 (N_9542,N_7132,N_6183);
nand U9543 (N_9543,N_6982,N_7747);
nor U9544 (N_9544,N_6081,N_6282);
or U9545 (N_9545,N_6360,N_7591);
or U9546 (N_9546,N_7977,N_6156);
and U9547 (N_9547,N_7773,N_7143);
nor U9548 (N_9548,N_7588,N_7320);
or U9549 (N_9549,N_6282,N_7523);
and U9550 (N_9550,N_6718,N_7790);
nor U9551 (N_9551,N_7997,N_7550);
xor U9552 (N_9552,N_6830,N_7448);
nand U9553 (N_9553,N_6598,N_7986);
and U9554 (N_9554,N_7374,N_6123);
and U9555 (N_9555,N_6706,N_6353);
nor U9556 (N_9556,N_7753,N_7327);
nand U9557 (N_9557,N_7365,N_6679);
nor U9558 (N_9558,N_6536,N_6272);
nand U9559 (N_9559,N_6925,N_6876);
nand U9560 (N_9560,N_6817,N_7473);
nand U9561 (N_9561,N_6611,N_7785);
or U9562 (N_9562,N_6798,N_6836);
nor U9563 (N_9563,N_6393,N_7556);
nor U9564 (N_9564,N_7132,N_6401);
nand U9565 (N_9565,N_7190,N_6365);
nand U9566 (N_9566,N_7466,N_6135);
nor U9567 (N_9567,N_6393,N_7108);
nor U9568 (N_9568,N_6320,N_6785);
or U9569 (N_9569,N_6418,N_6571);
nor U9570 (N_9570,N_7230,N_7452);
nand U9571 (N_9571,N_6991,N_6844);
nand U9572 (N_9572,N_7328,N_6409);
nand U9573 (N_9573,N_7642,N_6904);
nor U9574 (N_9574,N_6184,N_6533);
and U9575 (N_9575,N_7570,N_6287);
and U9576 (N_9576,N_7648,N_6298);
nand U9577 (N_9577,N_6306,N_7702);
and U9578 (N_9578,N_6037,N_7868);
nor U9579 (N_9579,N_7679,N_6017);
nand U9580 (N_9580,N_6025,N_7774);
and U9581 (N_9581,N_6714,N_7441);
nand U9582 (N_9582,N_7001,N_6303);
nor U9583 (N_9583,N_7437,N_6240);
nand U9584 (N_9584,N_7161,N_6159);
or U9585 (N_9585,N_7916,N_6963);
or U9586 (N_9586,N_6127,N_6377);
nand U9587 (N_9587,N_7677,N_7057);
nor U9588 (N_9588,N_6398,N_7132);
and U9589 (N_9589,N_6200,N_7710);
and U9590 (N_9590,N_7958,N_7032);
and U9591 (N_9591,N_7737,N_7970);
nand U9592 (N_9592,N_7572,N_7545);
or U9593 (N_9593,N_6554,N_7517);
nor U9594 (N_9594,N_7123,N_6102);
nand U9595 (N_9595,N_6656,N_6194);
and U9596 (N_9596,N_6388,N_7002);
nand U9597 (N_9597,N_6257,N_7961);
nor U9598 (N_9598,N_7159,N_6364);
nor U9599 (N_9599,N_6786,N_7372);
nor U9600 (N_9600,N_7664,N_6498);
or U9601 (N_9601,N_7938,N_6278);
nand U9602 (N_9602,N_6433,N_6863);
or U9603 (N_9603,N_6043,N_6948);
or U9604 (N_9604,N_6924,N_7617);
nor U9605 (N_9605,N_7870,N_7427);
and U9606 (N_9606,N_7379,N_7832);
and U9607 (N_9607,N_7509,N_7860);
or U9608 (N_9608,N_6299,N_6743);
or U9609 (N_9609,N_6582,N_7767);
nor U9610 (N_9610,N_6004,N_7752);
nand U9611 (N_9611,N_6241,N_6279);
or U9612 (N_9612,N_7321,N_7368);
and U9613 (N_9613,N_6011,N_7369);
nand U9614 (N_9614,N_7295,N_6113);
nand U9615 (N_9615,N_6668,N_6364);
nor U9616 (N_9616,N_7904,N_6509);
nand U9617 (N_9617,N_7237,N_6141);
and U9618 (N_9618,N_6710,N_6910);
nor U9619 (N_9619,N_7069,N_7056);
or U9620 (N_9620,N_6152,N_6552);
and U9621 (N_9621,N_7352,N_6122);
xor U9622 (N_9622,N_6212,N_6601);
and U9623 (N_9623,N_6017,N_6883);
and U9624 (N_9624,N_7922,N_6993);
and U9625 (N_9625,N_6824,N_7292);
nor U9626 (N_9626,N_6667,N_7594);
or U9627 (N_9627,N_7722,N_7932);
or U9628 (N_9628,N_7075,N_7678);
nand U9629 (N_9629,N_7423,N_6412);
or U9630 (N_9630,N_6865,N_6754);
nand U9631 (N_9631,N_7512,N_6894);
and U9632 (N_9632,N_7819,N_6232);
nand U9633 (N_9633,N_6455,N_6836);
nand U9634 (N_9634,N_6885,N_7263);
and U9635 (N_9635,N_7577,N_6867);
nor U9636 (N_9636,N_6367,N_7804);
or U9637 (N_9637,N_7601,N_7172);
nor U9638 (N_9638,N_7904,N_7951);
nand U9639 (N_9639,N_6480,N_6290);
and U9640 (N_9640,N_6264,N_6852);
and U9641 (N_9641,N_7954,N_7596);
xnor U9642 (N_9642,N_7741,N_7573);
nand U9643 (N_9643,N_7102,N_6851);
and U9644 (N_9644,N_7560,N_7485);
nor U9645 (N_9645,N_6158,N_7312);
and U9646 (N_9646,N_7754,N_6516);
nand U9647 (N_9647,N_6969,N_6736);
nor U9648 (N_9648,N_7068,N_6247);
xor U9649 (N_9649,N_6118,N_6710);
or U9650 (N_9650,N_6415,N_6380);
and U9651 (N_9651,N_7880,N_6424);
and U9652 (N_9652,N_7633,N_6833);
or U9653 (N_9653,N_6068,N_7181);
and U9654 (N_9654,N_7205,N_6608);
or U9655 (N_9655,N_6860,N_6513);
nor U9656 (N_9656,N_7498,N_7816);
and U9657 (N_9657,N_6526,N_7165);
or U9658 (N_9658,N_6233,N_6824);
and U9659 (N_9659,N_6676,N_7127);
nand U9660 (N_9660,N_7120,N_7642);
nor U9661 (N_9661,N_7274,N_7476);
or U9662 (N_9662,N_6019,N_7168);
or U9663 (N_9663,N_7152,N_6223);
nor U9664 (N_9664,N_6653,N_7191);
xor U9665 (N_9665,N_6861,N_7361);
or U9666 (N_9666,N_6534,N_6758);
or U9667 (N_9667,N_6348,N_7079);
or U9668 (N_9668,N_6748,N_7027);
xor U9669 (N_9669,N_7027,N_7911);
or U9670 (N_9670,N_7922,N_7322);
nand U9671 (N_9671,N_6622,N_6208);
or U9672 (N_9672,N_6027,N_6883);
nand U9673 (N_9673,N_7413,N_6212);
or U9674 (N_9674,N_7346,N_6525);
nand U9675 (N_9675,N_6107,N_7397);
nor U9676 (N_9676,N_6434,N_6291);
nand U9677 (N_9677,N_7425,N_6308);
or U9678 (N_9678,N_6779,N_7231);
nor U9679 (N_9679,N_7950,N_6796);
nor U9680 (N_9680,N_6024,N_6693);
nand U9681 (N_9681,N_6277,N_6760);
nand U9682 (N_9682,N_6821,N_6477);
or U9683 (N_9683,N_6065,N_7076);
and U9684 (N_9684,N_6767,N_6742);
or U9685 (N_9685,N_7964,N_7543);
nand U9686 (N_9686,N_6799,N_6570);
nor U9687 (N_9687,N_6048,N_6756);
or U9688 (N_9688,N_6732,N_7089);
or U9689 (N_9689,N_6324,N_6166);
nor U9690 (N_9690,N_7578,N_6111);
nor U9691 (N_9691,N_7749,N_7233);
nor U9692 (N_9692,N_7878,N_6054);
nand U9693 (N_9693,N_7948,N_6121);
nor U9694 (N_9694,N_7446,N_6806);
or U9695 (N_9695,N_7625,N_7196);
and U9696 (N_9696,N_6276,N_6013);
nand U9697 (N_9697,N_6889,N_6533);
and U9698 (N_9698,N_6602,N_7120);
nand U9699 (N_9699,N_7475,N_6996);
nand U9700 (N_9700,N_6342,N_7497);
or U9701 (N_9701,N_6267,N_6902);
and U9702 (N_9702,N_6470,N_7985);
and U9703 (N_9703,N_6845,N_6055);
nand U9704 (N_9704,N_7048,N_6265);
nor U9705 (N_9705,N_6883,N_7975);
nor U9706 (N_9706,N_7436,N_6637);
nand U9707 (N_9707,N_7385,N_6314);
or U9708 (N_9708,N_7100,N_6864);
nand U9709 (N_9709,N_6070,N_7454);
nor U9710 (N_9710,N_7431,N_6186);
and U9711 (N_9711,N_7216,N_6188);
and U9712 (N_9712,N_6592,N_6284);
nor U9713 (N_9713,N_6303,N_7235);
nand U9714 (N_9714,N_7380,N_7468);
and U9715 (N_9715,N_7505,N_6411);
nor U9716 (N_9716,N_7933,N_6544);
or U9717 (N_9717,N_6993,N_6592);
and U9718 (N_9718,N_7703,N_7591);
nor U9719 (N_9719,N_6945,N_6795);
and U9720 (N_9720,N_6963,N_7212);
or U9721 (N_9721,N_7340,N_6357);
and U9722 (N_9722,N_6520,N_6134);
nor U9723 (N_9723,N_6320,N_7727);
nand U9724 (N_9724,N_6076,N_7711);
or U9725 (N_9725,N_6331,N_6570);
and U9726 (N_9726,N_6466,N_6561);
and U9727 (N_9727,N_7501,N_6244);
and U9728 (N_9728,N_6416,N_7032);
or U9729 (N_9729,N_7816,N_7184);
or U9730 (N_9730,N_6258,N_6704);
nor U9731 (N_9731,N_6783,N_7759);
or U9732 (N_9732,N_7646,N_7991);
or U9733 (N_9733,N_6406,N_7949);
or U9734 (N_9734,N_6164,N_7566);
nand U9735 (N_9735,N_7559,N_7215);
or U9736 (N_9736,N_7028,N_7633);
nand U9737 (N_9737,N_7964,N_7412);
nor U9738 (N_9738,N_6539,N_6782);
or U9739 (N_9739,N_7371,N_6865);
and U9740 (N_9740,N_7794,N_7608);
and U9741 (N_9741,N_7477,N_7501);
or U9742 (N_9742,N_6223,N_7944);
nand U9743 (N_9743,N_7986,N_6917);
and U9744 (N_9744,N_6632,N_7084);
nor U9745 (N_9745,N_7572,N_7971);
nand U9746 (N_9746,N_7977,N_6408);
or U9747 (N_9747,N_6312,N_6512);
nor U9748 (N_9748,N_6340,N_7575);
nand U9749 (N_9749,N_7658,N_6827);
nor U9750 (N_9750,N_7457,N_6896);
or U9751 (N_9751,N_7375,N_7112);
nor U9752 (N_9752,N_7028,N_7484);
nor U9753 (N_9753,N_7457,N_6981);
xor U9754 (N_9754,N_7396,N_7551);
xor U9755 (N_9755,N_7515,N_7064);
nand U9756 (N_9756,N_7181,N_7240);
nand U9757 (N_9757,N_6652,N_6057);
nand U9758 (N_9758,N_7291,N_7726);
or U9759 (N_9759,N_7575,N_6493);
and U9760 (N_9760,N_7613,N_7679);
nand U9761 (N_9761,N_6072,N_6341);
and U9762 (N_9762,N_6168,N_7189);
nand U9763 (N_9763,N_6781,N_7712);
nand U9764 (N_9764,N_6954,N_6650);
nor U9765 (N_9765,N_7963,N_7872);
nand U9766 (N_9766,N_7113,N_7048);
and U9767 (N_9767,N_6370,N_6898);
nor U9768 (N_9768,N_6347,N_7766);
or U9769 (N_9769,N_7728,N_7358);
nand U9770 (N_9770,N_6155,N_7533);
or U9771 (N_9771,N_6493,N_6354);
or U9772 (N_9772,N_6606,N_7657);
nor U9773 (N_9773,N_6201,N_6142);
and U9774 (N_9774,N_6002,N_6225);
nor U9775 (N_9775,N_7413,N_7814);
or U9776 (N_9776,N_6368,N_6926);
or U9777 (N_9777,N_7593,N_6012);
nor U9778 (N_9778,N_6941,N_7175);
and U9779 (N_9779,N_6501,N_7663);
and U9780 (N_9780,N_6154,N_6668);
or U9781 (N_9781,N_6822,N_7266);
nor U9782 (N_9782,N_7914,N_7347);
nand U9783 (N_9783,N_7131,N_7797);
nand U9784 (N_9784,N_6577,N_6361);
or U9785 (N_9785,N_7084,N_6102);
and U9786 (N_9786,N_7032,N_6480);
nor U9787 (N_9787,N_7091,N_7666);
nor U9788 (N_9788,N_6828,N_7835);
and U9789 (N_9789,N_7122,N_7420);
nand U9790 (N_9790,N_6278,N_6748);
or U9791 (N_9791,N_6002,N_6273);
nand U9792 (N_9792,N_6332,N_6322);
nand U9793 (N_9793,N_7318,N_7303);
or U9794 (N_9794,N_6577,N_7071);
and U9795 (N_9795,N_7759,N_6942);
nand U9796 (N_9796,N_7187,N_6774);
nand U9797 (N_9797,N_6088,N_6116);
nand U9798 (N_9798,N_7768,N_7188);
and U9799 (N_9799,N_6361,N_7426);
and U9800 (N_9800,N_7635,N_7498);
nand U9801 (N_9801,N_6543,N_7235);
nand U9802 (N_9802,N_6862,N_6616);
or U9803 (N_9803,N_7502,N_7440);
nand U9804 (N_9804,N_6013,N_6839);
nand U9805 (N_9805,N_6717,N_6974);
nor U9806 (N_9806,N_7121,N_7106);
nor U9807 (N_9807,N_7349,N_6780);
or U9808 (N_9808,N_6167,N_7062);
and U9809 (N_9809,N_7213,N_7112);
and U9810 (N_9810,N_6198,N_6954);
or U9811 (N_9811,N_7542,N_6709);
or U9812 (N_9812,N_6861,N_7260);
nor U9813 (N_9813,N_6684,N_7004);
nand U9814 (N_9814,N_6212,N_6991);
nor U9815 (N_9815,N_6539,N_7777);
nor U9816 (N_9816,N_7308,N_7398);
or U9817 (N_9817,N_6396,N_7169);
nand U9818 (N_9818,N_6074,N_6537);
nor U9819 (N_9819,N_6756,N_6500);
nand U9820 (N_9820,N_6403,N_7530);
nor U9821 (N_9821,N_7526,N_6459);
nand U9822 (N_9822,N_6616,N_6515);
nor U9823 (N_9823,N_7073,N_6635);
nor U9824 (N_9824,N_6097,N_6662);
nor U9825 (N_9825,N_7361,N_7420);
or U9826 (N_9826,N_6702,N_6746);
nand U9827 (N_9827,N_6584,N_7377);
or U9828 (N_9828,N_7184,N_6577);
or U9829 (N_9829,N_6436,N_7197);
nand U9830 (N_9830,N_6381,N_6109);
and U9831 (N_9831,N_7069,N_6405);
nand U9832 (N_9832,N_6821,N_6651);
nand U9833 (N_9833,N_6608,N_7234);
and U9834 (N_9834,N_7984,N_7562);
nand U9835 (N_9835,N_6240,N_6280);
nor U9836 (N_9836,N_6225,N_7742);
and U9837 (N_9837,N_7163,N_7542);
or U9838 (N_9838,N_7505,N_6665);
nor U9839 (N_9839,N_7178,N_6882);
nand U9840 (N_9840,N_7726,N_6878);
nor U9841 (N_9841,N_7682,N_6901);
or U9842 (N_9842,N_6377,N_6856);
and U9843 (N_9843,N_7738,N_6980);
nor U9844 (N_9844,N_7748,N_7156);
nor U9845 (N_9845,N_6019,N_7375);
nand U9846 (N_9846,N_6952,N_6620);
nand U9847 (N_9847,N_7216,N_6487);
nor U9848 (N_9848,N_6721,N_6920);
nor U9849 (N_9849,N_6853,N_6502);
or U9850 (N_9850,N_6968,N_6760);
and U9851 (N_9851,N_7241,N_6210);
nand U9852 (N_9852,N_7129,N_7146);
and U9853 (N_9853,N_6774,N_6465);
or U9854 (N_9854,N_6908,N_7921);
or U9855 (N_9855,N_7675,N_6803);
and U9856 (N_9856,N_6286,N_7794);
or U9857 (N_9857,N_6156,N_7748);
or U9858 (N_9858,N_6556,N_6245);
or U9859 (N_9859,N_6599,N_6044);
and U9860 (N_9860,N_6101,N_7526);
and U9861 (N_9861,N_7542,N_6714);
and U9862 (N_9862,N_6927,N_6083);
and U9863 (N_9863,N_6823,N_7859);
and U9864 (N_9864,N_7337,N_6851);
nand U9865 (N_9865,N_7201,N_6176);
or U9866 (N_9866,N_7845,N_6684);
nor U9867 (N_9867,N_7172,N_7946);
nand U9868 (N_9868,N_7184,N_7230);
nor U9869 (N_9869,N_7501,N_6159);
and U9870 (N_9870,N_7191,N_7929);
or U9871 (N_9871,N_7358,N_7999);
nor U9872 (N_9872,N_6880,N_6953);
nand U9873 (N_9873,N_7141,N_6462);
nand U9874 (N_9874,N_7312,N_7249);
and U9875 (N_9875,N_7493,N_6200);
nor U9876 (N_9876,N_6915,N_6340);
nand U9877 (N_9877,N_7400,N_6795);
or U9878 (N_9878,N_7245,N_6760);
nor U9879 (N_9879,N_6415,N_7379);
and U9880 (N_9880,N_6756,N_7933);
nand U9881 (N_9881,N_7954,N_7750);
nand U9882 (N_9882,N_6030,N_6340);
or U9883 (N_9883,N_6878,N_7285);
or U9884 (N_9884,N_7681,N_6284);
or U9885 (N_9885,N_7181,N_7729);
nor U9886 (N_9886,N_7386,N_7414);
or U9887 (N_9887,N_6919,N_7867);
and U9888 (N_9888,N_7572,N_7575);
or U9889 (N_9889,N_7364,N_7716);
nor U9890 (N_9890,N_6358,N_6507);
nand U9891 (N_9891,N_7804,N_6696);
or U9892 (N_9892,N_7857,N_6584);
and U9893 (N_9893,N_6167,N_6288);
or U9894 (N_9894,N_7548,N_7709);
nor U9895 (N_9895,N_7646,N_7502);
or U9896 (N_9896,N_7769,N_6266);
and U9897 (N_9897,N_6525,N_6483);
nand U9898 (N_9898,N_6964,N_6987);
nand U9899 (N_9899,N_7389,N_7460);
and U9900 (N_9900,N_6760,N_6067);
or U9901 (N_9901,N_6576,N_7376);
and U9902 (N_9902,N_7064,N_6155);
and U9903 (N_9903,N_7765,N_7304);
or U9904 (N_9904,N_6716,N_7286);
xnor U9905 (N_9905,N_7865,N_6490);
or U9906 (N_9906,N_6709,N_7398);
or U9907 (N_9907,N_7773,N_6932);
nand U9908 (N_9908,N_6652,N_7310);
and U9909 (N_9909,N_7774,N_7432);
nor U9910 (N_9910,N_7848,N_6943);
or U9911 (N_9911,N_7861,N_7453);
or U9912 (N_9912,N_7981,N_6595);
and U9913 (N_9913,N_6382,N_6781);
or U9914 (N_9914,N_6350,N_6531);
or U9915 (N_9915,N_6625,N_7210);
or U9916 (N_9916,N_6168,N_7762);
or U9917 (N_9917,N_6506,N_7048);
nor U9918 (N_9918,N_6742,N_6143);
or U9919 (N_9919,N_6029,N_6931);
or U9920 (N_9920,N_7625,N_7265);
and U9921 (N_9921,N_6637,N_6474);
nand U9922 (N_9922,N_6313,N_6167);
or U9923 (N_9923,N_7473,N_6014);
or U9924 (N_9924,N_7226,N_7417);
nor U9925 (N_9925,N_7183,N_6627);
or U9926 (N_9926,N_7520,N_7505);
and U9927 (N_9927,N_7116,N_6737);
or U9928 (N_9928,N_6931,N_6047);
or U9929 (N_9929,N_7952,N_7250);
nand U9930 (N_9930,N_6630,N_6578);
or U9931 (N_9931,N_7019,N_7632);
and U9932 (N_9932,N_6469,N_7500);
and U9933 (N_9933,N_6496,N_7929);
and U9934 (N_9934,N_7603,N_7202);
and U9935 (N_9935,N_7434,N_7253);
nor U9936 (N_9936,N_6062,N_6829);
nand U9937 (N_9937,N_6195,N_6540);
and U9938 (N_9938,N_6898,N_6278);
or U9939 (N_9939,N_6991,N_6953);
or U9940 (N_9940,N_7239,N_7820);
nor U9941 (N_9941,N_7758,N_7195);
or U9942 (N_9942,N_7038,N_7007);
nor U9943 (N_9943,N_6713,N_7766);
nand U9944 (N_9944,N_6126,N_6019);
and U9945 (N_9945,N_7597,N_7992);
and U9946 (N_9946,N_7449,N_7671);
or U9947 (N_9947,N_6374,N_6839);
nor U9948 (N_9948,N_7439,N_7589);
or U9949 (N_9949,N_7493,N_7244);
nor U9950 (N_9950,N_6209,N_6703);
nor U9951 (N_9951,N_7453,N_6144);
nand U9952 (N_9952,N_6248,N_7325);
and U9953 (N_9953,N_7517,N_6988);
and U9954 (N_9954,N_6937,N_6051);
nor U9955 (N_9955,N_6840,N_6558);
nand U9956 (N_9956,N_6882,N_7775);
or U9957 (N_9957,N_7202,N_6937);
nand U9958 (N_9958,N_7678,N_7297);
or U9959 (N_9959,N_7532,N_6276);
or U9960 (N_9960,N_6149,N_7179);
or U9961 (N_9961,N_7264,N_6821);
nand U9962 (N_9962,N_6580,N_7827);
or U9963 (N_9963,N_7464,N_6128);
or U9964 (N_9964,N_6986,N_7593);
and U9965 (N_9965,N_7853,N_6256);
nor U9966 (N_9966,N_7546,N_6852);
xnor U9967 (N_9967,N_6298,N_6969);
and U9968 (N_9968,N_6620,N_6115);
nor U9969 (N_9969,N_7102,N_7541);
nand U9970 (N_9970,N_7716,N_6620);
nand U9971 (N_9971,N_7088,N_7220);
nand U9972 (N_9972,N_7577,N_7526);
or U9973 (N_9973,N_7481,N_6454);
or U9974 (N_9974,N_7344,N_6031);
nor U9975 (N_9975,N_6120,N_7050);
nand U9976 (N_9976,N_6769,N_6861);
or U9977 (N_9977,N_6534,N_6058);
nor U9978 (N_9978,N_7411,N_6604);
nand U9979 (N_9979,N_6578,N_6792);
nor U9980 (N_9980,N_6032,N_7658);
and U9981 (N_9981,N_7981,N_7324);
nand U9982 (N_9982,N_7247,N_7521);
and U9983 (N_9983,N_6607,N_7674);
or U9984 (N_9984,N_6410,N_6759);
or U9985 (N_9985,N_7674,N_6981);
nand U9986 (N_9986,N_6809,N_7560);
nand U9987 (N_9987,N_6344,N_6895);
and U9988 (N_9988,N_6164,N_6358);
nand U9989 (N_9989,N_6921,N_7106);
nand U9990 (N_9990,N_7126,N_7187);
or U9991 (N_9991,N_7688,N_6271);
and U9992 (N_9992,N_6102,N_6716);
or U9993 (N_9993,N_7888,N_6342);
nor U9994 (N_9994,N_6475,N_6457);
nor U9995 (N_9995,N_7085,N_7487);
nor U9996 (N_9996,N_7265,N_7550);
nor U9997 (N_9997,N_6318,N_7426);
nor U9998 (N_9998,N_7665,N_6413);
xnor U9999 (N_9999,N_7641,N_7132);
nor UO_0 (O_0,N_8542,N_9382);
or UO_1 (O_1,N_9410,N_9997);
and UO_2 (O_2,N_8691,N_8842);
or UO_3 (O_3,N_8917,N_9046);
nor UO_4 (O_4,N_8744,N_9883);
or UO_5 (O_5,N_9842,N_9537);
and UO_6 (O_6,N_8574,N_8406);
nand UO_7 (O_7,N_8086,N_9792);
or UO_8 (O_8,N_8258,N_9300);
and UO_9 (O_9,N_8056,N_8407);
and UO_10 (O_10,N_8064,N_9404);
nor UO_11 (O_11,N_8414,N_8921);
or UO_12 (O_12,N_9444,N_9192);
and UO_13 (O_13,N_9779,N_9712);
or UO_14 (O_14,N_9502,N_8468);
nand UO_15 (O_15,N_9500,N_8969);
nand UO_16 (O_16,N_8730,N_9752);
nand UO_17 (O_17,N_9324,N_9281);
nand UO_18 (O_18,N_8853,N_9298);
or UO_19 (O_19,N_9828,N_9598);
or UO_20 (O_20,N_9418,N_8888);
nand UO_21 (O_21,N_9062,N_8837);
nand UO_22 (O_22,N_8732,N_9222);
nand UO_23 (O_23,N_9727,N_8368);
nand UO_24 (O_24,N_9487,N_9831);
nor UO_25 (O_25,N_9987,N_9659);
nand UO_26 (O_26,N_9636,N_8022);
or UO_27 (O_27,N_9611,N_8235);
nand UO_28 (O_28,N_8668,N_8637);
or UO_29 (O_29,N_8321,N_8452);
and UO_30 (O_30,N_9888,N_8309);
or UO_31 (O_31,N_9314,N_8536);
nand UO_32 (O_32,N_9120,N_9640);
nand UO_33 (O_33,N_9207,N_9844);
or UO_34 (O_34,N_9993,N_9103);
and UO_35 (O_35,N_9913,N_9294);
and UO_36 (O_36,N_9946,N_9902);
nand UO_37 (O_37,N_8051,N_9377);
nor UO_38 (O_38,N_9244,N_9512);
nand UO_39 (O_39,N_8008,N_8314);
and UO_40 (O_40,N_8857,N_9199);
nor UO_41 (O_41,N_9544,N_8750);
nand UO_42 (O_42,N_8769,N_8598);
xor UO_43 (O_43,N_8654,N_9671);
nor UO_44 (O_44,N_9220,N_9525);
and UO_45 (O_45,N_9271,N_8793);
nand UO_46 (O_46,N_9647,N_9134);
and UO_47 (O_47,N_9650,N_9925);
or UO_48 (O_48,N_9540,N_8320);
or UO_49 (O_49,N_9680,N_9228);
or UO_50 (O_50,N_9509,N_9375);
nand UO_51 (O_51,N_8829,N_8119);
nor UO_52 (O_52,N_8566,N_8285);
nor UO_53 (O_53,N_8313,N_8603);
or UO_54 (O_54,N_8231,N_8679);
and UO_55 (O_55,N_8948,N_9567);
nor UO_56 (O_56,N_8813,N_9168);
and UO_57 (O_57,N_8931,N_9612);
nor UO_58 (O_58,N_9604,N_9012);
nand UO_59 (O_59,N_9847,N_8913);
and UO_60 (O_60,N_9864,N_8239);
and UO_61 (O_61,N_8173,N_8800);
nand UO_62 (O_62,N_8593,N_9610);
or UO_63 (O_63,N_9665,N_9743);
and UO_64 (O_64,N_9411,N_9579);
or UO_65 (O_65,N_8601,N_9110);
or UO_66 (O_66,N_9463,N_9440);
and UO_67 (O_67,N_8815,N_9584);
and UO_68 (O_68,N_8812,N_9710);
or UO_69 (O_69,N_9292,N_9084);
or UO_70 (O_70,N_8473,N_9148);
nor UO_71 (O_71,N_8791,N_8934);
nand UO_72 (O_72,N_9362,N_8332);
nand UO_73 (O_73,N_8415,N_9036);
and UO_74 (O_74,N_8977,N_9080);
and UO_75 (O_75,N_9623,N_9033);
or UO_76 (O_76,N_9170,N_9725);
xor UO_77 (O_77,N_9398,N_8804);
or UO_78 (O_78,N_8605,N_9204);
and UO_79 (O_79,N_8297,N_9976);
or UO_80 (O_80,N_9672,N_9620);
and UO_81 (O_81,N_8018,N_9180);
or UO_82 (O_82,N_9153,N_8349);
nor UO_83 (O_83,N_8648,N_9102);
nand UO_84 (O_84,N_8042,N_9554);
and UO_85 (O_85,N_8659,N_8789);
and UO_86 (O_86,N_9215,N_9403);
and UO_87 (O_87,N_9285,N_8990);
and UO_88 (O_88,N_9218,N_9332);
and UO_89 (O_89,N_9662,N_9510);
nand UO_90 (O_90,N_9124,N_8463);
nor UO_91 (O_91,N_9852,N_9826);
and UO_92 (O_92,N_8446,N_9159);
and UO_93 (O_93,N_8865,N_8792);
and UO_94 (O_94,N_9704,N_9132);
and UO_95 (O_95,N_9821,N_8295);
or UO_96 (O_96,N_9034,N_8839);
or UO_97 (O_97,N_9870,N_9953);
nor UO_98 (O_98,N_8786,N_8643);
and UO_99 (O_99,N_9916,N_9786);
or UO_100 (O_100,N_9200,N_9967);
or UO_101 (O_101,N_9459,N_8568);
or UO_102 (O_102,N_9532,N_8366);
or UO_103 (O_103,N_9566,N_8634);
nor UO_104 (O_104,N_8535,N_8227);
and UO_105 (O_105,N_9855,N_9342);
nor UO_106 (O_106,N_8021,N_9890);
nand UO_107 (O_107,N_9470,N_9293);
xnor UO_108 (O_108,N_9058,N_9906);
and UO_109 (O_109,N_8633,N_9982);
or UO_110 (O_110,N_9301,N_9923);
and UO_111 (O_111,N_9988,N_9734);
nand UO_112 (O_112,N_8044,N_8094);
or UO_113 (O_113,N_8998,N_8631);
and UO_114 (O_114,N_8110,N_8331);
nor UO_115 (O_115,N_9594,N_8095);
and UO_116 (O_116,N_8203,N_8009);
nand UO_117 (O_117,N_9358,N_8287);
and UO_118 (O_118,N_9094,N_8030);
nor UO_119 (O_119,N_9771,N_8555);
or UO_120 (O_120,N_8395,N_8382);
or UO_121 (O_121,N_8393,N_9565);
nor UO_122 (O_122,N_9551,N_8509);
and UO_123 (O_123,N_9631,N_8143);
nor UO_124 (O_124,N_9678,N_8392);
or UO_125 (O_125,N_9969,N_9092);
nor UO_126 (O_126,N_9827,N_8184);
nor UO_127 (O_127,N_8667,N_8438);
or UO_128 (O_128,N_9360,N_9056);
nor UO_129 (O_129,N_9260,N_8486);
nor UO_130 (O_130,N_9331,N_9151);
nor UO_131 (O_131,N_9165,N_9885);
nor UO_132 (O_132,N_9624,N_9927);
nand UO_133 (O_133,N_9235,N_8880);
and UO_134 (O_134,N_8749,N_9492);
or UO_135 (O_135,N_9157,N_8411);
and UO_136 (O_136,N_9942,N_9841);
nand UO_137 (O_137,N_9390,N_9087);
and UO_138 (O_138,N_8499,N_8088);
or UO_139 (O_139,N_9737,N_9529);
or UO_140 (O_140,N_8099,N_8380);
nand UO_141 (O_141,N_8284,N_9434);
nand UO_142 (O_142,N_8100,N_8511);
nand UO_143 (O_143,N_8255,N_9385);
and UO_144 (O_144,N_9937,N_9488);
nand UO_145 (O_145,N_8569,N_9716);
nand UO_146 (O_146,N_9736,N_8767);
nand UO_147 (O_147,N_8635,N_9085);
and UO_148 (O_148,N_8062,N_8361);
and UO_149 (O_149,N_8409,N_9055);
and UO_150 (O_150,N_8494,N_9769);
or UO_151 (O_151,N_9593,N_9649);
and UO_152 (O_152,N_8897,N_9871);
and UO_153 (O_153,N_8753,N_9107);
or UO_154 (O_154,N_9978,N_9547);
and UO_155 (O_155,N_9951,N_8307);
and UO_156 (O_156,N_8093,N_8656);
or UO_157 (O_157,N_9676,N_9854);
nand UO_158 (O_158,N_9641,N_8306);
or UO_159 (O_159,N_9315,N_9637);
nor UO_160 (O_160,N_8764,N_8134);
nor UO_161 (O_161,N_8132,N_9184);
and UO_162 (O_162,N_8770,N_9796);
nor UO_163 (O_163,N_8490,N_9920);
and UO_164 (O_164,N_9111,N_9130);
and UO_165 (O_165,N_9962,N_8903);
nor UO_166 (O_166,N_9353,N_8766);
and UO_167 (O_167,N_9867,N_8773);
or UO_168 (O_168,N_9202,N_8290);
nor UO_169 (O_169,N_8478,N_8629);
nor UO_170 (O_170,N_8076,N_9945);
nor UO_171 (O_171,N_9707,N_9368);
and UO_172 (O_172,N_8782,N_9364);
nand UO_173 (O_173,N_8618,N_9523);
nor UO_174 (O_174,N_8529,N_8015);
nor UO_175 (O_175,N_9424,N_9572);
or UO_176 (O_176,N_9017,N_9098);
xnor UO_177 (O_177,N_8780,N_9761);
nand UO_178 (O_178,N_8149,N_9476);
nand UO_179 (O_179,N_8836,N_8456);
nor UO_180 (O_180,N_8945,N_9802);
or UO_181 (O_181,N_8952,N_9318);
nor UO_182 (O_182,N_8279,N_9522);
or UO_183 (O_183,N_8704,N_8402);
nand UO_184 (O_184,N_8164,N_9198);
and UO_185 (O_185,N_8869,N_9044);
nor UO_186 (O_186,N_8822,N_8563);
and UO_187 (O_187,N_8199,N_8252);
and UO_188 (O_188,N_9327,N_8445);
and UO_189 (O_189,N_9995,N_9490);
nand UO_190 (O_190,N_9455,N_8647);
and UO_191 (O_191,N_8571,N_8984);
and UO_192 (O_192,N_9272,N_9477);
nand UO_193 (O_193,N_8167,N_9741);
nor UO_194 (O_194,N_9237,N_8216);
or UO_195 (O_195,N_9135,N_8066);
nor UO_196 (O_196,N_9086,N_9592);
nand UO_197 (O_197,N_8177,N_9820);
or UO_198 (O_198,N_9437,N_9503);
nand UO_199 (O_199,N_8703,N_9817);
nor UO_200 (O_200,N_8575,N_8814);
or UO_201 (O_201,N_8026,N_8615);
and UO_202 (O_202,N_9112,N_9048);
and UO_203 (O_203,N_8363,N_9001);
nor UO_204 (O_204,N_8096,N_8628);
nand UO_205 (O_205,N_9798,N_8055);
nor UO_206 (O_206,N_8747,N_9545);
or UO_207 (O_207,N_9429,N_8609);
or UO_208 (O_208,N_8882,N_9681);
or UO_209 (O_209,N_9694,N_9756);
and UO_210 (O_210,N_9775,N_9744);
nor UO_211 (O_211,N_8323,N_9378);
and UO_212 (O_212,N_8751,N_9699);
nor UO_213 (O_213,N_9250,N_8310);
and UO_214 (O_214,N_9471,N_8215);
and UO_215 (O_215,N_8233,N_9930);
nor UO_216 (O_216,N_8013,N_8818);
and UO_217 (O_217,N_8560,N_8492);
nor UO_218 (O_218,N_9663,N_9768);
and UO_219 (O_219,N_9685,N_8932);
xnor UO_220 (O_220,N_9507,N_8092);
and UO_221 (O_221,N_8480,N_9451);
or UO_222 (O_222,N_9465,N_9173);
nor UO_223 (O_223,N_8241,N_8288);
and UO_224 (O_224,N_9719,N_8613);
nand UO_225 (O_225,N_9999,N_8311);
nand UO_226 (O_226,N_8713,N_9117);
or UO_227 (O_227,N_9456,N_8895);
nor UO_228 (O_228,N_8627,N_8007);
nor UO_229 (O_229,N_9016,N_9628);
or UO_230 (O_230,N_9276,N_9878);
or UO_231 (O_231,N_8665,N_8678);
nand UO_232 (O_232,N_8501,N_9041);
and UO_233 (O_233,N_9797,N_8046);
nand UO_234 (O_234,N_9380,N_8212);
nand UO_235 (O_235,N_9050,N_9116);
nand UO_236 (O_236,N_9944,N_9642);
nand UO_237 (O_237,N_9328,N_9918);
nand UO_238 (O_238,N_8379,N_8541);
or UO_239 (O_239,N_9223,N_8193);
or UO_240 (O_240,N_9126,N_9865);
and UO_241 (O_241,N_8074,N_8250);
or UO_242 (O_242,N_9639,N_9341);
nor UO_243 (O_243,N_8978,N_9505);
nand UO_244 (O_244,N_8851,N_8127);
and UO_245 (O_245,N_9825,N_8675);
or UO_246 (O_246,N_9583,N_9635);
nor UO_247 (O_247,N_8114,N_8467);
nand UO_248 (O_248,N_9702,N_8709);
and UO_249 (O_249,N_8852,N_8386);
nor UO_250 (O_250,N_9216,N_8442);
or UO_251 (O_251,N_8028,N_8506);
and UO_252 (O_252,N_8611,N_9433);
nor UO_253 (O_253,N_8435,N_8372);
nand UO_254 (O_254,N_9959,N_9270);
nor UO_255 (O_255,N_9806,N_9316);
and UO_256 (O_256,N_8104,N_8690);
xnor UO_257 (O_257,N_9416,N_8632);
or UO_258 (O_258,N_9241,N_8449);
and UO_259 (O_259,N_9977,N_8440);
or UO_260 (O_260,N_8430,N_8500);
and UO_261 (O_261,N_9778,N_8784);
nor UO_262 (O_262,N_8810,N_9002);
nand UO_263 (O_263,N_8427,N_9196);
or UO_264 (O_264,N_9129,N_8357);
nand UO_265 (O_265,N_9032,N_9723);
nor UO_266 (O_266,N_9484,N_9305);
nand UO_267 (O_267,N_8182,N_9323);
or UO_268 (O_268,N_9549,N_8738);
nor UO_269 (O_269,N_9677,N_8148);
nand UO_270 (O_270,N_9210,N_9275);
and UO_271 (O_271,N_8752,N_8210);
or UO_272 (O_272,N_8020,N_8228);
and UO_273 (O_273,N_9560,N_8211);
nor UO_274 (O_274,N_8493,N_9162);
nor UO_275 (O_275,N_9577,N_8197);
or UO_276 (O_276,N_9861,N_8073);
or UO_277 (O_277,N_9109,N_8825);
nor UO_278 (O_278,N_9435,N_9115);
or UO_279 (O_279,N_9366,N_8065);
and UO_280 (O_280,N_9675,N_8619);
nand UO_281 (O_281,N_9167,N_9239);
or UO_282 (O_282,N_9057,N_8620);
nor UO_283 (O_283,N_8908,N_9422);
or UO_284 (O_284,N_8489,N_8701);
or UO_285 (O_285,N_9466,N_8685);
nand UO_286 (O_286,N_8354,N_9155);
nor UO_287 (O_287,N_9531,N_9794);
nor UO_288 (O_288,N_8968,N_9934);
and UO_289 (O_289,N_8399,N_9501);
or UO_290 (O_290,N_9100,N_9652);
or UO_291 (O_291,N_9591,N_8824);
and UO_292 (O_292,N_9968,N_9843);
nand UO_293 (O_293,N_8696,N_8973);
nand UO_294 (O_294,N_9766,N_9513);
nand UO_295 (O_295,N_9701,N_9759);
nor UO_296 (O_296,N_8756,N_8374);
or UO_297 (O_297,N_9691,N_9308);
nor UO_298 (O_298,N_8775,N_8036);
nor UO_299 (O_299,N_9339,N_9748);
and UO_300 (O_300,N_8892,N_9149);
and UO_301 (O_301,N_9892,N_9019);
nand UO_302 (O_302,N_9452,N_9622);
or UO_303 (O_303,N_9933,N_8133);
or UO_304 (O_304,N_9108,N_8873);
nand UO_305 (O_305,N_8835,N_8401);
nor UO_306 (O_306,N_9633,N_8123);
or UO_307 (O_307,N_9900,N_9013);
nand UO_308 (O_308,N_8006,N_9138);
and UO_309 (O_309,N_8229,N_8920);
and UO_310 (O_310,N_9897,N_9351);
and UO_311 (O_311,N_8264,N_9355);
nand UO_312 (O_312,N_8237,N_8953);
or UO_313 (O_313,N_9986,N_8847);
nand UO_314 (O_314,N_9372,N_8885);
and UO_315 (O_315,N_8146,N_9253);
and UO_316 (O_316,N_8849,N_9521);
nor UO_317 (O_317,N_9066,N_8845);
and UO_318 (O_318,N_9514,N_9346);
or UO_319 (O_319,N_9436,N_8596);
or UO_320 (O_320,N_8638,N_8544);
or UO_321 (O_321,N_9005,N_8400);
and UO_322 (O_322,N_9499,N_8875);
nor UO_323 (O_323,N_9072,N_8154);
nor UO_324 (O_324,N_8963,N_8622);
nand UO_325 (O_325,N_8448,N_8524);
or UO_326 (O_326,N_8650,N_8029);
nand UO_327 (O_327,N_8669,N_8023);
or UO_328 (O_328,N_9600,N_9834);
and UO_329 (O_329,N_9627,N_9373);
or UO_330 (O_330,N_8170,N_9582);
and UO_331 (O_331,N_9527,N_8011);
nor UO_332 (O_332,N_9618,N_9919);
nand UO_333 (O_333,N_8068,N_8341);
xor UO_334 (O_334,N_8682,N_9767);
nand UO_335 (O_335,N_9947,N_9585);
or UO_336 (O_336,N_9803,N_9143);
xnor UO_337 (O_337,N_9371,N_9230);
or UO_338 (O_338,N_9597,N_9142);
nand UO_339 (O_339,N_9217,N_8218);
nand UO_340 (O_340,N_8388,N_9257);
and UO_341 (O_341,N_9653,N_8653);
and UO_342 (O_342,N_9334,N_8808);
or UO_343 (O_343,N_9879,N_8526);
and UO_344 (O_344,N_9992,N_8491);
and UO_345 (O_345,N_9197,N_8190);
nor UO_346 (O_346,N_9007,N_8534);
or UO_347 (O_347,N_8707,N_9238);
or UO_348 (O_348,N_8941,N_9395);
and UO_349 (O_349,N_8298,N_9518);
or UO_350 (O_350,N_9485,N_8955);
nand UO_351 (O_351,N_8488,N_9697);
or UO_352 (O_352,N_9692,N_8168);
and UO_353 (O_353,N_8147,N_9077);
xor UO_354 (O_354,N_8772,N_8479);
nor UO_355 (O_355,N_8418,N_9886);
nand UO_356 (O_356,N_9833,N_9495);
nand UO_357 (O_357,N_8275,N_8302);
and UO_358 (O_358,N_8459,N_9709);
nor UO_359 (O_359,N_8369,N_9000);
nand UO_360 (O_360,N_8040,N_8666);
nand UO_361 (O_361,N_9823,N_9407);
nor UO_362 (O_362,N_9096,N_9164);
xor UO_363 (O_363,N_8512,N_9446);
or UO_364 (O_364,N_8305,N_9090);
nor UO_365 (O_365,N_8802,N_8597);
nor UO_366 (O_366,N_8602,N_8515);
or UO_367 (O_367,N_8408,N_9454);
and UO_368 (O_368,N_8985,N_8367);
nand UO_369 (O_369,N_8797,N_9790);
and UO_370 (O_370,N_8970,N_9895);
or UO_371 (O_371,N_8518,N_9348);
or UO_372 (O_372,N_9475,N_9935);
nor UO_373 (O_373,N_9860,N_9388);
and UO_374 (O_374,N_9483,N_8166);
and UO_375 (O_375,N_9189,N_8454);
nor UO_376 (O_376,N_8827,N_8943);
nor UO_377 (O_377,N_9065,N_8219);
and UO_378 (O_378,N_8412,N_9417);
and UO_379 (O_379,N_8991,N_9236);
and UO_380 (O_380,N_9857,N_8712);
and UO_381 (O_381,N_8201,N_8856);
and UO_382 (O_382,N_9787,N_9227);
and UO_383 (O_383,N_8942,N_9273);
nor UO_384 (O_384,N_8583,N_9800);
nor UO_385 (O_385,N_9357,N_9564);
or UO_386 (O_386,N_9249,N_9615);
nor UO_387 (O_387,N_8781,N_8987);
nand UO_388 (O_388,N_9088,N_8005);
or UO_389 (O_389,N_8353,N_8960);
or UO_390 (O_390,N_8922,N_9365);
and UO_391 (O_391,N_9391,N_9091);
and UO_392 (O_392,N_8975,N_8933);
nor UO_393 (O_393,N_8513,N_9783);
and UO_394 (O_394,N_8994,N_8540);
and UO_395 (O_395,N_9337,N_9464);
or UO_396 (O_396,N_8919,N_9333);
nand UO_397 (O_397,N_8063,N_8139);
nand UO_398 (O_398,N_8181,N_9506);
and UO_399 (O_399,N_9303,N_8872);
and UO_400 (O_400,N_9617,N_8537);
nor UO_401 (O_401,N_9536,N_8192);
or UO_402 (O_402,N_9147,N_8457);
and UO_403 (O_403,N_9040,N_9379);
nand UO_404 (O_404,N_9261,N_8672);
or UO_405 (O_405,N_9054,N_9609);
and UO_406 (O_406,N_9780,N_9114);
nor UO_407 (O_407,N_9875,N_8807);
and UO_408 (O_408,N_8102,N_8763);
nand UO_409 (O_409,N_9081,N_9634);
nand UO_410 (O_410,N_8131,N_8746);
and UO_411 (O_411,N_8276,N_8277);
nand UO_412 (O_412,N_8906,N_8539);
and UO_413 (O_413,N_9245,N_9309);
nor UO_414 (O_414,N_9426,N_8129);
and UO_415 (O_415,N_8204,N_9370);
nor UO_416 (O_416,N_8159,N_8900);
nand UO_417 (O_417,N_8652,N_9504);
or UO_418 (O_418,N_9174,N_9412);
nor UO_419 (O_419,N_9035,N_8120);
or UO_420 (O_420,N_8471,N_9047);
nor UO_421 (O_421,N_9750,N_9025);
nor UO_422 (O_422,N_8291,N_8081);
nor UO_423 (O_423,N_8683,N_8464);
and UO_424 (O_424,N_8308,N_9106);
nor UO_425 (O_425,N_8474,N_9630);
nand UO_426 (O_426,N_8498,N_8087);
nor UO_427 (O_427,N_9666,N_9568);
and UO_428 (O_428,N_8971,N_8833);
or UO_429 (O_429,N_9472,N_9127);
nand UO_430 (O_430,N_9928,N_9432);
or UO_431 (O_431,N_9955,N_9696);
and UO_432 (O_432,N_9254,N_8817);
or UO_433 (O_433,N_9284,N_8043);
and UO_434 (O_434,N_8124,N_8083);
nor UO_435 (O_435,N_9808,N_9311);
nor UO_436 (O_436,N_9439,N_9268);
and UO_437 (O_437,N_9904,N_9924);
and UO_438 (O_438,N_8315,N_8929);
and UO_439 (O_439,N_8424,N_9858);
nor UO_440 (O_440,N_9754,N_9690);
nor UO_441 (O_441,N_8947,N_8728);
nand UO_442 (O_442,N_9872,N_9247);
and UO_443 (O_443,N_8260,N_8118);
nand UO_444 (O_444,N_8719,N_8614);
and UO_445 (O_445,N_8834,N_9979);
and UO_446 (O_446,N_8779,N_9835);
nor UO_447 (O_447,N_9541,N_8097);
and UO_448 (O_448,N_8538,N_9882);
or UO_449 (O_449,N_9099,N_8333);
or UO_450 (O_450,N_9966,N_9064);
nor UO_451 (O_451,N_8034,N_9740);
or UO_452 (O_452,N_8286,N_8508);
or UO_453 (O_453,N_9201,N_8964);
and UO_454 (O_454,N_8737,N_9083);
or UO_455 (O_455,N_8937,N_9645);
nand UO_456 (O_456,N_9082,N_9816);
or UO_457 (O_457,N_9039,N_8562);
and UO_458 (O_458,N_9733,N_9981);
and UO_459 (O_459,N_8178,N_8577);
nand UO_460 (O_460,N_8886,N_8319);
or UO_461 (O_461,N_9729,N_9060);
or UO_462 (O_462,N_8925,N_8579);
nor UO_463 (O_463,N_9728,N_9289);
nor UO_464 (O_464,N_9557,N_9789);
nor UO_465 (O_465,N_9497,N_8995);
nand UO_466 (O_466,N_9508,N_9994);
or UO_467 (O_467,N_9730,N_8253);
or UO_468 (O_468,N_9608,N_8505);
and UO_469 (O_469,N_9809,N_9076);
nand UO_470 (O_470,N_9848,N_8581);
nor UO_471 (O_471,N_8265,N_9498);
nor UO_472 (O_472,N_9837,N_8225);
or UO_473 (O_473,N_8894,N_8684);
or UO_474 (O_474,N_9845,N_9688);
and UO_475 (O_475,N_9214,N_9449);
or UO_476 (O_476,N_8686,N_9213);
nand UO_477 (O_477,N_8365,N_8282);
nand UO_478 (O_478,N_8548,N_8887);
nand UO_479 (O_479,N_9310,N_8346);
nor UO_480 (O_480,N_8582,N_8608);
nor UO_481 (O_481,N_8816,N_9898);
and UO_482 (O_482,N_8930,N_9259);
and UO_483 (O_483,N_9069,N_9824);
nor UO_484 (O_484,N_8103,N_8202);
and UO_485 (O_485,N_8338,N_8263);
or UO_486 (O_486,N_9795,N_9003);
nor UO_487 (O_487,N_8050,N_8405);
nand UO_488 (O_488,N_8432,N_8715);
nor UO_489 (O_489,N_9191,N_9430);
nand UO_490 (O_490,N_8460,N_9063);
or UO_491 (O_491,N_9374,N_8722);
nor UO_492 (O_492,N_9491,N_9219);
nor UO_493 (O_493,N_9419,N_8496);
and UO_494 (O_494,N_8251,N_9695);
nor UO_495 (O_495,N_8893,N_8385);
and UO_496 (O_496,N_8868,N_9256);
and UO_497 (O_497,N_9793,N_8904);
nor UO_498 (O_498,N_8710,N_8735);
nor UO_499 (O_499,N_9190,N_9161);
nand UO_500 (O_500,N_9829,N_9045);
or UO_501 (O_501,N_9661,N_9776);
nor UO_502 (O_502,N_8604,N_8617);
or UO_503 (O_503,N_9105,N_8785);
or UO_504 (O_504,N_8391,N_9619);
nand UO_505 (O_505,N_8967,N_8370);
or UO_506 (O_506,N_9874,N_8232);
nand UO_507 (O_507,N_9458,N_9397);
and UO_508 (O_508,N_9093,N_9326);
nor UO_509 (O_509,N_8483,N_9799);
nor UO_510 (O_510,N_8281,N_8954);
and UO_511 (O_511,N_9877,N_9850);
and UO_512 (O_512,N_9648,N_8530);
nand UO_513 (O_513,N_8708,N_8101);
nor UO_514 (O_514,N_9839,N_9474);
nand UO_515 (O_515,N_8137,N_9345);
nor UO_516 (O_516,N_9914,N_9322);
nor UO_517 (O_517,N_8848,N_8245);
nor UO_518 (O_518,N_9866,N_8316);
or UO_519 (O_519,N_9071,N_8832);
nand UO_520 (O_520,N_9038,N_8413);
or UO_521 (O_521,N_8157,N_8152);
and UO_522 (O_522,N_9757,N_8729);
nor UO_523 (O_523,N_9542,N_9335);
nand UO_524 (O_524,N_8451,N_8578);
or UO_525 (O_525,N_9049,N_9177);
nor UO_526 (O_526,N_8600,N_9735);
nand UO_527 (O_527,N_8236,N_8128);
nand UO_528 (O_528,N_8038,N_9941);
nor UO_529 (O_529,N_8355,N_8126);
or UO_530 (O_530,N_9851,N_9359);
and UO_531 (O_531,N_8731,N_8165);
and UO_532 (O_532,N_8268,N_9873);
nor UO_533 (O_533,N_9957,N_9122);
xnor UO_534 (O_534,N_9515,N_8798);
nor UO_535 (O_535,N_9563,N_9943);
or UO_536 (O_536,N_8674,N_8156);
and UO_537 (O_537,N_8052,N_9317);
nand UO_538 (O_538,N_9280,N_8533);
nor UO_539 (O_539,N_9188,N_8783);
nor UO_540 (O_540,N_8561,N_8626);
and UO_541 (O_541,N_9654,N_9646);
xnor UO_542 (O_542,N_9657,N_9559);
and UO_543 (O_543,N_8976,N_9274);
and UO_544 (O_544,N_9814,N_9307);
nor UO_545 (O_545,N_8377,N_9312);
nor UO_546 (O_546,N_8663,N_8794);
nor UO_547 (O_547,N_9008,N_8909);
or UO_548 (O_548,N_9804,N_8455);
nor UO_549 (O_549,N_8951,N_8339);
and UO_550 (O_550,N_8012,N_9606);
or UO_551 (O_551,N_9014,N_9059);
nor UO_552 (O_552,N_9457,N_8257);
or UO_553 (O_553,N_9078,N_9128);
or UO_554 (O_554,N_9352,N_8191);
or UO_555 (O_555,N_8962,N_9186);
nand UO_556 (O_556,N_9629,N_8714);
and UO_557 (O_557,N_9175,N_9950);
or UO_558 (O_558,N_9313,N_8918);
and UO_559 (O_559,N_9277,N_8003);
or UO_560 (O_560,N_9121,N_8671);
nor UO_561 (O_561,N_8514,N_8249);
nand UO_562 (O_562,N_8843,N_8485);
nand UO_563 (O_563,N_9524,N_9031);
or UO_564 (O_564,N_8717,N_8304);
nand UO_565 (O_565,N_9880,N_9746);
nor UO_566 (O_566,N_9354,N_9468);
nand UO_567 (O_567,N_8507,N_9133);
and UO_568 (O_568,N_9427,N_8226);
or UO_569 (O_569,N_8422,N_8145);
and UO_570 (O_570,N_9493,N_9580);
or UO_571 (O_571,N_8079,N_9203);
and UO_572 (O_572,N_8826,N_9413);
nor UO_573 (O_573,N_9538,N_9516);
nand UO_574 (O_574,N_8702,N_8472);
or UO_575 (O_575,N_8841,N_9519);
or UO_576 (O_576,N_8718,N_8586);
and UO_577 (O_577,N_9569,N_8550);
or UO_578 (O_578,N_8844,N_8523);
nor UO_579 (O_579,N_8048,N_9123);
or UO_580 (O_580,N_8105,N_8248);
and UO_581 (O_581,N_8325,N_8337);
nand UO_582 (O_582,N_8244,N_9229);
nor UO_583 (O_583,N_9461,N_9325);
and UO_584 (O_584,N_8175,N_9231);
xnor UO_585 (O_585,N_9546,N_9722);
nand UO_586 (O_586,N_8246,N_8693);
and UO_587 (O_587,N_9183,N_8322);
and UO_588 (O_588,N_8878,N_9974);
nand UO_589 (O_589,N_9601,N_8838);
nor UO_590 (O_590,N_8521,N_8466);
nand UO_591 (O_591,N_8116,N_9755);
and UO_592 (O_592,N_8974,N_9079);
nor UO_593 (O_593,N_8796,N_8439);
xor UO_594 (O_594,N_9443,N_8564);
and UO_595 (O_595,N_8004,N_8720);
nor UO_596 (O_596,N_9896,N_9469);
nor UO_597 (O_597,N_8986,N_9840);
and UO_598 (O_598,N_8261,N_9813);
or UO_599 (O_599,N_8031,N_9179);
or UO_600 (O_600,N_9246,N_8419);
nand UO_601 (O_601,N_8240,N_8790);
nor UO_602 (O_602,N_9996,N_9899);
nor UO_603 (O_603,N_9023,N_9975);
nand UO_604 (O_604,N_9383,N_9660);
nor UO_605 (O_605,N_9983,N_8345);
nor UO_606 (O_606,N_9146,N_8274);
and UO_607 (O_607,N_9596,N_8864);
and UO_608 (O_608,N_8019,N_9494);
nand UO_609 (O_609,N_8222,N_9889);
nand UO_610 (O_610,N_8646,N_9042);
and UO_611 (O_611,N_8238,N_9903);
nand UO_612 (O_612,N_9949,N_9961);
nand UO_613 (O_613,N_8223,N_8269);
nor UO_614 (O_614,N_9024,N_8336);
nand UO_615 (O_615,N_8551,N_8883);
nand UO_616 (O_616,N_8795,N_8559);
or UO_617 (O_617,N_9344,N_9517);
nand UO_618 (O_618,N_9807,N_8877);
nand UO_619 (O_619,N_8636,N_8687);
nand UO_620 (O_620,N_9632,N_9528);
and UO_621 (O_621,N_8371,N_9113);
and UO_622 (O_622,N_8481,N_8450);
and UO_623 (O_623,N_8946,N_9486);
and UO_624 (O_624,N_9972,N_8329);
nor UO_625 (O_625,N_8935,N_9448);
nor UO_626 (O_626,N_8915,N_8090);
nor UO_627 (O_627,N_9269,N_9526);
nor UO_628 (O_628,N_9721,N_9467);
and UO_629 (O_629,N_9749,N_8944);
and UO_630 (O_630,N_8091,N_9539);
or UO_631 (O_631,N_8901,N_9760);
and UO_632 (O_632,N_8592,N_8740);
nor UO_633 (O_633,N_8607,N_9656);
or UO_634 (O_634,N_8961,N_8196);
or UO_635 (O_635,N_9363,N_8657);
nand UO_636 (O_636,N_8884,N_9751);
nand UO_637 (O_637,N_8169,N_8383);
nor UO_638 (O_638,N_8923,N_9396);
and UO_639 (O_639,N_9705,N_8205);
and UO_640 (O_640,N_9252,N_8358);
nor UO_641 (O_641,N_9673,N_8375);
or UO_642 (O_642,N_8256,N_9400);
nand UO_643 (O_643,N_9037,N_9753);
or UO_644 (O_644,N_8625,N_8138);
or UO_645 (O_645,N_9296,N_8661);
or UO_646 (O_646,N_9990,N_9052);
nor UO_647 (O_647,N_9602,N_8516);
nor UO_648 (O_648,N_8736,N_8610);
nor UO_649 (O_649,N_9420,N_8423);
nor UO_650 (O_650,N_8981,N_9674);
nand UO_651 (O_651,N_8373,N_9288);
nand UO_652 (O_652,N_8360,N_8080);
nand UO_653 (O_653,N_8172,N_8743);
and UO_654 (O_654,N_8343,N_9613);
and UO_655 (O_655,N_9511,N_9010);
or UO_656 (O_656,N_8378,N_8660);
nand UO_657 (O_657,N_9020,N_8972);
nor UO_658 (O_658,N_9938,N_9535);
or UO_659 (O_659,N_9952,N_9708);
or UO_660 (O_660,N_9243,N_8352);
or UO_661 (O_661,N_8224,N_8142);
or UO_662 (O_662,N_9915,N_8462);
nor UO_663 (O_663,N_9832,N_9070);
nor UO_664 (O_664,N_9616,N_8520);
and UO_665 (O_665,N_8185,N_9881);
and UO_666 (O_666,N_8905,N_8437);
xnor UO_667 (O_667,N_8153,N_9338);
and UO_668 (O_668,N_8059,N_8670);
nor UO_669 (O_669,N_8024,N_8698);
nand UO_670 (O_670,N_8344,N_8673);
and UO_671 (O_671,N_8823,N_8549);
nor UO_672 (O_672,N_8828,N_8999);
or UO_673 (O_673,N_8176,N_9208);
nand UO_674 (O_674,N_8624,N_9282);
or UO_675 (O_675,N_8727,N_8280);
and UO_676 (O_676,N_8692,N_8039);
or UO_677 (O_677,N_8996,N_9158);
or UO_678 (O_678,N_9773,N_9225);
nand UO_679 (O_679,N_8699,N_9682);
nor UO_680 (O_680,N_8570,N_9575);
nand UO_681 (O_681,N_8045,N_8655);
or UO_682 (O_682,N_9819,N_9340);
nand UO_683 (O_683,N_9711,N_9669);
nor UO_684 (O_684,N_9853,N_9450);
xnor UO_685 (O_685,N_8811,N_9815);
nor UO_686 (O_686,N_8957,N_9195);
or UO_687 (O_687,N_9932,N_8161);
xor UO_688 (O_688,N_9703,N_9131);
and UO_689 (O_689,N_9956,N_9462);
xor UO_690 (O_690,N_8262,N_9421);
nor UO_691 (O_691,N_8723,N_8347);
and UO_692 (O_692,N_9553,N_8547);
nor UO_693 (O_693,N_8950,N_8434);
nor UO_694 (O_694,N_9991,N_9520);
nor UO_695 (O_695,N_9777,N_8174);
nand UO_696 (O_696,N_8135,N_8207);
and UO_697 (O_697,N_8862,N_8444);
nor UO_698 (O_698,N_8136,N_8916);
nor UO_699 (O_699,N_9856,N_8041);
nor UO_700 (O_700,N_8989,N_8979);
nand UO_701 (O_701,N_9489,N_8889);
nand UO_702 (O_702,N_8303,N_8846);
nand UO_703 (O_703,N_8688,N_8928);
or UO_704 (O_704,N_8700,N_9306);
nand UO_705 (O_705,N_8077,N_9367);
nand UO_706 (O_706,N_8594,N_8495);
nor UO_707 (O_707,N_8876,N_8107);
and UO_708 (O_708,N_8469,N_9561);
nand UO_709 (O_709,N_8724,N_8595);
nand UO_710 (O_710,N_8641,N_9030);
nand UO_711 (O_711,N_9212,N_8141);
and UO_712 (O_712,N_8787,N_8587);
nor UO_713 (O_713,N_8503,N_8071);
nor UO_714 (O_714,N_8340,N_9205);
or UO_715 (O_715,N_8879,N_9399);
and UO_716 (O_716,N_8959,N_9970);
nand UO_717 (O_717,N_9810,N_9948);
or UO_718 (O_718,N_8863,N_8926);
nand UO_719 (O_719,N_8032,N_9304);
or UO_720 (O_720,N_9384,N_9251);
nand UO_721 (O_721,N_9791,N_8725);
and UO_722 (O_722,N_9801,N_9891);
nor UO_723 (O_723,N_9811,N_8384);
nor UO_724 (O_724,N_8206,N_8745);
and UO_725 (O_725,N_9176,N_8299);
nor UO_726 (O_726,N_8106,N_8881);
and UO_727 (O_727,N_9118,N_8082);
nor UO_728 (O_728,N_9785,N_9859);
and UO_729 (O_729,N_8482,N_9921);
and UO_730 (O_730,N_9361,N_9738);
nand UO_731 (O_731,N_8788,N_9964);
and UO_732 (O_732,N_8398,N_9726);
and UO_733 (O_733,N_8982,N_8630);
nor UO_734 (O_734,N_9607,N_8381);
or UO_735 (O_735,N_8531,N_8254);
or UO_736 (O_736,N_8758,N_8155);
nand UO_737 (O_737,N_8590,N_8588);
or UO_738 (O_738,N_9724,N_8000);
nor UO_739 (O_739,N_8294,N_9242);
nor UO_740 (O_740,N_8644,N_8390);
nor UO_741 (O_741,N_8754,N_9713);
nor UO_742 (O_742,N_9481,N_8896);
or UO_743 (O_743,N_8151,N_8376);
xnor UO_744 (O_744,N_9171,N_9764);
and UO_745 (O_745,N_9862,N_8639);
nor UO_746 (O_746,N_8072,N_9960);
or UO_747 (O_747,N_8522,N_9614);
or UO_748 (O_748,N_8558,N_8334);
nor UO_749 (O_749,N_9140,N_9043);
or UO_750 (O_750,N_9905,N_8272);
nand UO_751 (O_751,N_8187,N_9291);
nand UO_752 (O_752,N_9574,N_9387);
and UO_753 (O_753,N_8861,N_9912);
nand UO_754 (O_754,N_8760,N_8504);
xnor UO_755 (O_755,N_8160,N_9788);
and UO_756 (O_756,N_8651,N_8426);
nand UO_757 (O_757,N_9910,N_8867);
or UO_758 (O_758,N_9028,N_9772);
or UO_759 (O_759,N_9350,N_9248);
nand UO_760 (O_760,N_8676,N_9004);
nand UO_761 (O_761,N_9264,N_9295);
nor UO_762 (O_762,N_8121,N_8517);
nor UO_763 (O_763,N_9954,N_8112);
xnor UO_764 (O_764,N_8364,N_9731);
nand UO_765 (O_765,N_8397,N_8458);
nand UO_766 (O_766,N_8075,N_9530);
nor UO_767 (O_767,N_9152,N_9973);
nor UO_768 (O_768,N_9849,N_8198);
nand UO_769 (O_769,N_8125,N_9068);
nand UO_770 (O_770,N_8230,N_9922);
nor UO_771 (O_771,N_9985,N_9441);
and UO_772 (O_772,N_9226,N_9479);
and UO_773 (O_773,N_8716,N_8765);
or UO_774 (O_774,N_9438,N_9178);
nor UO_775 (O_775,N_8033,N_8525);
nor UO_776 (O_776,N_9144,N_8840);
nand UO_777 (O_777,N_8312,N_8993);
and UO_778 (O_778,N_9887,N_8585);
nand UO_779 (O_779,N_9145,N_8417);
nand UO_780 (O_780,N_9818,N_8425);
nand UO_781 (O_781,N_8980,N_9119);
nor UO_782 (O_782,N_8677,N_8858);
and UO_783 (O_783,N_9009,N_9550);
and UO_784 (O_784,N_8247,N_8572);
or UO_785 (O_785,N_9689,N_8351);
or UO_786 (O_786,N_8278,N_8270);
and UO_787 (O_787,N_9160,N_8850);
and UO_788 (O_788,N_8711,N_9187);
nor UO_789 (O_789,N_8326,N_8606);
or UO_790 (O_790,N_8940,N_9095);
or UO_791 (O_791,N_8002,N_8739);
and UO_792 (O_792,N_8318,N_9006);
nor UO_793 (O_793,N_8573,N_8774);
nor UO_794 (O_794,N_9139,N_9929);
or UO_795 (O_795,N_8645,N_9453);
nand UO_796 (O_796,N_9926,N_8527);
and UO_797 (O_797,N_8890,N_9822);
or UO_798 (O_798,N_9166,N_9320);
or UO_799 (O_799,N_9679,N_9343);
or UO_800 (O_800,N_9626,N_9869);
nand UO_801 (O_801,N_9473,N_9595);
nor UO_802 (O_802,N_8017,N_8117);
and UO_803 (O_803,N_8776,N_8556);
nand UO_804 (O_804,N_9774,N_9884);
and UO_805 (O_805,N_8273,N_9423);
or UO_806 (O_806,N_9431,N_8510);
and UO_807 (O_807,N_9067,N_9163);
nand UO_808 (O_808,N_9401,N_8983);
nor UO_809 (O_809,N_9812,N_9963);
or UO_810 (O_810,N_8209,N_8553);
and UO_811 (O_811,N_8591,N_8621);
and UO_812 (O_812,N_9533,N_9409);
and UO_813 (O_813,N_9784,N_8057);
nor UO_814 (O_814,N_8259,N_8662);
nand UO_815 (O_815,N_9425,N_8443);
or UO_816 (O_816,N_9715,N_8680);
nor UO_817 (O_817,N_8300,N_8266);
and UO_818 (O_818,N_8060,N_9209);
and UO_819 (O_819,N_8113,N_8911);
nor UO_820 (O_820,N_8733,N_8580);
or UO_821 (O_821,N_9836,N_8037);
nor UO_822 (O_822,N_8403,N_9369);
nor UO_823 (O_823,N_8144,N_9392);
and UO_824 (O_824,N_9555,N_9758);
nor UO_825 (O_825,N_9763,N_9909);
nand UO_826 (O_826,N_8778,N_9638);
nand UO_827 (O_827,N_9141,N_8870);
and UO_828 (O_828,N_9562,N_8956);
or UO_829 (O_829,N_8420,N_8476);
nand UO_830 (O_830,N_8047,N_8194);
and UO_831 (O_831,N_8025,N_9414);
or UO_832 (O_832,N_9347,N_8350);
nor UO_833 (O_833,N_8163,N_8871);
nor UO_834 (O_834,N_9125,N_8283);
nor UO_835 (O_835,N_9286,N_9053);
and UO_836 (O_836,N_8085,N_8465);
or UO_837 (O_837,N_8221,N_9686);
and UO_838 (O_838,N_8433,N_8949);
and UO_839 (O_839,N_9029,N_9745);
nor UO_840 (O_840,N_8208,N_9018);
and UO_841 (O_841,N_9684,N_9319);
or UO_842 (O_842,N_9302,N_9097);
xor UO_843 (O_843,N_9336,N_8557);
nor UO_844 (O_844,N_8234,N_8477);
or UO_845 (O_845,N_8327,N_8111);
or UO_846 (O_846,N_9643,N_9863);
nor UO_847 (O_847,N_9782,N_8394);
nand UO_848 (O_848,N_9266,N_8768);
and UO_849 (O_849,N_9221,N_8389);
and UO_850 (O_850,N_8035,N_9194);
or UO_851 (O_851,N_8958,N_9447);
and UO_852 (O_852,N_9011,N_9717);
and UO_853 (O_853,N_9876,N_8721);
nand UO_854 (O_854,N_8891,N_8965);
and UO_855 (O_855,N_9279,N_9206);
or UO_856 (O_856,N_8180,N_9931);
and UO_857 (O_857,N_9664,N_9805);
nand UO_858 (O_858,N_8658,N_9406);
xor UO_859 (O_859,N_8599,N_9781);
or UO_860 (O_860,N_9940,N_8301);
nand UO_861 (O_861,N_9998,N_9283);
or UO_862 (O_862,N_8734,N_8910);
xor UO_863 (O_863,N_8664,N_8820);
nor UO_864 (O_864,N_9578,N_8171);
or UO_865 (O_865,N_9234,N_8089);
nand UO_866 (O_866,N_9556,N_8855);
or UO_867 (O_867,N_9442,N_8084);
or UO_868 (O_868,N_9668,N_8183);
nand UO_869 (O_869,N_8356,N_9376);
and UO_870 (O_870,N_9936,N_8271);
or UO_871 (O_871,N_8328,N_8441);
nand UO_872 (O_872,N_8162,N_9480);
nand UO_873 (O_873,N_9573,N_9075);
nor UO_874 (O_874,N_8801,N_8330);
nand UO_875 (O_875,N_9590,N_9747);
nand UO_876 (O_876,N_8697,N_8289);
or UO_877 (O_877,N_8761,N_8200);
nor UO_878 (O_878,N_9074,N_8335);
or UO_879 (O_879,N_9136,N_8640);
nor UO_880 (O_880,N_9428,N_9408);
nor UO_881 (O_881,N_9073,N_9386);
or UO_882 (O_882,N_9389,N_8899);
or UO_883 (O_883,N_8189,N_8453);
nor UO_884 (O_884,N_9137,N_8924);
nor UO_885 (O_885,N_8649,N_9714);
and UO_886 (O_886,N_8576,N_8108);
nand UO_887 (O_887,N_8348,N_8296);
or UO_888 (O_888,N_8387,N_9742);
or UO_889 (O_889,N_8830,N_9290);
or UO_890 (O_890,N_8759,N_9478);
or UO_891 (O_891,N_9415,N_8806);
or UO_892 (O_892,N_8487,N_9907);
nor UO_893 (O_893,N_8914,N_8902);
or UO_894 (O_894,N_9989,N_9534);
nor UO_895 (O_895,N_9548,N_9706);
or UO_896 (O_896,N_9445,N_9330);
nand UO_897 (O_897,N_8001,N_8362);
and UO_898 (O_898,N_8528,N_8461);
nand UO_899 (O_899,N_9558,N_8421);
nor UO_900 (O_900,N_9182,N_9698);
and UO_901 (O_901,N_8324,N_8195);
or UO_902 (O_902,N_9460,N_9394);
and UO_903 (O_903,N_9846,N_9552);
nand UO_904 (O_904,N_8546,N_8938);
nor UO_905 (O_905,N_9625,N_8907);
nand UO_906 (O_906,N_8748,N_8242);
nor UO_907 (O_907,N_9255,N_9027);
nand UO_908 (O_908,N_8912,N_9868);
and UO_909 (O_909,N_9258,N_9621);
or UO_910 (O_910,N_8429,N_9224);
and UO_911 (O_911,N_8803,N_8058);
nand UO_912 (O_912,N_8809,N_8552);
nor UO_913 (O_913,N_9172,N_8431);
nor UO_914 (O_914,N_9381,N_9321);
nand UO_915 (O_915,N_8874,N_8027);
and UO_916 (O_916,N_9015,N_8267);
and UO_917 (O_917,N_9971,N_8543);
nor UO_918 (O_918,N_8049,N_9154);
and UO_919 (O_919,N_8519,N_9482);
and UO_920 (O_920,N_8939,N_8762);
nand UO_921 (O_921,N_9026,N_8612);
nand UO_922 (O_922,N_8689,N_8966);
nor UO_923 (O_923,N_8584,N_9263);
nor UO_924 (O_924,N_9297,N_8470);
and UO_925 (O_925,N_9687,N_8292);
and UO_926 (O_926,N_8416,N_9587);
nand UO_927 (O_927,N_9150,N_9732);
and UO_928 (O_928,N_9605,N_8706);
and UO_929 (O_929,N_9658,N_9588);
nand UO_930 (O_930,N_9939,N_9965);
and UO_931 (O_931,N_9356,N_9393);
nor UO_932 (O_932,N_8054,N_8150);
xnor UO_933 (O_933,N_9021,N_9667);
nand UO_934 (O_934,N_8565,N_9651);
and UO_935 (O_935,N_9911,N_9739);
or UO_936 (O_936,N_9917,N_9765);
or UO_937 (O_937,N_9980,N_8681);
or UO_938 (O_938,N_9232,N_8502);
xnor UO_939 (O_939,N_9299,N_8694);
nand UO_940 (O_940,N_9169,N_8061);
nand UO_941 (O_941,N_8293,N_9089);
or UO_942 (O_942,N_9958,N_9908);
or UO_943 (O_943,N_8396,N_9576);
or UO_944 (O_944,N_9693,N_9762);
or UO_945 (O_945,N_8410,N_8098);
and UO_946 (O_946,N_9670,N_9581);
nand UO_947 (O_947,N_8992,N_8122);
nand UO_948 (O_948,N_8115,N_9571);
nor UO_949 (O_949,N_9240,N_8927);
or UO_950 (O_950,N_8771,N_9830);
and UO_951 (O_951,N_8705,N_8070);
nor UO_952 (O_952,N_9181,N_8757);
and UO_953 (O_953,N_9349,N_8130);
nand UO_954 (O_954,N_9233,N_8821);
or UO_955 (O_955,N_8742,N_8532);
nand UO_956 (O_956,N_8859,N_9051);
and UO_957 (O_957,N_9267,N_8726);
nand UO_958 (O_958,N_8317,N_9104);
and UO_959 (O_959,N_8866,N_8214);
and UO_960 (O_960,N_9720,N_8589);
and UO_961 (O_961,N_8243,N_8616);
xnor UO_962 (O_962,N_9022,N_8436);
and UO_963 (O_963,N_8695,N_9405);
nor UO_964 (O_964,N_9599,N_8854);
nor UO_965 (O_965,N_8741,N_8069);
or UO_966 (O_966,N_9984,N_8831);
or UO_967 (O_967,N_8936,N_8213);
or UO_968 (O_968,N_8860,N_9655);
or UO_969 (O_969,N_8898,N_9278);
nor UO_970 (O_970,N_8404,N_8217);
nor UO_971 (O_971,N_9156,N_8428);
or UO_972 (O_972,N_9262,N_8220);
or UO_973 (O_973,N_8014,N_9718);
or UO_974 (O_974,N_8186,N_8567);
and UO_975 (O_975,N_8475,N_8010);
nor UO_976 (O_976,N_9644,N_8777);
nand UO_977 (O_977,N_8158,N_8078);
and UO_978 (O_978,N_8642,N_8188);
nor UO_979 (O_979,N_9894,N_8755);
nand UO_980 (O_980,N_8805,N_8988);
nor UO_981 (O_981,N_8016,N_9193);
or UO_982 (O_982,N_9901,N_9603);
and UO_983 (O_983,N_9543,N_8497);
nor UO_984 (O_984,N_9185,N_9329);
and UO_985 (O_985,N_8484,N_9101);
or UO_986 (O_986,N_8140,N_8545);
nand UO_987 (O_987,N_8342,N_8997);
and UO_988 (O_988,N_8819,N_8359);
or UO_989 (O_989,N_9586,N_9683);
and UO_990 (O_990,N_9700,N_9265);
nor UO_991 (O_991,N_8179,N_8053);
nor UO_992 (O_992,N_8623,N_9211);
nor UO_993 (O_993,N_8799,N_9287);
nand UO_994 (O_994,N_9061,N_9838);
nand UO_995 (O_995,N_9402,N_9496);
or UO_996 (O_996,N_9770,N_8067);
nand UO_997 (O_997,N_9893,N_9589);
or UO_998 (O_998,N_8109,N_8447);
nand UO_999 (O_999,N_8554,N_9570);
and UO_1000 (O_1000,N_8342,N_9548);
nand UO_1001 (O_1001,N_9798,N_9611);
or UO_1002 (O_1002,N_9630,N_9363);
or UO_1003 (O_1003,N_9468,N_9396);
and UO_1004 (O_1004,N_9517,N_8122);
nand UO_1005 (O_1005,N_8694,N_9987);
nand UO_1006 (O_1006,N_8216,N_9007);
nor UO_1007 (O_1007,N_9103,N_8748);
and UO_1008 (O_1008,N_9351,N_8704);
or UO_1009 (O_1009,N_8621,N_8631);
or UO_1010 (O_1010,N_9966,N_8996);
nor UO_1011 (O_1011,N_8532,N_8082);
nor UO_1012 (O_1012,N_9781,N_8676);
or UO_1013 (O_1013,N_8481,N_9476);
nand UO_1014 (O_1014,N_8579,N_9673);
nor UO_1015 (O_1015,N_9194,N_9583);
nand UO_1016 (O_1016,N_9627,N_8657);
nand UO_1017 (O_1017,N_9076,N_8378);
and UO_1018 (O_1018,N_9301,N_8052);
xnor UO_1019 (O_1019,N_9591,N_8934);
nor UO_1020 (O_1020,N_8629,N_9461);
nor UO_1021 (O_1021,N_8188,N_9392);
nand UO_1022 (O_1022,N_8725,N_8930);
or UO_1023 (O_1023,N_8177,N_8069);
nand UO_1024 (O_1024,N_9235,N_8056);
nand UO_1025 (O_1025,N_9716,N_8053);
nor UO_1026 (O_1026,N_9770,N_8882);
nor UO_1027 (O_1027,N_8019,N_9901);
and UO_1028 (O_1028,N_8424,N_8546);
nand UO_1029 (O_1029,N_8403,N_9093);
or UO_1030 (O_1030,N_8132,N_8153);
nor UO_1031 (O_1031,N_8734,N_8353);
or UO_1032 (O_1032,N_9309,N_8710);
nand UO_1033 (O_1033,N_8752,N_8039);
or UO_1034 (O_1034,N_8189,N_8788);
and UO_1035 (O_1035,N_9983,N_9930);
nor UO_1036 (O_1036,N_9106,N_9683);
or UO_1037 (O_1037,N_9336,N_9206);
nor UO_1038 (O_1038,N_9445,N_9579);
nor UO_1039 (O_1039,N_9706,N_8907);
and UO_1040 (O_1040,N_9408,N_9010);
nor UO_1041 (O_1041,N_8475,N_8999);
nor UO_1042 (O_1042,N_9261,N_9971);
or UO_1043 (O_1043,N_9013,N_9859);
and UO_1044 (O_1044,N_8604,N_8614);
or UO_1045 (O_1045,N_9812,N_9374);
nor UO_1046 (O_1046,N_9210,N_8836);
or UO_1047 (O_1047,N_8430,N_9826);
nand UO_1048 (O_1048,N_8294,N_9017);
or UO_1049 (O_1049,N_8632,N_8043);
nor UO_1050 (O_1050,N_9447,N_8750);
nand UO_1051 (O_1051,N_9277,N_9831);
nand UO_1052 (O_1052,N_8219,N_9790);
or UO_1053 (O_1053,N_9783,N_8585);
and UO_1054 (O_1054,N_9632,N_8361);
or UO_1055 (O_1055,N_8268,N_8398);
nor UO_1056 (O_1056,N_9471,N_8590);
nor UO_1057 (O_1057,N_9935,N_9323);
and UO_1058 (O_1058,N_8600,N_9425);
and UO_1059 (O_1059,N_9349,N_9382);
nor UO_1060 (O_1060,N_8473,N_9057);
and UO_1061 (O_1061,N_9847,N_9291);
or UO_1062 (O_1062,N_9709,N_9772);
and UO_1063 (O_1063,N_8711,N_9715);
and UO_1064 (O_1064,N_8139,N_8827);
and UO_1065 (O_1065,N_9337,N_8474);
nand UO_1066 (O_1066,N_8623,N_9402);
nor UO_1067 (O_1067,N_8381,N_8461);
nor UO_1068 (O_1068,N_9274,N_8890);
nand UO_1069 (O_1069,N_9505,N_9820);
nor UO_1070 (O_1070,N_8751,N_9482);
or UO_1071 (O_1071,N_9191,N_8886);
nor UO_1072 (O_1072,N_9380,N_9419);
nand UO_1073 (O_1073,N_9968,N_9849);
and UO_1074 (O_1074,N_8751,N_9095);
and UO_1075 (O_1075,N_8727,N_8889);
nand UO_1076 (O_1076,N_8773,N_8296);
or UO_1077 (O_1077,N_8848,N_9456);
or UO_1078 (O_1078,N_8598,N_8683);
or UO_1079 (O_1079,N_8718,N_9123);
nand UO_1080 (O_1080,N_8034,N_8004);
nor UO_1081 (O_1081,N_8523,N_9021);
nor UO_1082 (O_1082,N_9798,N_9362);
and UO_1083 (O_1083,N_9214,N_9270);
nor UO_1084 (O_1084,N_8851,N_9395);
or UO_1085 (O_1085,N_8318,N_9739);
nor UO_1086 (O_1086,N_8027,N_9309);
or UO_1087 (O_1087,N_8604,N_8881);
and UO_1088 (O_1088,N_9284,N_9251);
nor UO_1089 (O_1089,N_8697,N_9682);
and UO_1090 (O_1090,N_8361,N_8118);
and UO_1091 (O_1091,N_9565,N_9944);
or UO_1092 (O_1092,N_9131,N_9902);
nor UO_1093 (O_1093,N_9815,N_9688);
and UO_1094 (O_1094,N_9860,N_9967);
or UO_1095 (O_1095,N_9872,N_8802);
and UO_1096 (O_1096,N_8745,N_9254);
and UO_1097 (O_1097,N_8552,N_8766);
or UO_1098 (O_1098,N_9684,N_8298);
and UO_1099 (O_1099,N_9392,N_9579);
and UO_1100 (O_1100,N_8475,N_8217);
nand UO_1101 (O_1101,N_9142,N_9071);
and UO_1102 (O_1102,N_9795,N_8035);
or UO_1103 (O_1103,N_8947,N_8079);
or UO_1104 (O_1104,N_9103,N_8248);
nor UO_1105 (O_1105,N_8250,N_9828);
nor UO_1106 (O_1106,N_8325,N_8949);
and UO_1107 (O_1107,N_9362,N_9949);
xor UO_1108 (O_1108,N_8362,N_9218);
and UO_1109 (O_1109,N_8942,N_8879);
nor UO_1110 (O_1110,N_8335,N_8318);
nor UO_1111 (O_1111,N_9365,N_8406);
nand UO_1112 (O_1112,N_8312,N_9648);
nand UO_1113 (O_1113,N_8600,N_9351);
nor UO_1114 (O_1114,N_8768,N_9388);
nand UO_1115 (O_1115,N_9900,N_9068);
or UO_1116 (O_1116,N_8061,N_9372);
or UO_1117 (O_1117,N_8017,N_9397);
and UO_1118 (O_1118,N_9205,N_8219);
xor UO_1119 (O_1119,N_9395,N_9904);
nand UO_1120 (O_1120,N_9869,N_9562);
nand UO_1121 (O_1121,N_9986,N_8638);
xor UO_1122 (O_1122,N_9855,N_8893);
and UO_1123 (O_1123,N_8670,N_9334);
nand UO_1124 (O_1124,N_8044,N_9797);
nor UO_1125 (O_1125,N_8612,N_9054);
nand UO_1126 (O_1126,N_9399,N_9018);
or UO_1127 (O_1127,N_8309,N_8104);
nand UO_1128 (O_1128,N_8927,N_9102);
or UO_1129 (O_1129,N_8605,N_8181);
or UO_1130 (O_1130,N_9055,N_9045);
nor UO_1131 (O_1131,N_9698,N_8299);
nand UO_1132 (O_1132,N_8353,N_9130);
and UO_1133 (O_1133,N_9270,N_8988);
nor UO_1134 (O_1134,N_8604,N_8404);
or UO_1135 (O_1135,N_9966,N_9618);
nor UO_1136 (O_1136,N_9796,N_8794);
nor UO_1137 (O_1137,N_8174,N_8712);
or UO_1138 (O_1138,N_8847,N_8699);
nor UO_1139 (O_1139,N_8867,N_8116);
nand UO_1140 (O_1140,N_8454,N_8032);
and UO_1141 (O_1141,N_9865,N_9017);
nor UO_1142 (O_1142,N_8265,N_9419);
nand UO_1143 (O_1143,N_8188,N_8501);
and UO_1144 (O_1144,N_9712,N_8913);
and UO_1145 (O_1145,N_9702,N_8360);
nor UO_1146 (O_1146,N_9164,N_8528);
or UO_1147 (O_1147,N_8676,N_8251);
nor UO_1148 (O_1148,N_8192,N_8090);
and UO_1149 (O_1149,N_8430,N_9530);
nand UO_1150 (O_1150,N_9603,N_8592);
nand UO_1151 (O_1151,N_9981,N_8458);
and UO_1152 (O_1152,N_9346,N_9110);
or UO_1153 (O_1153,N_8879,N_9244);
and UO_1154 (O_1154,N_8586,N_9328);
nand UO_1155 (O_1155,N_8438,N_9397);
nor UO_1156 (O_1156,N_9255,N_8117);
nand UO_1157 (O_1157,N_9101,N_9319);
and UO_1158 (O_1158,N_9614,N_8753);
and UO_1159 (O_1159,N_8180,N_8852);
or UO_1160 (O_1160,N_8985,N_8322);
nand UO_1161 (O_1161,N_8300,N_8567);
nand UO_1162 (O_1162,N_8855,N_8561);
and UO_1163 (O_1163,N_8139,N_8169);
nand UO_1164 (O_1164,N_8740,N_8352);
and UO_1165 (O_1165,N_9965,N_9389);
nor UO_1166 (O_1166,N_8498,N_9502);
nor UO_1167 (O_1167,N_8294,N_8322);
or UO_1168 (O_1168,N_8588,N_9590);
nor UO_1169 (O_1169,N_8396,N_9113);
nand UO_1170 (O_1170,N_9135,N_8759);
or UO_1171 (O_1171,N_8426,N_8635);
nor UO_1172 (O_1172,N_8788,N_9250);
and UO_1173 (O_1173,N_9953,N_9003);
or UO_1174 (O_1174,N_9590,N_9596);
nor UO_1175 (O_1175,N_8380,N_9663);
or UO_1176 (O_1176,N_8608,N_8545);
or UO_1177 (O_1177,N_8035,N_9922);
or UO_1178 (O_1178,N_9614,N_9014);
and UO_1179 (O_1179,N_8418,N_9082);
and UO_1180 (O_1180,N_8841,N_8666);
and UO_1181 (O_1181,N_9402,N_8695);
or UO_1182 (O_1182,N_9877,N_8115);
or UO_1183 (O_1183,N_8248,N_9933);
nand UO_1184 (O_1184,N_8536,N_9111);
and UO_1185 (O_1185,N_9303,N_9330);
or UO_1186 (O_1186,N_8017,N_8085);
nor UO_1187 (O_1187,N_9330,N_8221);
nand UO_1188 (O_1188,N_9581,N_8468);
or UO_1189 (O_1189,N_9936,N_9102);
or UO_1190 (O_1190,N_8287,N_9252);
nand UO_1191 (O_1191,N_8289,N_9163);
and UO_1192 (O_1192,N_8606,N_8332);
nand UO_1193 (O_1193,N_8386,N_9319);
nor UO_1194 (O_1194,N_8964,N_9567);
or UO_1195 (O_1195,N_9687,N_9959);
or UO_1196 (O_1196,N_8366,N_9610);
or UO_1197 (O_1197,N_9234,N_8406);
or UO_1198 (O_1198,N_9762,N_8600);
and UO_1199 (O_1199,N_8232,N_9249);
nand UO_1200 (O_1200,N_9553,N_9496);
nor UO_1201 (O_1201,N_9118,N_9955);
or UO_1202 (O_1202,N_9952,N_9945);
xor UO_1203 (O_1203,N_8793,N_8316);
nor UO_1204 (O_1204,N_8103,N_9945);
and UO_1205 (O_1205,N_8394,N_9053);
or UO_1206 (O_1206,N_8006,N_9543);
or UO_1207 (O_1207,N_9441,N_8491);
nor UO_1208 (O_1208,N_8590,N_9925);
or UO_1209 (O_1209,N_9702,N_8937);
and UO_1210 (O_1210,N_8700,N_8124);
nor UO_1211 (O_1211,N_8248,N_8601);
nand UO_1212 (O_1212,N_8572,N_9835);
nand UO_1213 (O_1213,N_9432,N_8605);
nand UO_1214 (O_1214,N_8308,N_9426);
nor UO_1215 (O_1215,N_9082,N_8313);
nand UO_1216 (O_1216,N_9422,N_8330);
or UO_1217 (O_1217,N_9744,N_9880);
or UO_1218 (O_1218,N_9244,N_8968);
and UO_1219 (O_1219,N_8656,N_9978);
and UO_1220 (O_1220,N_9353,N_9011);
or UO_1221 (O_1221,N_8440,N_9536);
or UO_1222 (O_1222,N_8957,N_8463);
nand UO_1223 (O_1223,N_9124,N_8108);
and UO_1224 (O_1224,N_9186,N_9932);
nor UO_1225 (O_1225,N_9927,N_8898);
nor UO_1226 (O_1226,N_9567,N_9981);
or UO_1227 (O_1227,N_9936,N_9759);
and UO_1228 (O_1228,N_8320,N_8260);
nand UO_1229 (O_1229,N_8214,N_9984);
and UO_1230 (O_1230,N_8439,N_9021);
nor UO_1231 (O_1231,N_9197,N_9577);
nand UO_1232 (O_1232,N_8123,N_9811);
nand UO_1233 (O_1233,N_9732,N_8016);
and UO_1234 (O_1234,N_9082,N_8292);
or UO_1235 (O_1235,N_8200,N_9760);
or UO_1236 (O_1236,N_9983,N_8110);
and UO_1237 (O_1237,N_8579,N_9524);
and UO_1238 (O_1238,N_8704,N_8913);
nor UO_1239 (O_1239,N_8332,N_8780);
or UO_1240 (O_1240,N_8008,N_9981);
and UO_1241 (O_1241,N_9268,N_9827);
or UO_1242 (O_1242,N_9523,N_8235);
nand UO_1243 (O_1243,N_8667,N_8608);
or UO_1244 (O_1244,N_8605,N_9051);
and UO_1245 (O_1245,N_8873,N_8143);
or UO_1246 (O_1246,N_9322,N_8125);
or UO_1247 (O_1247,N_8417,N_8119);
nand UO_1248 (O_1248,N_8882,N_9010);
or UO_1249 (O_1249,N_9875,N_9637);
or UO_1250 (O_1250,N_8191,N_8862);
nor UO_1251 (O_1251,N_9553,N_8052);
or UO_1252 (O_1252,N_9322,N_8039);
or UO_1253 (O_1253,N_8780,N_8100);
or UO_1254 (O_1254,N_9524,N_9890);
and UO_1255 (O_1255,N_9353,N_9798);
or UO_1256 (O_1256,N_9190,N_8536);
nor UO_1257 (O_1257,N_8127,N_8785);
and UO_1258 (O_1258,N_9678,N_8984);
nand UO_1259 (O_1259,N_9662,N_9941);
and UO_1260 (O_1260,N_9663,N_8903);
and UO_1261 (O_1261,N_9602,N_9630);
or UO_1262 (O_1262,N_9574,N_9365);
and UO_1263 (O_1263,N_8337,N_8111);
and UO_1264 (O_1264,N_9695,N_8399);
nor UO_1265 (O_1265,N_9623,N_8867);
nand UO_1266 (O_1266,N_9463,N_8785);
nor UO_1267 (O_1267,N_9043,N_8430);
nand UO_1268 (O_1268,N_8764,N_8432);
nand UO_1269 (O_1269,N_9123,N_9149);
and UO_1270 (O_1270,N_8573,N_9299);
and UO_1271 (O_1271,N_8852,N_9711);
nor UO_1272 (O_1272,N_9624,N_9302);
nor UO_1273 (O_1273,N_9582,N_9197);
and UO_1274 (O_1274,N_9873,N_9417);
and UO_1275 (O_1275,N_9582,N_9475);
and UO_1276 (O_1276,N_8798,N_9242);
and UO_1277 (O_1277,N_8108,N_9513);
and UO_1278 (O_1278,N_8481,N_9391);
and UO_1279 (O_1279,N_9571,N_8492);
nand UO_1280 (O_1280,N_9611,N_9881);
nor UO_1281 (O_1281,N_9284,N_9253);
nor UO_1282 (O_1282,N_9688,N_8967);
xor UO_1283 (O_1283,N_9087,N_8105);
nand UO_1284 (O_1284,N_8678,N_9049);
and UO_1285 (O_1285,N_8173,N_9830);
xnor UO_1286 (O_1286,N_8051,N_8312);
nor UO_1287 (O_1287,N_9184,N_8652);
nor UO_1288 (O_1288,N_8041,N_9393);
nor UO_1289 (O_1289,N_8677,N_9395);
or UO_1290 (O_1290,N_8622,N_8309);
nor UO_1291 (O_1291,N_9390,N_9833);
or UO_1292 (O_1292,N_9056,N_8544);
nor UO_1293 (O_1293,N_8459,N_8561);
nand UO_1294 (O_1294,N_9925,N_8081);
nand UO_1295 (O_1295,N_8751,N_8597);
and UO_1296 (O_1296,N_9471,N_8772);
nor UO_1297 (O_1297,N_9516,N_8347);
nand UO_1298 (O_1298,N_9643,N_9389);
or UO_1299 (O_1299,N_8370,N_9201);
nand UO_1300 (O_1300,N_8541,N_9889);
nor UO_1301 (O_1301,N_8210,N_8713);
nand UO_1302 (O_1302,N_8109,N_8446);
and UO_1303 (O_1303,N_9980,N_9172);
or UO_1304 (O_1304,N_8349,N_9453);
nor UO_1305 (O_1305,N_9414,N_9032);
nand UO_1306 (O_1306,N_9311,N_8531);
nor UO_1307 (O_1307,N_9872,N_8211);
nor UO_1308 (O_1308,N_9225,N_8035);
or UO_1309 (O_1309,N_8394,N_9177);
and UO_1310 (O_1310,N_9434,N_9728);
nand UO_1311 (O_1311,N_9735,N_9060);
nand UO_1312 (O_1312,N_8422,N_8819);
nor UO_1313 (O_1313,N_8214,N_9509);
nor UO_1314 (O_1314,N_8272,N_8795);
nor UO_1315 (O_1315,N_8325,N_8333);
nand UO_1316 (O_1316,N_8701,N_8512);
nor UO_1317 (O_1317,N_8076,N_8271);
nor UO_1318 (O_1318,N_8934,N_8793);
and UO_1319 (O_1319,N_8430,N_9282);
and UO_1320 (O_1320,N_9330,N_9482);
nand UO_1321 (O_1321,N_8181,N_9150);
or UO_1322 (O_1322,N_9867,N_8214);
and UO_1323 (O_1323,N_8789,N_9003);
and UO_1324 (O_1324,N_9930,N_8606);
and UO_1325 (O_1325,N_8241,N_8908);
nor UO_1326 (O_1326,N_9614,N_9813);
nand UO_1327 (O_1327,N_9877,N_9470);
nand UO_1328 (O_1328,N_8569,N_9333);
and UO_1329 (O_1329,N_8203,N_9362);
and UO_1330 (O_1330,N_9665,N_9401);
nand UO_1331 (O_1331,N_8074,N_8168);
nand UO_1332 (O_1332,N_9610,N_8909);
nor UO_1333 (O_1333,N_8762,N_9891);
nand UO_1334 (O_1334,N_8951,N_9420);
or UO_1335 (O_1335,N_8810,N_8588);
and UO_1336 (O_1336,N_9592,N_9646);
nand UO_1337 (O_1337,N_8232,N_8013);
nor UO_1338 (O_1338,N_8458,N_8050);
nor UO_1339 (O_1339,N_8024,N_9739);
nor UO_1340 (O_1340,N_9900,N_8224);
and UO_1341 (O_1341,N_8324,N_8401);
and UO_1342 (O_1342,N_8265,N_9839);
and UO_1343 (O_1343,N_8992,N_8901);
nand UO_1344 (O_1344,N_9221,N_9512);
nor UO_1345 (O_1345,N_9775,N_9881);
nand UO_1346 (O_1346,N_8834,N_9443);
or UO_1347 (O_1347,N_8059,N_8334);
and UO_1348 (O_1348,N_9080,N_8482);
nand UO_1349 (O_1349,N_9041,N_8289);
nand UO_1350 (O_1350,N_8361,N_8274);
or UO_1351 (O_1351,N_8903,N_9812);
nand UO_1352 (O_1352,N_8596,N_9337);
and UO_1353 (O_1353,N_9345,N_8493);
or UO_1354 (O_1354,N_9965,N_8074);
nand UO_1355 (O_1355,N_8702,N_8815);
nor UO_1356 (O_1356,N_9219,N_8885);
nand UO_1357 (O_1357,N_9830,N_9539);
nand UO_1358 (O_1358,N_9683,N_9261);
nand UO_1359 (O_1359,N_8425,N_8779);
and UO_1360 (O_1360,N_8871,N_8598);
nor UO_1361 (O_1361,N_8752,N_9258);
and UO_1362 (O_1362,N_9033,N_8672);
and UO_1363 (O_1363,N_8047,N_9370);
nor UO_1364 (O_1364,N_8298,N_8170);
nor UO_1365 (O_1365,N_9330,N_8184);
and UO_1366 (O_1366,N_9293,N_9816);
and UO_1367 (O_1367,N_9063,N_9739);
or UO_1368 (O_1368,N_8971,N_9562);
nor UO_1369 (O_1369,N_9674,N_9206);
or UO_1370 (O_1370,N_8545,N_8943);
and UO_1371 (O_1371,N_9190,N_9243);
or UO_1372 (O_1372,N_8666,N_8105);
and UO_1373 (O_1373,N_8071,N_9459);
or UO_1374 (O_1374,N_9334,N_8604);
and UO_1375 (O_1375,N_8958,N_9670);
and UO_1376 (O_1376,N_8126,N_8400);
or UO_1377 (O_1377,N_8763,N_8131);
nand UO_1378 (O_1378,N_8147,N_9245);
and UO_1379 (O_1379,N_8315,N_9833);
or UO_1380 (O_1380,N_8556,N_8672);
nand UO_1381 (O_1381,N_9747,N_9865);
and UO_1382 (O_1382,N_8085,N_8646);
or UO_1383 (O_1383,N_9058,N_8000);
or UO_1384 (O_1384,N_9847,N_8488);
nand UO_1385 (O_1385,N_9913,N_8054);
nand UO_1386 (O_1386,N_8784,N_9542);
or UO_1387 (O_1387,N_8642,N_8846);
nor UO_1388 (O_1388,N_8735,N_8334);
nand UO_1389 (O_1389,N_8800,N_8181);
nand UO_1390 (O_1390,N_8191,N_8618);
nor UO_1391 (O_1391,N_8394,N_8531);
nand UO_1392 (O_1392,N_8260,N_9498);
nor UO_1393 (O_1393,N_8483,N_8060);
nand UO_1394 (O_1394,N_8294,N_8231);
nand UO_1395 (O_1395,N_9722,N_8505);
nor UO_1396 (O_1396,N_9290,N_8970);
nand UO_1397 (O_1397,N_8661,N_9415);
nor UO_1398 (O_1398,N_8692,N_9373);
and UO_1399 (O_1399,N_9086,N_8483);
nand UO_1400 (O_1400,N_8158,N_8497);
and UO_1401 (O_1401,N_9113,N_8348);
and UO_1402 (O_1402,N_8661,N_9557);
nor UO_1403 (O_1403,N_9153,N_9529);
nand UO_1404 (O_1404,N_8262,N_8440);
nor UO_1405 (O_1405,N_9215,N_9932);
and UO_1406 (O_1406,N_8167,N_8977);
or UO_1407 (O_1407,N_8203,N_9645);
nand UO_1408 (O_1408,N_8125,N_8443);
and UO_1409 (O_1409,N_8550,N_8382);
and UO_1410 (O_1410,N_9645,N_9694);
nand UO_1411 (O_1411,N_9910,N_8507);
nor UO_1412 (O_1412,N_8031,N_8877);
nor UO_1413 (O_1413,N_9810,N_8424);
or UO_1414 (O_1414,N_9064,N_9759);
and UO_1415 (O_1415,N_9598,N_9929);
nand UO_1416 (O_1416,N_8464,N_9663);
and UO_1417 (O_1417,N_8428,N_9577);
or UO_1418 (O_1418,N_9108,N_9189);
nor UO_1419 (O_1419,N_8575,N_8441);
nand UO_1420 (O_1420,N_8748,N_8721);
nor UO_1421 (O_1421,N_9829,N_9654);
and UO_1422 (O_1422,N_9841,N_9807);
and UO_1423 (O_1423,N_8386,N_9897);
and UO_1424 (O_1424,N_8688,N_9693);
nor UO_1425 (O_1425,N_8736,N_9782);
nor UO_1426 (O_1426,N_8085,N_9034);
nor UO_1427 (O_1427,N_9454,N_8860);
nor UO_1428 (O_1428,N_8606,N_8302);
nor UO_1429 (O_1429,N_8894,N_8570);
nand UO_1430 (O_1430,N_8237,N_8902);
nor UO_1431 (O_1431,N_9562,N_8245);
nand UO_1432 (O_1432,N_8363,N_8289);
nand UO_1433 (O_1433,N_8592,N_8182);
and UO_1434 (O_1434,N_9877,N_8720);
and UO_1435 (O_1435,N_8538,N_9610);
xor UO_1436 (O_1436,N_9642,N_9265);
nand UO_1437 (O_1437,N_8223,N_9196);
nand UO_1438 (O_1438,N_8039,N_8586);
nor UO_1439 (O_1439,N_8895,N_9822);
and UO_1440 (O_1440,N_9416,N_8465);
nand UO_1441 (O_1441,N_8909,N_9387);
nor UO_1442 (O_1442,N_9137,N_8656);
and UO_1443 (O_1443,N_8716,N_8382);
or UO_1444 (O_1444,N_9931,N_8619);
nand UO_1445 (O_1445,N_9243,N_8379);
nor UO_1446 (O_1446,N_8951,N_8024);
nand UO_1447 (O_1447,N_8201,N_9562);
and UO_1448 (O_1448,N_9674,N_8706);
or UO_1449 (O_1449,N_9540,N_9508);
or UO_1450 (O_1450,N_8522,N_8710);
or UO_1451 (O_1451,N_9868,N_8132);
and UO_1452 (O_1452,N_8347,N_8194);
nand UO_1453 (O_1453,N_9124,N_9126);
nor UO_1454 (O_1454,N_9343,N_8759);
nor UO_1455 (O_1455,N_8141,N_8790);
nor UO_1456 (O_1456,N_9639,N_8393);
or UO_1457 (O_1457,N_8911,N_8634);
nand UO_1458 (O_1458,N_8459,N_8598);
or UO_1459 (O_1459,N_8979,N_8845);
nand UO_1460 (O_1460,N_9030,N_9444);
nor UO_1461 (O_1461,N_8398,N_8921);
and UO_1462 (O_1462,N_8496,N_9192);
nand UO_1463 (O_1463,N_8593,N_9361);
or UO_1464 (O_1464,N_8215,N_8871);
nor UO_1465 (O_1465,N_8411,N_9796);
nand UO_1466 (O_1466,N_9566,N_9856);
or UO_1467 (O_1467,N_9338,N_9937);
or UO_1468 (O_1468,N_8969,N_8828);
and UO_1469 (O_1469,N_9047,N_8124);
or UO_1470 (O_1470,N_9761,N_8721);
nor UO_1471 (O_1471,N_8819,N_8519);
xor UO_1472 (O_1472,N_8600,N_8263);
or UO_1473 (O_1473,N_8996,N_8171);
or UO_1474 (O_1474,N_8789,N_8145);
or UO_1475 (O_1475,N_9354,N_8278);
nor UO_1476 (O_1476,N_8447,N_8278);
nand UO_1477 (O_1477,N_8891,N_9053);
and UO_1478 (O_1478,N_8948,N_9779);
or UO_1479 (O_1479,N_8290,N_9076);
nand UO_1480 (O_1480,N_9125,N_8308);
nand UO_1481 (O_1481,N_9217,N_9726);
nand UO_1482 (O_1482,N_8197,N_8530);
nand UO_1483 (O_1483,N_8419,N_9513);
or UO_1484 (O_1484,N_8122,N_8372);
or UO_1485 (O_1485,N_9540,N_9394);
and UO_1486 (O_1486,N_9136,N_8076);
or UO_1487 (O_1487,N_8721,N_8203);
nor UO_1488 (O_1488,N_8451,N_9326);
nand UO_1489 (O_1489,N_8752,N_8203);
or UO_1490 (O_1490,N_9740,N_9062);
and UO_1491 (O_1491,N_9438,N_9173);
or UO_1492 (O_1492,N_9432,N_8832);
or UO_1493 (O_1493,N_8141,N_8221);
and UO_1494 (O_1494,N_8951,N_9997);
and UO_1495 (O_1495,N_9302,N_9233);
nor UO_1496 (O_1496,N_8467,N_8768);
or UO_1497 (O_1497,N_9822,N_8049);
or UO_1498 (O_1498,N_9604,N_9629);
nand UO_1499 (O_1499,N_8384,N_8413);
endmodule