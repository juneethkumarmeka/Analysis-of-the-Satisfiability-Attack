module basic_5000_50000_5000_25_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_2214,In_4576);
nor U1 (N_1,In_3200,In_4172);
nor U2 (N_2,In_2847,In_450);
and U3 (N_3,In_2608,In_146);
and U4 (N_4,In_4622,In_335);
xnor U5 (N_5,In_4814,In_2171);
and U6 (N_6,In_2488,In_1400);
nor U7 (N_7,In_3800,In_3240);
or U8 (N_8,In_1461,In_2117);
nand U9 (N_9,In_4104,In_2668);
xnor U10 (N_10,In_769,In_2567);
and U11 (N_11,In_2445,In_4951);
nand U12 (N_12,In_457,In_3688);
nand U13 (N_13,In_1862,In_3958);
and U14 (N_14,In_4584,In_339);
and U15 (N_15,In_3488,In_4975);
or U16 (N_16,In_1677,In_4707);
nand U17 (N_17,In_2890,In_3032);
xor U18 (N_18,In_4564,In_4846);
nand U19 (N_19,In_3299,In_3636);
xnor U20 (N_20,In_4596,In_4363);
nand U21 (N_21,In_3565,In_4725);
or U22 (N_22,In_1494,In_2741);
xor U23 (N_23,In_2,In_3214);
and U24 (N_24,In_3450,In_1625);
or U25 (N_25,In_2589,In_662);
nor U26 (N_26,In_2563,In_117);
nor U27 (N_27,In_3393,In_3180);
nor U28 (N_28,In_2813,In_4991);
nor U29 (N_29,In_2732,In_434);
and U30 (N_30,In_1323,In_3763);
nor U31 (N_31,In_4849,In_3655);
and U32 (N_32,In_3169,In_2487);
nor U33 (N_33,In_578,In_137);
xnor U34 (N_34,In_559,In_3802);
nor U35 (N_35,In_475,In_3713);
xnor U36 (N_36,In_888,In_3796);
nand U37 (N_37,In_665,In_639);
or U38 (N_38,In_1420,In_3339);
nor U39 (N_39,In_4842,In_1962);
or U40 (N_40,In_1208,In_69);
and U41 (N_41,In_4890,In_4536);
or U42 (N_42,In_1104,In_1140);
nor U43 (N_43,In_4010,In_1412);
xor U44 (N_44,In_2226,In_3257);
and U45 (N_45,In_4838,In_2225);
nor U46 (N_46,In_4482,In_1541);
xor U47 (N_47,In_325,In_1610);
xnor U48 (N_48,In_4452,In_677);
xnor U49 (N_49,In_2158,In_2256);
xor U50 (N_50,In_937,In_98);
or U51 (N_51,In_245,In_4784);
nand U52 (N_52,In_1313,In_2235);
and U53 (N_53,In_3203,In_142);
and U54 (N_54,In_2877,In_3593);
xor U55 (N_55,In_566,In_1266);
nand U56 (N_56,In_4278,In_984);
nor U57 (N_57,In_3185,In_957);
nand U58 (N_58,In_2764,In_3624);
or U59 (N_59,In_1711,In_4261);
or U60 (N_60,In_1054,In_2245);
and U61 (N_61,In_3657,In_2830);
or U62 (N_62,In_1404,In_220);
and U63 (N_63,In_3569,In_3972);
nor U64 (N_64,In_1315,In_827);
or U65 (N_65,In_2963,In_261);
or U66 (N_66,In_4511,In_1675);
xnor U67 (N_67,In_2693,In_3838);
nand U68 (N_68,In_2818,In_1828);
nand U69 (N_69,In_1339,In_4603);
or U70 (N_70,In_3816,In_3403);
xnor U71 (N_71,In_3392,In_2377);
and U72 (N_72,In_2882,In_4309);
and U73 (N_73,In_1361,In_2146);
or U74 (N_74,In_4444,In_1952);
xnor U75 (N_75,In_4978,In_648);
nor U76 (N_76,In_2585,In_1255);
and U77 (N_77,In_4754,In_417);
and U78 (N_78,In_4762,In_2701);
and U79 (N_79,In_4864,In_2035);
xnor U80 (N_80,In_49,In_2573);
and U81 (N_81,In_1394,In_2466);
xnor U82 (N_82,In_3464,In_176);
or U83 (N_83,In_2221,In_2948);
and U84 (N_84,In_3093,In_3253);
and U85 (N_85,In_4717,In_2874);
and U86 (N_86,In_3060,In_343);
xor U87 (N_87,In_2926,In_4569);
or U88 (N_88,In_2736,In_4456);
and U89 (N_89,In_3276,In_2189);
or U90 (N_90,In_3009,In_4001);
xnor U91 (N_91,In_3415,In_3159);
and U92 (N_92,In_4225,In_519);
and U93 (N_93,In_787,In_851);
nand U94 (N_94,In_740,In_4934);
or U95 (N_95,In_1654,In_697);
nand U96 (N_96,In_2233,In_3505);
nor U97 (N_97,In_37,In_3387);
or U98 (N_98,In_3806,In_3943);
and U99 (N_99,In_2938,In_2443);
or U100 (N_100,In_359,In_35);
or U101 (N_101,In_702,In_3601);
nor U102 (N_102,In_4961,In_100);
and U103 (N_103,In_3422,In_4562);
nand U104 (N_104,In_268,In_1396);
nand U105 (N_105,In_1892,In_2496);
xnor U106 (N_106,In_4966,In_338);
nor U107 (N_107,In_938,In_3735);
and U108 (N_108,In_4906,In_2160);
nor U109 (N_109,In_599,In_1035);
or U110 (N_110,In_90,In_4165);
nor U111 (N_111,In_3150,In_1919);
or U112 (N_112,In_2578,In_4559);
nand U113 (N_113,In_2424,In_3099);
or U114 (N_114,In_2248,In_2694);
and U115 (N_115,In_1101,In_4072);
nand U116 (N_116,In_3467,In_4310);
nand U117 (N_117,In_4221,In_4874);
nor U118 (N_118,In_131,In_4568);
nor U119 (N_119,In_2678,In_308);
and U120 (N_120,In_4630,In_1572);
nor U121 (N_121,In_1302,In_1940);
and U122 (N_122,In_1434,In_357);
xor U123 (N_123,In_3506,In_4346);
nor U124 (N_124,In_2329,In_2744);
and U125 (N_125,In_206,In_3518);
or U126 (N_126,In_2613,In_201);
or U127 (N_127,In_111,In_1145);
xor U128 (N_128,In_3545,In_1126);
and U129 (N_129,In_1188,In_4818);
and U130 (N_130,In_1656,In_4583);
nor U131 (N_131,In_4698,In_22);
xor U132 (N_132,In_74,In_4997);
and U133 (N_133,In_813,In_3237);
xnor U134 (N_134,In_2902,In_4872);
or U135 (N_135,In_996,In_208);
and U136 (N_136,In_1578,In_4429);
and U137 (N_137,In_3566,In_977);
xor U138 (N_138,In_700,In_372);
xnor U139 (N_139,In_604,In_3373);
nand U140 (N_140,In_2116,In_66);
or U141 (N_141,In_2331,In_4548);
nor U142 (N_142,In_4572,In_2104);
nor U143 (N_143,In_4254,In_2522);
and U144 (N_144,In_4915,In_3644);
nand U145 (N_145,In_4718,In_3001);
xor U146 (N_146,In_3508,In_4445);
xor U147 (N_147,In_1866,In_632);
or U148 (N_148,In_1148,In_480);
or U149 (N_149,In_687,In_3496);
xor U150 (N_150,In_3535,In_961);
nor U151 (N_151,In_377,In_3143);
and U152 (N_152,In_635,In_1053);
nor U153 (N_153,In_1813,In_3115);
nor U154 (N_154,In_1336,In_1926);
and U155 (N_155,In_307,In_570);
and U156 (N_156,In_2346,In_257);
nor U157 (N_157,In_751,In_2727);
or U158 (N_158,In_316,In_4777);
nor U159 (N_159,In_336,In_1069);
or U160 (N_160,In_2760,In_4831);
xnor U161 (N_161,In_1128,In_3628);
nor U162 (N_162,In_4637,In_2971);
nand U163 (N_163,In_2396,In_1679);
or U164 (N_164,In_1614,In_2807);
xor U165 (N_165,In_724,In_3707);
xor U166 (N_166,In_3483,In_3348);
and U167 (N_167,In_25,In_2539);
xnor U168 (N_168,In_2577,In_2389);
and U169 (N_169,In_215,In_302);
and U170 (N_170,In_3604,In_1523);
nand U171 (N_171,In_4928,In_2211);
nor U172 (N_172,In_3794,In_1582);
nor U173 (N_173,In_1213,In_2754);
or U174 (N_174,In_972,In_3942);
and U175 (N_175,In_3853,In_2328);
nand U176 (N_176,In_1534,In_1110);
xnor U177 (N_177,In_513,In_591);
xor U178 (N_178,In_534,In_3005);
nor U179 (N_179,In_4329,In_4667);
nor U180 (N_180,In_561,In_4832);
nor U181 (N_181,In_1540,In_706);
and U182 (N_182,In_2497,In_2817);
and U183 (N_183,In_4744,In_1489);
nor U184 (N_184,In_4401,In_3105);
and U185 (N_185,In_2936,In_1059);
and U186 (N_186,In_3771,In_2870);
and U187 (N_187,In_24,In_1560);
nor U188 (N_188,In_4813,In_4780);
nand U189 (N_189,In_1267,In_2651);
xnor U190 (N_190,In_4192,In_1611);
nand U191 (N_191,In_3044,In_2940);
or U192 (N_192,In_2291,In_4294);
xor U193 (N_193,In_1387,In_4478);
or U194 (N_194,In_1165,In_3663);
or U195 (N_195,In_4407,In_4328);
or U196 (N_196,In_2342,In_330);
and U197 (N_197,In_2683,In_4626);
nor U198 (N_198,In_3848,In_3936);
xnor U199 (N_199,In_4948,In_1229);
xnor U200 (N_200,In_3772,In_3017);
and U201 (N_201,In_766,In_3109);
xor U202 (N_202,In_444,In_3474);
xor U203 (N_203,In_3256,In_1997);
nand U204 (N_204,In_2460,In_1383);
or U205 (N_205,In_4235,In_471);
or U206 (N_206,In_4674,In_1485);
and U207 (N_207,In_1057,In_3858);
nor U208 (N_208,In_1401,In_56);
or U209 (N_209,In_2878,In_2257);
nand U210 (N_210,In_1080,In_1143);
or U211 (N_211,In_2663,In_1009);
or U212 (N_212,In_3343,In_2723);
xnor U213 (N_213,In_2274,In_212);
xnor U214 (N_214,In_3807,In_4435);
and U215 (N_215,In_2849,In_1586);
nand U216 (N_216,In_4306,In_224);
or U217 (N_217,In_4402,In_4681);
nand U218 (N_218,In_4161,In_3291);
and U219 (N_219,In_3597,In_2434);
nand U220 (N_220,In_28,In_3964);
or U221 (N_221,In_1472,In_4140);
xnor U222 (N_222,In_1773,In_1929);
nor U223 (N_223,In_1694,In_2250);
nand U224 (N_224,In_1884,In_4910);
nor U225 (N_225,In_637,In_4312);
or U226 (N_226,In_895,In_2333);
and U227 (N_227,In_4947,In_2494);
nand U228 (N_228,In_843,In_3426);
nand U229 (N_229,In_2929,In_2476);
xnor U230 (N_230,In_1024,In_3420);
nand U231 (N_231,In_2832,In_4038);
xor U232 (N_232,In_699,In_4246);
or U233 (N_233,In_1139,In_3578);
xnor U234 (N_234,In_3114,In_2699);
xnor U235 (N_235,In_3304,In_1349);
nand U236 (N_236,In_4544,In_1294);
nor U237 (N_237,In_182,In_2096);
or U238 (N_238,In_1506,In_2144);
nand U239 (N_239,In_4214,In_499);
and U240 (N_240,In_2360,In_1214);
nor U241 (N_241,In_725,In_850);
xor U242 (N_242,In_1844,In_2889);
and U243 (N_243,In_2822,In_3768);
or U244 (N_244,In_4411,In_68);
nor U245 (N_245,In_1580,In_776);
and U246 (N_246,In_4446,In_2408);
nor U247 (N_247,In_1777,In_2587);
nor U248 (N_248,In_1367,In_1298);
nand U249 (N_249,In_1486,In_2285);
xor U250 (N_250,In_1971,In_4183);
nand U251 (N_251,In_1525,In_4169);
nor U252 (N_252,In_1236,In_1549);
or U253 (N_253,In_4336,In_3736);
nor U254 (N_254,In_3085,In_3079);
xnor U255 (N_255,In_2196,In_1303);
xnor U256 (N_256,In_775,In_2569);
and U257 (N_257,In_833,In_3012);
nand U258 (N_258,In_1920,In_4537);
and U259 (N_259,In_1835,In_1175);
and U260 (N_260,In_2630,In_2247);
or U261 (N_261,In_3424,In_3011);
xor U262 (N_262,In_3481,In_2195);
nand U263 (N_263,In_4281,In_3619);
and U264 (N_264,In_600,In_3504);
xnor U265 (N_265,In_2486,In_232);
xor U266 (N_266,In_3473,In_1766);
xnor U267 (N_267,In_3466,In_2553);
nor U268 (N_268,In_4403,In_3478);
xnor U269 (N_269,In_3544,In_4956);
and U270 (N_270,In_183,In_4260);
xor U271 (N_271,In_2307,In_3219);
nand U272 (N_272,In_3563,In_4550);
nor U273 (N_273,In_1855,In_2115);
nand U274 (N_274,In_3808,In_2136);
and U275 (N_275,In_289,In_862);
xnor U276 (N_276,In_4413,In_321);
nand U277 (N_277,In_2323,In_1697);
and U278 (N_278,In_713,In_408);
and U279 (N_279,In_3446,In_2781);
and U280 (N_280,In_2062,In_180);
or U281 (N_281,In_219,In_1);
or U282 (N_282,In_2498,In_1391);
nand U283 (N_283,In_4676,In_1762);
nor U284 (N_284,In_741,In_3674);
nand U285 (N_285,In_3318,In_463);
nand U286 (N_286,In_2384,In_3133);
and U287 (N_287,In_4259,In_145);
and U288 (N_288,In_4468,In_489);
and U289 (N_289,In_4922,In_4936);
xor U290 (N_290,In_2427,In_4073);
and U291 (N_291,In_1842,In_4206);
nor U292 (N_292,In_4783,In_3618);
nor U293 (N_293,In_358,In_4076);
xnor U294 (N_294,In_4412,In_1763);
nor U295 (N_295,In_571,In_4766);
nor U296 (N_296,In_3698,In_4641);
xor U297 (N_297,In_4332,In_1025);
xnor U298 (N_298,In_314,In_233);
xnor U299 (N_299,In_428,In_750);
and U300 (N_300,In_33,In_2834);
xor U301 (N_301,In_2441,In_2049);
xnor U302 (N_302,In_2395,In_1512);
xor U303 (N_303,In_3208,In_1853);
xnor U304 (N_304,In_1969,In_798);
or U305 (N_305,In_1160,In_642);
or U306 (N_306,In_732,In_1871);
xor U307 (N_307,In_1681,In_3377);
and U308 (N_308,In_555,In_2432);
nand U309 (N_309,In_2960,In_1432);
nor U310 (N_310,In_4670,In_2737);
or U311 (N_311,In_3340,In_3465);
and U312 (N_312,In_2875,In_2511);
and U313 (N_313,In_4409,In_4949);
nand U314 (N_314,In_1219,In_2230);
or U315 (N_315,In_905,In_1822);
xor U316 (N_316,In_1861,In_3441);
xnor U317 (N_317,In_254,In_3658);
nor U318 (N_318,In_326,In_3090);
or U319 (N_319,In_3234,In_3595);
and U320 (N_320,In_4355,In_4252);
nand U321 (N_321,In_617,In_3551);
nor U322 (N_322,In_2249,In_2201);
nor U323 (N_323,In_2504,In_2893);
nor U324 (N_324,In_834,In_2625);
xor U325 (N_325,In_2583,In_4597);
nand U326 (N_326,In_527,In_3954);
or U327 (N_327,In_4437,In_535);
and U328 (N_328,In_2361,In_3919);
nand U329 (N_329,In_2648,In_3194);
and U330 (N_330,In_1498,In_3306);
xnor U331 (N_331,In_2021,In_1501);
and U332 (N_332,In_2510,In_3730);
nor U333 (N_333,In_1370,In_2927);
nor U334 (N_334,In_46,In_2658);
and U335 (N_335,In_2961,In_3589);
nand U336 (N_336,In_4048,In_3137);
and U337 (N_337,In_970,In_2854);
xnor U338 (N_338,In_1173,In_3096);
nor U339 (N_339,In_3696,In_1182);
nand U340 (N_340,In_237,In_2362);
nand U341 (N_341,In_3358,In_1118);
xnor U342 (N_342,In_2205,In_4022);
xnor U343 (N_343,In_3899,In_890);
xor U344 (N_344,In_1860,In_3100);
and U345 (N_345,In_3705,In_2685);
xor U346 (N_346,In_1598,In_1450);
nand U347 (N_347,In_3434,In_2857);
and U348 (N_348,In_1123,In_2707);
nand U349 (N_349,In_4506,In_3372);
nand U350 (N_350,In_2325,In_4602);
nand U351 (N_351,In_4615,In_1590);
and U352 (N_352,In_2976,In_2002);
xnor U353 (N_353,In_1975,In_2916);
and U354 (N_354,In_3469,In_759);
nand U355 (N_355,In_1960,In_1588);
xnor U356 (N_356,In_1648,In_3832);
or U357 (N_357,In_2197,In_501);
or U358 (N_358,In_3877,In_4428);
nor U359 (N_359,In_1505,In_2763);
nand U360 (N_360,In_200,In_2458);
xnor U361 (N_361,In_4067,In_2442);
nand U362 (N_362,In_4954,In_2808);
and U363 (N_363,In_1904,In_3245);
and U364 (N_364,In_3228,In_2789);
or U365 (N_365,In_2611,In_2646);
or U366 (N_366,In_3065,In_4202);
xor U367 (N_367,In_3632,In_1639);
or U368 (N_368,In_2311,In_3834);
and U369 (N_369,In_4111,In_1829);
nand U370 (N_370,In_3052,In_3945);
xor U371 (N_371,In_299,In_854);
nor U372 (N_372,In_2181,In_2097);
xnor U373 (N_373,In_4496,In_135);
nor U374 (N_374,In_891,In_332);
nor U375 (N_375,In_1493,In_3725);
nand U376 (N_376,In_576,In_4440);
and U377 (N_377,In_1528,In_2549);
nor U378 (N_378,In_3436,In_4491);
nor U379 (N_379,In_72,In_3210);
xnor U380 (N_380,In_835,In_1942);
nor U381 (N_381,In_2503,In_4099);
and U382 (N_382,In_2066,In_2556);
xor U383 (N_383,In_3334,In_805);
and U384 (N_384,In_2239,In_3748);
xor U385 (N_385,In_1655,In_719);
xnor U386 (N_386,In_853,In_2572);
nor U387 (N_387,In_2244,In_4231);
nand U388 (N_388,In_2977,In_1778);
nand U389 (N_389,In_2842,In_2526);
or U390 (N_390,In_4899,In_1760);
nor U391 (N_391,In_3171,In_446);
or U392 (N_392,In_696,In_2751);
and U393 (N_393,In_1562,In_2785);
nor U394 (N_394,In_3879,In_156);
xor U395 (N_395,In_4772,In_898);
xnor U396 (N_396,In_4387,In_3692);
or U397 (N_397,In_3991,In_2345);
xor U398 (N_398,In_1637,In_288);
nand U399 (N_399,In_4493,In_2406);
nor U400 (N_400,In_491,In_3579);
and U401 (N_401,In_3388,In_985);
and U402 (N_402,In_2644,In_2080);
xnor U403 (N_403,In_558,In_2538);
or U404 (N_404,In_1407,In_4663);
nor U405 (N_405,In_4366,In_881);
and U406 (N_406,In_3611,In_3835);
xnor U407 (N_407,In_1807,In_3330);
and U408 (N_408,In_1972,In_3775);
nor U409 (N_409,In_419,In_778);
nor U410 (N_410,In_4,In_3801);
or U411 (N_411,In_4324,In_3074);
or U412 (N_412,In_974,In_1288);
or U413 (N_413,In_2680,In_794);
xor U414 (N_414,In_351,In_2018);
xor U415 (N_415,In_3984,In_1487);
nand U416 (N_416,In_2617,In_4530);
or U417 (N_417,In_2622,In_1774);
xor U418 (N_418,In_185,In_4664);
nand U419 (N_419,In_2547,In_3867);
xor U420 (N_420,In_2495,In_3831);
or U421 (N_421,In_2895,In_1153);
nor U422 (N_422,In_2787,In_2672);
or U423 (N_423,In_2967,In_2453);
nand U424 (N_424,In_560,In_384);
nand U425 (N_425,In_1812,In_966);
or U426 (N_426,In_2816,In_3917);
or U427 (N_427,In_1682,In_949);
nor U428 (N_428,In_388,In_3587);
and U429 (N_429,In_102,In_986);
or U430 (N_430,In_2480,In_777);
nand U431 (N_431,In_2966,In_3026);
nor U432 (N_432,In_1470,In_2492);
and U433 (N_433,In_1047,In_3818);
xor U434 (N_434,In_540,In_4694);
and U435 (N_435,In_4495,In_4981);
or U436 (N_436,In_2861,In_598);
nand U437 (N_437,In_2845,In_3108);
and U438 (N_438,In_2319,In_1845);
or U439 (N_439,In_3347,In_3195);
or U440 (N_440,In_93,In_1410);
or U441 (N_441,In_3212,In_3070);
nand U442 (N_442,In_2083,In_187);
or U443 (N_443,In_1547,In_4416);
and U444 (N_444,In_4893,In_508);
xor U445 (N_445,In_886,In_2555);
and U446 (N_446,In_1692,In_2054);
nand U447 (N_447,In_3091,In_2521);
xnor U448 (N_448,In_3843,In_2414);
or U449 (N_449,In_1631,In_1877);
nor U450 (N_450,In_95,In_2700);
xnor U451 (N_451,In_1245,In_4904);
xor U452 (N_452,In_659,In_375);
and U453 (N_453,In_407,In_3718);
and U454 (N_454,In_4012,In_935);
or U455 (N_455,In_4251,In_3670);
or U456 (N_456,In_4984,In_1258);
nor U457 (N_457,In_147,In_4770);
or U458 (N_458,In_4205,In_2720);
nand U459 (N_459,In_189,In_171);
and U460 (N_460,In_2695,In_1851);
nand U461 (N_461,In_4529,In_4851);
and U462 (N_462,In_1089,In_251);
nor U463 (N_463,In_3847,In_235);
nor U464 (N_464,In_4662,In_1604);
xnor U465 (N_465,In_1981,In_1429);
or U466 (N_466,In_4425,In_1193);
or U467 (N_467,In_4862,In_2184);
and U468 (N_468,In_3264,In_4937);
or U469 (N_469,In_4273,In_3815);
and U470 (N_470,In_3897,In_1242);
and U471 (N_471,In_1841,In_3191);
nand U472 (N_472,In_2517,In_3173);
or U473 (N_473,In_3432,In_476);
and U474 (N_474,In_4907,In_3872);
xnor U475 (N_475,In_1244,In_3206);
xor U476 (N_476,In_4215,In_4656);
nand U477 (N_477,In_1990,In_1748);
xor U478 (N_478,In_109,In_4642);
and U479 (N_479,In_202,In_337);
nor U480 (N_480,In_2490,In_1230);
and U481 (N_481,In_158,In_686);
nand U482 (N_482,In_2766,In_1696);
or U483 (N_483,In_4586,In_4480);
nor U484 (N_484,In_928,In_2381);
xnor U485 (N_485,In_2440,In_3665);
xor U486 (N_486,In_2979,In_4066);
nor U487 (N_487,In_2472,In_1462);
nor U488 (N_488,In_4341,In_356);
nand U489 (N_489,In_1466,In_1559);
or U490 (N_490,In_1911,In_2600);
nand U491 (N_491,In_4392,In_317);
nor U492 (N_492,In_4088,In_2429);
nand U493 (N_493,In_141,In_1949);
or U494 (N_494,In_4349,In_892);
nand U495 (N_495,In_4953,In_4512);
nand U496 (N_496,In_4634,In_4730);
nor U497 (N_497,In_4905,In_367);
nand U498 (N_498,In_4521,In_1521);
nand U499 (N_499,In_1815,In_4386);
and U500 (N_500,In_3939,In_2161);
and U501 (N_501,In_2717,In_216);
and U502 (N_502,In_4684,In_4016);
nor U503 (N_503,In_899,In_4645);
nor U504 (N_504,In_2987,In_1986);
xor U505 (N_505,In_1366,In_3561);
or U506 (N_506,In_646,In_2118);
or U507 (N_507,In_2959,In_3425);
and U508 (N_508,In_1715,In_1318);
xnor U509 (N_509,In_4086,In_2657);
xnor U510 (N_510,In_2964,In_4398);
nand U511 (N_511,In_3856,In_1418);
nand U512 (N_512,In_2641,In_295);
or U513 (N_513,In_4234,In_3476);
xnor U514 (N_514,In_2298,In_2173);
or U515 (N_515,In_3321,In_2283);
nor U516 (N_516,In_2778,In_81);
xnor U517 (N_517,In_1371,In_2532);
or U518 (N_518,In_1710,In_1174);
xnor U519 (N_519,In_4857,In_1129);
nand U520 (N_520,In_3814,In_4296);
or U521 (N_521,In_2838,In_3397);
xnor U522 (N_522,In_3533,In_2452);
xor U523 (N_523,In_4973,In_398);
or U524 (N_524,In_4219,In_3072);
or U525 (N_525,In_3331,In_586);
nor U526 (N_526,In_4515,In_3221);
xor U527 (N_527,In_3523,In_2343);
nor U528 (N_528,In_3937,In_3746);
and U529 (N_529,In_2322,In_3129);
or U530 (N_530,In_4131,In_1909);
xnor U531 (N_531,In_1082,In_4728);
and U532 (N_532,In_4058,In_3706);
nor U533 (N_533,In_551,In_2380);
nor U534 (N_534,In_4554,In_80);
xor U535 (N_535,In_2299,In_3147);
nand U536 (N_536,In_3944,In_875);
nand U537 (N_537,In_1482,In_4224);
or U538 (N_538,In_121,In_2885);
and U539 (N_539,In_2227,In_4958);
nor U540 (N_540,In_3592,In_211);
xnor U541 (N_541,In_4049,In_2293);
nor U542 (N_542,In_3435,In_4701);
and U543 (N_543,In_1617,In_2484);
or U544 (N_544,In_1901,In_2590);
and U545 (N_545,In_3837,In_8);
xor U546 (N_546,In_2475,In_58);
or U547 (N_547,In_3830,In_4077);
nor U548 (N_548,In_1848,In_4926);
and U549 (N_549,In_574,In_3679);
and U550 (N_550,In_675,In_4360);
and U551 (N_551,In_1234,In_4271);
xnor U552 (N_552,In_3289,In_376);
xnor U553 (N_553,In_839,In_1978);
nand U554 (N_554,In_3172,In_887);
xnor U555 (N_555,In_333,In_310);
and U556 (N_556,In_1719,In_3226);
or U557 (N_557,In_2518,In_4527);
and U558 (N_558,In_4117,In_4280);
xnor U559 (N_559,In_567,In_2788);
nand U560 (N_560,In_3056,In_1448);
nor U561 (N_561,In_3993,In_175);
nor U562 (N_562,In_4244,In_999);
or U563 (N_563,In_96,In_402);
nor U564 (N_564,In_1212,In_3341);
nor U565 (N_565,In_4249,In_296);
nand U566 (N_566,In_2614,In_2631);
and U567 (N_567,In_4031,In_4319);
nand U568 (N_568,In_2072,In_59);
nand U569 (N_569,In_60,In_381);
or U570 (N_570,In_1091,In_3826);
or U571 (N_571,In_1613,In_3183);
nand U572 (N_572,In_1832,In_4475);
and U573 (N_573,In_4704,In_4870);
and U574 (N_574,In_1379,In_1061);
and U575 (N_575,In_1417,In_2679);
nor U576 (N_576,In_2190,In_1085);
nor U577 (N_577,In_3440,In_3000);
and U578 (N_578,In_3697,In_4778);
nor U579 (N_579,In_3727,In_3087);
nor U580 (N_580,In_1456,In_238);
nor U581 (N_581,In_4321,In_4052);
or U582 (N_582,In_679,In_461);
and U583 (N_583,In_1713,In_4253);
and U584 (N_584,In_91,In_167);
nor U585 (N_585,In_653,In_1704);
nor U586 (N_586,In_3482,In_277);
xnor U587 (N_587,In_3038,In_99);
xor U588 (N_588,In_4798,In_3468);
xnor U589 (N_589,In_163,In_4085);
nor U590 (N_590,In_579,In_4391);
nand U591 (N_591,In_1729,In_4287);
nor U592 (N_592,In_3591,In_2702);
or U593 (N_593,In_4123,In_2864);
xnor U594 (N_594,In_1413,In_4174);
and U595 (N_595,In_2336,In_4566);
or U596 (N_596,In_1051,In_1532);
xnor U597 (N_597,In_2046,In_4064);
and U598 (N_598,In_723,In_772);
or U599 (N_599,In_1914,In_2310);
and U600 (N_600,In_4025,In_4348);
and U601 (N_601,In_2457,In_3132);
nand U602 (N_602,In_3548,In_3092);
nand U603 (N_603,In_569,In_1312);
or U604 (N_604,In_1759,In_618);
xnor U605 (N_605,In_248,In_4079);
nor U606 (N_606,In_3607,In_3462);
or U607 (N_607,In_1159,In_2958);
nand U608 (N_608,In_549,In_4142);
and U609 (N_609,In_3213,In_3841);
nor U610 (N_610,In_4320,In_3168);
xor U611 (N_611,In_783,In_5);
or U612 (N_612,In_573,In_3873);
nor U613 (N_613,In_3614,In_4087);
nand U614 (N_614,In_855,In_260);
or U615 (N_615,In_3277,In_934);
and U616 (N_616,In_0,In_1957);
nand U617 (N_617,In_2326,In_2655);
xor U618 (N_618,In_1439,In_4264);
nand U619 (N_619,In_1181,In_16);
and U620 (N_620,In_42,In_4649);
nor U621 (N_621,In_4033,In_3300);
nor U622 (N_622,In_4466,In_941);
xor U623 (N_623,In_3479,In_2444);
xor U624 (N_624,In_340,In_1150);
and U625 (N_625,In_2945,In_676);
and U626 (N_626,In_1596,In_2092);
xor U627 (N_627,In_1566,In_3715);
or U628 (N_628,In_705,In_1261);
and U629 (N_629,In_1131,In_1595);
nor U630 (N_630,In_2748,In_2493);
nor U631 (N_631,In_3652,In_4394);
and U632 (N_632,In_2186,In_154);
xor U633 (N_633,In_4775,In_149);
and U634 (N_634,In_455,In_1615);
nand U635 (N_635,In_4697,In_791);
nand U636 (N_636,In_4354,In_26);
or U637 (N_637,In_4107,In_1825);
or U638 (N_638,In_3828,In_1752);
or U639 (N_639,In_3777,In_2253);
xnor U640 (N_640,In_1636,In_1157);
and U641 (N_641,In_1468,In_1108);
nand U642 (N_642,In_3948,In_3555);
and U643 (N_643,In_1431,In_3145);
nor U644 (N_644,In_878,In_1907);
or U645 (N_645,In_256,In_3448);
nand U646 (N_646,In_3024,In_322);
xnor U647 (N_647,In_2623,In_1938);
and U648 (N_648,In_1747,In_286);
nor U649 (N_649,In_2388,In_2757);
nor U650 (N_650,In_19,In_4914);
nor U651 (N_651,In_2943,In_4116);
xnor U652 (N_652,In_1691,In_2576);
xnor U653 (N_653,In_4361,In_2897);
xnor U654 (N_654,In_4614,In_2393);
and U655 (N_655,In_3493,In_4828);
nor U656 (N_656,In_873,In_3540);
and U657 (N_657,In_2447,In_4528);
nor U658 (N_658,In_3878,In_3238);
or U659 (N_659,In_1358,In_1570);
nor U660 (N_660,In_3524,In_4836);
and U661 (N_661,In_2348,In_988);
or U662 (N_662,In_1194,In_4539);
or U663 (N_663,In_3231,In_630);
and U664 (N_664,In_2898,In_4742);
xnor U665 (N_665,In_1965,In_1751);
nor U666 (N_666,In_3492,In_1973);
or U667 (N_667,In_3881,In_2918);
nor U668 (N_668,In_806,In_2662);
and U669 (N_669,In_1013,In_221);
nor U670 (N_670,In_2193,In_3320);
or U671 (N_671,In_1137,In_488);
nand U672 (N_672,In_2375,In_4218);
and U673 (N_673,In_1520,In_864);
nor U674 (N_674,In_210,In_369);
nand U675 (N_675,In_729,In_4136);
and U676 (N_676,In_3556,In_1502);
nand U677 (N_677,In_4620,In_971);
nor U678 (N_678,In_4485,In_2934);
nor U679 (N_679,In_3385,In_1481);
or U680 (N_680,In_3016,In_1296);
nor U681 (N_681,In_3282,In_2917);
xor U682 (N_682,In_842,In_913);
xor U683 (N_683,In_3297,In_3825);
nor U684 (N_684,In_3410,In_2185);
or U685 (N_685,In_1423,In_1231);
nand U686 (N_686,In_4228,In_1666);
or U687 (N_687,In_1628,In_1690);
nand U688 (N_688,In_908,In_4610);
and U689 (N_689,In_4063,In_1223);
xor U690 (N_690,In_234,In_3849);
and U691 (N_691,In_1269,In_1600);
nand U692 (N_692,In_32,In_2752);
nor U693 (N_693,In_2629,In_2957);
xor U694 (N_694,In_979,In_1289);
xor U695 (N_695,In_1026,In_2351);
xor U696 (N_696,In_2863,In_2901);
or U697 (N_697,In_4459,In_4331);
nand U698 (N_698,In_1970,In_2284);
nor U699 (N_699,In_4643,In_1178);
nand U700 (N_700,In_2636,In_2437);
nand U701 (N_701,In_2015,In_2581);
nor U702 (N_702,In_2131,In_385);
nor U703 (N_703,In_3014,In_821);
nor U704 (N_704,In_1720,In_1341);
and U705 (N_705,In_738,In_4604);
nand U706 (N_706,In_1698,In_2514);
nor U707 (N_707,In_2411,In_3649);
and U708 (N_708,In_884,In_4103);
nand U709 (N_709,In_657,In_2597);
and U710 (N_710,In_1818,In_2304);
or U711 (N_711,In_2876,In_4473);
xor U712 (N_712,In_2837,In_2252);
and U713 (N_713,In_3871,In_485);
nor U714 (N_714,In_1142,In_2223);
nand U715 (N_715,In_511,In_722);
and U716 (N_716,In_4333,In_2251);
or U717 (N_717,In_258,In_4494);
nor U718 (N_718,In_139,In_2564);
xnor U719 (N_719,In_3668,In_247);
xor U720 (N_720,In_1622,In_2318);
xor U721 (N_721,In_3230,In_733);
xnor U722 (N_722,In_3973,In_231);
nor U723 (N_723,In_3033,In_848);
nand U724 (N_724,In_390,In_490);
and U725 (N_725,In_658,In_1237);
xor U726 (N_726,In_4167,In_2673);
nor U727 (N_727,In_3577,In_1517);
nor U728 (N_728,In_3411,In_3760);
and U729 (N_729,In_2095,In_917);
xnor U730 (N_730,In_159,In_582);
and U731 (N_731,In_1116,In_2594);
nor U732 (N_732,In_4567,In_2933);
or U733 (N_733,In_1620,In_4977);
nand U734 (N_734,In_4892,In_1601);
or U735 (N_735,In_2919,In_1310);
nand U736 (N_736,In_373,In_1088);
nand U737 (N_737,In_2143,In_487);
nor U738 (N_738,In_1438,In_3724);
or U739 (N_739,In_3491,In_846);
nand U740 (N_740,In_3225,In_3684);
and U741 (N_741,In_2905,In_300);
and U742 (N_742,In_2833,In_868);
xor U743 (N_743,In_198,In_990);
xnor U744 (N_744,In_2855,In_817);
or U745 (N_745,In_1279,In_1317);
or U746 (N_746,In_76,In_4120);
nand U747 (N_747,In_533,In_3804);
xnor U748 (N_748,In_4547,In_1838);
nor U749 (N_749,In_1473,In_2664);
nor U750 (N_750,In_1757,In_306);
and U751 (N_751,In_3490,In_482);
nand U752 (N_752,In_1638,In_4942);
nor U753 (N_753,In_1623,In_3559);
and U754 (N_754,In_2014,In_1442);
and U755 (N_755,In_2768,In_4029);
nor U756 (N_756,In_4210,In_2236);
and U757 (N_757,In_3733,In_4184);
xnor U758 (N_758,In_1643,In_4969);
nor U759 (N_759,In_3274,In_2011);
nand U760 (N_760,In_2174,In_2881);
nor U761 (N_761,In_1044,In_3259);
and U762 (N_762,In_1700,In_939);
nor U763 (N_763,In_1898,In_39);
nor U764 (N_764,In_3193,In_919);
and U765 (N_765,In_4703,In_3840);
or U766 (N_766,In_1568,In_902);
and U767 (N_767,In_3547,In_2779);
nor U768 (N_768,In_502,In_437);
nand U769 (N_769,In_2286,In_2975);
nor U770 (N_770,In_716,In_4767);
nand U771 (N_771,In_3709,In_1395);
nor U772 (N_772,In_1663,In_803);
or U773 (N_773,In_2006,In_3295);
and U774 (N_774,In_831,In_2109);
nand U775 (N_775,In_3266,In_3181);
xor U776 (N_776,In_4523,In_2191);
or U777 (N_777,In_2423,In_4648);
nor U778 (N_778,In_2029,In_1355);
xor U779 (N_779,In_795,In_3081);
or U780 (N_780,In_4158,In_4431);
nor U781 (N_781,In_153,In_4855);
or U782 (N_782,In_460,In_4255);
nor U783 (N_783,In_2281,In_1021);
nor U784 (N_784,In_399,In_2735);
and U785 (N_785,In_3623,In_987);
and U786 (N_786,In_2199,In_3992);
xnor U787 (N_787,In_1465,In_624);
or U788 (N_788,In_4458,In_3418);
nor U789 (N_789,In_53,In_2810);
or U790 (N_790,In_962,In_4900);
nand U791 (N_791,In_521,In_701);
xnor U792 (N_792,In_2397,In_1081);
and U793 (N_793,In_3451,In_3058);
nand U794 (N_794,In_341,In_3537);
and U795 (N_795,In_368,In_3204);
and U796 (N_796,In_1854,In_2262);
nand U797 (N_797,In_4555,In_4414);
nor U798 (N_798,In_3638,In_1510);
or U799 (N_799,In_3738,In_2012);
and U800 (N_800,In_964,In_1183);
xor U801 (N_801,In_1954,In_108);
nor U802 (N_802,In_4434,In_132);
and U803 (N_803,In_3015,In_1368);
nor U804 (N_804,In_581,In_3910);
or U805 (N_805,In_2666,In_4146);
and U806 (N_806,In_517,In_3439);
nand U807 (N_807,In_4600,In_3606);
nand U808 (N_808,In_1220,In_3511);
xor U809 (N_809,In_3626,In_2991);
nand U810 (N_810,In_168,In_4848);
and U811 (N_811,In_4678,In_2907);
nand U812 (N_812,In_1944,In_2231);
xnor U813 (N_813,In_1736,In_2370);
and U814 (N_814,In_315,In_4081);
and U815 (N_815,In_4791,In_4941);
xnor U816 (N_816,In_829,In_323);
xnor U817 (N_817,In_1603,In_4878);
nor U818 (N_818,In_4118,In_3627);
and U819 (N_819,In_2659,In_2835);
nand U820 (N_820,In_2061,In_4430);
nand U821 (N_821,In_4171,In_4712);
and U822 (N_822,In_4923,In_682);
and U823 (N_823,In_1504,In_3258);
nand U824 (N_824,In_4896,In_529);
nor U825 (N_825,In_1933,In_4359);
or U826 (N_826,In_2797,In_2825);
nand U827 (N_827,In_3723,In_404);
and U828 (N_828,In_3543,In_2033);
and U829 (N_829,In_799,In_4746);
nand U830 (N_830,In_3702,In_3549);
xor U831 (N_831,In_2982,In_727);
nand U832 (N_832,In_3030,In_4112);
xnor U833 (N_833,In_4901,In_3243);
nand U834 (N_834,In_267,In_2132);
and U835 (N_835,In_2401,In_4657);
nand U836 (N_836,In_2405,In_1066);
and U837 (N_837,In_4222,In_3722);
or U838 (N_838,In_4563,In_2942);
and U839 (N_839,In_1529,In_3077);
nand U840 (N_840,In_4190,In_178);
nand U841 (N_841,In_2776,In_1295);
nand U842 (N_842,In_3811,In_746);
nor U843 (N_843,In_3322,In_2268);
and U844 (N_844,In_3803,In_619);
nor U845 (N_845,In_3309,In_3217);
nand U846 (N_846,In_933,In_1718);
and U847 (N_847,In_2391,In_4432);
and U848 (N_848,In_1561,In_4124);
nor U849 (N_849,In_2912,In_3516);
nand U850 (N_850,In_2228,In_1007);
nand U851 (N_851,In_2769,In_4763);
or U852 (N_852,In_3960,In_967);
xnor U853 (N_853,In_2366,In_918);
nand U854 (N_854,In_2390,In_3980);
nor U855 (N_855,In_3884,In_2712);
and U856 (N_856,In_4272,In_2824);
xor U857 (N_857,In_1107,In_896);
nand U858 (N_858,In_383,In_4499);
or U859 (N_859,In_2169,In_4628);
or U860 (N_860,In_4788,In_4599);
xor U861 (N_861,In_3552,In_1186);
xnor U862 (N_862,In_4113,In_2034);
and U863 (N_863,In_3758,In_3765);
or U864 (N_864,In_3743,In_4965);
nor U865 (N_865,In_3154,In_1741);
nor U866 (N_866,In_1430,In_1156);
and U867 (N_867,In_1687,In_65);
nor U868 (N_868,In_3766,In_882);
xor U869 (N_869,In_353,In_4028);
or U870 (N_870,In_2467,In_669);
and U871 (N_871,In_2219,In_462);
xnor U872 (N_872,In_2058,In_698);
nor U873 (N_873,In_4820,In_3430);
or U874 (N_874,In_2241,In_4817);
or U875 (N_875,In_2840,In_2653);
and U876 (N_876,In_2022,In_4122);
nor U877 (N_877,In_4050,In_4030);
nand U878 (N_878,In_423,In_4719);
nor U879 (N_879,In_4835,In_4508);
or U880 (N_880,In_204,In_4837);
xnor U881 (N_881,In_2288,In_4976);
and U882 (N_882,In_1806,In_3603);
xor U883 (N_883,In_2347,In_1354);
nand U884 (N_884,In_3965,In_6);
and U885 (N_885,In_1321,In_1075);
or U886 (N_886,In_1052,In_2418);
nor U887 (N_887,In_3793,In_1837);
xnor U888 (N_888,In_3981,In_507);
nor U889 (N_889,In_3662,In_4047);
nor U890 (N_890,In_1921,In_2120);
nand U891 (N_891,In_3602,In_920);
xor U892 (N_892,In_1084,In_2264);
or U893 (N_893,In_2119,In_2294);
and U894 (N_894,In_4789,In_3938);
nor U895 (N_895,In_2485,In_1895);
and U896 (N_896,In_3693,In_768);
and U897 (N_897,In_3820,In_4687);
nand U898 (N_898,In_3701,In_4105);
and U899 (N_899,In_3390,In_3211);
or U900 (N_900,In_3622,In_1014);
or U901 (N_901,In_4776,In_1513);
and U902 (N_902,In_1735,In_4236);
nand U903 (N_903,In_4316,In_4062);
xnor U904 (N_904,In_656,In_4739);
nand U905 (N_905,In_3113,In_505);
nand U906 (N_906,In_3394,In_2170);
nor U907 (N_907,In_1252,In_2166);
nor U908 (N_908,In_4702,In_1330);
or U909 (N_909,In_414,In_1019);
or U910 (N_910,In_625,In_3514);
and U911 (N_911,In_3633,In_4178);
nor U912 (N_912,In_683,In_1707);
and U913 (N_913,In_4275,In_2860);
nor U914 (N_914,In_552,In_453);
or U915 (N_915,In_3095,In_3164);
nand U916 (N_916,In_1873,In_3836);
xor U917 (N_917,In_3656,In_3599);
or U918 (N_918,In_2745,In_3971);
xor U919 (N_919,In_2303,In_845);
and U920 (N_920,In_2935,In_3216);
nor U921 (N_921,In_4990,In_3507);
nand U922 (N_922,In_866,In_4292);
and U923 (N_923,In_2155,In_2266);
xnor U924 (N_924,In_2570,In_3059);
xor U925 (N_925,In_4985,In_4541);
nand U926 (N_926,In_4303,In_1991);
xor U927 (N_927,In_3761,In_2770);
nor U928 (N_928,In_2542,In_4241);
xor U929 (N_929,In_4089,In_782);
or U930 (N_930,In_1397,In_524);
or U931 (N_931,In_284,In_1115);
nor U932 (N_932,In_2402,In_161);
nand U933 (N_933,In_1437,In_708);
nor U934 (N_934,In_4731,In_4295);
or U935 (N_935,In_2338,In_2544);
nand U936 (N_936,In_1268,In_1012);
or U937 (N_937,In_1702,In_1632);
and U938 (N_938,In_1055,In_4526);
xnor U939 (N_939,In_2337,In_1287);
and U940 (N_940,In_3918,In_2952);
nor U941 (N_941,In_1556,In_13);
and U942 (N_942,In_4175,In_580);
and U943 (N_943,In_3127,In_3710);
xnor U944 (N_944,In_2154,In_1928);
nand U945 (N_945,In_4276,In_3025);
xnor U946 (N_946,In_771,In_41);
nor U947 (N_947,In_4654,In_2473);
and U948 (N_948,In_1392,In_3323);
or U949 (N_949,In_4034,In_1352);
or U950 (N_950,In_3845,In_4196);
nand U951 (N_951,In_1071,In_2156);
or U952 (N_952,In_3893,In_301);
nor U953 (N_953,In_584,In_670);
nand U954 (N_954,In_4743,In_3104);
and U955 (N_955,In_2026,In_334);
and U956 (N_956,In_2584,In_730);
nand U957 (N_957,In_500,In_874);
xnor U958 (N_958,In_2149,In_633);
nor U959 (N_959,In_2640,In_3177);
xnor U960 (N_960,In_3959,In_4785);
or U961 (N_961,In_4757,In_4621);
nor U962 (N_962,In_3088,In_2175);
nor U963 (N_963,In_2565,In_4672);
and U964 (N_964,In_1659,In_2150);
nor U965 (N_965,In_1939,In_1114);
or U966 (N_966,In_2660,In_3554);
nand U967 (N_967,In_194,In_2043);
or U968 (N_968,In_1761,In_1271);
or U969 (N_969,In_1618,In_728);
and U970 (N_970,In_2134,In_4369);
and U971 (N_971,In_2846,In_948);
nor U972 (N_972,In_4115,In_4781);
and U973 (N_973,In_4601,In_2462);
nand U974 (N_974,In_2039,In_947);
nand U975 (N_975,In_4338,In_609);
or U976 (N_976,In_832,In_226);
nor U977 (N_977,In_3859,In_3497);
and U978 (N_978,In_86,In_1712);
or U979 (N_979,In_1201,In_3255);
nor U980 (N_980,In_1514,In_4151);
or U981 (N_981,In_3608,In_464);
or U982 (N_982,In_3156,In_4774);
nand U983 (N_983,In_431,In_1558);
nor U984 (N_984,In_4420,In_1206);
and U985 (N_985,In_4185,In_4722);
nand U986 (N_986,In_3359,In_4365);
nand U987 (N_987,In_3963,In_826);
xor U988 (N_988,In_3708,In_1591);
and U989 (N_989,In_18,In_4585);
nand U990 (N_990,In_188,In_4139);
nand U991 (N_991,In_4623,In_3947);
nand U992 (N_992,In_2969,In_4269);
nand U993 (N_993,In_2880,In_2051);
nor U994 (N_994,In_4417,In_223);
or U995 (N_995,In_3442,In_2474);
or U996 (N_996,In_3279,In_4004);
or U997 (N_997,In_3634,In_3500);
nor U998 (N_998,In_3188,In_1644);
nand U999 (N_999,In_1452,In_747);
nand U1000 (N_1000,In_1730,In_459);
nor U1001 (N_1001,In_1239,In_1974);
nand U1002 (N_1002,In_2410,In_1027);
xnor U1003 (N_1003,In_3503,In_426);
xnor U1004 (N_1004,In_3637,In_1994);
nand U1005 (N_1005,In_144,In_4852);
nand U1006 (N_1006,In_877,In_3824);
and U1007 (N_1007,In_610,In_4998);
and U1008 (N_1008,In_4517,In_523);
xnor U1009 (N_1009,In_1040,In_3344);
nor U1010 (N_1010,In_424,In_134);
or U1011 (N_1011,In_3227,In_2030);
nor U1012 (N_1012,In_1475,In_1665);
xor U1013 (N_1013,In_380,In_2984);
nand U1014 (N_1014,In_3117,In_4723);
and U1015 (N_1015,In_4422,In_1935);
and U1016 (N_1016,In_83,In_1017);
nand U1017 (N_1017,In_994,In_2290);
nand U1018 (N_1018,In_3262,In_2168);
and U1019 (N_1019,In_3055,In_2147);
nand U1020 (N_1020,In_3744,In_4607);
xnor U1021 (N_1021,In_4971,In_328);
or U1022 (N_1022,In_3712,In_2661);
nor U1023 (N_1023,In_4368,In_3988);
nor U1024 (N_1024,In_4551,In_3041);
nand U1025 (N_1025,In_1416,In_1454);
and U1026 (N_1026,In_3677,In_514);
and U1027 (N_1027,In_1519,In_4737);
and U1028 (N_1028,In_2282,In_2690);
or U1029 (N_1029,In_3073,In_3986);
xor U1030 (N_1030,In_1727,In_1380);
nor U1031 (N_1031,In_4760,In_3912);
and U1032 (N_1032,In_1184,In_963);
xnor U1033 (N_1033,In_525,In_2260);
nand U1034 (N_1034,In_3094,In_54);
nand U1035 (N_1035,In_3290,In_1210);
or U1036 (N_1036,In_1553,In_2020);
nor U1037 (N_1037,In_4751,In_1096);
nand U1038 (N_1038,In_89,In_3023);
or U1039 (N_1039,In_2040,In_3376);
xnor U1040 (N_1040,In_3889,In_2364);
xor U1041 (N_1041,In_663,In_3337);
or U1042 (N_1042,In_2378,In_3929);
nand U1043 (N_1043,In_2954,In_2604);
or U1044 (N_1044,In_757,In_1754);
xnor U1045 (N_1045,In_3957,In_1399);
and U1046 (N_1046,In_1527,In_2896);
nand U1047 (N_1047,In_2130,In_1215);
xor U1048 (N_1048,In_2470,In_3671);
nand U1049 (N_1049,In_800,In_3542);
nor U1050 (N_1050,In_2041,In_4886);
nand U1051 (N_1051,In_3809,In_2607);
nand U1052 (N_1052,In_4448,In_229);
or U1053 (N_1053,In_506,In_1875);
xor U1054 (N_1054,In_4700,In_2771);
nand U1055 (N_1055,In_718,In_1037);
nor U1056 (N_1056,In_2603,In_3646);
nor U1057 (N_1057,In_1880,In_196);
nor U1058 (N_1058,In_11,In_4690);
and U1059 (N_1059,In_3764,In_4617);
nor U1060 (N_1060,In_1946,In_1867);
or U1061 (N_1061,In_4301,In_1924);
xnor U1062 (N_1062,In_959,In_94);
xnor U1063 (N_1063,In_3648,In_84);
xor U1064 (N_1064,In_3682,In_3750);
xnor U1065 (N_1065,In_2320,In_70);
nand U1066 (N_1066,In_4484,In_3103);
and U1067 (N_1067,In_115,In_3333);
or U1068 (N_1068,In_1440,In_2862);
or U1069 (N_1069,In_3431,In_3311);
nor U1070 (N_1070,In_4741,In_1070);
or U1071 (N_1071,In_546,In_1683);
or U1072 (N_1072,In_21,In_2525);
and U1073 (N_1073,In_1676,In_1634);
nor U1074 (N_1074,In_3997,In_4582);
xor U1075 (N_1075,In_4752,In_2983);
or U1076 (N_1076,In_3572,In_3629);
nor U1077 (N_1077,In_1121,In_4377);
nand U1078 (N_1078,In_2407,In_3484);
or U1079 (N_1079,In_4194,In_1780);
nor U1080 (N_1080,In_2946,In_809);
or U1081 (N_1081,In_1122,In_1947);
nor U1082 (N_1082,In_1948,In_1608);
and U1083 (N_1083,In_1585,In_3184);
and U1084 (N_1084,In_2359,In_4808);
xor U1085 (N_1085,In_4830,In_1124);
nand U1086 (N_1086,In_1776,In_3931);
and U1087 (N_1087,In_1474,In_345);
or U1088 (N_1088,In_4472,In_541);
xor U1089 (N_1089,In_2024,In_4177);
nand U1090 (N_1090,In_1078,In_4347);
nand U1091 (N_1091,In_3427,In_4390);
or U1092 (N_1092,In_1005,In_1447);
nand U1093 (N_1093,In_4683,In_1033);
nand U1094 (N_1094,In_4362,In_1817);
and U1095 (N_1095,In_1202,In_3261);
nand U1096 (N_1096,In_3128,In_3449);
and U1097 (N_1097,In_1927,In_1424);
nand U1098 (N_1098,In_23,In_2048);
and U1099 (N_1099,In_4520,In_4925);
nor U1100 (N_1100,In_4285,In_2172);
xor U1101 (N_1101,In_82,In_1262);
and U1102 (N_1102,In_2124,In_2101);
nor U1103 (N_1103,In_449,In_927);
nor U1104 (N_1104,In_3409,In_3987);
xor U1105 (N_1105,In_4658,In_4593);
nor U1106 (N_1106,In_2385,In_611);
nand U1107 (N_1107,In_4833,In_4795);
and U1108 (N_1108,In_4883,In_1619);
nand U1109 (N_1109,In_4633,In_396);
xor U1110 (N_1110,In_2188,In_1624);
xnor U1111 (N_1111,In_2710,In_3134);
or U1112 (N_1112,In_3019,In_4176);
and U1113 (N_1113,In_225,In_1495);
xor U1114 (N_1114,In_2540,In_4581);
nand U1115 (N_1115,In_3531,In_793);
nand U1116 (N_1116,In_2996,In_2358);
or U1117 (N_1117,In_4121,In_4540);
nand U1118 (N_1118,In_1923,In_1046);
nand U1119 (N_1119,In_4930,In_477);
nor U1120 (N_1120,In_397,In_4858);
or U1121 (N_1121,In_1917,In_2708);
nand U1122 (N_1122,In_930,In_4068);
xnor U1123 (N_1123,In_3327,In_503);
nand U1124 (N_1124,In_1823,In_2413);
xor U1125 (N_1125,In_4322,In_3371);
and U1126 (N_1126,In_29,In_3866);
or U1127 (N_1127,In_3374,In_672);
xor U1128 (N_1128,In_3570,In_418);
or U1129 (N_1129,In_1363,In_982);
or U1130 (N_1130,In_179,In_1900);
nor U1131 (N_1131,In_2371,In_2254);
or U1132 (N_1132,In_1373,In_3135);
nor U1133 (N_1133,In_1889,In_1311);
nand U1134 (N_1134,In_2968,In_3370);
nor U1135 (N_1135,In_1457,In_2007);
or U1136 (N_1136,In_1187,In_3842);
or U1137 (N_1137,In_2561,In_123);
nor U1138 (N_1138,In_1886,In_4909);
xnor U1139 (N_1139,In_4096,In_1992);
xnor U1140 (N_1140,In_870,In_2017);
or U1141 (N_1141,In_1686,In_3653);
xnor U1142 (N_1142,In_3641,In_4382);
nand U1143 (N_1143,In_1925,In_103);
and U1144 (N_1144,In_409,In_1189);
or U1145 (N_1145,In_3280,In_1740);
nor U1146 (N_1146,In_2915,In_4065);
xor U1147 (N_1147,In_2568,In_4946);
xor U1148 (N_1148,In_422,In_3486);
or U1149 (N_1149,In_2669,In_236);
or U1150 (N_1150,In_3250,In_4374);
xor U1151 (N_1151,In_2821,In_3082);
nor U1152 (N_1152,In_4082,In_3166);
nor U1153 (N_1153,In_4924,In_1945);
nor U1154 (N_1154,In_4265,In_4823);
nand U1155 (N_1155,In_2543,In_2215);
xnor U1156 (N_1156,In_4199,In_3704);
nor U1157 (N_1157,In_3283,In_1095);
and U1158 (N_1158,In_4298,In_3882);
or U1159 (N_1159,In_4574,In_654);
nor U1160 (N_1160,In_2222,In_2894);
xnor U1161 (N_1161,In_1708,In_1565);
nand U1162 (N_1162,In_628,In_2010);
xor U1163 (N_1163,In_3833,In_411);
nand U1164 (N_1164,In_230,In_849);
and U1165 (N_1165,In_2598,In_3244);
xor U1166 (N_1166,In_4282,In_4470);
xnor U1167 (N_1167,In_4410,In_3433);
xor U1168 (N_1168,In_4546,In_2479);
nand U1169 (N_1169,In_3084,In_1406);
nor U1170 (N_1170,In_1388,In_2758);
and U1171 (N_1171,In_2780,In_4159);
and U1172 (N_1172,In_1545,In_1733);
nand U1173 (N_1173,In_3405,In_655);
nor U1174 (N_1174,In_965,In_4427);
nand U1175 (N_1175,In_4844,In_4498);
nor U1176 (N_1176,In_2422,In_3475);
and U1177 (N_1177,In_3066,In_1910);
and U1178 (N_1178,In_3900,In_1166);
xor U1179 (N_1179,In_3398,In_797);
or U1180 (N_1180,In_1293,In_4580);
nor U1181 (N_1181,In_1627,In_4327);
nand U1182 (N_1182,In_2853,In_2605);
or U1183 (N_1183,In_3020,In_550);
or U1184 (N_1184,In_4279,In_3286);
and U1185 (N_1185,In_1499,In_4357);
or U1186 (N_1186,In_2151,In_1453);
xnor U1187 (N_1187,In_3532,In_4532);
nor U1188 (N_1188,In_789,In_1802);
and U1189 (N_1189,In_3316,In_4182);
nor U1190 (N_1190,In_4132,In_4804);
xnor U1191 (N_1191,In_1781,In_4453);
nor U1192 (N_1192,In_2107,In_3798);
or U1193 (N_1193,In_1350,In_2733);
nand U1194 (N_1194,In_3661,In_360);
or U1195 (N_1195,In_1796,In_4589);
nor U1196 (N_1196,In_64,In_2430);
nand U1197 (N_1197,In_2993,In_1238);
xnor U1198 (N_1198,In_859,In_1966);
and U1199 (N_1199,In_3610,In_602);
nor U1200 (N_1200,In_4441,In_4286);
nand U1201 (N_1201,In_1805,In_1351);
nor U1202 (N_1202,In_4765,In_1204);
or U1203 (N_1203,In_4595,In_2795);
nor U1204 (N_1204,In_2729,In_3412);
xor U1205 (N_1205,In_4913,In_754);
or U1206 (N_1206,In_1260,In_1874);
nand U1207 (N_1207,In_2044,In_1934);
nor U1208 (N_1208,In_2962,In_861);
and U1209 (N_1209,In_51,In_4987);
and U1210 (N_1210,In_2053,In_320);
xnor U1211 (N_1211,In_3921,In_4212);
nand U1212 (N_1212,In_1536,In_1240);
or U1213 (N_1213,In_2696,In_1789);
xor U1214 (N_1214,In_1094,In_4609);
nor U1215 (N_1215,In_405,In_1090);
and U1216 (N_1216,In_3994,In_4376);
or U1217 (N_1217,In_1218,In_4810);
nand U1218 (N_1218,In_4093,In_4972);
xor U1219 (N_1219,In_2509,In_3251);
or U1220 (N_1220,In_2865,In_2557);
xor U1221 (N_1221,In_3911,In_1200);
xnor U1222 (N_1222,In_3247,In_1277);
nor U1223 (N_1223,In_3525,In_3294);
nand U1224 (N_1224,In_4570,In_792);
nor U1225 (N_1225,In_2709,In_496);
nand U1226 (N_1226,In_612,In_1668);
or U1227 (N_1227,In_3903,In_3998);
and U1228 (N_1228,In_1881,In_3558);
and U1229 (N_1229,In_1170,In_3163);
and U1230 (N_1230,In_1836,In_1301);
or U1231 (N_1231,In_298,In_4091);
xnor U1232 (N_1232,In_925,In_2688);
and U1233 (N_1233,In_4471,In_2140);
nor U1234 (N_1234,In_3119,In_1569);
xor U1235 (N_1235,In_4404,In_4026);
nor U1236 (N_1236,In_2756,In_36);
or U1237 (N_1237,In_1272,In_2740);
nor U1238 (N_1238,In_4740,In_2560);
or U1239 (N_1239,In_1325,In_4738);
nor U1240 (N_1240,In_1819,In_4734);
nand U1241 (N_1241,In_926,In_1584);
and U1242 (N_1242,In_309,In_931);
xor U1243 (N_1243,In_575,In_4525);
and U1244 (N_1244,In_371,In_2084);
nor U1245 (N_1245,In_2777,In_4483);
nand U1246 (N_1246,In_2812,In_4661);
or U1247 (N_1247,In_4974,In_3378);
or U1248 (N_1248,In_3062,In_2240);
xor U1249 (N_1249,In_3273,In_160);
nor U1250 (N_1250,In_852,In_2505);
nand U1251 (N_1251,In_1743,In_1888);
and U1252 (N_1252,In_1689,In_2306);
xor U1253 (N_1253,In_2923,In_30);
and U1254 (N_1254,In_1385,In_3401);
or U1255 (N_1255,In_4960,In_804);
xor U1256 (N_1256,In_4556,In_532);
nand U1257 (N_1257,In_2182,In_2027);
nor U1258 (N_1258,In_3749,In_2259);
or U1259 (N_1259,In_2731,In_4535);
xnor U1260 (N_1260,In_2312,In_2513);
nor U1261 (N_1261,In_1563,In_4284);
xor U1262 (N_1262,In_3061,In_361);
xnor U1263 (N_1263,In_615,In_2949);
nand U1264 (N_1264,In_1594,In_433);
or U1265 (N_1265,In_1551,In_3864);
nand U1266 (N_1266,In_3529,In_1419);
nor U1267 (N_1267,In_4699,In_4227);
xor U1268 (N_1268,In_4023,In_2986);
and U1269 (N_1269,In_1988,In_3190);
and U1270 (N_1270,In_4565,In_841);
xor U1271 (N_1271,In_605,In_4270);
or U1272 (N_1272,In_3883,In_2883);
and U1273 (N_1273,In_509,In_2990);
nand U1274 (N_1274,In_3513,In_1606);
and U1275 (N_1275,In_1299,In_4419);
nor U1276 (N_1276,In_1445,In_2367);
nor U1277 (N_1277,In_1031,In_4339);
nor U1278 (N_1278,In_1753,In_2209);
nand U1279 (N_1279,In_1488,In_3360);
xor U1280 (N_1280,In_4764,In_2355);
xor U1281 (N_1281,In_4935,In_2692);
or U1282 (N_1282,In_3270,In_542);
or U1283 (N_1283,In_246,In_1076);
nand U1284 (N_1284,In_3178,In_743);
nor U1285 (N_1285,In_2951,In_1386);
or U1286 (N_1286,In_2045,In_3367);
or U1287 (N_1287,In_2258,In_2301);
xnor U1288 (N_1288,In_4796,In_1967);
and U1289 (N_1289,In_1248,In_4608);
or U1290 (N_1290,In_1334,In_3053);
xor U1291 (N_1291,In_1134,In_1961);
nand U1292 (N_1292,In_3983,In_614);
nor U1293 (N_1293,In_4881,In_1422);
xnor U1294 (N_1294,In_3035,In_3239);
and U1295 (N_1295,In_1629,In_4853);
nor U1296 (N_1296,In_681,In_113);
nand U1297 (N_1297,In_583,In_3039);
nor U1298 (N_1298,In_2309,In_1041);
or U1299 (N_1299,In_1931,In_2500);
or U1300 (N_1300,In_2767,In_1381);
nor U1301 (N_1301,In_395,In_4226);
nor U1302 (N_1302,In_3999,In_3447);
nand U1303 (N_1303,In_1745,In_4800);
nand U1304 (N_1304,In_4871,In_2784);
and U1305 (N_1305,In_2098,In_3850);
xnor U1306 (N_1306,In_4042,In_3389);
or U1307 (N_1307,In_2988,In_1958);
xor U1308 (N_1308,In_3975,In_2924);
and U1309 (N_1309,In_3138,In_4152);
xor U1310 (N_1310,In_911,In_1086);
nor U1311 (N_1311,In_3538,In_2400);
xnor U1312 (N_1312,In_960,In_4577);
nor U1313 (N_1313,In_38,In_1135);
or U1314 (N_1314,In_2713,In_50);
or U1315 (N_1315,In_1721,In_174);
or U1316 (N_1316,In_1068,In_1376);
and U1317 (N_1317,In_4216,In_244);
nand U1318 (N_1318,In_2232,In_4198);
or U1319 (N_1319,In_1427,In_692);
or U1320 (N_1320,In_1405,In_2085);
nand U1321 (N_1321,In_721,In_4467);
and U1322 (N_1322,In_3862,In_4400);
nor U1323 (N_1323,In_4335,In_3452);
and U1324 (N_1324,In_4616,In_4060);
nor U1325 (N_1325,In_1273,In_273);
nor U1326 (N_1326,In_2459,In_2261);
xor U1327 (N_1327,In_4932,In_3769);
or U1328 (N_1328,In_2277,In_3721);
and U1329 (N_1329,In_1508,In_1408);
xnor U1330 (N_1330,In_4841,In_2552);
and U1331 (N_1331,In_3805,In_3519);
nand U1332 (N_1332,In_1464,In_2368);
and U1333 (N_1333,In_3616,In_392);
xnor U1334 (N_1334,In_1552,In_1463);
or U1335 (N_1335,In_1833,In_1709);
xnor U1336 (N_1336,In_956,In_324);
nor U1337 (N_1337,In_4490,In_4358);
or U1338 (N_1338,In_4465,In_2332);
xnor U1339 (N_1339,In_4075,In_671);
xnor U1340 (N_1340,In_4488,In_2535);
or U1341 (N_1341,In_4618,In_992);
and U1342 (N_1342,In_1377,In_4542);
nor U1343 (N_1343,In_1161,In_218);
xor U1344 (N_1344,In_3148,In_1768);
nand U1345 (N_1345,In_3196,In_707);
or U1346 (N_1346,In_2804,In_2208);
nor U1347 (N_1347,In_1191,In_4588);
nor U1348 (N_1348,In_1980,In_486);
and U1349 (N_1349,In_2634,In_4963);
nand U1350 (N_1350,In_263,In_4057);
nor U1351 (N_1351,In_483,In_4711);
or U1352 (N_1352,In_3787,In_3362);
xnor U1353 (N_1353,In_1415,In_2844);
or U1354 (N_1354,In_4514,In_481);
and U1355 (N_1355,In_2431,In_4691);
xnor U1356 (N_1356,In_4070,In_4999);
nor U1357 (N_1357,In_4170,In_318);
nand U1358 (N_1358,In_761,In_749);
xor U1359 (N_1359,In_2899,In_2063);
xor U1360 (N_1360,In_1891,In_7);
nor U1361 (N_1361,In_4141,In_530);
or U1362 (N_1362,In_4647,In_3681);
xor U1363 (N_1363,In_2353,In_1734);
or U1364 (N_1364,In_1099,In_4787);
nor U1365 (N_1365,In_3647,In_2800);
xor U1366 (N_1366,In_3586,In_2465);
and U1367 (N_1367,In_265,In_3315);
and U1368 (N_1368,In_2213,In_4451);
and U1369 (N_1369,In_4538,In_365);
and U1370 (N_1370,In_1375,In_2892);
or U1371 (N_1371,In_4821,In_4035);
and U1372 (N_1372,In_2914,In_1511);
and U1373 (N_1373,In_621,In_3189);
and U1374 (N_1374,In_4659,In_4207);
xor U1375 (N_1375,In_3069,In_1198);
nand U1376 (N_1376,In_3536,In_3182);
nor U1377 (N_1377,In_2159,In_2327);
and U1378 (N_1378,In_4024,In_3812);
nor U1379 (N_1379,In_1573,In_1362);
or U1380 (N_1380,In_294,In_1653);
nor U1381 (N_1381,In_4518,In_1203);
and U1382 (N_1382,In_4302,In_2005);
xor U1383 (N_1383,In_901,In_2858);
and U1384 (N_1384,In_1571,In_1783);
and U1385 (N_1385,In_2519,In_2676);
and U1386 (N_1386,In_4861,In_4912);
nor U1387 (N_1387,In_1998,In_1820);
and U1388 (N_1388,In_2373,In_980);
or U1389 (N_1389,In_4334,In_1004);
xnor U1390 (N_1390,In_3666,In_3651);
or U1391 (N_1391,In_4891,In_4455);
and U1392 (N_1392,In_4927,In_3174);
xnor U1393 (N_1393,In_537,In_856);
or U1394 (N_1394,In_1788,In_1103);
or U1395 (N_1395,In_2032,In_2618);
and U1396 (N_1396,In_2595,In_4979);
and U1397 (N_1397,In_650,In_4415);
nor U1398 (N_1398,In_1435,In_3906);
nor U1399 (N_1399,In_2141,In_2643);
nor U1400 (N_1400,In_1821,In_3404);
or U1401 (N_1401,In_2137,In_192);
nand U1402 (N_1402,In_3950,In_165);
nor U1403 (N_1403,In_2850,In_1849);
or U1404 (N_1404,In_243,In_954);
and U1405 (N_1405,In_1179,In_3932);
nor U1406 (N_1406,In_2970,In_1799);
nor U1407 (N_1407,In_1642,In_1196);
nand U1408 (N_1408,In_4729,In_969);
and U1409 (N_1409,In_1524,In_4308);
nor U1410 (N_1410,In_4750,In_3142);
xor U1411 (N_1411,In_1964,In_2999);
nand U1412 (N_1412,In_266,In_1887);
nand U1413 (N_1413,In_1127,In_4474);
nand U1414 (N_1414,In_3600,In_720);
nand U1415 (N_1415,In_2491,In_2300);
nand U1416 (N_1416,In_3335,In_900);
nor U1417 (N_1417,In_1353,In_1804);
and U1418 (N_1418,In_773,In_2105);
or U1419 (N_1419,In_4462,In_1963);
xor U1420 (N_1420,In_2722,In_3928);
xor U1421 (N_1421,In_3515,In_3795);
and U1422 (N_1422,In_2068,In_2903);
or U1423 (N_1423,In_1913,In_4163);
xnor U1424 (N_1424,In_3345,In_2324);
and U1425 (N_1425,In_440,In_4130);
xor U1426 (N_1426,In_2019,In_3799);
nand U1427 (N_1427,In_4213,In_2386);
nand U1428 (N_1428,In_2512,In_4919);
nor U1429 (N_1429,In_4644,In_1332);
nor U1430 (N_1430,In_2523,In_1726);
xnor U1431 (N_1431,In_1451,In_203);
xor U1432 (N_1432,In_2978,In_2356);
nand U1433 (N_1433,In_1039,In_3199);
or U1434 (N_1434,In_27,In_3887);
and U1435 (N_1435,In_4424,In_2435);
nand U1436 (N_1436,In_3526,In_1516);
nand U1437 (N_1437,In_879,In_3396);
nand U1438 (N_1438,In_3534,In_4173);
nand U1439 (N_1439,In_1285,In_3925);
nor U1440 (N_1440,In_4606,In_1790);
or U1441 (N_1441,In_2652,In_2198);
xnor U1442 (N_1442,In_825,In_1060);
xor U1443 (N_1443,In_2667,In_4879);
nand U1444 (N_1444,In_847,In_3827);
xnor U1445 (N_1445,In_2050,In_3457);
xor U1446 (N_1446,In_1322,In_1567);
nor U1447 (N_1447,In_355,In_170);
nor U1448 (N_1448,In_1426,In_2278);
nor U1449 (N_1449,In_2093,In_4880);
nand U1450 (N_1450,In_3977,In_1471);
nand U1451 (N_1451,In_1635,In_1257);
nor U1452 (N_1452,In_4938,In_3729);
or U1453 (N_1453,In_946,In_2111);
nor U1454 (N_1454,In_1374,In_1950);
nor U1455 (N_1455,In_1125,In_2481);
or U1456 (N_1456,In_953,In_4013);
nand U1457 (N_1457,In_1673,In_1467);
nor U1458 (N_1458,In_736,In_55);
nor U1459 (N_1459,In_3902,In_1879);
nor U1460 (N_1460,In_2363,In_2743);
nand U1461 (N_1461,In_3870,In_2110);
nand U1462 (N_1462,In_3342,In_2217);
or U1463 (N_1463,In_1576,In_280);
xnor U1464 (N_1464,In_4102,In_1722);
nand U1465 (N_1465,In_1956,In_2730);
nor U1466 (N_1466,In_3654,In_2374);
and U1467 (N_1467,In_4492,In_1764);
and U1468 (N_1468,In_3625,In_4533);
or U1469 (N_1469,In_143,In_3272);
and U1470 (N_1470,In_3581,In_1036);
and U1471 (N_1471,In_1797,In_3363);
xnor U1472 (N_1472,In_4343,In_4373);
or U1473 (N_1473,In_3444,In_4745);
and U1474 (N_1474,In_1333,In_3686);
xnor U1475 (N_1475,In_631,In_3908);
or U1476 (N_1476,In_282,In_3753);
nand U1477 (N_1477,In_4352,In_1357);
or U1478 (N_1478,In_2069,In_2801);
or U1479 (N_1479,In_3445,In_2183);
nand U1480 (N_1480,In_3366,In_3460);
xnor U1481 (N_1481,In_4150,In_3197);
xnor U1482 (N_1482,In_3176,In_2297);
and U1483 (N_1483,In_4078,In_3368);
nor U1484 (N_1484,In_1347,In_2715);
or U1485 (N_1485,In_1633,In_1548);
nand U1486 (N_1486,In_1785,In_885);
nand U1487 (N_1487,In_4888,In_126);
or U1488 (N_1488,In_3905,In_1149);
nand U1489 (N_1489,In_2869,In_3382);
nor U1490 (N_1490,In_3006,In_2403);
nor U1491 (N_1491,In_2099,In_4002);
nand U1492 (N_1492,In_4128,In_1141);
nor U1493 (N_1493,In_2554,In_528);
nand U1494 (N_1494,In_4300,In_1827);
nor U1495 (N_1495,In_4727,In_748);
xor U1496 (N_1496,In_3031,In_3615);
and U1497 (N_1497,In_4381,In_4500);
nand U1498 (N_1498,In_1284,In_4268);
xor U1499 (N_1499,In_3786,In_2973);
and U1500 (N_1500,In_3741,In_2953);
nand U1501 (N_1501,In_711,In_406);
or U1502 (N_1502,In_844,In_52);
and U1503 (N_1503,In_689,In_1130);
or U1504 (N_1504,In_2551,In_1359);
or U1505 (N_1505,In_2433,In_4815);
or U1506 (N_1506,In_4510,In_2665);
nor U1507 (N_1507,In_3101,In_1369);
nand U1508 (N_1508,In_1856,In_152);
nand U1509 (N_1509,In_2714,In_31);
xnor U1510 (N_1510,In_1436,In_1180);
nor U1511 (N_1511,In_1058,In_1169);
or U1512 (N_1512,In_4043,In_2421);
nand U1513 (N_1513,In_1959,In_2350);
and U1514 (N_1514,In_1389,In_1767);
nor U1515 (N_1515,In_430,In_2031);
nor U1516 (N_1516,In_1433,In_2075);
and U1517 (N_1517,In_4996,In_3680);
nand U1518 (N_1518,In_61,In_822);
and U1519 (N_1519,In_1286,In_978);
nand U1520 (N_1520,In_4110,In_3896);
or U1521 (N_1521,In_1340,In_1999);
nor U1522 (N_1522,In_3583,In_3955);
nand U1523 (N_1523,In_2610,In_4220);
nor U1524 (N_1524,In_770,In_3265);
nand U1525 (N_1525,In_1093,In_3890);
xor U1526 (N_1526,In_493,In_755);
xor U1527 (N_1527,In_1067,In_2689);
xnor U1528 (N_1528,In_3782,In_2009);
xnor U1529 (N_1529,In_3416,In_401);
or U1530 (N_1530,In_4011,In_347);
or U1531 (N_1531,In_3673,In_3594);
nand U1532 (N_1532,In_2203,In_249);
nor U1533 (N_1533,In_2836,In_2997);
xor U1534 (N_1534,In_4442,In_3487);
or U1535 (N_1535,In_764,In_4356);
xor U1536 (N_1536,In_4164,In_3588);
nand U1537 (N_1537,In_1337,In_2772);
nand U1538 (N_1538,In_2152,In_2704);
or U1539 (N_1539,In_3876,In_279);
or U1540 (N_1540,In_2428,In_2315);
xnor U1541 (N_1541,In_1065,In_903);
and U1542 (N_1542,In_867,In_1022);
or U1543 (N_1543,In_2383,In_4267);
nor U1544 (N_1544,In_538,In_3495);
xor U1545 (N_1545,In_382,In_2891);
nand U1546 (N_1546,In_3892,In_3546);
xor U1547 (N_1547,In_2079,In_2828);
or U1548 (N_1548,In_942,In_3110);
or U1549 (N_1549,In_828,In_1226);
nor U1550 (N_1550,In_3456,In_1045);
nand U1551 (N_1551,In_3823,In_4384);
or U1552 (N_1552,In_2650,In_3454);
xor U1553 (N_1553,In_1839,In_350);
nor U1554 (N_1554,In_3267,In_3813);
nand U1555 (N_1555,In_2089,In_554);
and U1556 (N_1556,In_3967,In_1167);
or U1557 (N_1557,In_1172,In_2582);
and U1558 (N_1558,In_2357,In_3004);
nand U1559 (N_1559,In_4866,In_151);
xnor U1560 (N_1560,In_3201,In_1739);
xor U1561 (N_1561,In_2204,In_688);
nor U1562 (N_1562,In_120,In_1779);
nand U1563 (N_1563,In_1824,In_2354);
xnor U1564 (N_1564,In_3402,In_1011);
nor U1565 (N_1565,In_3120,In_3155);
nor U1566 (N_1566,In_2113,In_4229);
or U1567 (N_1567,In_824,In_3186);
or U1568 (N_1568,In_3969,In_4720);
or U1569 (N_1569,In_1784,In_4680);
and U1570 (N_1570,In_2706,In_2989);
or U1571 (N_1571,In_75,In_4450);
nor U1572 (N_1572,In_1503,In_693);
nor U1573 (N_1573,In_1106,In_4545);
and U1574 (N_1574,In_3232,In_128);
nand U1575 (N_1575,In_1023,In_4782);
and U1576 (N_1576,In_2995,In_1006);
xnor U1577 (N_1577,In_227,In_1985);
xor U1578 (N_1578,In_2212,In_1098);
or U1579 (N_1579,In_2645,In_2477);
or U1580 (N_1580,In_2087,In_3209);
and U1581 (N_1581,In_726,In_3920);
nor U1582 (N_1582,In_3907,In_3922);
or U1583 (N_1583,In_3687,In_4631);
nand U1584 (N_1584,In_4439,In_2060);
nand U1585 (N_1585,In_3028,In_504);
xor U1586 (N_1586,In_4036,In_293);
and U1587 (N_1587,In_239,In_3913);
nor U1588 (N_1588,In_4933,In_4827);
xnor U1589 (N_1589,In_3755,In_4673);
nor U1590 (N_1590,In_2042,In_4418);
xnor U1591 (N_1591,In_2823,In_2317);
nor U1592 (N_1592,In_1772,In_3047);
xor U1593 (N_1593,In_2094,In_3242);
and U1594 (N_1594,In_4639,In_2280);
and U1595 (N_1595,In_1162,In_1232);
or U1596 (N_1596,In_3472,In_2724);
and U1597 (N_1597,In_4232,In_4726);
xnor U1598 (N_1598,In_2210,In_785);
nor U1599 (N_1599,In_1609,In_3550);
xor U1600 (N_1600,In_2091,In_981);
nor U1601 (N_1601,In_472,In_660);
and U1602 (N_1602,In_4008,In_1840);
and U1603 (N_1603,In_1414,In_3246);
nor U1604 (N_1604,In_494,In_3140);
xnor U1605 (N_1605,In_1535,In_3567);
xnor U1606 (N_1606,In_1491,In_3562);
and U1607 (N_1607,In_1530,In_2177);
xor U1608 (N_1608,In_1803,In_3419);
and U1609 (N_1609,In_1221,In_2941);
xor U1610 (N_1610,In_4822,In_2802);
xor U1611 (N_1611,In_1348,In_2586);
or U1612 (N_1612,In_4943,In_3915);
nand U1613 (N_1613,In_104,In_4619);
xnor U1614 (N_1614,In_3288,In_2734);
nand U1615 (N_1615,In_1449,In_2352);
nor U1616 (N_1616,In_1409,In_1478);
nand U1617 (N_1617,In_3083,In_3220);
xnor U1618 (N_1618,In_3027,In_788);
or U1619 (N_1619,In_2508,In_467);
nand U1620 (N_1620,In_2076,In_1254);
xor U1621 (N_1621,In_2591,In_3609);
or U1622 (N_1622,In_2416,In_4877);
or U1623 (N_1623,In_3541,In_3499);
nand U1624 (N_1624,In_1597,In_4200);
and U1625 (N_1625,In_2167,In_3480);
nor U1626 (N_1626,In_4903,In_2308);
or U1627 (N_1627,In_2911,In_2612);
nand U1628 (N_1628,In_1050,In_4317);
nand U1629 (N_1629,In_3865,In_4902);
or U1630 (N_1630,In_3029,In_836);
xnor U1631 (N_1631,In_780,In_4988);
xor U1632 (N_1632,In_4612,In_2534);
xor U1633 (N_1633,In_4147,In_4395);
nand U1634 (N_1634,In_1834,In_4037);
or U1635 (N_1635,In_661,In_2528);
xnor U1636 (N_1636,In_164,In_2588);
nand U1637 (N_1637,In_3312,In_2436);
or U1638 (N_1638,In_4397,In_1338);
xor U1639 (N_1639,In_2404,In_3585);
xnor U1640 (N_1640,In_4364,In_3118);
or U1641 (N_1641,In_1769,In_3784);
nand U1642 (N_1642,In_3406,In_1652);
nand U1643 (N_1643,In_3990,In_2859);
or U1644 (N_1644,In_1360,In_1792);
xnor U1645 (N_1645,In_3924,In_2546);
or U1646 (N_1646,In_3202,In_3198);
xor U1647 (N_1647,In_3218,In_1225);
and U1648 (N_1648,In_1968,In_3313);
nor U1649 (N_1649,In_1577,In_4095);
nor U1650 (N_1650,In_4209,In_976);
xnor U1651 (N_1651,In_515,In_291);
xor U1652 (N_1652,In_592,In_4168);
and U1653 (N_1653,In_3131,In_3810);
nor U1654 (N_1654,In_3791,In_762);
and U1655 (N_1655,In_3453,In_3170);
xnor U1656 (N_1656,In_3160,In_1002);
xnor U1657 (N_1657,In_4005,In_4307);
nor U1658 (N_1658,In_865,In_87);
and U1659 (N_1659,In_1932,In_2139);
and U1660 (N_1660,In_983,In_4262);
xnor U1661 (N_1661,In_1885,In_4389);
nor U1662 (N_1662,In_2344,In_2305);
and U1663 (N_1663,In_2220,In_148);
nand U1664 (N_1664,In_4201,In_4671);
nor U1665 (N_1665,In_1171,In_3909);
xnor U1666 (N_1666,In_3459,In_2930);
nand U1667 (N_1667,In_4479,In_1826);
xor U1668 (N_1668,In_2023,In_1937);
xnor U1669 (N_1669,In_2471,In_522);
xnor U1670 (N_1670,In_3571,In_1787);
nand U1671 (N_1671,In_3946,In_3324);
nand U1672 (N_1672,In_2775,In_1020);
and U1673 (N_1673,In_1372,In_2806);
or U1674 (N_1674,In_191,In_3121);
and U1675 (N_1675,In_4156,In_815);
and U1676 (N_1676,In_4114,In_391);
or U1677 (N_1677,In_4054,In_4887);
and U1678 (N_1678,In_3260,In_2206);
nand U1679 (N_1679,In_3063,In_645);
xnor U1680 (N_1680,In_1650,In_348);
and U1681 (N_1681,In_2765,In_4137);
or U1682 (N_1682,In_3175,In_2349);
and U1683 (N_1683,In_3051,In_4371);
nand U1684 (N_1684,In_742,In_3613);
nand U1685 (N_1685,In_2376,In_2677);
nand U1686 (N_1686,In_2939,In_4378);
or U1687 (N_1687,In_1073,In_2164);
xor U1688 (N_1688,In_2287,In_2783);
xnor U1689 (N_1689,In_1222,In_4819);
nand U1690 (N_1690,In_1731,In_4421);
and U1691 (N_1691,In_1446,In_2670);
nand U1692 (N_1692,In_3539,In_1250);
xor U1693 (N_1693,In_3380,In_904);
nor U1694 (N_1694,In_4646,In_3292);
and U1695 (N_1695,In_3080,In_1507);
and U1696 (N_1696,In_1185,In_3790);
and U1697 (N_1697,In_807,In_4895);
nor U1698 (N_1698,In_4370,In_3303);
nor U1699 (N_1699,In_114,In_2122);
xor U1700 (N_1700,In_4501,In_3379);
nand U1701 (N_1701,In_3759,In_760);
or U1702 (N_1702,In_668,In_15);
nor U1703 (N_1703,In_3,In_1798);
or U1704 (N_1704,In_3582,In_4399);
and U1705 (N_1705,In_2738,In_2574);
nand U1706 (N_1706,In_1209,In_2128);
nand U1707 (N_1707,In_2809,In_4531);
xnor U1708 (N_1708,In_1158,In_756);
and U1709 (N_1709,In_4959,In_3553);
or U1710 (N_1710,In_4921,In_2506);
nor U1711 (N_1711,In_4108,In_2379);
or U1712 (N_1712,In_416,In_4299);
nand U1713 (N_1713,In_1869,In_2163);
xor U1714 (N_1714,In_4486,In_1744);
nand U1715 (N_1715,In_1936,In_577);
xor U1716 (N_1716,In_547,In_1575);
xnor U1717 (N_1717,In_3353,In_3302);
nand U1718 (N_1718,In_4153,In_3463);
nand U1719 (N_1719,In_73,In_4721);
and U1720 (N_1720,In_2218,In_4653);
or U1721 (N_1721,In_1211,In_819);
xor U1722 (N_1722,In_4290,In_4083);
nand U1723 (N_1723,In_3961,In_1749);
nor U1724 (N_1724,In_2482,In_4611);
nand U1725 (N_1725,In_3935,In_3694);
xor U1726 (N_1726,In_704,In_1074);
or U1727 (N_1727,In_1793,In_1119);
or U1728 (N_1728,In_1484,In_1308);
and U1729 (N_1729,In_312,In_3319);
nand U1730 (N_1730,In_3557,In_810);
nor U1731 (N_1731,In_4350,In_363);
xor U1732 (N_1732,In_1192,In_4675);
nand U1733 (N_1733,In_3517,In_1331);
xnor U1734 (N_1734,In_563,In_4433);
and U1735 (N_1735,In_3328,In_4447);
and U1736 (N_1736,In_1878,In_2950);
and U1737 (N_1737,In_4940,In_2792);
nand U1738 (N_1738,In_4040,In_1072);
nand U1739 (N_1739,In_271,In_3951);
nand U1740 (N_1740,In_4469,In_1555);
nand U1741 (N_1741,In_520,In_3672);
nand U1742 (N_1742,In_4457,In_2873);
xnor U1743 (N_1743,In_3489,In_228);
nor U1744 (N_1744,In_1544,In_801);
and U1745 (N_1745,In_4688,In_4385);
or U1746 (N_1746,In_2719,In_4845);
xor U1747 (N_1747,In_441,In_1015);
nor U1748 (N_1748,In_2255,In_622);
nand U1749 (N_1749,In_2886,In_3754);
nand U1750 (N_1750,In_2839,In_837);
xor U1751 (N_1751,In_3875,In_667);
xnor U1752 (N_1752,In_3888,In_1227);
or U1753 (N_1753,In_4885,In_4850);
nor U1754 (N_1754,In_1270,In_998);
or U1755 (N_1755,In_2238,In_2750);
nand U1756 (N_1756,In_936,In_2142);
xor U1757 (N_1757,In_2382,In_3573);
and U1758 (N_1758,In_4868,In_2592);
and U1759 (N_1759,In_2647,In_1132);
or U1760 (N_1760,In_3576,In_2316);
xnor U1761 (N_1761,In_1852,In_2831);
and U1762 (N_1762,In_2815,In_3349);
nand U1763 (N_1763,In_1276,In_544);
xnor U1764 (N_1764,In_1112,In_3049);
and U1765 (N_1765,In_3222,In_943);
nand U1766 (N_1766,In_2932,In_4867);
or U1767 (N_1767,In_4709,In_649);
xor U1768 (N_1768,In_2037,In_2399);
nor U1769 (N_1769,In_4046,In_1770);
or U1770 (N_1770,In_2794,In_3739);
xor U1771 (N_1771,In_478,In_4092);
or U1772 (N_1772,In_4477,In_1699);
and U1773 (N_1773,In_3098,In_2980);
nand U1774 (N_1774,In_2279,In_3631);
or U1775 (N_1775,In_2074,In_281);
xnor U1776 (N_1776,In_155,In_1000);
nor U1777 (N_1777,In_2602,In_448);
nor U1778 (N_1778,In_2856,In_97);
or U1779 (N_1779,In_3067,In_2114);
nor U1780 (N_1780,In_57,In_4513);
nor U1781 (N_1781,In_1460,In_1816);
and U1782 (N_1782,In_4090,In_3125);
nand U1783 (N_1783,In_1309,In_2121);
nor U1784 (N_1784,In_4186,In_3018);
nand U1785 (N_1785,In_1616,In_3940);
xnor U1786 (N_1786,In_2868,In_1701);
nor U1787 (N_1787,In_603,In_4126);
nand U1788 (N_1788,In_4769,In_1120);
or U1789 (N_1789,In_2562,In_4799);
or U1790 (N_1790,In_906,In_3350);
nand U1791 (N_1791,In_4685,In_447);
xnor U1792 (N_1792,In_1083,In_1249);
or U1793 (N_1793,In_2871,In_3455);
and U1794 (N_1794,In_4449,In_1111);
nor U1795 (N_1795,In_3757,In_2675);
and U1796 (N_1796,In_3689,In_4534);
nand U1797 (N_1797,In_125,In_2726);
or U1798 (N_1798,In_2739,In_2369);
nor U1799 (N_1799,In_3742,In_1593);
nor U1800 (N_1800,In_587,In_4989);
xor U1801 (N_1801,In_4367,In_1459);
nor U1802 (N_1802,In_2550,In_3863);
xor U1803 (N_1803,In_4689,In_694);
xor U1804 (N_1804,In_1742,In_1868);
nand U1805 (N_1805,In_1384,In_564);
xnor U1806 (N_1806,In_1378,In_2108);
xor U1807 (N_1807,In_1297,In_4502);
nand U1808 (N_1808,In_2524,In_991);
or U1809 (N_1809,In_863,In_739);
xnor U1810 (N_1810,In_2559,In_209);
and U1811 (N_1811,In_3470,In_1444);
xnor U1812 (N_1812,In_1092,In_3407);
xnor U1813 (N_1813,In_3111,In_2502);
and U1814 (N_1814,In_4283,In_1987);
xnor U1815 (N_1815,In_264,In_250);
nor U1816 (N_1816,In_811,In_647);
xnor U1817 (N_1817,In_4594,In_2867);
and U1818 (N_1818,In_627,In_3136);
or U1819 (N_1819,In_2271,In_3007);
nor U1820 (N_1820,In_2302,In_2848);
or U1821 (N_1821,In_4460,In_4575);
xnor U1822 (N_1822,In_2425,In_1038);
xnor U1823 (N_1823,In_3332,In_4293);
xnor U1824 (N_1824,In_3568,In_1531);
nand U1825 (N_1825,In_278,In_2499);
nand U1826 (N_1826,In_3747,In_4573);
or U1827 (N_1827,In_3819,In_2599);
nand U1828 (N_1828,In_3075,In_370);
nand U1829 (N_1829,In_4277,In_4968);
or U1830 (N_1830,In_950,In_403);
and U1831 (N_1831,In_4790,In_2626);
and U1832 (N_1832,In_62,In_2000);
nor U1833 (N_1833,In_4967,In_4344);
and U1834 (N_1834,In_1897,In_3669);
or U1835 (N_1835,In_1795,In_2157);
and U1836 (N_1836,In_1539,In_838);
or U1837 (N_1837,In_2773,In_4127);
and U1838 (N_1838,In_3949,In_1345);
or U1839 (N_1839,In_303,In_3660);
nor U1840 (N_1840,In_820,In_2820);
xor U1841 (N_1841,In_1810,In_2129);
or U1842 (N_1842,In_3395,In_626);
or U1843 (N_1843,In_2243,In_425);
nand U1844 (N_1844,In_1393,In_4436);
nor U1845 (N_1845,In_1307,In_1304);
xor U1846 (N_1846,In_342,In_2879);
nand U1847 (N_1847,In_3165,In_2798);
nor U1848 (N_1848,In_636,In_2501);
xor U1849 (N_1849,In_3355,In_944);
nor U1850 (N_1850,In_1105,In_4801);
nand U1851 (N_1851,In_9,In_543);
and U1852 (N_1852,In_872,In_4982);
or U1853 (N_1853,In_1079,In_2439);
and U1854 (N_1854,In_4666,In_2409);
xnor U1855 (N_1855,In_1876,In_4682);
or U1856 (N_1856,In_269,In_3010);
or U1857 (N_1857,In_4195,In_3650);
nand U1858 (N_1858,In_3734,In_3281);
and U1859 (N_1859,In_2270,In_2086);
or U1860 (N_1860,In_2913,In_2721);
or U1861 (N_1861,In_3895,In_2819);
xor U1862 (N_1862,In_1228,In_1291);
nor U1863 (N_1863,In_2483,In_3752);
or U1864 (N_1864,In_3271,In_3822);
nor U1865 (N_1865,In_3580,In_1328);
nor U1866 (N_1866,In_1989,In_695);
xnor U1867 (N_1867,In_127,In_744);
nand U1868 (N_1868,In_2088,In_781);
xor U1869 (N_1869,In_4557,In_3933);
xnor U1870 (N_1870,In_3894,In_1235);
or U1871 (N_1871,In_4824,In_1283);
xor U1872 (N_1872,In_2449,In_3699);
and U1873 (N_1873,In_4706,In_3241);
and U1874 (N_1874,In_3498,In_1915);
or U1875 (N_1875,In_1282,In_1583);
nor U1876 (N_1876,In_830,In_710);
nor U1877 (N_1877,In_1680,In_1049);
or U1878 (N_1878,In_4558,In_2003);
nor U1879 (N_1879,In_3953,In_3414);
xor U1880 (N_1880,In_3112,In_173);
nor U1881 (N_1881,In_3364,In_1669);
nor U1882 (N_1882,In_3361,In_1064);
and U1883 (N_1883,In_410,In_3351);
nand U1884 (N_1884,In_4955,In_2922);
nor U1885 (N_1885,In_140,In_3891);
nor U1886 (N_1886,In_613,In_3630);
nand U1887 (N_1887,In_1077,In_1883);
and U1888 (N_1888,In_3728,In_1870);
xnor U1889 (N_1889,In_2671,In_3043);
or U1890 (N_1890,In_276,In_4342);
nand U1891 (N_1891,In_468,In_765);
and U1892 (N_1892,In_4705,In_1190);
and U1893 (N_1893,In_2047,In_814);
nor U1894 (N_1894,In_2620,In_3683);
or U1895 (N_1895,In_177,In_63);
and U1896 (N_1896,In_4166,In_924);
nor U1897 (N_1897,In_737,In_4211);
nor U1898 (N_1898,In_4516,In_1402);
nand U1899 (N_1899,In_344,In_3162);
nor U1900 (N_1900,In_666,In_4856);
xnor U1901 (N_1901,In_4669,In_456);
nor U1902 (N_1902,In_3417,In_4489);
xnor U1903 (N_1903,In_3774,In_1737);
nand U1904 (N_1904,In_4860,In_1916);
and U1905 (N_1905,In_2718,In_1983);
and U1906 (N_1906,In_4759,In_4372);
nand U1907 (N_1907,In_2638,In_808);
or U1908 (N_1908,In_3215,In_673);
nand U1909 (N_1909,In_4406,In_3783);
xor U1910 (N_1910,In_2786,In_1097);
xor U1911 (N_1911,In_1557,In_2827);
or U1912 (N_1912,In_2392,In_2269);
nor U1913 (N_1913,In_4957,In_2082);
xnor U1914 (N_1914,In_4632,In_674);
nor U1915 (N_1915,In_2272,In_2615);
xnor U1916 (N_1916,In_172,In_4003);
nor U1917 (N_1917,In_907,In_3821);
nor U1918 (N_1918,In_2081,In_3846);
xor U1919 (N_1919,In_1703,In_43);
nand U1920 (N_1920,In_3788,In_1684);
and U1921 (N_1921,In_1850,In_3356);
and U1922 (N_1922,In_4553,In_2412);
or U1923 (N_1923,In_2888,In_3248);
and U1924 (N_1924,In_2415,In_1163);
or U1925 (N_1925,In_4843,In_860);
or U1926 (N_1926,In_466,In_4345);
nor U1927 (N_1927,In_4109,In_4983);
nor U1928 (N_1928,In_973,In_1843);
nor U1929 (N_1929,In_858,In_4379);
nand U1930 (N_1930,In_545,In_3785);
xnor U1931 (N_1931,In_2028,In_2762);
nor U1932 (N_1932,In_1872,In_3923);
and U1933 (N_1933,In_1265,In_2639);
nand U1934 (N_1934,In_4724,In_4145);
nor U1935 (N_1935,In_283,In_3978);
and U1936 (N_1936,In_4007,In_2426);
nor U1937 (N_1937,In_1109,In_4106);
and U1938 (N_1938,In_2755,In_3574);
nor U1939 (N_1939,In_2705,In_4203);
and U1940 (N_1940,In_1048,In_327);
nor U1941 (N_1941,In_1688,In_2920);
xnor U1942 (N_1942,In_1951,In_1207);
nand U1943 (N_1943,In_4463,In_374);
xor U1944 (N_1944,In_2008,In_112);
nor U1945 (N_1945,In_319,In_2468);
or U1946 (N_1946,In_474,In_4098);
nor U1947 (N_1947,In_1018,In_3116);
nand U1948 (N_1948,In_2947,In_157);
xnor U1949 (N_1949,In_4592,In_4994);
and U1950 (N_1950,In_3384,In_3071);
xor U1951 (N_1951,In_3278,In_1168);
nand U1952 (N_1952,In_1724,In_105);
nand U1953 (N_1953,In_1251,In_952);
xnor U1954 (N_1954,In_3751,In_473);
nand U1955 (N_1955,In_4716,In_2419);
nand U1956 (N_1956,In_608,In_562);
nand U1957 (N_1957,In_3346,In_4561);
nor U1958 (N_1958,In_3645,In_3123);
xor U1959 (N_1959,In_4044,In_4340);
xnor U1960 (N_1960,In_4889,In_4238);
xnor U1961 (N_1961,In_4829,In_2529);
or U1962 (N_1962,In_3485,In_955);
nand U1963 (N_1963,In_14,In_2001);
nand U1964 (N_1964,In_2965,In_1016);
nor U1965 (N_1965,In_2016,In_2627);
or U1966 (N_1966,In_4019,In_620);
and U1967 (N_1967,In_2013,In_1859);
nand U1968 (N_1968,In_1390,In_1661);
nand U1969 (N_1969,In_2649,In_536);
or U1970 (N_1970,In_2126,In_4847);
or U1971 (N_1971,In_3399,In_10);
and U1972 (N_1972,In_1195,In_997);
and U1973 (N_1973,In_2910,In_3040);
or U1974 (N_1974,In_1001,In_2200);
nand U1975 (N_1975,In_3598,In_129);
xor U1976 (N_1976,In_362,In_1630);
xor U1977 (N_1977,In_4454,In_1728);
xnor U1978 (N_1978,In_3008,In_3296);
or U1979 (N_1979,In_469,In_1771);
and U1980 (N_1980,In_413,In_1421);
and U1981 (N_1981,In_2814,In_386);
and U1982 (N_1982,In_3046,In_2703);
nor U1983 (N_1983,In_1246,In_2656);
or U1984 (N_1984,In_1995,In_3512);
nand U1985 (N_1985,In_4408,In_2004);
nand U1986 (N_1986,In_3428,In_275);
xor U1987 (N_1987,In_1755,In_3659);
nand U1988 (N_1988,In_4304,In_2900);
or U1989 (N_1989,In_4443,In_1670);
nand U1990 (N_1990,In_1908,In_2276);
and U1991 (N_1991,In_2642,In_2112);
nand U1992 (N_1992,In_1671,In_4289);
or U1993 (N_1993,In_4426,In_3013);
nor U1994 (N_1994,In_2985,In_4793);
nand U1995 (N_1995,In_2790,In_1984);
nor U1996 (N_1996,In_880,In_4188);
or U1997 (N_1997,In_4756,In_1658);
nor U1998 (N_1998,In_2624,In_1564);
or U1999 (N_1999,In_2067,In_1274);
xor U2000 (N_2000,N_353,In_3762);
nand U2001 (N_2001,N_336,N_629);
nand U2002 (N_2002,In_1993,N_425);
xnor U2003 (N_2003,In_329,N_860);
and U2004 (N_2004,N_391,In_4794);
or U2005 (N_2005,N_1891,In_4464);
nor U2006 (N_2006,In_3861,In_2127);
and U2007 (N_2007,N_879,N_190);
nor U2008 (N_2008,N_1944,N_750);
nand U2009 (N_2009,In_3429,In_1003);
nor U2010 (N_2010,In_2162,N_1419);
nor U2011 (N_2011,N_568,N_1083);
nand U2012 (N_2012,N_706,N_450);
or U2013 (N_2013,N_1899,N_683);
and U2014 (N_2014,N_1388,N_922);
nor U2015 (N_2015,N_1410,N_1465);
xor U2016 (N_2016,N_1670,N_1371);
or U2017 (N_2017,N_853,N_501);
nand U2018 (N_2018,N_420,N_1653);
or U2019 (N_2019,N_1876,N_1213);
or U2020 (N_2020,N_1523,N_1771);
or U2021 (N_2021,N_671,N_592);
nand U2022 (N_2022,N_614,N_475);
nor U2023 (N_2023,N_153,N_1350);
and U2024 (N_2024,N_221,N_1763);
or U2025 (N_2025,N_998,In_3596);
or U2026 (N_2026,In_1197,In_1292);
nor U2027 (N_2027,In_3161,N_345);
or U2028 (N_2028,N_1813,N_1571);
or U2029 (N_2029,N_115,N_1013);
or U2030 (N_2030,N_318,In_3086);
or U2031 (N_2031,N_847,N_1355);
nor U2032 (N_2032,N_183,In_107);
nand U2033 (N_2033,N_1158,In_4181);
nand U2034 (N_2034,N_536,In_1056);
or U2035 (N_2035,N_1930,In_4587);
or U2036 (N_2036,N_409,N_1703);
or U2037 (N_2037,N_1495,N_308);
and U2038 (N_2038,N_796,N_1940);
xnor U2039 (N_2039,In_3621,N_1259);
nand U2040 (N_2040,N_1545,In_4237);
nand U2041 (N_2041,In_3869,In_2908);
and U2042 (N_2042,N_1391,In_4590);
and U2043 (N_2043,N_322,N_1016);
nor U2044 (N_2044,N_901,In_2059);
nand U2045 (N_2045,In_4160,N_1509);
or U2046 (N_2046,In_4041,In_3854);
and U2047 (N_2047,N_1305,In_415);
nor U2048 (N_2048,N_538,In_3229);
xnor U2049 (N_2049,In_2628,In_3477);
or U2050 (N_2050,In_4768,N_1555);
xor U2051 (N_2051,In_590,In_181);
nor U2052 (N_2052,N_622,N_258);
and U2053 (N_2053,N_703,N_1534);
xor U2054 (N_2054,N_745,N_1423);
nor U2055 (N_2055,N_201,N_333);
nor U2056 (N_2056,N_1962,In_199);
and U2057 (N_2057,In_4138,N_1089);
or U2058 (N_2058,In_2077,N_1774);
and U2059 (N_2059,N_545,N_95);
and U2060 (N_2060,N_1889,In_3308);
or U2061 (N_2061,N_342,N_1945);
nor U2062 (N_2062,In_4315,N_828);
or U2063 (N_2063,In_3502,N_1407);
and U2064 (N_2064,N_1828,In_4258);
or U2065 (N_2065,In_3745,In_3314);
and U2066 (N_2066,N_194,N_1927);
or U2067 (N_2067,N_1119,N_1268);
or U2068 (N_2068,N_598,N_1466);
nand U2069 (N_2069,In_607,In_2937);
nor U2070 (N_2070,N_532,In_3298);
xor U2071 (N_2071,In_432,In_3792);
nand U2072 (N_2072,N_1875,N_707);
and U2073 (N_2073,In_2711,N_1185);
or U2074 (N_2074,N_1149,N_1117);
nand U2075 (N_2075,In_2566,In_2464);
or U2076 (N_2076,N_1124,In_1518);
or U2077 (N_2077,N_539,N_404);
and U2078 (N_2078,In_4325,N_1363);
nor U2079 (N_2079,N_543,N_1404);
nand U2080 (N_2080,In_1278,N_231);
xnor U2081 (N_2081,N_615,N_1972);
and U2082 (N_2082,N_714,In_1327);
nor U2083 (N_2083,In_3612,N_1074);
and U2084 (N_2084,N_804,N_1910);
or U2085 (N_2085,N_136,In_1865);
or U2086 (N_2086,N_429,N_1924);
or U2087 (N_2087,N_1338,N_952);
or U2088 (N_2088,N_1137,N_718);
xor U2089 (N_2089,N_659,N_163);
nand U2090 (N_2090,N_1221,N_11);
nor U2091 (N_2091,In_3089,In_779);
or U2092 (N_2092,N_436,In_4758);
and U2093 (N_2093,In_3714,N_1282);
nand U2094 (N_2094,In_1705,N_760);
nor U2095 (N_2095,N_214,N_1939);
xnor U2096 (N_2096,In_4149,In_518);
nand U2097 (N_2097,N_1236,N_1114);
nand U2098 (N_2098,N_127,N_1848);
and U2099 (N_2099,In_2637,N_579);
nand U2100 (N_2100,N_132,In_3868);
xor U2101 (N_2101,In_897,N_573);
or U2102 (N_2102,N_1691,N_1251);
xor U2103 (N_2103,N_1739,N_1845);
or U2104 (N_2104,N_1665,In_3124);
nand U2105 (N_2105,N_64,N_1269);
or U2106 (N_2106,N_1559,N_1579);
nand U2107 (N_2107,N_56,N_1973);
or U2108 (N_2108,N_42,N_1515);
nand U2109 (N_2109,N_1377,N_477);
and U2110 (N_2110,In_1509,N_516);
nor U2111 (N_2111,N_1053,N_1867);
nand U2112 (N_2112,N_164,N_57);
nand U2113 (N_2113,In_2455,In_4245);
nor U2114 (N_2114,N_1120,In_3284);
and U2115 (N_2115,N_789,In_3391);
xnor U2116 (N_2116,In_4736,N_1617);
nand U2117 (N_2117,N_1796,N_628);
nand U2118 (N_2118,N_1462,In_4613);
or U2119 (N_2119,In_4505,N_1646);
xnor U2120 (N_2120,N_222,N_641);
nand U2121 (N_2121,In_4330,In_916);
and U2122 (N_2122,N_871,N_111);
nor U2123 (N_2123,In_1647,N_1521);
or U2124 (N_2124,N_925,In_387);
xor U2125 (N_2125,N_206,In_4918);
and U2126 (N_2126,N_1065,N_1912);
and U2127 (N_2127,N_443,In_3179);
or U2128 (N_2128,N_470,N_1473);
nor U2129 (N_2129,In_4375,In_593);
and U2130 (N_2130,In_1738,N_1731);
nor U2131 (N_2131,In_3797,N_1205);
or U2132 (N_2132,In_3639,N_1548);
and U2133 (N_2133,N_645,N_77);
xor U2134 (N_2134,In_4250,N_514);
nor U2135 (N_2135,N_1490,N_1309);
and U2136 (N_2136,N_910,N_492);
xor U2137 (N_2137,In_4180,In_1364);
and U2138 (N_2138,N_1109,In_3048);
or U2139 (N_2139,N_229,N_987);
xnor U2140 (N_2140,In_470,N_148);
and U2141 (N_2141,In_3461,N_1822);
nor U2142 (N_2142,N_1264,N_416);
and U2143 (N_2143,N_47,N_1513);
xnor U2144 (N_2144,In_4939,N_1683);
and U2145 (N_2145,In_162,N_1582);
or U2146 (N_2146,In_2826,N_1814);
nor U2147 (N_2147,In_3564,N_1233);
or U2148 (N_2148,N_1488,N_923);
nand U2149 (N_2149,In_2609,N_1202);
xor U2150 (N_2150,N_1428,N_455);
nand U2151 (N_2151,In_4811,In_4931);
nor U2152 (N_2152,In_1809,N_1411);
or U2153 (N_2153,N_1788,N_1306);
nand U2154 (N_2154,N_1865,N_1911);
nand U2155 (N_2155,In_3152,In_745);
nand U2156 (N_2156,N_66,N_7);
xor U2157 (N_2157,N_872,In_1716);
nand U2158 (N_2158,In_305,N_302);
and U2159 (N_2159,N_1971,In_2194);
or U2160 (N_2160,N_881,In_2036);
nand U2161 (N_2161,N_819,N_1589);
xor U2162 (N_2162,N_877,N_432);
nor U2163 (N_2163,In_1319,N_176);
and U2164 (N_2164,N_70,In_2056);
xor U2165 (N_2165,N_1553,In_3740);
nand U2166 (N_2166,N_1575,N_1914);
nand U2167 (N_2167,N_1435,N_794);
nand U2168 (N_2168,N_1935,N_711);
xnor U2169 (N_2169,N_1574,N_239);
nand U2170 (N_2170,N_669,In_4208);
nand U2171 (N_2171,N_1655,N_780);
nor U2172 (N_2172,In_2621,N_1864);
nor U2173 (N_2173,N_521,In_1382);
and U2174 (N_2174,In_1685,N_1007);
xor U2175 (N_2175,N_1386,N_1879);
or U2176 (N_2176,N_8,N_627);
and U2177 (N_2177,N_1200,In_3383);
and U2178 (N_2178,In_136,N_1923);
and U2179 (N_2179,In_4944,N_1805);
nand U2180 (N_2180,N_220,N_387);
xor U2181 (N_2181,N_1764,N_252);
or U2182 (N_2182,N_788,N_1044);
xor U2183 (N_2183,N_1223,In_346);
nor U2184 (N_2184,In_4405,N_966);
or U2185 (N_2185,N_1012,N_1499);
and U2186 (N_2186,In_4695,N_565);
nor U2187 (N_2187,N_1692,In_4297);
nand U2188 (N_2188,In_3381,N_1754);
or U2189 (N_2189,N_1281,N_1232);
nand U2190 (N_2190,N_981,In_3719);
nor U2191 (N_2191,In_4061,N_1084);
nor U2192 (N_2192,In_4006,In_4911);
nand U2193 (N_2193,N_765,N_307);
and U2194 (N_2194,In_311,N_972);
and U2195 (N_2195,In_1469,N_1847);
and U2196 (N_2196,In_2749,In_1177);
nor U2197 (N_2197,In_1589,N_1897);
or U2198 (N_2198,N_1227,N_827);
or U2199 (N_2199,In_4242,N_1031);
or U2200 (N_2200,In_1443,N_482);
xor U2201 (N_2201,N_1174,N_341);
nand U2202 (N_2202,N_1562,N_374);
nand U2203 (N_2203,N_1,In_616);
xnor U2204 (N_2204,N_106,In_4509);
or U2205 (N_2205,In_1247,N_1165);
and U2206 (N_2206,In_1765,In_1857);
and U2207 (N_2207,N_1037,N_1270);
and U2208 (N_2208,N_664,N_1427);
nor U2209 (N_2209,In_2246,In_4423);
nand U2210 (N_2210,N_334,In_3421);
and U2211 (N_2211,N_1284,In_4840);
nor U2212 (N_2212,In_4771,In_691);
nor U2213 (N_2213,N_850,N_559);
nand U2214 (N_2214,In_3106,N_655);
nand U2215 (N_2215,N_1095,In_421);
nand U2216 (N_2216,N_30,N_159);
xor U2217 (N_2217,N_1131,N_735);
nor U2218 (N_2218,In_2365,N_1453);
or U2219 (N_2219,In_1791,N_1140);
and U2220 (N_2220,In_4191,In_1695);
or U2221 (N_2221,N_888,N_26);
or U2222 (N_2222,N_1367,N_1424);
and U2223 (N_2223,N_1105,N_287);
xor U2224 (N_2224,N_911,In_1579);
nand U2225 (N_2225,In_2691,In_4080);
nor U2226 (N_2226,N_1516,N_1396);
and U2227 (N_2227,N_1167,N_701);
nor U2228 (N_2228,N_1999,N_1003);
or U2229 (N_2229,In_436,N_580);
nand U2230 (N_2230,In_1010,N_1654);
xnor U2231 (N_2231,In_262,N_1838);
or U2232 (N_2232,N_1815,N_1981);
xor U2233 (N_2233,N_1792,N_338);
nor U2234 (N_2234,N_1359,N_1021);
nand U2235 (N_2235,N_63,N_616);
nor U2236 (N_2236,In_78,In_3130);
and U2237 (N_2237,N_10,N_314);
xor U2238 (N_2238,N_945,N_192);
nand U2239 (N_2239,N_1573,In_3527);
and U2240 (N_2240,N_566,In_2292);
and U2241 (N_2241,In_1314,N_1491);
or U2242 (N_2242,N_893,In_3146);
or U2243 (N_2243,In_184,N_526);
or U2244 (N_2244,N_1725,In_259);
nand U2245 (N_2245,N_1958,N_688);
nor U2246 (N_2246,In_869,In_4497);
and U2247 (N_2247,N_1368,N_460);
and U2248 (N_2248,In_2334,N_332);
xnor U2249 (N_2249,In_4839,In_3310);
xor U2250 (N_2250,N_984,N_831);
nor U2251 (N_2251,In_1087,N_1379);
nand U2252 (N_2252,N_676,In_4383);
and U2253 (N_2253,N_535,N_976);
and U2254 (N_2254,N_1773,In_1906);
xor U2255 (N_2255,In_680,In_2052);
and U2256 (N_2256,N_1769,In_712);
xnor U2257 (N_2257,In_3829,N_1479);
xnor U2258 (N_2258,In_510,In_1660);
and U2259 (N_2259,N_1634,N_1014);
and U2260 (N_2260,N_719,In_1649);
or U2261 (N_2261,In_3857,N_34);
nand U2262 (N_2262,In_3325,In_2635);
or U2263 (N_2263,In_4964,N_863);
xnor U2264 (N_2264,In_4223,N_1965);
nor U2265 (N_2265,N_1730,In_958);
or U2266 (N_2266,N_6,In_124);
nor U2267 (N_2267,N_509,N_1470);
nand U2268 (N_2268,N_1237,In_2791);
xor U2269 (N_2269,N_1000,In_1714);
and U2270 (N_2270,N_433,N_1934);
nand U2271 (N_2271,In_914,N_609);
nor U2272 (N_2272,N_962,N_130);
xnor U2273 (N_2273,N_253,In_2981);
xor U2274 (N_2274,N_424,In_588);
and U2275 (N_2275,N_1403,In_539);
or U2276 (N_2276,N_67,N_694);
or U2277 (N_2277,N_1426,In_3471);
and U2278 (N_2278,N_563,In_1922);
nor U2279 (N_2279,N_1255,N_1782);
or U2280 (N_2280,N_1810,In_1515);
xor U2281 (N_2281,N_1833,N_232);
or U2282 (N_2282,N_360,N_1842);
and U2283 (N_2283,In_4247,N_1153);
and U2284 (N_2284,N_200,N_895);
and U2285 (N_2285,N_1330,N_493);
or U2286 (N_2286,N_1852,N_961);
nor U2287 (N_2287,N_84,N_1229);
nand U2288 (N_2288,N_1599,N_663);
nand U2289 (N_2289,N_1493,N_403);
or U2290 (N_2290,N_1178,In_3956);
nor U2291 (N_2291,N_1855,N_857);
or U2292 (N_2292,N_1787,In_4021);
nand U2293 (N_2293,N_657,N_205);
or U2294 (N_2294,N_454,N_1262);
or U2295 (N_2295,N_574,In_2887);
xor U2296 (N_2296,N_273,N_1890);
or U2297 (N_2297,N_523,N_241);
or U2298 (N_2298,N_330,N_752);
or U2299 (N_2299,In_894,N_1314);
or U2300 (N_2300,N_1551,In_2456);
nand U2301 (N_2301,In_4187,N_916);
nand U2302 (N_2302,N_269,In_1199);
xor U2303 (N_2303,In_4217,N_430);
or U2304 (N_2304,N_1866,N_806);
nor U2305 (N_2305,N_558,In_1758);
nand U2306 (N_2306,N_1334,In_2469);
and U2307 (N_2307,In_4337,In_3640);
xor U2308 (N_2308,N_1613,In_1479);
or U2309 (N_2309,N_354,In_3590);
xor U2310 (N_2310,N_388,N_1895);
xnor U2311 (N_2311,In_1903,N_1706);
xor U2312 (N_2312,N_704,In_993);
or U2313 (N_2313,N_1331,In_1441);
and U2314 (N_2314,N_684,In_3400);
nor U2315 (N_2315,N_1452,N_186);
xor U2316 (N_2316,N_255,N_1840);
nand U2317 (N_2317,N_68,N_1008);
nand U2318 (N_2318,In_734,N_1871);
nand U2319 (N_2319,N_917,N_1100);
and U2320 (N_2320,N_298,N_634);
or U2321 (N_2321,In_3097,In_1542);
nor U2322 (N_2322,N_94,In_4802);
xnor U2323 (N_2323,In_1899,In_3914);
xor U2324 (N_2324,In_1428,N_135);
or U2325 (N_2325,In_1151,In_3438);
nand U2326 (N_2326,N_1627,N_165);
nor U2327 (N_2327,N_208,N_1561);
or U2328 (N_2328,N_774,In_4318);
and U2329 (N_2329,In_4579,In_3737);
nand U2330 (N_2330,In_909,In_1693);
nor U2331 (N_2331,In_1458,In_4692);
nor U2332 (N_2332,N_1402,N_744);
or U2333 (N_2333,N_767,N_1795);
nor U2334 (N_2334,N_1418,N_502);
xor U2335 (N_2335,N_1444,N_1503);
or U2336 (N_2336,N_818,In_427);
nand U2337 (N_2337,N_264,In_2684);
nor U2338 (N_2338,N_1618,N_71);
nor U2339 (N_2339,N_1621,N_1721);
nor U2340 (N_2340,In_3691,N_55);
xor U2341 (N_2341,In_2071,N_891);
nor U2342 (N_2342,In_634,In_290);
nor U2343 (N_2343,In_1896,In_2654);
xor U2344 (N_2344,N_1430,N_1337);
nor U2345 (N_2345,In_2448,N_227);
or U2346 (N_2346,In_1280,N_555);
or U2347 (N_2347,In_1144,In_1243);
and U2348 (N_2348,N_1738,In_1133);
and U2349 (N_2349,In_4045,N_300);
nand U2350 (N_2350,N_447,N_81);
nor U2351 (N_2351,N_824,N_1888);
or U2352 (N_2352,N_365,In_753);
nand U2353 (N_2353,N_1915,In_4715);
xnor U2354 (N_2354,N_1819,In_4101);
or U2355 (N_2355,N_400,In_3605);
or U2356 (N_2356,In_3501,N_1032);
or U2357 (N_2357,N_38,N_621);
and U2358 (N_2358,In_439,N_129);
xor U2359 (N_2359,N_665,N_53);
xor U2360 (N_2360,N_1041,N_1790);
nor U2361 (N_2361,N_5,N_1317);
and U2362 (N_2362,N_1979,N_949);
nor U2363 (N_2363,N_904,N_121);
or U2364 (N_2364,N_1702,N_1145);
nor U2365 (N_2365,N_444,N_995);
and U2366 (N_2366,N_597,N_1989);
xnor U2367 (N_2367,N_412,N_1241);
nand U2368 (N_2368,N_9,In_4638);
nand U2369 (N_2369,In_349,N_1917);
nand U2370 (N_2370,N_1287,In_3057);
nor U2371 (N_2371,In_548,N_936);
and U2372 (N_2372,In_2545,N_723);
or U2373 (N_2373,N_1583,N_1794);
or U2374 (N_2374,In_4571,N_1936);
nor U2375 (N_2375,N_803,N_1841);
xnor U2376 (N_2376,N_1751,In_4243);
or U2377 (N_2377,N_1986,In_4134);
and U2378 (N_2378,N_78,In_1253);
nand U2379 (N_2379,N_285,N_414);
xnor U2380 (N_2380,In_3904,N_670);
nor U2381 (N_2381,N_690,In_910);
nand U2382 (N_2382,N_1786,N_797);
xor U2383 (N_2383,N_739,In_1062);
and U2384 (N_2384,In_1723,N_1296);
or U2385 (N_2385,N_1849,N_1946);
nand U2386 (N_2386,N_491,N_1686);
and U2387 (N_2387,N_1957,In_989);
xnor U2388 (N_2388,N_1481,N_1762);
nand U2389 (N_2389,In_3336,In_3307);
or U2390 (N_2390,N_1492,N_1189);
and U2391 (N_2391,In_4549,N_982);
nand U2392 (N_2392,In_3022,In_3851);
nand U2393 (N_2393,N_356,N_779);
nand U2394 (N_2394,In_366,In_812);
or U2395 (N_2395,N_1015,N_1460);
or U2396 (N_2396,N_1443,N_1125);
nand U2397 (N_2397,N_1791,N_1349);
xnor U2398 (N_2398,N_699,N_364);
or U2399 (N_2399,N_866,In_4875);
xor U2400 (N_2400,N_954,In_4155);
or U2401 (N_2401,N_1705,N_1345);
nor U2402 (N_2402,In_2921,N_1950);
and U2403 (N_2403,In_106,In_2843);
xor U2404 (N_2404,N_340,N_1887);
nand U2405 (N_2405,In_270,N_459);
xor U2406 (N_2406,N_1238,In_3962);
nor U2407 (N_2407,In_4503,N_1184);
xnor U2408 (N_2408,In_1882,N_715);
nor U2409 (N_2409,N_1722,N_1123);
xor U2410 (N_2410,In_3898,N_503);
nand U2411 (N_2411,In_3982,In_1574);
nor U2412 (N_2412,N_1687,In_4710);
or U2413 (N_2413,N_654,N_604);
xor U2414 (N_2414,In_1864,In_3927);
nand U2415 (N_2415,In_3732,N_61);
nor U2416 (N_2416,N_1129,N_997);
and U2417 (N_2417,N_845,N_14);
or U2418 (N_2418,N_73,N_920);
nor U2419 (N_2419,In_1953,N_329);
nand U2420 (N_2420,N_1802,N_237);
xnor U2421 (N_2421,In_2596,In_3776);
nor U2422 (N_2422,N_487,N_1056);
xor U2423 (N_2423,N_41,In_1746);
nor U2424 (N_2424,N_1464,N_197);
or U2425 (N_2425,In_3233,N_1803);
nand U2426 (N_2426,N_1156,N_107);
nand U2427 (N_2427,N_326,N_887);
or U2428 (N_2428,N_286,N_1461);
nand U2429 (N_2429,N_1995,N_1707);
or U2430 (N_2430,In_1533,In_1725);
and U2431 (N_2431,N_1079,N_396);
nand U2432 (N_2432,N_1169,N_147);
nand U2433 (N_2433,N_80,N_1072);
and U2434 (N_2434,N_561,In_3703);
and U2435 (N_2435,N_110,N_631);
and U2436 (N_2436,N_986,N_607);
nand U2437 (N_2437,In_2616,N_1421);
xor U2438 (N_2438,In_2579,In_2974);
or U2439 (N_2439,In_1008,In_4652);
xnor U2440 (N_2440,N_1242,N_829);
xnor U2441 (N_2441,N_1508,N_1004);
nor U2442 (N_2442,N_964,N_1442);
nand U2443 (N_2443,In_1976,N_17);
xor U2444 (N_2444,N_584,N_1533);
xor U2445 (N_2445,In_921,N_1514);
or U2446 (N_2446,N_422,N_303);
and U2447 (N_2447,N_1226,N_24);
xor U2448 (N_2448,N_272,In_4055);
and U2449 (N_2449,N_1299,N_1148);
and U2450 (N_2450,N_1907,N_1173);
xor U2451 (N_2451,In_638,In_297);
or U2452 (N_2452,N_281,In_4481);
nor U2453 (N_2453,In_3144,N_295);
xnor U2454 (N_2454,In_3352,In_3305);
or U2455 (N_2455,In_252,In_1621);
nand U2456 (N_2456,N_288,N_452);
and U2457 (N_2457,N_716,N_1637);
and U2458 (N_2458,In_4625,N_524);
and U2459 (N_2459,In_678,N_85);
nor U2460 (N_2460,In_3952,N_1001);
and U2461 (N_2461,N_594,N_1035);
or U2462 (N_2462,N_463,N_1458);
and U2463 (N_2463,N_697,N_823);
xor U2464 (N_2464,N_661,N_1478);
nand U2465 (N_2465,N_417,In_2619);
or U2466 (N_2466,N_1603,N_1285);
nand U2467 (N_2467,N_1456,In_1672);
or U2468 (N_2468,N_835,N_930);
nand U2469 (N_2469,N_1554,N_116);
nor U2470 (N_2470,N_1526,In_1667);
xor U2471 (N_2471,N_1565,N_1179);
xnor U2472 (N_2472,N_1812,N_126);
and U2473 (N_2473,N_1087,N_906);
or U2474 (N_2474,N_1057,N_1220);
nand U2475 (N_2475,In_640,In_2148);
or U2476 (N_2476,N_79,N_468);
nor U2477 (N_2477,In_304,In_1233);
nor U2478 (N_2478,N_742,N_1199);
xor U2479 (N_2479,N_1075,N_1183);
and U2480 (N_2480,N_440,N_1502);
and U2481 (N_2481,In_4263,N_1715);
nor U2482 (N_2482,In_664,In_643);
and U2483 (N_2483,In_12,N_786);
and U2484 (N_2484,N_1365,In_2055);
nand U2485 (N_2485,N_709,N_1506);
and U2486 (N_2486,N_23,N_1454);
nand U2487 (N_2487,In_3102,N_48);
and U2488 (N_2488,N_884,N_1801);
nor U2489 (N_2489,In_2994,In_1811);
nand U2490 (N_2490,In_2106,N_1085);
xnor U2491 (N_2491,In_3885,In_1344);
nor U2492 (N_2492,N_1869,N_851);
nand U2493 (N_2493,N_182,In_3205);
and U2494 (N_2494,In_3530,N_88);
and U2495 (N_2495,In_4732,N_951);
and U2496 (N_2496,N_1279,N_1716);
nand U2497 (N_2497,N_1984,In_4826);
nor U2498 (N_2498,N_1542,N_91);
xnor U2499 (N_2499,N_572,N_383);
nor U2500 (N_2500,N_1530,In_2537);
xor U2501 (N_2501,N_1441,N_1532);
and U2502 (N_2502,N_638,N_1918);
xor U2503 (N_2503,N_1856,N_875);
or U2504 (N_2504,N_462,N_98);
and U2505 (N_2505,In_394,In_4543);
xor U2506 (N_2506,In_130,In_465);
xnor U2507 (N_2507,N_1050,N_1382);
xnor U2508 (N_2508,N_682,N_1612);
xnor U2509 (N_2509,N_637,In_915);
nand U2510 (N_2510,In_4380,In_945);
and U2511 (N_2511,N_1664,N_1295);
nor U2512 (N_2512,In_3620,N_1952);
xor U2513 (N_2513,N_247,N_114);
or U2514 (N_2514,In_4733,N_211);
nand U2515 (N_2515,N_321,N_1422);
nor U2516 (N_2516,N_1324,In_4917);
and U2517 (N_2517,N_497,N_1699);
or U2518 (N_2518,In_400,N_1289);
and U2519 (N_2519,In_3509,N_1688);
nor U2520 (N_2520,N_1425,N_155);
nand U2521 (N_2521,N_927,N_761);
or U2522 (N_2522,In_4992,N_1298);
xnor U2523 (N_2523,In_3789,N_1440);
or U2524 (N_2524,In_3716,N_1552);
or U2525 (N_2525,N_1340,N_974);
or U2526 (N_2526,N_395,In_594);
or U2527 (N_2527,N_978,In_2558);
nor U2528 (N_2528,N_152,N_1009);
nand U2529 (N_2529,N_1431,In_2782);
nand U2530 (N_2530,In_1483,N_219);
xor U2531 (N_2531,N_710,In_4873);
or U2532 (N_2532,In_2237,N_1101);
nand U2533 (N_2533,N_510,In_3365);
and U2534 (N_2534,N_1619,In_651);
or U2535 (N_2535,N_1415,N_1128);
xor U2536 (N_2536,N_800,N_1230);
nand U2537 (N_2537,N_1384,N_1712);
xor U2538 (N_2538,N_1861,N_1868);
xnor U2539 (N_2539,N_245,N_1040);
nand U2540 (N_2540,N_202,N_442);
or U2541 (N_2541,N_1528,N_118);
or U2542 (N_2542,In_1425,N_1970);
xor U2543 (N_2543,N_900,N_1445);
xnor U2544 (N_2544,N_859,N_569);
or U2545 (N_2545,N_1327,In_3916);
and U2546 (N_2546,N_1273,N_305);
or U2547 (N_2547,N_1217,N_35);
or U2548 (N_2548,N_428,N_613);
or U2549 (N_2549,In_889,In_1996);
or U2550 (N_2550,In_4014,N_1272);
nand U2551 (N_2551,In_4438,In_2102);
nor U2552 (N_2552,In_4522,N_963);
nand U2553 (N_2553,N_988,In_3329);
nor U2554 (N_2554,N_674,In_3695);
and U2555 (N_2555,N_1373,In_2176);
nand U2556 (N_2556,In_2536,In_292);
or U2557 (N_2557,N_1248,In_2478);
xor U2558 (N_2558,N_515,In_1706);
xnor U2559 (N_2559,N_758,N_1993);
xor U2560 (N_2560,In_379,In_4854);
xnor U2561 (N_2561,N_977,N_1118);
nand U2562 (N_2562,In_4313,In_1217);
or U2563 (N_2563,In_169,N_1726);
nor U2564 (N_2564,N_134,N_1094);
nand U2565 (N_2565,In_1587,In_3263);
or U2566 (N_2566,N_1188,N_1322);
or U2567 (N_2567,N_1231,In_1342);
and U2568 (N_2568,In_3996,N_1759);
or U2569 (N_2569,N_1604,In_4162);
or U2570 (N_2570,In_1830,N_1420);
or U2571 (N_2571,In_703,N_1160);
xor U2572 (N_2572,N_193,N_1071);
and U2573 (N_2573,N_1905,N_4);
or U2574 (N_2574,In_715,N_145);
nor U2575 (N_2575,In_1335,N_1097);
xor U2576 (N_2576,N_743,N_979);
or U2577 (N_2577,In_3667,N_626);
nand U2578 (N_2578,In_3989,In_3778);
and U2579 (N_2579,N_1804,N_907);
xnor U2580 (N_2580,N_672,In_3369);
xor U2581 (N_2581,N_461,N_801);
or U2582 (N_2582,N_1385,N_950);
xnor U2583 (N_2583,N_612,N_1477);
xor U2584 (N_2584,N_1585,N_1409);
or U2585 (N_2585,N_1313,In_4560);
and U2586 (N_2586,N_1099,N_1312);
nor U2587 (N_2587,N_1406,N_1954);
or U2588 (N_2588,N_466,N_1744);
xor U2589 (N_2589,In_3664,N_1467);
and U2590 (N_2590,N_1076,N_1736);
nand U2591 (N_2591,N_1894,N_1288);
and U2592 (N_2592,N_39,N_291);
xnor U2593 (N_2593,N_1648,In_484);
xor U2594 (N_2594,In_1612,N_833);
or U2595 (N_2595,In_3522,N_234);
nor U2596 (N_2596,N_1693,In_4749);
xnor U2597 (N_2597,In_110,N_407);
nand U2598 (N_2598,In_2341,In_4071);
or U2599 (N_2599,N_1283,N_858);
or U2600 (N_2600,N_1577,In_3852);
xor U2601 (N_2601,N_1615,N_1874);
nor U2602 (N_2602,N_1629,N_316);
and U2603 (N_2603,N_46,N_802);
or U2604 (N_2604,N_762,N_358);
and U2605 (N_2605,In_195,N_290);
nand U2606 (N_2606,In_3767,In_2242);
and U2607 (N_2607,N_366,N_1320);
xnor U2608 (N_2608,N_1329,N_1609);
and U2609 (N_2609,N_1066,N_1510);
and U2610 (N_2610,N_1246,N_878);
and U2611 (N_2611,N_437,N_1181);
nor U2612 (N_2612,N_199,N_1155);
or U2613 (N_2613,N_1092,N_821);
nor U2614 (N_2614,In_763,N_692);
and U2615 (N_2615,N_1608,N_99);
and U2616 (N_2616,In_4256,In_4920);
or U2617 (N_2617,N_1741,N_1820);
nand U2618 (N_2618,In_2180,N_1310);
xnor U2619 (N_2619,N_278,In_2531);
nand U2620 (N_2620,In_585,In_4898);
and U2621 (N_2621,In_3685,In_4629);
nand U2622 (N_2622,N_686,N_1742);
and U2623 (N_2623,N_1500,N_339);
and U2624 (N_2624,N_177,N_1463);
nor U2625 (N_2625,In_253,In_1326);
nor U2626 (N_2626,N_849,In_3979);
nor U2627 (N_2627,N_1161,In_4761);
or U2628 (N_2628,N_235,N_1392);
xnor U2629 (N_2629,In_1678,In_2296);
xor U2630 (N_2630,N_620,N_1517);
nand U2631 (N_2631,N_498,N_1991);
nand U2632 (N_2632,N_277,N_1832);
nand U2633 (N_2633,N_656,N_652);
or U2634 (N_2634,N_257,N_938);
nand U2635 (N_2635,N_1186,N_113);
nand U2636 (N_2636,In_4125,N_1381);
and U2637 (N_2637,N_1225,N_973);
nor U2638 (N_2638,In_4779,In_4894);
xor U2639 (N_2639,N_1916,In_1592);
xor U2640 (N_2640,In_3042,In_3675);
and U2641 (N_2641,N_1449,N_212);
and U2642 (N_2642,N_441,N_1150);
nor U2643 (N_2643,N_1151,In_4797);
xnor U2644 (N_2644,N_160,N_1536);
and U2645 (N_2645,N_1550,In_4884);
xor U2646 (N_2646,N_588,In_1264);
xnor U2647 (N_2647,In_1538,In_3050);
nand U2648 (N_2648,N_274,In_1546);
nor U2649 (N_2649,N_1067,In_3711);
nor U2650 (N_2650,N_1750,In_4708);
xnor U2651 (N_2651,N_1042,N_1765);
nor U2652 (N_2652,N_1343,In_2138);
and U2653 (N_2653,In_951,N_149);
nand U2654 (N_2654,N_784,N_226);
and U2655 (N_2655,N_1323,In_3268);
xnor U2656 (N_2656,N_1194,N_867);
and U2657 (N_2657,N_1512,N_1354);
and U2658 (N_2658,N_1469,In_3642);
nor U2659 (N_2659,N_386,In_922);
nand U2660 (N_2660,N_1372,In_443);
nor U2661 (N_2661,N_1696,N_553);
xnor U2662 (N_2662,N_1353,In_4056);
xnor U2663 (N_2663,In_4189,N_1732);
xnor U2664 (N_2664,N_1942,N_695);
xnor U2665 (N_2665,N_903,In_1136);
and U2666 (N_2666,N_489,In_1662);
xor U2667 (N_2667,In_4816,In_1943);
or U2668 (N_2668,N_1374,In_1490);
nor U2669 (N_2669,In_438,N_1854);
xor U2670 (N_2670,N_352,In_4015);
xnor U2671 (N_2671,N_1197,In_4803);
nand U2672 (N_2672,N_1839,In_3064);
nand U2673 (N_2673,N_522,N_259);
and U2674 (N_2674,N_1527,N_1260);
xnor U2675 (N_2675,In_2103,In_3443);
nor U2676 (N_2676,N_680,N_248);
or U2677 (N_2677,N_381,N_713);
or U2678 (N_2678,In_3301,In_857);
xor U2679 (N_2679,N_283,In_1102);
and U2680 (N_2680,N_1520,In_20);
and U2681 (N_2681,N_1093,N_1663);
or U2682 (N_2682,N_1034,N_830);
or U2683 (N_2683,N_1318,N_282);
nor U2684 (N_2684,N_304,N_371);
xnor U2685 (N_2685,N_476,In_4039);
nor U2686 (N_2686,In_2100,In_4980);
or U2687 (N_2687,N_1695,N_1824);
or U2688 (N_2688,In_629,In_1607);
nand U2689 (N_2689,In_3860,N_431);
nor U2690 (N_2690,In_4053,In_150);
nor U2691 (N_2691,In_442,In_118);
or U2692 (N_2692,In_1155,In_1113);
nor U2693 (N_2693,In_3386,In_3037);
and U2694 (N_2694,In_1526,N_547);
or U2695 (N_2695,N_590,In_3275);
nor U2696 (N_2696,N_228,N_834);
nor U2697 (N_2697,In_3773,N_1201);
and U2698 (N_2698,N_576,N_1727);
xnor U2699 (N_2699,N_512,In_3149);
nand U2700 (N_2700,N_1051,N_178);
xor U2701 (N_2701,In_4640,N_753);
nand U2702 (N_2702,N_1341,In_2606);
nand U2703 (N_2703,In_644,In_3968);
nand U2704 (N_2704,N_1581,In_77);
nand U2705 (N_2705,In_3690,In_1537);
or U2706 (N_2706,N_944,N_438);
or U2707 (N_2707,In_4773,N_1632);
or U2708 (N_2708,N_1058,In_498);
and U2709 (N_2709,In_1863,N_1781);
xor U2710 (N_2710,N_1844,N_1280);
nand U2711 (N_2711,N_840,In_2575);
xor U2712 (N_2712,N_423,N_1955);
nor U2713 (N_2713,In_2202,N_1734);
nand U2714 (N_2714,In_4144,N_1723);
xnor U2715 (N_2715,N_1992,N_1214);
and U2716 (N_2716,N_1990,N_519);
xnor U2717 (N_2717,N_1953,N_1212);
and U2718 (N_2718,In_2998,In_3326);
or U2719 (N_2719,In_1732,N_1684);
nor U2720 (N_2720,In_1154,N_75);
or U2721 (N_2721,In_3036,N_1525);
and U2722 (N_2722,In_2728,N_397);
nor U2723 (N_2723,In_2884,N_1476);
nand U2724 (N_2724,N_1682,N_18);
or U2725 (N_2725,N_36,N_726);
xnor U2726 (N_2726,In_3839,In_3510);
nor U2727 (N_2727,In_2571,In_1794);
or U2728 (N_2728,N_549,N_864);
nand U2729 (N_2729,In_2811,In_4792);
xor U2730 (N_2730,N_112,In_1801);
and U2731 (N_2731,N_1321,In_684);
nand U2732 (N_2732,N_419,N_93);
xnor U2733 (N_2733,In_568,N_473);
xnor U2734 (N_2734,In_48,In_4696);
nand U2735 (N_2735,In_1100,N_1448);
xor U2736 (N_2736,N_846,N_729);
xnor U2737 (N_2737,In_4605,N_1030);
nor U2738 (N_2738,N_1286,N_822);
nand U2739 (N_2739,N_1086,N_1351);
xnor U2740 (N_2740,N_1902,N_389);
nor U2741 (N_2741,In_205,N_1204);
nor U2742 (N_2742,In_4807,N_554);
and U2743 (N_2743,In_709,N_167);
and U2744 (N_2744,In_2507,In_3187);
nor U2745 (N_2745,N_861,In_1224);
nor U2746 (N_2746,N_985,In_2681);
or U2747 (N_2747,N_319,In_4995);
nor U2748 (N_2748,N_527,N_691);
nand U2749 (N_2749,N_343,In_1042);
or U2750 (N_2750,N_1496,N_595);
nand U2751 (N_2751,N_143,N_757);
nand U2752 (N_2752,N_600,N_1457);
and U2753 (N_2753,N_1018,N_826);
or U2754 (N_2754,N_260,N_908);
nor U2755 (N_2755,N_1275,N_1250);
and U2756 (N_2756,In_4660,N_1398);
and U2757 (N_2757,N_89,N_1835);
or U2758 (N_2758,N_1146,In_2289);
nor U2759 (N_2759,N_1416,N_138);
and U2760 (N_2760,N_764,N_792);
nand U2761 (N_2761,N_967,N_25);
nand U2762 (N_2762,In_4693,In_2925);
nor U2763 (N_2763,N_151,In_3780);
or U2764 (N_2764,N_1394,In_2135);
nand U2765 (N_2765,In_2516,N_1297);
or U2766 (N_2766,N_496,In_2541);
nor U2767 (N_2767,In_2451,N_119);
or U2768 (N_2768,N_392,N_1922);
and U2769 (N_2769,N_1966,In_1651);
and U2770 (N_2770,N_1900,N_1584);
and U2771 (N_2771,In_3700,In_3458);
nand U2772 (N_2772,N_1913,N_736);
nor U2773 (N_2773,In_2725,In_840);
or U2774 (N_2774,N_82,In_2841);
and U2775 (N_2775,In_1982,N_1881);
and U2776 (N_2776,N_751,In_1543);
nor U2777 (N_2777,N_924,In_2387);
nand U2778 (N_2778,In_4119,N_250);
and U2779 (N_2779,N_312,N_599);
and U2780 (N_2780,N_49,N_1951);
and U2781 (N_2781,N_1768,N_1829);
xor U2782 (N_2782,N_54,N_1636);
and U2783 (N_2783,N_267,In_2398);
nor U2784 (N_2784,In_2394,N_1669);
xnor U2785 (N_2785,In_2224,In_287);
or U2786 (N_2786,N_97,N_678);
xnor U2787 (N_2787,In_454,N_1713);
nor U2788 (N_2788,N_1809,In_1522);
or U2789 (N_2789,N_965,N_1274);
xor U2790 (N_2790,N_1010,In_2686);
nor U2791 (N_2791,In_1847,In_1329);
xor U2792 (N_2792,N_813,In_4651);
or U2793 (N_2793,In_3034,N_1588);
or U2794 (N_2794,N_783,N_1896);
nand U2795 (N_2795,N_1641,N_1586);
nor U2796 (N_2796,In_4094,In_3720);
nor U2797 (N_2797,In_2955,N_1267);
or U2798 (N_2798,N_1644,N_708);
and U2799 (N_2799,N_725,N_836);
nor U2800 (N_2800,In_4179,N_105);
nor U2801 (N_2801,N_28,N_21);
and U2802 (N_2802,In_1346,In_1554);
nand U2803 (N_2803,N_1154,N_586);
nand U2804 (N_2804,N_90,N_376);
xor U2805 (N_2805,N_1633,N_591);
or U2806 (N_2806,N_1429,N_1772);
and U2807 (N_2807,N_1138,In_2829);
or U2808 (N_2808,N_896,N_348);
xnor U2809 (N_2809,N_1348,In_1476);
nor U2810 (N_2810,N_346,N_837);
and U2811 (N_2811,N_766,N_1689);
or U2812 (N_2812,In_3985,In_1480);
nand U2813 (N_2813,In_4747,N_1361);
and U2814 (N_2814,N_991,In_3678);
nor U2815 (N_2815,N_1052,N_480);
xnor U2816 (N_2816,In_3078,N_1113);
nor U2817 (N_2817,In_4897,In_3617);
or U2818 (N_2818,In_3966,N_210);
or U2819 (N_2819,In_3926,N_215);
or U2820 (N_2820,N_1587,N_1834);
nor U2821 (N_2821,N_1254,N_540);
nand U2822 (N_2822,N_230,N_544);
nor U2823 (N_2823,N_379,N_1580);
or U2824 (N_2824,N_530,N_941);
nand U2825 (N_2825,N_905,In_2687);
nor U2826 (N_2826,In_133,N_484);
and U2827 (N_2827,N_1218,N_1497);
nor U2828 (N_2828,In_4100,N_1346);
xnor U2829 (N_2829,In_1941,N_1244);
nand U2830 (N_2830,N_1261,N_653);
nor U2831 (N_2831,N_1412,In_3584);
or U2832 (N_2832,N_724,In_3317);
nor U2833 (N_2833,N_902,N_297);
and U2834 (N_2834,N_1937,In_1281);
nor U2835 (N_2835,In_929,N_968);
nor U2836 (N_2836,N_483,In_4859);
xor U2837 (N_2837,N_179,N_882);
and U2838 (N_2838,N_755,In_1263);
or U2839 (N_2839,N_1694,N_582);
nand U2840 (N_2840,N_141,N_781);
xnor U2841 (N_2841,N_855,N_943);
or U2842 (N_2842,N_256,N_469);
or U2843 (N_2843,N_618,N_402);
nand U2844 (N_2844,N_1336,In_685);
and U2845 (N_2845,In_1030,N_1249);
and U2846 (N_2846,In_2295,N_1026);
xor U2847 (N_2847,In_3643,N_40);
nand U2848 (N_2848,N_185,N_310);
xnor U2849 (N_2849,N_72,N_1366);
or U2850 (N_2850,In_893,N_439);
nand U2851 (N_2851,N_1302,In_3054);
nand U2852 (N_2852,N_1872,N_1484);
nand U2853 (N_2853,In_2489,N_292);
nor U2854 (N_2854,N_1294,In_2454);
nor U2855 (N_2855,N_890,N_919);
nor U2856 (N_2856,N_1784,N_971);
nor U2857 (N_2857,In_3021,In_2747);
nor U2858 (N_2858,In_4487,N_505);
xor U2859 (N_2859,N_104,In_4714);
xor U2860 (N_2860,In_193,N_1652);
nor U2861 (N_2861,N_733,N_1048);
nor U2862 (N_2862,N_1968,In_119);
or U2863 (N_2863,In_138,N_372);
nand U2864 (N_2864,In_2533,In_714);
or U2865 (N_2865,In_823,N_1880);
nand U2866 (N_2866,N_123,N_294);
nand U2867 (N_2867,In_1411,N_1745);
xnor U2868 (N_2868,In_3003,In_2450);
or U2869 (N_2869,N_1628,N_1159);
nand U2870 (N_2870,N_1878,In_1775);
nor U2871 (N_2871,N_1126,N_1326);
or U2872 (N_2872,In_4288,N_897);
and U2873 (N_2873,N_1643,In_4962);
xnor U2874 (N_2874,In_565,N_848);
and U2875 (N_2875,N_453,In_1977);
nand U2876 (N_2876,N_1027,N_337);
nand U2877 (N_2877,N_1756,In_4636);
and U2878 (N_2878,N_1208,N_541);
xor U2879 (N_2879,In_2682,In_2153);
nand U2880 (N_2880,N_1256,N_947);
or U2881 (N_2881,N_393,N_1808);
or U2882 (N_2882,N_32,In_2548);
nand U2883 (N_2883,N_50,N_662);
and U2884 (N_2884,N_1339,N_150);
xor U2885 (N_2885,N_1610,N_1626);
or U2886 (N_2886,N_458,N_769);
or U2887 (N_2887,In_3974,N_1258);
xor U2888 (N_2888,N_799,N_842);
nor U2889 (N_2889,In_2774,N_746);
xnor U2890 (N_2890,N_777,N_1023);
xnor U2891 (N_2891,N_605,N_1570);
nor U2892 (N_2892,N_1413,N_1566);
or U2893 (N_2893,In_3770,N_350);
and U2894 (N_2894,In_45,In_1164);
nor U2895 (N_2895,N_1209,N_970);
nor U2896 (N_2896,N_1193,N_1078);
nand U2897 (N_2897,N_198,N_894);
or U2898 (N_2898,In_4863,N_1080);
nand U2899 (N_2899,In_802,N_642);
nand U2900 (N_2900,In_4230,In_2125);
nor U2901 (N_2901,In_3122,N_131);
or U2902 (N_2902,N_1928,In_2852);
nand U2903 (N_2903,N_275,N_1446);
and U2904 (N_2904,N_651,In_4233);
and U2905 (N_2905,N_1674,N_158);
xnor U2906 (N_2906,N_15,In_2805);
xnor U2907 (N_2907,N_1672,N_1519);
nand U2908 (N_2908,In_883,N_1060);
xnor U2909 (N_2909,N_325,N_1196);
xor U2910 (N_2910,N_798,In_3192);
or U2911 (N_2911,N_1837,N_1240);
nor U2912 (N_2912,N_717,N_992);
nand U2913 (N_2913,N_993,N_1235);
nand U2914 (N_2914,N_1567,N_589);
and U2915 (N_2915,N_1811,N_20);
xor U2916 (N_2916,N_1405,N_537);
or U2917 (N_2917,N_874,N_1714);
or U2918 (N_2918,N_1622,N_1700);
or U2919 (N_2919,N_117,In_1717);
or U2920 (N_2920,N_69,In_1063);
and U2921 (N_2921,N_1011,N_1592);
xnor U2922 (N_2922,N_415,N_1369);
xor U2923 (N_2923,N_1886,N_474);
or U2924 (N_2924,In_207,N_1779);
and U2925 (N_2925,In_17,N_1827);
and U2926 (N_2926,In_4027,N_156);
and U2927 (N_2927,N_317,N_1678);
xnor U2928 (N_2928,In_596,N_1483);
xor U2929 (N_2929,N_608,N_1311);
nand U2930 (N_2930,In_4020,N_1143);
or U2931 (N_2931,N_1432,N_518);
nor U2932 (N_2932,N_399,N_1451);
xnor U2933 (N_2933,N_1002,N_1399);
nor U2934 (N_2934,N_1982,N_486);
xor U2935 (N_2935,N_1657,In_4812);
and U2936 (N_2936,N_478,N_529);
and U2937 (N_2937,N_1920,N_1006);
nor U2938 (N_2938,N_571,N_807);
nand U2939 (N_2939,N_1414,In_352);
nand U2940 (N_2940,In_4133,In_2372);
and U2941 (N_2941,N_912,In_516);
and U2942 (N_2942,N_1328,N_188);
xnor U2943 (N_2943,In_526,In_1455);
or U2944 (N_2944,N_1068,N_915);
and U2945 (N_2945,N_1046,In_2057);
nand U2946 (N_2946,N_668,In_4353);
and U2947 (N_2947,N_1977,In_85);
or U2948 (N_2948,N_1224,N_1142);
and U2949 (N_2949,N_382,In_595);
nor U2950 (N_2950,N_92,N_1724);
or U2951 (N_2951,N_876,In_1477);
nor U2952 (N_2952,In_606,In_1497);
and U2953 (N_2953,N_1091,In_2872);
and U2954 (N_2954,N_196,In_4950);
or U2955 (N_2955,In_3252,In_1918);
nor U2956 (N_2956,N_1308,N_625);
and U2957 (N_2957,N_280,N_1925);
nor U2958 (N_2958,N_1059,N_1785);
or U2959 (N_2959,N_76,In_1305);
nor U2960 (N_2960,N_1293,N_983);
nand U2961 (N_2961,N_513,N_1625);
or U2962 (N_2962,N_667,In_4735);
xor U2963 (N_2963,N_225,N_1591);
nand U2964 (N_2964,N_748,N_1088);
or U2965 (N_2965,N_323,In_4679);
and U2966 (N_2966,N_405,N_1504);
nand U2967 (N_2967,In_2909,N_166);
and U2968 (N_2968,N_331,N_1767);
nor U2969 (N_2969,N_782,In_553);
nand U2970 (N_2970,N_644,N_181);
nand U2971 (N_2971,N_1486,N_31);
and U2972 (N_2972,In_731,N_832);
nor U2973 (N_2973,N_1325,N_606);
or U2974 (N_2974,N_630,In_3076);
and U2975 (N_2975,N_1569,In_2674);
nand U2976 (N_2976,In_92,In_3941);
xnor U2977 (N_2977,N_464,In_2321);
and U2978 (N_2978,In_4993,N_811);
nand U2979 (N_2979,N_1662,In_2339);
xor U2980 (N_2980,N_1969,In_597);
nor U2981 (N_2981,In_4524,N_839);
or U2982 (N_2982,In_4311,N_1719);
xor U2983 (N_2983,N_649,N_1315);
xnor U2984 (N_2984,In_4882,In_1605);
xnor U2985 (N_2985,In_1117,N_1747);
nor U2986 (N_2986,N_1522,N_759);
and U2987 (N_2987,N_596,In_1674);
or U2988 (N_2988,In_4507,N_154);
and U2989 (N_2989,N_1798,In_2632);
nand U2990 (N_2990,N_1401,N_1926);
and U2991 (N_2991,N_1606,N_1998);
and U2992 (N_2992,N_1659,N_367);
nand U2993 (N_2993,N_1364,In_116);
nand U2994 (N_2994,N_602,In_3223);
nand U2995 (N_2995,In_3254,N_1133);
and U2996 (N_2996,N_1362,In_2746);
and U2997 (N_2997,In_641,In_3408);
and U2998 (N_2998,N_1843,N_1959);
and U2999 (N_2999,N_1300,N_721);
or U3000 (N_3000,N_1127,N_320);
or U3001 (N_3001,N_1436,N_344);
and U3002 (N_3002,N_370,N_1620);
or U3003 (N_3003,In_717,N_1245);
nor U3004 (N_3004,N_1081,N_1475);
and U3005 (N_3005,N_1980,In_1320);
nand U3006 (N_3006,N_1624,N_1540);
nor U3007 (N_3007,N_611,N_1112);
nor U3008 (N_3008,In_4396,In_458);
and U3009 (N_3009,In_4239,In_4598);
nor U3010 (N_3010,N_1877,In_3886);
or U3011 (N_3011,N_1685,N_373);
nor U3012 (N_3012,In_3560,N_687);
nand U3013 (N_3013,N_648,In_1930);
xor U3014 (N_3014,N_1758,N_22);
nor U3015 (N_3015,N_747,N_673);
or U3016 (N_3016,N_1851,N_1728);
nand U3017 (N_3017,N_862,N_457);
nor U3018 (N_3018,In_4806,N_1518);
or U3019 (N_3019,In_274,N_1539);
and U3020 (N_3020,N_1045,N_361);
xnor U3021 (N_3021,N_1360,N_1135);
nor U3022 (N_3022,N_1383,N_1544);
nor U3023 (N_3023,In_1365,N_2);
nand U3024 (N_3024,N_1873,N_1332);
xnor U3025 (N_3025,N_1190,N_720);
nand U3026 (N_3026,N_1417,In_2078);
or U3027 (N_3027,In_4143,N_1978);
or U3028 (N_3028,N_465,N_1152);
and U3029 (N_3029,In_3235,N_650);
nor U3030 (N_3030,N_1831,N_1775);
xor U3031 (N_3031,N_1853,N_1028);
and U3032 (N_3032,N_1863,N_994);
or U3033 (N_3033,In_4193,In_3375);
and U3034 (N_3034,N_1941,In_1290);
nand U3035 (N_3035,N_1557,In_67);
xor U3036 (N_3036,N_276,N_187);
nor U3037 (N_3037,N_1679,N_1893);
xnor U3038 (N_3038,N_1746,In_1756);
and U3039 (N_3039,N_172,N_1611);
and U3040 (N_3040,In_3354,N_969);
or U3041 (N_3041,In_4135,N_1598);
and U3042 (N_3042,N_162,N_1252);
nor U3043 (N_3043,N_1600,In_2580);
xor U3044 (N_3044,N_1639,In_44);
xnor U3045 (N_3045,N_520,N_899);
or U3046 (N_3046,In_1581,N_581);
nor U3047 (N_3047,In_1858,N_223);
or U3048 (N_3048,In_3413,N_1823);
nand U3049 (N_3049,N_1748,N_772);
xnor U3050 (N_3050,N_1708,N_62);
nand U3051 (N_3051,In_497,N_929);
xor U3052 (N_3052,N_1961,N_533);
xnor U3053 (N_3053,In_4266,In_4970);
or U3054 (N_3054,In_1028,N_1883);
nand U3055 (N_3055,N_996,N_1985);
xor U3056 (N_3056,N_1568,N_1666);
nor U3057 (N_3057,In_4834,In_4686);
xor U3058 (N_3058,N_313,N_880);
xor U3059 (N_3059,In_932,In_4668);
nand U3060 (N_3060,In_2273,N_1903);
nor U3061 (N_3061,In_4552,N_1234);
xnor U3062 (N_3062,N_980,N_550);
nor U3063 (N_3063,N_1017,N_562);
nand U3064 (N_3064,N_1601,N_660);
or U3065 (N_3065,N_168,In_1808);
xnor U3066 (N_3066,N_1983,In_3676);
nand U3067 (N_3067,N_1033,N_52);
xnor U3068 (N_3068,In_3249,N_534);
xnor U3069 (N_3069,N_139,N_820);
nor U3070 (N_3070,N_1661,N_1210);
nor U3071 (N_3071,In_774,N_1069);
nand U3072 (N_3072,In_2265,N_869);
nor U3073 (N_3073,N_411,N_741);
or U3074 (N_3074,N_1352,In_2463);
xor U3075 (N_3075,N_265,N_427);
or U3076 (N_3076,N_773,N_791);
nor U3077 (N_3077,In_1626,N_27);
and U3078 (N_3078,N_271,N_698);
xor U3079 (N_3079,In_3287,In_2742);
xnor U3080 (N_3080,In_2593,In_1043);
and U3081 (N_3081,In_4665,In_3731);
nand U3082 (N_3082,N_937,N_1157);
and U3083 (N_3083,N_1761,N_1656);
nand U3084 (N_3084,N_1602,In_2716);
and U3085 (N_3085,In_240,N_1203);
nand U3086 (N_3086,N_956,In_1205);
xor U3087 (N_3087,N_13,In_1029);
and U3088 (N_3088,N_587,In_1912);
nand U3089 (N_3089,N_349,N_421);
nand U3090 (N_3090,In_2275,N_102);
and U3091 (N_3091,N_426,N_418);
and U3092 (N_3092,In_3167,N_1884);
and U3093 (N_3093,In_101,In_479);
and U3094 (N_3094,N_731,N_1547);
nand U3095 (N_3095,In_40,N_1974);
nand U3096 (N_3096,N_1106,In_4157);
xor U3097 (N_3097,N_1291,In_2972);
nand U3098 (N_3098,N_120,N_1698);
and U3099 (N_3099,N_1770,N_467);
and U3100 (N_3100,In_4274,N_633);
nand U3101 (N_3101,N_567,In_4051);
and U3102 (N_3102,In_2520,In_378);
and U3103 (N_3103,In_1152,In_445);
and U3104 (N_3104,In_4351,N_1111);
xor U3105 (N_3105,N_268,N_1395);
xor U3106 (N_3106,N_844,In_190);
and U3107 (N_3107,In_4069,N_808);
nor U3108 (N_3108,N_369,In_4627);
and U3109 (N_3109,N_125,In_4032);
nor U3110 (N_3110,N_1163,N_1480);
or U3111 (N_3111,In_4876,In_197);
nand U3112 (N_3112,N_1766,In_3995);
nand U3113 (N_3113,N_1717,N_359);
xnor U3114 (N_3114,N_86,N_1450);
nor U3115 (N_3115,N_1121,In_4154);
and U3116 (N_3116,N_1676,N_1271);
nor U3117 (N_3117,N_108,N_1247);
and U3118 (N_3118,In_186,N_180);
nor U3119 (N_3119,N_1729,N_1631);
nand U3120 (N_3120,N_666,N_1029);
or U3121 (N_3121,N_1677,N_301);
nor U3122 (N_3122,N_647,N_852);
xor U3123 (N_3123,N_1956,N_1933);
or U3124 (N_3124,N_517,In_4018);
nor U3125 (N_3125,N_511,N_3);
or U3126 (N_3126,N_1806,N_100);
nor U3127 (N_3127,N_1333,N_1472);
nand U3128 (N_3128,N_128,N_355);
and U3129 (N_3129,N_1857,In_784);
xor U3130 (N_3130,N_681,N_1743);
xor U3131 (N_3131,In_4257,N_1645);
nand U3132 (N_3132,N_236,N_1215);
nand U3133 (N_3133,In_2234,In_4000);
xor U3134 (N_3134,N_1437,N_868);
xnor U3135 (N_3135,N_451,N_1020);
nand U3136 (N_3136,N_1711,N_1850);
and U3137 (N_3137,N_362,N_270);
or U3138 (N_3138,N_1776,N_948);
xnor U3139 (N_3139,N_1036,N_1594);
nor U3140 (N_3140,N_209,N_1860);
nor U3141 (N_3141,In_2515,In_1893);
or U3142 (N_3142,N_1605,N_19);
xnor U3143 (N_3143,In_2803,In_786);
and U3144 (N_3144,N_1616,In_492);
and U3145 (N_3145,N_1651,In_2931);
or U3146 (N_3146,N_242,In_3224);
or U3147 (N_3147,In_3141,N_1909);
or U3148 (N_3148,N_398,N_471);
nand U3149 (N_3149,In_4323,N_677);
and U3150 (N_3150,N_1960,N_1375);
and U3151 (N_3151,N_932,N_1947);
and U3152 (N_3152,N_1817,N_1304);
nor U3153 (N_3153,N_700,N_1108);
or U3154 (N_3154,In_1356,N_169);
or U3155 (N_3155,N_564,N_603);
or U3156 (N_3156,N_161,N_1104);
or U3157 (N_3157,N_1780,N_1563);
and U3158 (N_3158,In_2192,N_689);
nand U3159 (N_3159,N_548,N_1797);
nor U3160 (N_3160,In_2633,In_2313);
nand U3161 (N_3161,N_109,N_140);
and U3162 (N_3162,N_500,N_33);
nand U3163 (N_3163,N_1507,N_560);
or U3164 (N_3164,N_1596,In_2420);
nor U3165 (N_3165,In_3139,N_1658);
xnor U3166 (N_3166,In_412,N_1560);
xor U3167 (N_3167,N_261,N_83);
nand U3168 (N_3168,In_4865,N_734);
xnor U3169 (N_3169,In_1138,N_1710);
or U3170 (N_3170,In_2335,N_1191);
nand U3171 (N_3171,In_3844,In_122);
xnor U3172 (N_3172,N_1239,N_37);
or U3173 (N_3173,In_2697,N_528);
or U3174 (N_3174,N_1468,N_1709);
nor U3175 (N_3175,N_1901,N_1623);
and U3176 (N_3176,N_1649,In_690);
or U3177 (N_3177,N_1195,In_4326);
nor U3178 (N_3178,N_934,N_490);
or U3179 (N_3179,N_1301,N_406);
or U3180 (N_3180,In_531,In_3874);
and U3181 (N_3181,N_737,N_508);
nand U3182 (N_3182,N_1433,N_898);
nor U3183 (N_3183,In_4009,N_913);
or U3184 (N_3184,N_175,N_1755);
and U3185 (N_3185,In_2090,In_4677);
nand U3186 (N_3186,N_1147,In_623);
xnor U3187 (N_3187,N_885,In_1814);
and U3188 (N_3188,N_551,N_1038);
nand U3189 (N_3189,In_4809,N_311);
and U3190 (N_3190,In_752,N_585);
xor U3191 (N_3191,In_4059,N_556);
or U3192 (N_3192,N_1904,N_507);
nand U3193 (N_3193,In_557,In_3717);
nand U3194 (N_3194,N_1531,In_735);
nor U3195 (N_3195,N_45,N_619);
nor U3196 (N_3196,N_1278,In_3494);
xor U3197 (N_3197,N_1116,In_3520);
nand U3198 (N_3198,In_1324,N_610);
or U3199 (N_3199,N_263,N_1130);
or U3200 (N_3200,In_4916,In_3934);
nand U3201 (N_3201,N_999,N_1640);
or U3202 (N_3202,N_1122,N_1022);
and U3203 (N_3203,In_451,In_3002);
xor U3204 (N_3204,In_2793,N_1821);
nor U3205 (N_3205,N_1943,N_1882);
nand U3206 (N_3206,N_1277,N_218);
xor U3207 (N_3207,In_1831,In_1602);
nand U3208 (N_3208,In_975,N_1439);
nor U3209 (N_3209,N_479,N_1595);
nor U3210 (N_3210,N_1597,In_2038);
nor U3211 (N_3211,N_646,N_1777);
xnor U3212 (N_3212,N_933,N_1760);
and U3213 (N_3213,In_1955,N_495);
nor U3214 (N_3214,N_1025,In_4786);
and U3215 (N_3215,In_393,N_133);
and U3216 (N_3216,N_1438,N_1718);
xor U3217 (N_3217,In_2698,N_1171);
nand U3218 (N_3218,N_531,N_1474);
nand U3219 (N_3219,N_815,N_506);
xnor U3220 (N_3220,N_1487,N_1132);
nand U3221 (N_3221,In_2866,N_171);
and U3222 (N_3222,N_1347,N_1043);
nor U3223 (N_3223,N_103,N_262);
xnor U3224 (N_3224,In_4240,N_1222);
nor U3225 (N_3225,N_1524,N_926);
nor U3226 (N_3226,N_146,N_390);
nand U3227 (N_3227,N_59,N_1668);
or U3228 (N_3228,In_4291,In_940);
and U3229 (N_3229,In_3528,In_2133);
xor U3230 (N_3230,N_1830,N_722);
nand U3231 (N_3231,N_1671,In_1657);
nor U3232 (N_3232,In_556,In_1645);
nand U3233 (N_3233,N_485,N_1793);
nand U3234 (N_3234,In_217,In_2446);
and U3235 (N_3235,N_1207,In_2179);
and U3236 (N_3236,N_309,N_65);
xor U3237 (N_3237,N_570,N_583);
or U3238 (N_3238,N_170,N_1921);
nand U3239 (N_3239,In_4017,N_504);
or U3240 (N_3240,In_3068,N_1390);
or U3241 (N_3241,N_1387,N_1175);
or U3242 (N_3242,N_754,N_1988);
nand U3243 (N_3243,N_1614,N_1019);
nand U3244 (N_3244,N_1735,In_3151);
nor U3245 (N_3245,N_1964,N_892);
and U3246 (N_3246,N_96,In_1786);
nor U3247 (N_3247,N_1172,In_512);
and U3248 (N_3248,N_1908,In_3285);
and U3249 (N_3249,N_456,In_1034);
xnor U3250 (N_3250,N_1630,N_1192);
xnor U3251 (N_3251,N_770,N_357);
nand U3252 (N_3252,N_790,In_4986);
or U3253 (N_3253,N_137,N_601);
and U3254 (N_3254,N_1996,N_243);
xor U3255 (N_3255,N_542,N_173);
nand U3256 (N_3256,N_1342,N_1090);
or U3257 (N_3257,N_1650,In_4635);
nand U3258 (N_3258,N_959,In_452);
xor U3259 (N_3259,N_810,N_1862);
nor U3260 (N_3260,N_377,N_347);
or U3261 (N_3261,In_995,N_315);
xnor U3262 (N_3262,N_1168,In_313);
xnor U3263 (N_3263,N_1408,In_4805);
and U3264 (N_3264,N_1139,In_1259);
and U3265 (N_3265,In_3158,N_775);
and U3266 (N_3266,In_2527,In_2761);
and U3267 (N_3267,In_213,N_1303);
and U3268 (N_3268,N_195,N_60);
nor U3269 (N_3269,In_758,N_435);
xnor U3270 (N_3270,N_1976,In_2065);
nand U3271 (N_3271,N_1141,In_1256);
or U3272 (N_3272,N_408,In_2207);
or U3273 (N_3273,N_577,In_364);
xnor U3274 (N_3274,N_1690,In_876);
xnor U3275 (N_3275,In_1902,In_2906);
or U3276 (N_3276,N_957,In_1300);
or U3277 (N_3277,In_3357,N_335);
or U3278 (N_3278,In_4825,In_331);
xnor U3279 (N_3279,In_2216,In_4908);
nor U3280 (N_3280,In_3107,In_4650);
nand U3281 (N_3281,In_2438,N_1967);
nor U3282 (N_3282,In_1846,N_1660);
nand U3283 (N_3283,N_1228,N_756);
nor U3284 (N_3284,In_4305,N_289);
and U3285 (N_3285,In_4624,N_1358);
and U3286 (N_3286,N_1816,In_2340);
or U3287 (N_3287,N_693,N_204);
and U3288 (N_3288,In_389,N_1211);
or U3289 (N_3289,N_960,N_184);
or U3290 (N_3290,N_351,N_838);
and U3291 (N_3291,N_1266,N_1647);
xor U3292 (N_3292,N_1389,In_2314);
nor U3293 (N_3293,N_1593,N_1063);
or U3294 (N_3294,N_224,N_16);
xor U3295 (N_3295,In_241,N_378);
and U3296 (N_3296,N_1720,N_1489);
and U3297 (N_3297,In_1750,N_1110);
nand U3298 (N_3298,In_435,N_51);
xor U3299 (N_3299,N_1482,N_266);
or U3300 (N_3300,N_284,N_216);
and U3301 (N_3301,N_1177,N_1098);
xnor U3302 (N_3302,N_931,N_639);
nor U3303 (N_3303,N_1494,In_3521);
xor U3304 (N_3304,In_1275,N_293);
and U3305 (N_3305,N_1024,N_675);
or U3306 (N_3306,N_124,In_912);
nor U3307 (N_3307,N_1455,N_732);
and U3308 (N_3308,In_2759,N_946);
and U3309 (N_3309,In_3045,In_601);
xor U3310 (N_3310,N_101,N_843);
nand U3311 (N_3311,In_4504,N_1162);
xor U3312 (N_3312,In_4074,N_1471);
xor U3313 (N_3313,N_1697,In_2601);
nor U3314 (N_3314,In_1640,In_2928);
or U3315 (N_3315,In_354,N_217);
and U3316 (N_3316,N_1107,In_2851);
xnor U3317 (N_3317,N_1219,N_1319);
nand U3318 (N_3318,N_1836,In_1641);
and U3319 (N_3319,N_702,N_1216);
and U3320 (N_3320,N_1607,N_1198);
nand U3321 (N_3321,In_4753,N_12);
nor U3322 (N_3322,In_4655,N_74);
nor U3323 (N_3323,N_856,In_3575);
or U3324 (N_3324,N_1062,N_213);
nand U3325 (N_3325,N_488,N_324);
and U3326 (N_3326,N_1858,N_246);
and U3327 (N_3327,N_1825,N_728);
or U3328 (N_3328,N_1799,N_763);
nand U3329 (N_3329,In_3880,In_2530);
nor U3330 (N_3330,In_3157,N_955);
nand U3331 (N_3331,N_958,N_975);
or U3332 (N_3332,In_1905,In_4084);
or U3333 (N_3333,N_1103,N_1590);
xor U3334 (N_3334,N_593,In_3236);
xor U3335 (N_3335,N_1800,In_3635);
nor U3336 (N_3336,N_1134,N_1807);
nor U3337 (N_3337,N_1393,N_157);
or U3338 (N_3338,In_2944,N_1397);
nor U3339 (N_3339,In_1147,N_1870);
xor U3340 (N_3340,N_785,N_1054);
and U3341 (N_3341,N_174,In_420);
or U3342 (N_3342,N_989,N_705);
nor U3343 (N_3343,In_1979,N_251);
xor U3344 (N_3344,In_923,In_3207);
xnor U3345 (N_3345,N_1558,N_1077);
or U3346 (N_3346,N_635,N_249);
nor U3347 (N_3347,N_1316,N_1064);
nor U3348 (N_3348,N_1749,In_3126);
nand U3349 (N_3349,N_1290,In_4476);
nand U3350 (N_3350,N_380,N_44);
nand U3351 (N_3351,In_47,In_767);
nand U3352 (N_3352,N_525,N_1541);
and U3353 (N_3353,N_939,In_4748);
nand U3354 (N_3354,N_472,N_401);
or U3355 (N_3355,N_854,N_883);
xor U3356 (N_3356,N_816,In_4929);
or U3357 (N_3357,N_679,In_4393);
nand U3358 (N_3358,N_1485,In_1403);
or U3359 (N_3359,N_909,In_1550);
xnor U3360 (N_3360,N_793,N_1265);
xor U3361 (N_3361,N_557,N_870);
or U3362 (N_3362,N_203,N_1789);
nand U3363 (N_3363,N_738,In_1216);
or U3364 (N_3364,N_1370,N_1535);
nand U3365 (N_3365,N_552,In_2064);
nand U3366 (N_3366,N_1701,N_1704);
and U3367 (N_3367,N_1376,N_1556);
and U3368 (N_3368,N_375,N_1938);
or U3369 (N_3369,In_4148,N_632);
nor U3370 (N_3370,N_306,N_1538);
or U3371 (N_3371,In_1894,N_1102);
nand U3372 (N_3372,N_1892,N_1906);
xor U3373 (N_3373,In_3269,N_914);
nor U3374 (N_3374,In_1646,N_1826);
nor U3375 (N_3375,N_1164,N_1675);
xor U3376 (N_3376,N_1929,N_889);
nand U3377 (N_3377,In_4591,N_189);
xnor U3378 (N_3378,N_1859,N_244);
or U3379 (N_3379,N_1434,In_589);
nand U3380 (N_3380,N_233,In_4097);
nand U3381 (N_3381,In_3293,N_1740);
nor U3382 (N_3382,N_712,N_279);
xor U3383 (N_3383,N_385,N_1932);
nor U3384 (N_3384,In_4519,N_696);
nor U3385 (N_3385,In_1496,N_144);
or U3386 (N_3386,N_499,In_2992);
and U3387 (N_3387,In_796,In_4713);
and U3388 (N_3388,In_2123,In_4945);
nand U3389 (N_3389,N_575,N_812);
and U3390 (N_3390,In_4388,In_1241);
xor U3391 (N_3391,N_327,N_1180);
or U3392 (N_3392,N_990,N_1564);
xnor U3393 (N_3393,N_1546,In_4869);
or U3394 (N_3394,N_617,N_1176);
and U3395 (N_3395,In_4129,N_1257);
nor U3396 (N_3396,N_1498,In_4952);
nor U3397 (N_3397,N_1576,N_1949);
nand U3398 (N_3398,N_1898,In_1032);
nand U3399 (N_3399,In_3756,In_2070);
or U3400 (N_3400,In_2956,N_636);
or U3401 (N_3401,N_953,N_1511);
or U3402 (N_3402,N_1378,N_1166);
or U3403 (N_3403,N_394,In_71);
xor U3404 (N_3404,In_2229,In_2904);
xor U3405 (N_3405,N_873,N_1243);
and U3406 (N_3406,In_3726,N_1752);
or U3407 (N_3407,N_1635,N_445);
nor U3408 (N_3408,In_968,In_429);
and U3409 (N_3409,In_1800,N_1400);
nor U3410 (N_3410,N_1276,N_481);
and U3411 (N_3411,N_935,In_3970);
nor U3412 (N_3412,N_207,In_2417);
or U3413 (N_3413,N_809,N_1753);
xnor U3414 (N_3414,N_1919,In_1176);
and U3415 (N_3415,N_1987,N_1115);
nor U3416 (N_3416,In_1500,N_1144);
nor U3417 (N_3417,N_1206,In_790);
xor U3418 (N_3418,In_1146,N_1047);
nand U3419 (N_3419,N_328,N_1357);
nand U3420 (N_3420,N_1885,N_778);
nor U3421 (N_3421,N_449,In_34);
nand U3422 (N_3422,N_413,N_841);
nand U3423 (N_3423,N_1136,In_2187);
and U3424 (N_3424,N_1667,N_940);
or U3425 (N_3425,N_624,In_3976);
nor U3426 (N_3426,N_1380,In_1398);
xor U3427 (N_3427,N_1335,N_1975);
or U3428 (N_3428,N_1039,In_2799);
and U3429 (N_3429,N_1757,N_1997);
xnor U3430 (N_3430,In_79,N_296);
xor U3431 (N_3431,N_191,N_1356);
nand U3432 (N_3432,N_0,N_1505);
xor U3433 (N_3433,N_434,N_1737);
xnor U3434 (N_3434,In_4314,N_1459);
nand U3435 (N_3435,In_3930,N_1501);
nand U3436 (N_3436,N_1187,N_865);
xor U3437 (N_3437,N_299,N_122);
and U3438 (N_3438,In_2796,N_1673);
and U3439 (N_3439,N_825,N_1073);
xnor U3440 (N_3440,In_285,In_1664);
xor U3441 (N_3441,In_652,In_3779);
nand U3442 (N_3442,In_1343,In_214);
nand U3443 (N_3443,N_928,N_1578);
and U3444 (N_3444,In_3901,N_921);
nor U3445 (N_3445,N_1253,In_1890);
nor U3446 (N_3446,N_1263,N_1344);
xor U3447 (N_3447,N_410,N_142);
nor U3448 (N_3448,In_1782,N_918);
and U3449 (N_3449,N_942,N_1529);
or U3450 (N_3450,In_242,N_1931);
nor U3451 (N_3451,N_1543,In_88);
and U3452 (N_3452,N_446,In_2461);
nand U3453 (N_3453,N_363,N_805);
nand U3454 (N_3454,N_29,N_1778);
and U3455 (N_3455,N_640,N_727);
and U3456 (N_3456,N_1733,In_4197);
nor U3457 (N_3457,In_255,N_1681);
xor U3458 (N_3458,N_1783,N_749);
xnor U3459 (N_3459,N_817,In_2263);
and U3460 (N_3460,In_4755,In_818);
and U3461 (N_3461,In_4461,In_166);
nand U3462 (N_3462,In_2753,N_254);
xnor U3463 (N_3463,N_1055,N_240);
and U3464 (N_3464,N_1070,N_1307);
xnor U3465 (N_3465,In_2025,N_1638);
xnor U3466 (N_3466,In_816,N_87);
xnor U3467 (N_3467,N_740,N_448);
xnor U3468 (N_3468,N_643,In_3153);
and U3469 (N_3469,N_384,N_685);
and U3470 (N_3470,N_795,N_1182);
and U3471 (N_3471,N_1642,In_3817);
nand U3472 (N_3472,N_730,N_1963);
xor U3473 (N_3473,N_1096,N_787);
xnor U3474 (N_3474,In_3437,N_1061);
xnor U3475 (N_3475,In_572,N_1680);
and U3476 (N_3476,In_1599,In_2145);
xnor U3477 (N_3477,In_4578,N_578);
nor U3478 (N_3478,N_1948,N_43);
nor U3479 (N_3479,N_1846,N_886);
nor U3480 (N_3480,N_1170,In_222);
and U3481 (N_3481,In_2165,N_771);
xnor U3482 (N_3482,N_623,N_1994);
and U3483 (N_3483,N_1049,In_2073);
or U3484 (N_3484,In_2178,N_1005);
or U3485 (N_3485,In_4204,N_814);
nand U3486 (N_3486,N_776,N_658);
nor U3487 (N_3487,N_494,N_1818);
or U3488 (N_3488,N_1292,In_3781);
xnor U3489 (N_3489,N_238,N_1537);
and U3490 (N_3490,N_368,In_1306);
nand U3491 (N_3491,N_1572,N_1082);
nor U3492 (N_3492,In_495,In_272);
xor U3493 (N_3493,In_1316,N_1549);
xor U3494 (N_3494,In_2267,N_1447);
nand U3495 (N_3495,In_3423,N_58);
or U3496 (N_3496,In_3338,N_546);
and U3497 (N_3497,In_2330,N_768);
and U3498 (N_3498,In_871,In_1492);
or U3499 (N_3499,In_4248,In_3855);
or U3500 (N_3500,In_1814,N_476);
nand U3501 (N_3501,N_785,N_1676);
nor U3502 (N_3502,In_664,N_1285);
or U3503 (N_3503,In_240,N_73);
or U3504 (N_3504,N_865,In_389);
nor U3505 (N_3505,N_1148,N_1062);
or U3506 (N_3506,In_436,In_454);
or U3507 (N_3507,N_1923,N_728);
xor U3508 (N_3508,N_525,N_1090);
xnor U3509 (N_3509,In_2609,N_1328);
and U3510 (N_3510,In_1660,N_56);
nand U3511 (N_3511,N_1167,N_1725);
and U3512 (N_3512,In_3767,N_1938);
nor U3513 (N_3513,In_2314,N_1262);
and U3514 (N_3514,In_150,N_803);
and U3515 (N_3515,In_2759,In_4884);
xor U3516 (N_3516,N_1166,N_741);
xor U3517 (N_3517,In_1146,N_1219);
and U3518 (N_3518,N_439,N_1275);
nor U3519 (N_3519,In_2192,In_4375);
nor U3520 (N_3520,N_1911,In_4256);
nand U3521 (N_3521,N_1890,N_804);
nor U3522 (N_3522,N_577,In_1497);
or U3523 (N_3523,N_91,In_2566);
nand U3524 (N_3524,N_883,In_4041);
nand U3525 (N_3525,In_3861,N_336);
or U3526 (N_3526,In_2263,N_284);
xor U3527 (N_3527,N_1122,N_1072);
xnor U3528 (N_3528,N_860,N_688);
nand U3529 (N_3529,N_1598,N_983);
nand U3530 (N_3530,N_997,N_1710);
and U3531 (N_3531,N_1918,N_1562);
and U3532 (N_3532,N_459,N_1594);
nand U3533 (N_3533,In_4768,N_1909);
or U3534 (N_3534,N_1968,N_868);
xnor U3535 (N_3535,In_3732,N_715);
and U3536 (N_3536,N_1302,N_760);
nand U3537 (N_3537,In_2237,N_527);
and U3538 (N_3538,N_1809,N_488);
or U3539 (N_3539,N_47,N_1518);
nand U3540 (N_3540,N_817,N_923);
and U3541 (N_3541,N_989,N_1074);
nor U3542 (N_3542,In_1941,N_970);
and U3543 (N_3543,In_1102,N_1062);
xor U3544 (N_3544,N_1543,N_590);
and U3545 (N_3545,N_759,In_240);
and U3546 (N_3546,N_1086,N_793);
and U3547 (N_3547,N_1262,N_497);
nand U3548 (N_3548,In_3285,N_1594);
nand U3549 (N_3549,N_1174,N_1800);
xnor U3550 (N_3550,N_1066,N_1052);
and U3551 (N_3551,N_2,N_1278);
and U3552 (N_3552,N_773,N_431);
nor U3553 (N_3553,N_1192,In_2263);
nor U3554 (N_3554,N_994,In_1863);
nand U3555 (N_3555,N_163,N_1211);
xnor U3556 (N_3556,In_1155,N_1676);
nor U3557 (N_3557,N_930,N_700);
and U3558 (N_3558,N_899,N_1078);
xnor U3559 (N_3559,N_553,N_1541);
xnor U3560 (N_3560,N_420,In_4375);
nor U3561 (N_3561,In_3187,N_1960);
and U3562 (N_3562,N_1131,N_440);
nand U3563 (N_3563,In_921,N_1234);
nor U3564 (N_3564,N_913,N_712);
nand U3565 (N_3565,In_4006,In_3930);
or U3566 (N_3566,N_779,N_967);
nor U3567 (N_3567,In_779,In_1278);
nand U3568 (N_3568,N_362,In_912);
nand U3569 (N_3569,N_1622,N_1171);
xnor U3570 (N_3570,N_545,N_401);
or U3571 (N_3571,N_1564,N_396);
and U3572 (N_3572,In_4522,In_3995);
or U3573 (N_3573,N_615,In_3635);
nand U3574 (N_3574,N_1631,In_1010);
nand U3575 (N_3575,N_11,N_1692);
xnor U3576 (N_3576,N_1657,N_1244);
and U3577 (N_3577,In_349,N_1141);
and U3578 (N_3578,N_1160,N_775);
and U3579 (N_3579,In_2339,N_1567);
or U3580 (N_3580,N_1494,In_1714);
and U3581 (N_3581,N_1488,N_1025);
nor U3582 (N_3582,N_1233,In_1574);
nand U3583 (N_3583,In_4970,In_4217);
xnor U3584 (N_3584,N_1140,In_1542);
or U3585 (N_3585,N_919,In_4805);
nand U3586 (N_3586,N_1143,N_742);
nand U3587 (N_3587,N_1936,N_1152);
xor U3588 (N_3588,In_4193,N_1347);
and U3589 (N_3589,N_549,N_1463);
nand U3590 (N_3590,N_1640,N_1984);
xnor U3591 (N_3591,N_570,N_197);
nand U3592 (N_3592,In_452,In_2799);
and U3593 (N_3593,N_1150,N_665);
xor U3594 (N_3594,N_414,N_60);
nor U3595 (N_3595,N_1337,N_1114);
and U3596 (N_3596,N_920,In_2537);
xnor U3597 (N_3597,N_303,In_1662);
nor U3598 (N_3598,N_600,In_596);
xnor U3599 (N_3599,N_155,N_1931);
nor U3600 (N_3600,In_1830,In_4313);
and U3601 (N_3601,N_657,In_4074);
and U3602 (N_3602,N_1848,N_1297);
nor U3603 (N_3603,In_4017,N_239);
nand U3604 (N_3604,N_80,N_1932);
or U3605 (N_3605,In_1316,In_3617);
nor U3606 (N_3606,In_3408,In_3621);
and U3607 (N_3607,In_3855,In_47);
and U3608 (N_3608,In_2263,N_304);
nor U3609 (N_3609,N_1937,N_378);
or U3610 (N_3610,N_1652,In_1801);
nand U3611 (N_3611,N_1078,In_638);
or U3612 (N_3612,N_579,N_412);
nand U3613 (N_3613,N_1499,N_1719);
and U3614 (N_3614,N_341,N_1180);
nand U3615 (N_3615,N_577,N_1085);
and U3616 (N_3616,In_4816,In_2593);
or U3617 (N_3617,In_389,In_1403);
nand U3618 (N_3618,In_387,N_263);
nand U3619 (N_3619,In_993,N_1424);
and U3620 (N_3620,In_2803,N_961);
nand U3621 (N_3621,In_4708,N_1836);
or U3622 (N_3622,In_2025,N_801);
nand U3623 (N_3623,In_242,In_1723);
nor U3624 (N_3624,N_211,In_3740);
or U3625 (N_3625,N_1846,N_12);
and U3626 (N_3626,N_391,N_763);
nor U3627 (N_3627,N_247,N_816);
nor U3628 (N_3628,N_181,N_1057);
nor U3629 (N_3629,In_3620,In_3021);
nor U3630 (N_3630,N_178,N_176);
or U3631 (N_3631,N_1768,N_1673);
and U3632 (N_3632,N_350,N_1227);
and U3633 (N_3633,In_4053,N_768);
nand U3634 (N_3634,N_854,N_426);
nand U3635 (N_3635,N_1891,N_217);
nor U3636 (N_3636,In_1758,N_737);
xnor U3637 (N_3637,N_259,N_203);
nand U3638 (N_3638,N_233,N_1691);
xor U3639 (N_3639,N_1474,N_1173);
nor U3640 (N_3640,N_1214,N_1724);
or U3641 (N_3641,N_1404,N_1056);
or U3642 (N_3642,N_270,N_1269);
nor U3643 (N_3643,N_617,N_514);
xnor U3644 (N_3644,N_904,N_780);
xor U3645 (N_3645,N_1108,In_2981);
nor U3646 (N_3646,N_468,In_3391);
xor U3647 (N_3647,N_1621,N_1576);
or U3648 (N_3648,In_4041,N_1221);
nor U3649 (N_3649,N_941,In_432);
and U3650 (N_3650,N_853,N_1657);
or U3651 (N_3651,N_964,N_176);
or U3652 (N_3652,N_969,N_824);
nor U3653 (N_3653,N_1044,N_1754);
and U3654 (N_3654,In_2981,N_480);
nand U3655 (N_3655,N_312,N_1054);
and U3656 (N_3656,N_1044,In_4898);
nand U3657 (N_3657,In_4055,N_1885);
or U3658 (N_3658,N_1119,N_1015);
or U3659 (N_3659,N_1438,N_365);
or U3660 (N_3660,N_718,N_1002);
and U3661 (N_3661,In_429,N_1347);
xnor U3662 (N_3662,N_8,In_4651);
or U3663 (N_3663,N_274,N_1);
or U3664 (N_3664,N_771,N_874);
xor U3665 (N_3665,In_1324,N_998);
and U3666 (N_3666,In_1918,In_181);
or U3667 (N_3667,N_743,N_1161);
nand U3668 (N_3668,N_1275,In_1102);
xor U3669 (N_3669,N_413,In_588);
or U3670 (N_3670,N_1824,N_1201);
xnor U3671 (N_3671,N_595,N_353);
xnor U3672 (N_3672,In_1102,N_1035);
nor U3673 (N_3673,N_1143,In_2843);
nand U3674 (N_3674,N_267,N_1403);
nor U3675 (N_3675,N_791,N_433);
and U3676 (N_3676,In_4519,N_871);
nor U3677 (N_3677,In_585,N_313);
nand U3678 (N_3678,In_4149,N_1693);
xnor U3679 (N_3679,N_1600,N_1678);
nand U3680 (N_3680,N_24,N_486);
nor U3681 (N_3681,In_492,In_3443);
xnor U3682 (N_3682,N_1409,In_4811);
nor U3683 (N_3683,N_1929,N_323);
nor U3684 (N_3684,In_1912,In_717);
nor U3685 (N_3685,N_665,N_1746);
xor U3686 (N_3686,N_979,N_1232);
nor U3687 (N_3687,N_1600,N_8);
and U3688 (N_3688,In_3676,N_1392);
xor U3689 (N_3689,N_367,In_1626);
nor U3690 (N_3690,In_2928,In_3719);
nand U3691 (N_3691,N_783,N_445);
nor U3692 (N_3692,N_1913,N_1926);
or U3693 (N_3693,In_4908,N_1969);
xor U3694 (N_3694,N_630,In_1133);
or U3695 (N_3695,In_484,N_455);
or U3696 (N_3696,N_448,In_4635);
nor U3697 (N_3697,In_2937,In_4571);
xnor U3698 (N_3698,N_382,In_2537);
xnor U3699 (N_3699,N_1009,N_606);
and U3700 (N_3700,N_823,In_1335);
xnor U3701 (N_3701,N_1429,N_148);
and U3702 (N_3702,In_1791,In_4732);
nand U3703 (N_3703,N_750,In_2944);
nor U3704 (N_3704,In_2464,N_891);
or U3705 (N_3705,N_1136,N_1028);
and U3706 (N_3706,N_1129,N_1310);
nand U3707 (N_3707,In_3773,In_412);
or U3708 (N_3708,N_1115,In_4160);
nor U3709 (N_3709,N_1963,N_1406);
xnor U3710 (N_3710,In_4590,N_63);
xnor U3711 (N_3711,N_1620,N_1653);
and U3712 (N_3712,In_1010,N_951);
nor U3713 (N_3713,In_4138,In_4650);
and U3714 (N_3714,N_1653,N_529);
nor U3715 (N_3715,In_585,N_1561);
xnor U3716 (N_3716,N_1434,N_1709);
or U3717 (N_3717,In_1425,N_609);
nor U3718 (N_3718,N_958,N_1161);
or U3719 (N_3719,N_923,In_389);
nand U3720 (N_3720,N_367,N_1612);
or U3721 (N_3721,N_1394,N_1710);
and U3722 (N_3722,N_1473,N_778);
nand U3723 (N_3723,N_1200,N_378);
and U3724 (N_3724,In_3560,In_4605);
and U3725 (N_3725,N_1310,N_1895);
nand U3726 (N_3726,In_2579,N_1000);
nand U3727 (N_3727,N_1484,In_4375);
xor U3728 (N_3728,N_1008,N_662);
xor U3729 (N_3729,N_295,N_567);
and U3730 (N_3730,In_205,In_3770);
xor U3731 (N_3731,N_1992,In_993);
xor U3732 (N_3732,N_1609,In_1953);
nor U3733 (N_3733,In_4021,N_138);
nand U3734 (N_3734,In_3726,N_1210);
nor U3735 (N_3735,In_1133,N_1490);
nor U3736 (N_3736,N_1959,In_2805);
nand U3737 (N_3737,N_1702,N_425);
or U3738 (N_3738,N_781,N_1092);
and U3739 (N_3739,N_988,N_581);
xor U3740 (N_3740,In_3852,In_767);
nand U3741 (N_3741,N_1503,N_605);
or U3742 (N_3742,N_938,N_1430);
or U3743 (N_3743,N_29,N_1974);
or U3744 (N_3744,N_1605,In_1903);
xor U3745 (N_3745,N_1800,N_368);
nor U3746 (N_3746,In_3501,In_4715);
nand U3747 (N_3747,N_1186,N_1950);
nor U3748 (N_3748,In_1515,N_626);
nand U3749 (N_3749,N_1750,In_595);
nand U3750 (N_3750,N_494,N_366);
nor U3751 (N_3751,N_272,In_3901);
nor U3752 (N_3752,In_2956,N_1230);
or U3753 (N_3753,N_1170,In_1831);
and U3754 (N_3754,N_682,N_1376);
nor U3755 (N_3755,N_615,N_1622);
nand U3756 (N_3756,In_2687,In_400);
xor U3757 (N_3757,N_1698,In_2056);
and U3758 (N_3758,N_1722,N_407);
xor U3759 (N_3759,N_786,In_3310);
and U3760 (N_3760,In_393,In_2981);
or U3761 (N_3761,N_167,In_2687);
nand U3762 (N_3762,In_3383,N_1802);
xor U3763 (N_3763,N_1663,N_1318);
nor U3764 (N_3764,N_1385,N_674);
xnor U3765 (N_3765,N_1104,In_2162);
xor U3766 (N_3766,In_2998,N_158);
or U3767 (N_3767,N_1971,In_3956);
xor U3768 (N_3768,In_3167,N_1348);
nor U3769 (N_3769,N_1256,N_80);
and U3770 (N_3770,N_367,In_1403);
or U3771 (N_3771,In_4323,N_595);
and U3772 (N_3772,N_162,N_346);
nor U3773 (N_3773,In_4625,In_122);
or U3774 (N_3774,In_3703,In_1858);
nand U3775 (N_3775,In_4859,In_3106);
nand U3776 (N_3776,N_766,N_1208);
or U3777 (N_3777,In_4242,N_962);
nand U3778 (N_3778,N_1438,N_1103);
xor U3779 (N_3779,N_1951,N_902);
and U3780 (N_3780,N_919,N_857);
nor U3781 (N_3781,In_2956,In_3797);
xnor U3782 (N_3782,N_659,N_103);
or U3783 (N_3783,N_1385,N_937);
nor U3784 (N_3784,N_1232,N_1536);
or U3785 (N_3785,N_667,N_148);
xor U3786 (N_3786,In_1657,In_4039);
nor U3787 (N_3787,In_2202,N_281);
or U3788 (N_3788,In_1581,N_987);
or U3789 (N_3789,N_479,N_1621);
nor U3790 (N_3790,N_1342,N_71);
or U3791 (N_3791,In_2148,N_1398);
and U3792 (N_3792,N_661,N_272);
or U3793 (N_3793,In_4266,In_3413);
nand U3794 (N_3794,N_1018,N_1734);
nor U3795 (N_3795,In_3676,In_3717);
xnor U3796 (N_3796,N_1045,In_784);
nor U3797 (N_3797,In_818,N_234);
nor U3798 (N_3798,In_1411,In_4834);
nor U3799 (N_3799,N_596,N_1829);
or U3800 (N_3800,N_1223,N_1540);
and U3801 (N_3801,N_1124,In_3695);
or U3802 (N_3802,In_2295,N_1238);
and U3803 (N_3803,In_731,N_861);
nor U3804 (N_3804,N_22,In_3996);
nor U3805 (N_3805,In_1808,N_1157);
nand U3806 (N_3806,In_4797,N_669);
nor U3807 (N_3807,In_3076,N_541);
nor U3808 (N_3808,In_763,In_3868);
nand U3809 (N_3809,N_751,N_1953);
nor U3810 (N_3810,N_1168,N_382);
or U3811 (N_3811,N_1739,In_3068);
and U3812 (N_3812,N_1679,In_2516);
or U3813 (N_3813,N_1386,N_132);
xnor U3814 (N_3814,N_791,N_1387);
nand U3815 (N_3815,N_1406,N_1845);
nand U3816 (N_3816,N_1608,In_2057);
xnor U3817 (N_3817,N_96,N_304);
and U3818 (N_3818,N_432,In_3057);
and U3819 (N_3819,N_238,N_99);
nand U3820 (N_3820,In_4834,In_1509);
nand U3821 (N_3821,N_509,N_1779);
and U3822 (N_3822,In_2100,In_2246);
nor U3823 (N_3823,N_161,In_4911);
nor U3824 (N_3824,N_732,N_991);
or U3825 (N_3825,In_3691,In_3437);
or U3826 (N_3826,N_955,In_3855);
nand U3827 (N_3827,In_3620,N_335);
and U3828 (N_3828,In_2811,N_1919);
nor U3829 (N_3829,In_4749,N_1877);
nand U3830 (N_3830,N_100,N_1576);
xor U3831 (N_3831,N_1118,N_1311);
nand U3832 (N_3832,N_1758,In_4605);
or U3833 (N_3833,N_5,In_3413);
nor U3834 (N_3834,In_593,N_1472);
nand U3835 (N_3835,N_1097,N_981);
xnor U3836 (N_3836,N_1453,N_872);
nand U3837 (N_3837,N_1494,N_1840);
or U3838 (N_3838,N_208,N_1335);
nor U3839 (N_3839,N_1731,N_1251);
or U3840 (N_3840,In_869,N_541);
or U3841 (N_3841,N_1693,N_1976);
or U3842 (N_3842,N_661,N_978);
or U3843 (N_3843,N_907,In_712);
xnor U3844 (N_3844,In_329,N_561);
or U3845 (N_3845,In_3254,N_1907);
nand U3846 (N_3846,In_889,N_897);
and U3847 (N_3847,In_651,N_1159);
nor U3848 (N_3848,In_2059,N_1146);
nand U3849 (N_3849,N_1178,N_789);
xor U3850 (N_3850,N_138,N_1414);
nor U3851 (N_3851,N_619,N_1561);
nand U3852 (N_3852,N_519,N_562);
or U3853 (N_3853,N_1809,N_1629);
or U3854 (N_3854,N_156,N_311);
nor U3855 (N_3855,N_1977,N_603);
nor U3856 (N_3856,In_4247,N_1590);
and U3857 (N_3857,N_717,N_500);
and U3858 (N_3858,In_3974,In_1146);
xor U3859 (N_3859,N_678,In_4908);
or U3860 (N_3860,In_2761,N_841);
and U3861 (N_3861,N_221,N_967);
nor U3862 (N_3862,N_560,N_43);
xnor U3863 (N_3863,N_105,N_505);
and U3864 (N_3864,N_1185,N_1030);
xor U3865 (N_3865,N_1893,In_3780);
or U3866 (N_3866,N_1691,In_4297);
or U3867 (N_3867,In_3254,N_676);
nand U3868 (N_3868,N_1155,N_1302);
nor U3869 (N_3869,N_314,In_557);
nor U3870 (N_3870,N_974,In_4069);
nand U3871 (N_3871,N_1507,N_20);
or U3872 (N_3872,In_492,N_1598);
nor U3873 (N_3873,N_1470,In_4405);
or U3874 (N_3874,N_1780,In_1003);
xor U3875 (N_3875,N_694,N_43);
and U3876 (N_3876,N_469,In_2448);
xnor U3877 (N_3877,N_944,N_1309);
and U3878 (N_3878,In_34,N_722);
nor U3879 (N_3879,N_317,In_454);
and U3880 (N_3880,In_4323,In_2937);
or U3881 (N_3881,N_411,In_1490);
nand U3882 (N_3882,In_1649,N_923);
and U3883 (N_3883,N_296,In_2747);
and U3884 (N_3884,In_2133,N_871);
nor U3885 (N_3885,In_242,N_1005);
nor U3886 (N_3886,N_1995,N_433);
and U3887 (N_3887,In_2725,In_2841);
xor U3888 (N_3888,N_492,N_1685);
nand U3889 (N_3889,N_735,N_819);
or U3890 (N_3890,In_4125,N_1193);
xnor U3891 (N_3891,N_783,In_3149);
or U3892 (N_3892,N_1647,N_1207);
or U3893 (N_3893,N_4,N_922);
or U3894 (N_3894,N_1436,N_1981);
or U3895 (N_3895,N_715,In_1589);
or U3896 (N_3896,N_1312,N_832);
xor U3897 (N_3897,N_1781,In_2759);
nand U3898 (N_3898,N_895,In_241);
nand U3899 (N_3899,N_1585,N_1261);
nand U3900 (N_3900,In_262,N_1627);
nor U3901 (N_3901,In_1275,N_1923);
nor U3902 (N_3902,N_255,N_534);
or U3903 (N_3903,N_1480,In_2537);
nand U3904 (N_3904,N_1379,In_3107);
xor U3905 (N_3905,In_1403,N_59);
or U3906 (N_3906,In_85,N_1210);
xnor U3907 (N_3907,N_1128,N_103);
xor U3908 (N_3908,N_33,In_2446);
nor U3909 (N_3909,N_766,N_1316);
and U3910 (N_3910,N_1879,N_862);
nand U3911 (N_3911,N_1482,In_1480);
nand U3912 (N_3912,In_4840,N_1047);
and U3913 (N_3913,In_3502,N_1537);
nand U3914 (N_3914,N_1327,N_131);
xor U3915 (N_3915,N_1443,N_1137);
nand U3916 (N_3916,N_1641,N_1002);
and U3917 (N_3917,N_846,In_1647);
nor U3918 (N_3918,In_4911,N_1774);
nor U3919 (N_3919,N_679,N_1656);
or U3920 (N_3920,N_1358,N_1178);
and U3921 (N_3921,In_4423,N_111);
or U3922 (N_3922,In_349,N_356);
and U3923 (N_3923,In_3904,N_1542);
nand U3924 (N_3924,N_1690,In_4204);
xor U3925 (N_3925,N_577,In_1693);
xor U3926 (N_3926,N_1024,N_872);
xor U3927 (N_3927,N_765,N_52);
nor U3928 (N_3928,N_210,N_1246);
nand U3929 (N_3929,N_1074,N_950);
and U3930 (N_3930,N_779,In_1197);
and U3931 (N_3931,In_4898,N_365);
xnor U3932 (N_3932,N_1278,N_1081);
nor U3933 (N_3933,In_2267,N_1915);
xnor U3934 (N_3934,In_4624,N_504);
and U3935 (N_3935,In_2796,N_1945);
nor U3936 (N_3936,N_641,In_758);
nor U3937 (N_3937,N_1292,N_224);
and U3938 (N_3938,N_400,In_2635);
xnor U3939 (N_3939,In_1791,In_916);
or U3940 (N_3940,N_246,N_693);
nor U3941 (N_3941,N_118,N_1863);
nand U3942 (N_3942,N_930,In_4652);
nor U3943 (N_3943,N_118,N_1713);
nand U3944 (N_3944,N_1507,In_4629);
nor U3945 (N_3945,In_4710,In_910);
and U3946 (N_3946,N_436,In_3386);
xor U3947 (N_3947,N_1099,In_4713);
or U3948 (N_3948,N_1969,In_364);
and U3949 (N_3949,N_1993,In_893);
xor U3950 (N_3950,N_1386,In_3141);
nand U3951 (N_3951,In_2339,N_217);
xnor U3952 (N_3952,N_1852,In_4080);
nor U3953 (N_3953,In_2716,N_1195);
xor U3954 (N_3954,N_1394,In_709);
xor U3955 (N_3955,N_490,N_1244);
or U3956 (N_3956,N_532,N_1181);
nor U3957 (N_3957,N_1733,N_1642);
nor U3958 (N_3958,N_1680,In_2202);
xnor U3959 (N_3959,N_1252,N_1407);
xor U3960 (N_3960,N_297,N_482);
nor U3961 (N_3961,N_1020,N_1693);
nor U3962 (N_3962,N_1622,N_1763);
xnor U3963 (N_3963,N_1305,N_298);
nor U3964 (N_3964,N_383,N_816);
xor U3965 (N_3965,N_1043,In_3584);
and U3966 (N_3966,N_300,N_209);
nand U3967 (N_3967,N_134,N_705);
nand U3968 (N_3968,N_160,In_712);
or U3969 (N_3969,N_1348,N_1233);
xnor U3970 (N_3970,N_988,N_910);
and U3971 (N_3971,N_359,N_745);
or U3972 (N_3972,N_1228,N_1991);
xor U3973 (N_3973,N_902,In_3126);
nor U3974 (N_3974,N_966,In_1176);
nand U3975 (N_3975,N_88,In_4056);
nor U3976 (N_3976,N_832,N_1720);
nor U3977 (N_3977,In_479,In_3130);
nor U3978 (N_3978,In_3310,N_195);
nand U3979 (N_3979,In_678,In_2621);
or U3980 (N_3980,N_37,In_4243);
and U3981 (N_3981,N_1961,In_4613);
and U3982 (N_3982,N_1115,In_2179);
nor U3983 (N_3983,N_1971,In_3857);
and U3984 (N_3984,In_2654,N_361);
and U3985 (N_3985,In_352,N_966);
or U3986 (N_3986,N_295,In_3966);
and U3987 (N_3987,N_755,N_1711);
nand U3988 (N_3988,N_227,In_1259);
nor U3989 (N_3989,In_1365,N_1794);
and U3990 (N_3990,In_2533,N_1395);
nor U3991 (N_3991,N_1669,N_1328);
and U3992 (N_3992,N_198,N_14);
xnor U3993 (N_3993,N_1564,N_1373);
and U3994 (N_3994,N_766,N_354);
nor U3995 (N_3995,In_136,In_3789);
or U3996 (N_3996,N_1210,N_967);
nand U3997 (N_3997,N_1860,N_1755);
nand U3998 (N_3998,N_713,N_822);
nand U3999 (N_3999,In_17,N_1120);
nor U4000 (N_4000,N_2863,N_3935);
xor U4001 (N_4001,N_2245,N_3807);
nor U4002 (N_4002,N_3901,N_2335);
or U4003 (N_4003,N_2744,N_2944);
nand U4004 (N_4004,N_3898,N_2295);
or U4005 (N_4005,N_2745,N_2782);
or U4006 (N_4006,N_2401,N_3179);
and U4007 (N_4007,N_2681,N_3512);
nor U4008 (N_4008,N_2708,N_3309);
or U4009 (N_4009,N_2942,N_2317);
and U4010 (N_4010,N_2717,N_2080);
and U4011 (N_4011,N_3742,N_2904);
nand U4012 (N_4012,N_3975,N_2582);
or U4013 (N_4013,N_2957,N_3596);
and U4014 (N_4014,N_3516,N_2491);
and U4015 (N_4015,N_3958,N_2680);
nor U4016 (N_4016,N_2148,N_3577);
or U4017 (N_4017,N_3295,N_2751);
xnor U4018 (N_4018,N_3024,N_2369);
or U4019 (N_4019,N_2253,N_2059);
xor U4020 (N_4020,N_2410,N_3598);
nand U4021 (N_4021,N_2959,N_2179);
nor U4022 (N_4022,N_3730,N_2884);
nand U4023 (N_4023,N_3037,N_2125);
and U4024 (N_4024,N_2504,N_3484);
nand U4025 (N_4025,N_2409,N_2799);
or U4026 (N_4026,N_2083,N_3360);
and U4027 (N_4027,N_2065,N_2828);
and U4028 (N_4028,N_3877,N_3305);
xor U4029 (N_4029,N_2063,N_3056);
nor U4030 (N_4030,N_3226,N_3897);
and U4031 (N_4031,N_3814,N_2399);
and U4032 (N_4032,N_3448,N_2336);
nor U4033 (N_4033,N_3550,N_3185);
xnor U4034 (N_4034,N_3077,N_2593);
nand U4035 (N_4035,N_2263,N_2524);
nand U4036 (N_4036,N_3950,N_2881);
or U4037 (N_4037,N_2784,N_2662);
nand U4038 (N_4038,N_2756,N_2290);
and U4039 (N_4039,N_3416,N_3803);
nand U4040 (N_4040,N_2580,N_2071);
nand U4041 (N_4041,N_3228,N_2286);
nor U4042 (N_4042,N_2511,N_3816);
or U4043 (N_4043,N_3049,N_3015);
and U4044 (N_4044,N_3674,N_3621);
nand U4045 (N_4045,N_3557,N_3172);
and U4046 (N_4046,N_3451,N_2872);
nand U4047 (N_4047,N_3833,N_3836);
and U4048 (N_4048,N_2643,N_2352);
or U4049 (N_4049,N_2636,N_2014);
or U4050 (N_4050,N_3963,N_2283);
and U4051 (N_4051,N_3311,N_2720);
and U4052 (N_4052,N_2984,N_3107);
and U4053 (N_4053,N_2417,N_3834);
or U4054 (N_4054,N_3194,N_3640);
xnor U4055 (N_4055,N_2671,N_2235);
xor U4056 (N_4056,N_2246,N_2448);
and U4057 (N_4057,N_2172,N_2537);
xor U4058 (N_4058,N_3424,N_3671);
xor U4059 (N_4059,N_3708,N_3143);
xor U4060 (N_4060,N_3246,N_3085);
and U4061 (N_4061,N_3623,N_3321);
or U4062 (N_4062,N_2595,N_3337);
and U4063 (N_4063,N_3458,N_2338);
nand U4064 (N_4064,N_2199,N_3619);
or U4065 (N_4065,N_2534,N_3693);
xor U4066 (N_4066,N_2015,N_3526);
and U4067 (N_4067,N_2356,N_2438);
or U4068 (N_4068,N_2652,N_3464);
nand U4069 (N_4069,N_3601,N_2358);
and U4070 (N_4070,N_2702,N_2189);
or U4071 (N_4071,N_3747,N_2215);
nor U4072 (N_4072,N_2300,N_2182);
nand U4073 (N_4073,N_2735,N_3639);
xnor U4074 (N_4074,N_2510,N_3251);
or U4075 (N_4075,N_3072,N_2326);
xor U4076 (N_4076,N_3564,N_2183);
nor U4077 (N_4077,N_2441,N_2332);
or U4078 (N_4078,N_3993,N_2343);
xor U4079 (N_4079,N_2716,N_3213);
and U4080 (N_4080,N_2459,N_3981);
or U4081 (N_4081,N_3168,N_2700);
and U4082 (N_4082,N_2777,N_3644);
nand U4083 (N_4083,N_2827,N_3676);
xnor U4084 (N_4084,N_2365,N_2414);
and U4085 (N_4085,N_2536,N_2293);
nand U4086 (N_4086,N_2561,N_2411);
and U4087 (N_4087,N_3007,N_2073);
and U4088 (N_4088,N_2377,N_2210);
and U4089 (N_4089,N_3500,N_2242);
xnor U4090 (N_4090,N_2655,N_3068);
or U4091 (N_4091,N_2370,N_3414);
xor U4092 (N_4092,N_2668,N_2673);
nor U4093 (N_4093,N_2820,N_2113);
nor U4094 (N_4094,N_3805,N_2875);
xnor U4095 (N_4095,N_3562,N_2017);
or U4096 (N_4096,N_3064,N_3374);
nand U4097 (N_4097,N_2806,N_3934);
nand U4098 (N_4098,N_2496,N_3095);
and U4099 (N_4099,N_3438,N_2021);
xor U4100 (N_4100,N_2824,N_3849);
nand U4101 (N_4101,N_3983,N_2546);
xor U4102 (N_4102,N_2223,N_2285);
or U4103 (N_4103,N_3631,N_3535);
nor U4104 (N_4104,N_3613,N_3061);
nand U4105 (N_4105,N_2505,N_3120);
nand U4106 (N_4106,N_3405,N_2667);
and U4107 (N_4107,N_2575,N_2353);
xor U4108 (N_4108,N_2938,N_3561);
nor U4109 (N_4109,N_3112,N_3752);
or U4110 (N_4110,N_3231,N_2030);
or U4111 (N_4111,N_3300,N_3731);
xor U4112 (N_4112,N_2978,N_3522);
xor U4113 (N_4113,N_3303,N_3127);
or U4114 (N_4114,N_2960,N_3216);
or U4115 (N_4115,N_2882,N_3724);
and U4116 (N_4116,N_2614,N_3200);
or U4117 (N_4117,N_2874,N_2712);
or U4118 (N_4118,N_3971,N_3973);
or U4119 (N_4119,N_3253,N_3883);
or U4120 (N_4120,N_3060,N_3802);
or U4121 (N_4121,N_3402,N_2616);
xor U4122 (N_4122,N_2980,N_2856);
nor U4123 (N_4123,N_3086,N_2936);
or U4124 (N_4124,N_3835,N_2967);
or U4125 (N_4125,N_3543,N_2398);
nor U4126 (N_4126,N_2306,N_2109);
and U4127 (N_4127,N_3141,N_3385);
nor U4128 (N_4128,N_2328,N_2986);
and U4129 (N_4129,N_2547,N_3741);
or U4130 (N_4130,N_2452,N_3738);
or U4131 (N_4131,N_2044,N_2344);
and U4132 (N_4132,N_3480,N_2259);
and U4133 (N_4133,N_2832,N_3444);
and U4134 (N_4134,N_3383,N_2810);
nand U4135 (N_4135,N_2964,N_3767);
and U4136 (N_4136,N_3240,N_3599);
nand U4137 (N_4137,N_2270,N_2323);
nor U4138 (N_4138,N_3230,N_2072);
nand U4139 (N_4139,N_2633,N_2990);
and U4140 (N_4140,N_2579,N_2724);
or U4141 (N_4141,N_3638,N_2236);
xor U4142 (N_4142,N_3186,N_2418);
and U4143 (N_4143,N_3398,N_2953);
and U4144 (N_4144,N_3870,N_2238);
nor U4145 (N_4145,N_3361,N_2212);
xnor U4146 (N_4146,N_3207,N_2552);
xnor U4147 (N_4147,N_3697,N_2996);
or U4148 (N_4148,N_2887,N_2195);
and U4149 (N_4149,N_3918,N_3197);
nor U4150 (N_4150,N_3256,N_2256);
nand U4151 (N_4151,N_3652,N_2391);
nand U4152 (N_4152,N_3274,N_3495);
or U4153 (N_4153,N_3750,N_3600);
and U4154 (N_4154,N_3699,N_3084);
nor U4155 (N_4155,N_3616,N_3387);
nor U4156 (N_4156,N_2773,N_3225);
or U4157 (N_4157,N_2798,N_3316);
or U4158 (N_4158,N_2842,N_2097);
and U4159 (N_4159,N_3555,N_3649);
nand U4160 (N_4160,N_2704,N_3946);
xnor U4161 (N_4161,N_3536,N_3351);
nand U4162 (N_4162,N_3293,N_2831);
and U4163 (N_4163,N_2730,N_2787);
nand U4164 (N_4164,N_2280,N_2137);
nor U4165 (N_4165,N_3005,N_3714);
and U4166 (N_4166,N_3866,N_2495);
nand U4167 (N_4167,N_3733,N_3502);
nand U4168 (N_4168,N_3889,N_2781);
xnor U4169 (N_4169,N_2891,N_2185);
and U4170 (N_4170,N_3769,N_2443);
xor U4171 (N_4171,N_2146,N_2870);
and U4172 (N_4172,N_3931,N_3111);
and U4173 (N_4173,N_3146,N_3916);
xnor U4174 (N_4174,N_2892,N_3857);
nand U4175 (N_4175,N_2272,N_3915);
and U4176 (N_4176,N_2050,N_3521);
nand U4177 (N_4177,N_3284,N_2260);
xnor U4178 (N_4178,N_2927,N_2829);
or U4179 (N_4179,N_2718,N_3409);
and U4180 (N_4180,N_3426,N_2094);
nor U4181 (N_4181,N_3149,N_3882);
or U4182 (N_4182,N_3034,N_2309);
nor U4183 (N_4183,N_3909,N_2543);
and U4184 (N_4184,N_3356,N_3924);
xor U4185 (N_4185,N_2472,N_3030);
and U4186 (N_4186,N_3335,N_2732);
nor U4187 (N_4187,N_2170,N_2298);
and U4188 (N_4188,N_2991,N_2572);
xnor U4189 (N_4189,N_3578,N_3990);
nor U4190 (N_4190,N_2308,N_2115);
nand U4191 (N_4191,N_3250,N_3673);
and U4192 (N_4192,N_3195,N_3055);
or U4193 (N_4193,N_3887,N_2877);
and U4194 (N_4194,N_3142,N_2425);
xor U4195 (N_4195,N_2001,N_2808);
nand U4196 (N_4196,N_2248,N_2455);
nor U4197 (N_4197,N_3804,N_3080);
xnor U4198 (N_4198,N_3132,N_3991);
or U4199 (N_4199,N_3265,N_3144);
nor U4200 (N_4200,N_3393,N_2741);
xnor U4201 (N_4201,N_3192,N_3936);
and U4202 (N_4202,N_2368,N_2794);
xor U4203 (N_4203,N_2731,N_3945);
and U4204 (N_4204,N_2811,N_3241);
nand U4205 (N_4205,N_2049,N_2596);
or U4206 (N_4206,N_2427,N_3223);
nand U4207 (N_4207,N_3545,N_2861);
and U4208 (N_4208,N_3243,N_2802);
nand U4209 (N_4209,N_2167,N_3709);
nor U4210 (N_4210,N_3302,N_3252);
nand U4211 (N_4211,N_2121,N_2337);
nor U4212 (N_4212,N_2760,N_3329);
xor U4213 (N_4213,N_3419,N_3105);
xor U4214 (N_4214,N_3281,N_2618);
or U4215 (N_4215,N_2895,N_3988);
and U4216 (N_4216,N_2836,N_3394);
or U4217 (N_4217,N_3150,N_3319);
and U4218 (N_4218,N_3523,N_2150);
and U4219 (N_4219,N_2478,N_3560);
nor U4220 (N_4220,N_3841,N_3418);
or U4221 (N_4221,N_2713,N_3443);
nand U4222 (N_4222,N_2064,N_3129);
and U4223 (N_4223,N_2463,N_3460);
xnor U4224 (N_4224,N_2519,N_2181);
and U4225 (N_4225,N_2267,N_3538);
and U4226 (N_4226,N_2683,N_2051);
xnor U4227 (N_4227,N_2746,N_2650);
nand U4228 (N_4228,N_3683,N_2127);
nand U4229 (N_4229,N_2555,N_2645);
or U4230 (N_4230,N_3196,N_2800);
xnor U4231 (N_4231,N_2666,N_3271);
or U4232 (N_4232,N_3212,N_3905);
and U4233 (N_4233,N_3786,N_2322);
nand U4234 (N_4234,N_3908,N_3290);
nor U4235 (N_4235,N_2193,N_3382);
xor U4236 (N_4236,N_3239,N_3904);
or U4237 (N_4237,N_3357,N_3728);
and U4238 (N_4238,N_3862,N_2747);
or U4239 (N_4239,N_2405,N_2415);
and U4240 (N_4240,N_3907,N_2481);
nand U4241 (N_4241,N_3547,N_2845);
xor U4242 (N_4242,N_2494,N_3655);
and U4243 (N_4243,N_3315,N_3874);
or U4244 (N_4244,N_3900,N_2627);
or U4245 (N_4245,N_2940,N_2446);
and U4246 (N_4246,N_3336,N_2816);
nand U4247 (N_4247,N_3462,N_3258);
and U4248 (N_4248,N_3014,N_2641);
xor U4249 (N_4249,N_2319,N_3978);
nor U4250 (N_4250,N_2303,N_2779);
nand U4251 (N_4251,N_3853,N_3955);
nor U4252 (N_4252,N_2854,N_3592);
xnor U4253 (N_4253,N_2725,N_3411);
nor U4254 (N_4254,N_2048,N_3434);
nand U4255 (N_4255,N_2331,N_2682);
xnor U4256 (N_4256,N_2970,N_3746);
xor U4257 (N_4257,N_3646,N_2801);
nor U4258 (N_4258,N_2905,N_3020);
xor U4259 (N_4259,N_3466,N_3603);
or U4260 (N_4260,N_3622,N_3135);
or U4261 (N_4261,N_3039,N_3287);
nand U4262 (N_4262,N_2982,N_2684);
xnor U4263 (N_4263,N_3940,N_2227);
or U4264 (N_4264,N_3249,N_3997);
nor U4265 (N_4265,N_2363,N_2912);
or U4266 (N_4266,N_3795,N_3137);
nor U4267 (N_4267,N_3399,N_3735);
xnor U4268 (N_4268,N_2301,N_3827);
nor U4269 (N_4269,N_2602,N_3333);
nand U4270 (N_4270,N_3618,N_3110);
and U4271 (N_4271,N_3108,N_3620);
or U4272 (N_4272,N_2705,N_3670);
and U4273 (N_4273,N_2975,N_3777);
nor U4274 (N_4274,N_2287,N_2710);
nand U4275 (N_4275,N_2515,N_3776);
or U4276 (N_4276,N_2659,N_2771);
nor U4277 (N_4277,N_2512,N_3169);
and U4278 (N_4278,N_3152,N_2130);
and U4279 (N_4279,N_2623,N_3605);
or U4280 (N_4280,N_2216,N_3497);
nand U4281 (N_4281,N_3681,N_2722);
nand U4282 (N_4282,N_3867,N_2390);
or U4283 (N_4283,N_2089,N_3100);
nor U4284 (N_4284,N_3970,N_3962);
or U4285 (N_4285,N_3575,N_2145);
and U4286 (N_4286,N_2903,N_2734);
nand U4287 (N_4287,N_3275,N_2657);
xor U4288 (N_4288,N_2407,N_3856);
nand U4289 (N_4289,N_2429,N_3760);
xor U4290 (N_4290,N_2202,N_3001);
or U4291 (N_4291,N_3595,N_2442);
xnor U4292 (N_4292,N_3677,N_2841);
and U4293 (N_4293,N_2597,N_2979);
nor U4294 (N_4294,N_2209,N_2857);
xor U4295 (N_4295,N_3793,N_2554);
or U4296 (N_4296,N_3552,N_3762);
nor U4297 (N_4297,N_3939,N_2133);
xnor U4298 (N_4298,N_2120,N_2325);
xor U4299 (N_4299,N_3203,N_2822);
nand U4300 (N_4300,N_3477,N_3698);
nand U4301 (N_4301,N_2062,N_2578);
nor U4302 (N_4302,N_3685,N_2464);
nor U4303 (N_4303,N_2985,N_3604);
nor U4304 (N_4304,N_2240,N_3773);
nor U4305 (N_4305,N_3063,N_2630);
xnor U4306 (N_4306,N_3019,N_2016);
or U4307 (N_4307,N_2817,N_2833);
and U4308 (N_4308,N_2592,N_2013);
nor U4309 (N_4309,N_2250,N_3972);
and U4310 (N_4310,N_3178,N_3774);
nor U4311 (N_4311,N_2693,N_2826);
nor U4312 (N_4312,N_3042,N_3864);
and U4313 (N_4313,N_3554,N_2503);
or U4314 (N_4314,N_2526,N_3808);
nor U4315 (N_4315,N_3840,N_3820);
xor U4316 (N_4316,N_2428,N_2606);
and U4317 (N_4317,N_3288,N_2204);
xnor U4318 (N_4318,N_2469,N_3345);
and U4319 (N_4319,N_3224,N_3496);
xnor U4320 (N_4320,N_3283,N_2974);
and U4321 (N_4321,N_3513,N_2232);
nand U4322 (N_4322,N_2351,N_2729);
or U4323 (N_4323,N_2739,N_3974);
and U4324 (N_4324,N_3352,N_3279);
xnor U4325 (N_4325,N_3753,N_3104);
xnor U4326 (N_4326,N_2507,N_2753);
xnor U4327 (N_4327,N_3453,N_3199);
xnor U4328 (N_4328,N_2647,N_2525);
xor U4329 (N_4329,N_3667,N_2186);
and U4330 (N_4330,N_2562,N_3749);
and U4331 (N_4331,N_3420,N_3317);
nand U4332 (N_4332,N_3074,N_2333);
xor U4333 (N_4333,N_3184,N_3614);
xor U4334 (N_4334,N_3175,N_3891);
nand U4335 (N_4335,N_2114,N_2493);
xor U4336 (N_4336,N_3067,N_2689);
and U4337 (N_4337,N_2457,N_3524);
nand U4338 (N_4338,N_2925,N_3482);
nand U4339 (N_4339,N_2989,N_2359);
or U4340 (N_4340,N_3233,N_2141);
nor U4341 (N_4341,N_2255,N_3587);
nand U4342 (N_4342,N_3151,N_3177);
nand U4343 (N_4343,N_3126,N_3682);
or U4344 (N_4344,N_2347,N_2103);
nor U4345 (N_4345,N_2003,N_2733);
or U4346 (N_4346,N_2797,N_2023);
nand U4347 (N_4347,N_3826,N_3396);
or U4348 (N_4348,N_3914,N_3678);
or U4349 (N_4349,N_2169,N_2153);
xnor U4350 (N_4350,N_2589,N_3610);
nor U4351 (N_4351,N_2714,N_2497);
and U4352 (N_4352,N_3011,N_3308);
or U4353 (N_4353,N_2586,N_2803);
or U4354 (N_4354,N_3201,N_2297);
xor U4355 (N_4355,N_3162,N_3445);
nor U4356 (N_4356,N_2514,N_3320);
nor U4357 (N_4357,N_2913,N_3326);
or U4358 (N_4358,N_3291,N_2653);
and U4359 (N_4359,N_3851,N_3478);
or U4360 (N_4360,N_3625,N_2965);
and U4361 (N_4361,N_2381,N_3579);
nor U4362 (N_4362,N_2483,N_3036);
nand U4363 (N_4363,N_2180,N_3799);
nor U4364 (N_4364,N_3929,N_2581);
and U4365 (N_4365,N_2971,N_3517);
nor U4366 (N_4366,N_3789,N_3860);
xor U4367 (N_4367,N_2539,N_2585);
nand U4368 (N_4368,N_3245,N_3428);
xnor U4369 (N_4369,N_2921,N_2864);
and U4370 (N_4370,N_3781,N_2228);
nand U4371 (N_4371,N_2548,N_3875);
and U4372 (N_4372,N_3363,N_2897);
xor U4373 (N_4373,N_2421,N_3696);
or U4374 (N_4374,N_2609,N_2068);
nand U4375 (N_4375,N_2302,N_2403);
or U4376 (N_4376,N_3529,N_3318);
or U4377 (N_4377,N_2941,N_3541);
nand U4378 (N_4378,N_2885,N_3675);
and U4379 (N_4379,N_2406,N_2691);
xnor U4380 (N_4380,N_3757,N_2943);
nand U4381 (N_4381,N_2299,N_3995);
and U4382 (N_4382,N_3367,N_3871);
or U4383 (N_4383,N_3879,N_2530);
xnor U4384 (N_4384,N_3650,N_3761);
nand U4385 (N_4385,N_2375,N_3221);
nand U4386 (N_4386,N_2192,N_2624);
and U4387 (N_4387,N_2101,N_3285);
and U4388 (N_4388,N_2819,N_3485);
xor U4389 (N_4389,N_2709,N_3558);
xnor U4390 (N_4390,N_3691,N_3327);
xor U4391 (N_4391,N_3641,N_2092);
nor U4392 (N_4392,N_3611,N_3818);
nor U4393 (N_4393,N_3627,N_2136);
nand U4394 (N_4394,N_3312,N_2587);
xor U4395 (N_4395,N_3492,N_2855);
xor U4396 (N_4396,N_2262,N_3313);
xor U4397 (N_4397,N_3046,N_2191);
xor U4398 (N_4398,N_2273,N_3648);
nand U4399 (N_4399,N_2551,N_3029);
and U4400 (N_4400,N_3133,N_2635);
nand U4401 (N_4401,N_3645,N_2310);
nor U4402 (N_4402,N_3948,N_3532);
and U4403 (N_4403,N_3912,N_3830);
and U4404 (N_4404,N_3082,N_2674);
nor U4405 (N_4405,N_2574,N_3404);
nand U4406 (N_4406,N_3027,N_2266);
and U4407 (N_4407,N_3324,N_3260);
or U4408 (N_4408,N_2340,N_2763);
nand U4409 (N_4409,N_2339,N_2707);
or U4410 (N_4410,N_2727,N_2764);
xnor U4411 (N_4411,N_3941,N_3885);
nor U4412 (N_4412,N_3896,N_2203);
nor U4413 (N_4413,N_3938,N_2588);
nand U4414 (N_4414,N_2922,N_3032);
or U4415 (N_4415,N_3906,N_2171);
xnor U4416 (N_4416,N_3788,N_2294);
or U4417 (N_4417,N_3076,N_3264);
and U4418 (N_4418,N_2523,N_2631);
and U4419 (N_4419,N_2499,N_2008);
nand U4420 (N_4420,N_3825,N_3154);
xor U4421 (N_4421,N_2106,N_2037);
xnor U4422 (N_4422,N_2977,N_2498);
or U4423 (N_4423,N_2004,N_3736);
nor U4424 (N_4424,N_2976,N_3395);
and U4425 (N_4425,N_3109,N_3819);
nor U4426 (N_4426,N_3415,N_3280);
or U4427 (N_4427,N_2118,N_2814);
and U4428 (N_4428,N_3388,N_3937);
or U4429 (N_4429,N_2663,N_2159);
or U4430 (N_4430,N_3494,N_2994);
or U4431 (N_4431,N_2221,N_3134);
xnor U4432 (N_4432,N_2924,N_3968);
nor U4433 (N_4433,N_3989,N_3525);
nand U4434 (N_4434,N_2416,N_3801);
nand U4435 (N_4435,N_3106,N_2901);
and U4436 (N_4436,N_2615,N_2656);
and U4437 (N_4437,N_3455,N_3689);
or U4438 (N_4438,N_2096,N_2465);
or U4439 (N_4439,N_3515,N_3176);
nor U4440 (N_4440,N_2057,N_2919);
nor U4441 (N_4441,N_2433,N_3607);
xor U4442 (N_4442,N_2239,N_3071);
nor U4443 (N_4443,N_2762,N_3573);
or U4444 (N_4444,N_2754,N_2583);
nor U4445 (N_4445,N_2284,N_3986);
nor U4446 (N_4446,N_2541,N_3672);
nand U4447 (N_4447,N_3922,N_2649);
xor U4448 (N_4448,N_3089,N_2371);
nor U4449 (N_4449,N_2876,N_3124);
xnor U4450 (N_4450,N_2550,N_3191);
or U4451 (N_4451,N_3222,N_2557);
nor U4452 (N_4452,N_2231,N_3858);
nor U4453 (N_4453,N_2521,N_3759);
nor U4454 (N_4454,N_3406,N_3328);
nor U4455 (N_4455,N_2026,N_3704);
nand U4456 (N_4456,N_2669,N_2091);
and U4457 (N_4457,N_2038,N_2690);
xor U4458 (N_4458,N_3261,N_3439);
xnor U4459 (N_4459,N_3961,N_2968);
nor U4460 (N_4460,N_3943,N_3118);
nand U4461 (N_4461,N_2395,N_2642);
or U4462 (N_4462,N_2422,N_3121);
or U4463 (N_4463,N_2198,N_3182);
nand U4464 (N_4464,N_2312,N_2074);
nand U4465 (N_4465,N_2571,N_2998);
or U4466 (N_4466,N_3379,N_2156);
xnor U4467 (N_4467,N_3364,N_2840);
nor U4468 (N_4468,N_2098,N_2423);
or U4469 (N_4469,N_2608,N_3967);
nor U4470 (N_4470,N_3694,N_3227);
xnor U4471 (N_4471,N_2501,N_3421);
nand U4472 (N_4472,N_2871,N_2522);
nor U4473 (N_4473,N_3559,N_3911);
nand U4474 (N_4474,N_2402,N_2009);
and U4475 (N_4475,N_3433,N_2275);
or U4476 (N_4476,N_2379,N_2129);
nor U4477 (N_4477,N_2950,N_2878);
nand U4478 (N_4478,N_3873,N_3966);
nor U4479 (N_4479,N_2565,N_3574);
xor U4480 (N_4480,N_2629,N_3520);
and U4481 (N_4481,N_3998,N_2818);
nand U4482 (N_4482,N_3633,N_2676);
xor U4483 (N_4483,N_2229,N_2175);
xor U4484 (N_4484,N_3519,N_3702);
nand U4485 (N_4485,N_3066,N_3307);
nand U4486 (N_4486,N_3701,N_2226);
or U4487 (N_4487,N_3952,N_3727);
and U4488 (N_4488,N_2807,N_3982);
and U4489 (N_4489,N_3490,N_3145);
and U4490 (N_4490,N_2658,N_3476);
and U4491 (N_4491,N_2426,N_2830);
nand U4492 (N_4492,N_2424,N_3719);
xor U4493 (N_4493,N_2697,N_3050);
nor U4494 (N_4494,N_2850,N_3796);
nor U4495 (N_4495,N_2780,N_3729);
nor U4496 (N_4496,N_3242,N_3669);
and U4497 (N_4497,N_3472,N_3637);
xnor U4498 (N_4498,N_2999,N_2007);
and U4499 (N_4499,N_2222,N_2626);
nand U4500 (N_4500,N_3706,N_3430);
nor U4501 (N_4501,N_2462,N_2983);
nand U4502 (N_4502,N_2451,N_3344);
nand U4503 (N_4503,N_3768,N_3951);
or U4504 (N_4504,N_3365,N_2617);
xor U4505 (N_4505,N_3965,N_3498);
and U4506 (N_4506,N_3930,N_3778);
nand U4507 (N_4507,N_3254,N_3392);
nor U4508 (N_4508,N_3653,N_3359);
xnor U4509 (N_4509,N_3743,N_3954);
or U4510 (N_4510,N_3236,N_3028);
xor U4511 (N_4511,N_2492,N_3016);
nor U4512 (N_4512,N_3289,N_2364);
or U4513 (N_4513,N_3128,N_2440);
nor U4514 (N_4514,N_2349,N_3892);
xor U4515 (N_4515,N_3872,N_3259);
nor U4516 (N_4516,N_3407,N_2584);
and U4517 (N_4517,N_3045,N_2058);
xnor U4518 (N_4518,N_3563,N_3859);
xor U4519 (N_4519,N_3048,N_2138);
nor U4520 (N_4520,N_2894,N_2930);
and U4521 (N_4521,N_2566,N_3174);
nor U4522 (N_4522,N_2104,N_3278);
nand U4523 (N_4523,N_2549,N_3985);
xor U4524 (N_4524,N_2564,N_2789);
or U4525 (N_4525,N_2963,N_2374);
and U4526 (N_4526,N_3435,N_2292);
or U4527 (N_4527,N_3155,N_2450);
and U4528 (N_4528,N_3052,N_3488);
nor U4529 (N_4529,N_3957,N_2117);
nor U4530 (N_4530,N_3210,N_3716);
or U4531 (N_4531,N_2010,N_3659);
nor U4532 (N_4532,N_2908,N_3635);
nand U4533 (N_4533,N_2553,N_3572);
xnor U4534 (N_4534,N_3441,N_3098);
nand U4535 (N_4535,N_3220,N_3131);
and U4536 (N_4536,N_3597,N_3267);
xor U4537 (N_4537,N_2664,N_2460);
or U4538 (N_4538,N_3585,N_2721);
and U4539 (N_4539,N_3479,N_2776);
xnor U4540 (N_4540,N_2929,N_2314);
nand U4541 (N_4541,N_2765,N_3540);
nor U4542 (N_4542,N_3722,N_2470);
nor U4543 (N_4543,N_2973,N_3272);
and U4544 (N_4544,N_2520,N_2577);
or U4545 (N_4545,N_2914,N_3507);
nor U4546 (N_4546,N_2540,N_3553);
nand U4547 (N_4547,N_3923,N_3286);
xor U4548 (N_4548,N_3615,N_2207);
or U4549 (N_4549,N_3339,N_2563);
or U4550 (N_4550,N_3979,N_3764);
nand U4551 (N_4551,N_3390,N_2155);
nor U4552 (N_4552,N_2208,N_2567);
nand U4553 (N_4553,N_3606,N_3205);
or U4554 (N_4554,N_2093,N_2821);
or U4555 (N_4555,N_3880,N_3878);
xnor U4556 (N_4556,N_2196,N_2654);
nand U4557 (N_4557,N_3787,N_2726);
and U4558 (N_4558,N_2218,N_3403);
nor U4559 (N_4559,N_3581,N_2034);
xnor U4560 (N_4560,N_3070,N_3211);
or U4561 (N_4561,N_2509,N_2157);
and U4562 (N_4562,N_3589,N_2916);
nand U4563 (N_4563,N_3977,N_3431);
nand U4564 (N_4564,N_2320,N_3765);
and U4565 (N_4565,N_2889,N_3602);
nor U4566 (N_4566,N_3202,N_3457);
nor U4567 (N_4567,N_2706,N_3903);
nor U4568 (N_4568,N_3628,N_3349);
xor U4569 (N_4569,N_2482,N_2392);
nor U4570 (N_4570,N_2069,N_3831);
xor U4571 (N_4571,N_3821,N_2703);
or U4572 (N_4572,N_2603,N_2362);
xor U4573 (N_4573,N_3999,N_2445);
nor U4574 (N_4574,N_2237,N_2933);
and U4575 (N_4575,N_2688,N_2786);
nand U4576 (N_4576,N_2917,N_3008);
or U4577 (N_4577,N_2513,N_3139);
nor U4578 (N_4578,N_2134,N_2178);
nor U4579 (N_4579,N_3734,N_3703);
and U4580 (N_4580,N_2568,N_3330);
and U4581 (N_4581,N_3876,N_2467);
and U4582 (N_4582,N_2162,N_2860);
or U4583 (N_4583,N_2350,N_3437);
xor U4584 (N_4584,N_3782,N_2477);
nor U4585 (N_4585,N_3463,N_2728);
xor U4586 (N_4586,N_3350,N_3097);
or U4587 (N_4587,N_3475,N_3078);
xnor U4588 (N_4588,N_2981,N_2573);
nor U4589 (N_4589,N_3362,N_3823);
and U4590 (N_4590,N_3094,N_3688);
nor U4591 (N_4591,N_2961,N_3665);
xor U4592 (N_4592,N_2453,N_2838);
and U4593 (N_4593,N_3456,N_3075);
xnor U4594 (N_4594,N_2902,N_2958);
nor U4595 (N_4595,N_3854,N_2002);
nand U4596 (N_4596,N_2006,N_3371);
xnor U4597 (N_4597,N_2151,N_2378);
nand U4598 (N_4598,N_2533,N_3717);
or U4599 (N_4599,N_2995,N_2386);
nand U4600 (N_4600,N_3775,N_3377);
and U4601 (N_4601,N_2217,N_3422);
and U4602 (N_4602,N_3721,N_3461);
nor U4603 (N_4603,N_2373,N_3546);
and U4604 (N_4604,N_2011,N_2893);
or U4605 (N_4605,N_3413,N_3624);
nor U4606 (N_4606,N_2154,N_2695);
xnor U4607 (N_4607,N_2686,N_3474);
or U4608 (N_4608,N_3634,N_3294);
or U4609 (N_4609,N_3163,N_2147);
and U4610 (N_4610,N_2084,N_3235);
xor U4611 (N_4611,N_3680,N_3528);
xnor U4612 (N_4612,N_3338,N_2767);
xnor U4613 (N_4613,N_2022,N_2761);
nand U4614 (N_4614,N_3006,N_2675);
nand U4615 (N_4615,N_3331,N_3755);
or U4616 (N_4616,N_2434,N_3031);
xnor U4617 (N_4617,N_2354,N_2698);
xor U4618 (N_4618,N_2173,N_3248);
xnor U4619 (N_4619,N_2243,N_2862);
nor U4620 (N_4620,N_3041,N_2435);
or U4621 (N_4621,N_2318,N_2040);
and U4622 (N_4622,N_2075,N_2947);
or U4623 (N_4623,N_2920,N_2397);
xor U4624 (N_4624,N_2738,N_3486);
nand U4625 (N_4625,N_3165,N_3797);
nor U4626 (N_4626,N_3499,N_2060);
and U4627 (N_4627,N_2648,N_2997);
and U4628 (N_4628,N_2139,N_3266);
and U4629 (N_4629,N_3888,N_3206);
or U4630 (N_4630,N_3469,N_2324);
xnor U4631 (N_4631,N_3173,N_3832);
or U4632 (N_4632,N_2082,N_3964);
or U4633 (N_4633,N_3565,N_3187);
xnor U4634 (N_4634,N_2570,N_3744);
and U4635 (N_4635,N_2188,N_2644);
and U4636 (N_4636,N_3189,N_2949);
and U4637 (N_4637,N_3798,N_3810);
xor U4638 (N_4638,N_3695,N_2041);
nand U4639 (N_4639,N_2601,N_2785);
and U4640 (N_4640,N_2788,N_2711);
xor U4641 (N_4641,N_3153,N_2490);
nand U4642 (N_4642,N_2907,N_2031);
nand U4643 (N_4643,N_2969,N_3270);
or U4644 (N_4644,N_3454,N_2201);
nor U4645 (N_4645,N_2890,N_2883);
or U4646 (N_4646,N_2694,N_3921);
and U4647 (N_4647,N_2843,N_2687);
nand U4648 (N_4648,N_2219,N_2254);
and U4649 (N_4649,N_2951,N_3158);
nor U4650 (N_4650,N_2899,N_3257);
and U4651 (N_4651,N_2054,N_3160);
and U4652 (N_4652,N_3660,N_2791);
or U4653 (N_4653,N_3425,N_2956);
and U4654 (N_4654,N_3022,N_3489);
and U4655 (N_4655,N_2278,N_2111);
or U4656 (N_4656,N_2679,N_2865);
nand U4657 (N_4657,N_3247,N_3380);
nor U4658 (N_4658,N_3920,N_3612);
or U4659 (N_4659,N_2419,N_2955);
and U4660 (N_4660,N_2622,N_3737);
or U4661 (N_4661,N_2620,N_3058);
and U4662 (N_4662,N_3549,N_3643);
xor U4663 (N_4663,N_3237,N_3800);
and U4664 (N_4664,N_3232,N_2105);
xnor U4665 (N_4665,N_3378,N_2305);
or U4666 (N_4666,N_3471,N_2685);
and U4667 (N_4667,N_2327,N_2056);
xnor U4668 (N_4668,N_3171,N_2500);
nor U4669 (N_4669,N_3863,N_3090);
xnor U4670 (N_4670,N_3663,N_3370);
nor U4671 (N_4671,N_3933,N_3447);
nand U4672 (N_4672,N_3065,N_3386);
nor U4673 (N_4673,N_3666,N_2431);
nand U4674 (N_4674,N_3346,N_2265);
xor U4675 (N_4675,N_2079,N_2122);
or U4676 (N_4676,N_3657,N_3570);
and U4677 (N_4677,N_2258,N_3059);
xnor U4678 (N_4678,N_2108,N_3310);
or U4679 (N_4679,N_3511,N_3229);
or U4680 (N_4680,N_2244,N_2852);
nor U4681 (N_4681,N_3298,N_3452);
nand U4682 (N_4682,N_2665,N_3238);
xor U4683 (N_4683,N_2382,N_3720);
and U4684 (N_4684,N_2087,N_2758);
or U4685 (N_4685,N_2000,N_2282);
xor U4686 (N_4686,N_2099,N_3987);
or U4687 (N_4687,N_2479,N_2909);
and U4688 (N_4688,N_3130,N_2027);
xor U4689 (N_4689,N_3282,N_3269);
xnor U4690 (N_4690,N_2915,N_3944);
or U4691 (N_4691,N_3292,N_2321);
nand U4692 (N_4692,N_3035,N_3004);
nor U4693 (N_4693,N_2165,N_3984);
nand U4694 (N_4694,N_3783,N_3459);
nand U4695 (N_4695,N_2772,N_3824);
nand U4696 (N_4696,N_3865,N_2367);
xnor U4697 (N_4697,N_3580,N_3372);
or U4698 (N_4698,N_2923,N_3758);
nand U4699 (N_4699,N_3481,N_3884);
nor U4700 (N_4700,N_2289,N_2061);
and U4701 (N_4701,N_3113,N_3530);
and U4702 (N_4702,N_2778,N_2307);
xor U4703 (N_4703,N_2931,N_3341);
nor U4704 (N_4704,N_3852,N_2535);
or U4705 (N_4705,N_2848,N_2660);
and U4706 (N_4706,N_3140,N_3503);
nor U4707 (N_4707,N_3446,N_3114);
nand U4708 (N_4708,N_3895,N_3391);
or U4709 (N_4709,N_2792,N_3375);
or U4710 (N_4710,N_3018,N_3043);
nand U4711 (N_4711,N_2610,N_3725);
and U4712 (N_4712,N_2430,N_3427);
nor U4713 (N_4713,N_2187,N_3534);
nand U4714 (N_4714,N_3166,N_2184);
or U4715 (N_4715,N_2723,N_3408);
nor U4716 (N_4716,N_2110,N_3009);
or U4717 (N_4717,N_2388,N_3568);
or U4718 (N_4718,N_2911,N_3073);
or U4719 (N_4719,N_2594,N_3299);
or U4720 (N_4720,N_2357,N_2444);
nand U4721 (N_4721,N_2640,N_2432);
and U4722 (N_4722,N_3608,N_3493);
and U4723 (N_4723,N_3103,N_2851);
xnor U4724 (N_4724,N_2088,N_2315);
nand U4725 (N_4725,N_3491,N_2055);
or U4726 (N_4726,N_2032,N_3548);
xnor U4727 (N_4727,N_2839,N_3062);
and U4728 (N_4728,N_3473,N_3510);
and U4729 (N_4729,N_3822,N_3183);
or U4730 (N_4730,N_3000,N_2783);
or U4731 (N_4731,N_3843,N_3167);
or U4732 (N_4732,N_2625,N_2928);
nand U4733 (N_4733,N_3845,N_2166);
nand U4734 (N_4734,N_2484,N_3518);
xor U4735 (N_4735,N_2045,N_2888);
nor U4736 (N_4736,N_2396,N_2487);
nand U4737 (N_4737,N_2449,N_2420);
nor U4738 (N_4738,N_2692,N_2311);
nor U4739 (N_4739,N_3590,N_3136);
nand U4740 (N_4740,N_3850,N_3180);
nor U4741 (N_4741,N_3739,N_2458);
nand U4742 (N_4742,N_3204,N_2859);
or U4743 (N_4743,N_2342,N_2412);
nand U4744 (N_4744,N_3583,N_2355);
nand U4745 (N_4745,N_2126,N_3772);
nand U4746 (N_4746,N_2591,N_2646);
xnor U4747 (N_4747,N_3710,N_3322);
and U4748 (N_4748,N_2067,N_2288);
nand U4749 (N_4749,N_3894,N_3122);
nand U4750 (N_4750,N_2556,N_2932);
nor U4751 (N_4751,N_3994,N_3686);
nor U4752 (N_4752,N_3651,N_2132);
nor U4753 (N_4753,N_3959,N_3809);
or U4754 (N_4754,N_3846,N_3244);
or U4755 (N_4755,N_3751,N_2176);
xor U4756 (N_4756,N_2740,N_2634);
or U4757 (N_4757,N_3842,N_2880);
or U4758 (N_4758,N_3432,N_2241);
and U4759 (N_4759,N_2281,N_2439);
xor U4760 (N_4760,N_2028,N_2158);
xnor U4761 (N_4761,N_3038,N_3869);
nand U4762 (N_4762,N_2719,N_3839);
nor U4763 (N_4763,N_2488,N_2993);
and U4764 (N_4764,N_3569,N_3101);
nand U4765 (N_4765,N_3219,N_3044);
or U4766 (N_4766,N_3092,N_3726);
nand U4767 (N_4767,N_2847,N_3069);
or U4768 (N_4768,N_3218,N_2102);
and U4769 (N_4769,N_2858,N_3053);
nand U4770 (N_4770,N_3397,N_3417);
nand U4771 (N_4771,N_2269,N_2225);
nand U4772 (N_4772,N_2715,N_2205);
nor U4773 (N_4773,N_3609,N_3487);
and U4774 (N_4774,N_2385,N_3763);
or U4775 (N_4775,N_2077,N_3465);
and U4776 (N_4776,N_2793,N_3332);
and U4777 (N_4777,N_3571,N_3700);
nor U4778 (N_4778,N_2394,N_2447);
xnor U4779 (N_4779,N_3847,N_2639);
and U4780 (N_4780,N_2095,N_2769);
or U4781 (N_4781,N_3713,N_3156);
nand U4782 (N_4782,N_2140,N_2174);
or U4783 (N_4783,N_2768,N_3301);
nand U4784 (N_4784,N_3617,N_3784);
or U4785 (N_4785,N_3263,N_3684);
nand U4786 (N_4786,N_3692,N_3013);
nor U4787 (N_4787,N_3806,N_2770);
and U4788 (N_4788,N_2569,N_2119);
nor U4789 (N_4789,N_2197,N_3890);
xor U4790 (N_4790,N_2164,N_3647);
or U4791 (N_4791,N_2200,N_3754);
nand U4792 (N_4792,N_2220,N_3591);
nor U4793 (N_4793,N_2612,N_2613);
and U4794 (N_4794,N_2867,N_3687);
nand U4795 (N_4795,N_2825,N_3868);
and U4796 (N_4796,N_2873,N_3188);
or U4797 (N_4797,N_2454,N_3088);
xnor U4798 (N_4798,N_3412,N_3707);
and U4799 (N_4799,N_3147,N_3566);
or U4800 (N_4800,N_2844,N_3658);
nor U4801 (N_4801,N_3325,N_2837);
nor U4802 (N_4802,N_3366,N_3848);
xnor U4803 (N_4803,N_2123,N_3779);
or U4804 (N_4804,N_3190,N_2766);
and U4805 (N_4805,N_2701,N_2085);
nand U4806 (N_4806,N_2475,N_2638);
or U4807 (N_4807,N_3040,N_2755);
nor U4808 (N_4808,N_2532,N_2143);
nor U4809 (N_4809,N_3116,N_2853);
xnor U4810 (N_4810,N_2906,N_2972);
and U4811 (N_4811,N_3026,N_2835);
nand U4812 (N_4812,N_3273,N_3992);
xor U4813 (N_4813,N_2508,N_2946);
nand U4814 (N_4814,N_2211,N_2619);
nand U4815 (N_4815,N_3304,N_2966);
nand U4816 (N_4816,N_2380,N_2486);
and U4817 (N_4817,N_3551,N_3323);
or U4818 (N_4818,N_3125,N_2053);
or U4819 (N_4819,N_2468,N_3679);
and U4820 (N_4820,N_3093,N_3021);
and U4821 (N_4821,N_2934,N_3504);
nor U4822 (N_4822,N_2670,N_2036);
or U4823 (N_4823,N_3662,N_3715);
or U4824 (N_4824,N_3588,N_2752);
or U4825 (N_4825,N_2012,N_2213);
nor U4826 (N_4826,N_3718,N_3664);
nor U4827 (N_4827,N_2538,N_3861);
xor U4828 (N_4828,N_3969,N_3373);
nand U4829 (N_4829,N_2952,N_3567);
nor U4830 (N_4830,N_2316,N_3881);
and U4831 (N_4831,N_3514,N_3811);
and U4832 (N_4832,N_3358,N_3429);
or U4833 (N_4833,N_2948,N_2516);
and U4834 (N_4834,N_2276,N_3838);
and U4835 (N_4835,N_3083,N_3436);
xnor U4836 (N_4836,N_2372,N_3193);
or U4837 (N_4837,N_3668,N_3342);
or U4838 (N_4838,N_3947,N_3470);
nand U4839 (N_4839,N_2559,N_3533);
nor U4840 (N_4840,N_3340,N_3629);
and U4841 (N_4841,N_2360,N_2076);
nor U4842 (N_4842,N_2304,N_2019);
or U4843 (N_4843,N_2206,N_2558);
xnor U4844 (N_4844,N_2529,N_2345);
or U4845 (N_4845,N_3369,N_2361);
and U4846 (N_4846,N_3790,N_2161);
xnor U4847 (N_4847,N_2268,N_3501);
nor U4848 (N_4848,N_2607,N_2604);
nor U4849 (N_4849,N_2329,N_2474);
nand U4850 (N_4850,N_2230,N_3910);
xnor U4851 (N_4851,N_2502,N_3376);
or U4852 (N_4852,N_2461,N_2090);
xor U4853 (N_4853,N_3927,N_2264);
nand U4854 (N_4854,N_3096,N_3584);
and U4855 (N_4855,N_3712,N_3732);
and U4856 (N_4856,N_3593,N_3928);
and U4857 (N_4857,N_3306,N_2812);
xor U4858 (N_4858,N_2466,N_2896);
nor U4859 (N_4859,N_3576,N_3047);
nor U4860 (N_4860,N_3010,N_3012);
xor U4861 (N_4861,N_2632,N_3913);
xor U4862 (N_4862,N_3661,N_2249);
xnor U4863 (N_4863,N_3942,N_3748);
nand U4864 (N_4864,N_3844,N_2939);
nor U4865 (N_4865,N_2506,N_2029);
and U4866 (N_4866,N_2485,N_2590);
or U4867 (N_4867,N_3949,N_3023);
xor U4868 (N_4868,N_3960,N_3505);
xor U4869 (N_4869,N_2834,N_2987);
xnor U4870 (N_4870,N_3410,N_3556);
and U4871 (N_4871,N_2757,N_2177);
nor U4872 (N_4872,N_3384,N_2346);
nand U4873 (N_4873,N_3117,N_2918);
nor U4874 (N_4874,N_2383,N_3334);
or U4875 (N_4875,N_2749,N_3277);
xnor U4876 (N_4876,N_3527,N_2194);
or U4877 (N_4877,N_3081,N_2279);
nor U4878 (N_4878,N_2480,N_3157);
xnor U4879 (N_4879,N_2805,N_3723);
xor U4880 (N_4880,N_3449,N_2809);
or U4881 (N_4881,N_3198,N_2910);
and U4882 (N_4882,N_3771,N_3381);
or U4883 (N_4883,N_3953,N_2677);
xnor U4884 (N_4884,N_3780,N_3483);
and U4885 (N_4885,N_2066,N_3812);
nor U4886 (N_4886,N_2823,N_3791);
and U4887 (N_4887,N_3355,N_2025);
xnor U4888 (N_4888,N_2988,N_2070);
or U4889 (N_4889,N_2868,N_3148);
or U4890 (N_4890,N_2436,N_3976);
or U4891 (N_4891,N_3813,N_2945);
and U4892 (N_4892,N_3506,N_3138);
xnor U4893 (N_4893,N_2116,N_2039);
nand U4894 (N_4894,N_2043,N_3017);
xnor U4895 (N_4895,N_2804,N_3626);
and U4896 (N_4896,N_2869,N_2341);
nor U4897 (N_4897,N_2135,N_2737);
nor U4898 (N_4898,N_3051,N_2404);
and U4899 (N_4899,N_3508,N_3509);
xnor U4900 (N_4900,N_2775,N_3002);
nand U4901 (N_4901,N_2437,N_2962);
xor U4902 (N_4902,N_2384,N_2408);
and U4903 (N_4903,N_3925,N_3542);
xnor U4904 (N_4904,N_3099,N_2100);
nand U4905 (N_4905,N_2128,N_2560);
nand U4906 (N_4906,N_3057,N_3917);
nor U4907 (N_4907,N_2886,N_2846);
xor U4908 (N_4908,N_2898,N_2748);
and U4909 (N_4909,N_3181,N_3539);
or U4910 (N_4910,N_3531,N_3033);
or U4911 (N_4911,N_3855,N_3314);
and U4912 (N_4912,N_3087,N_2296);
and U4913 (N_4913,N_2393,N_3214);
xor U4914 (N_4914,N_2598,N_2528);
xor U4915 (N_4915,N_3902,N_3815);
and U4916 (N_4916,N_2736,N_3268);
and U4917 (N_4917,N_2935,N_2035);
xor U4918 (N_4918,N_2168,N_2291);
or U4919 (N_4919,N_2813,N_2545);
and U4920 (N_4920,N_3234,N_3450);
or U4921 (N_4921,N_2992,N_3690);
xnor U4922 (N_4922,N_2018,N_3745);
nor U4923 (N_4923,N_3003,N_3956);
nand U4924 (N_4924,N_2046,N_3354);
nor U4925 (N_4925,N_2400,N_2672);
xnor U4926 (N_4926,N_3586,N_3400);
nor U4927 (N_4927,N_3785,N_2678);
nor U4928 (N_4928,N_3467,N_3794);
nor U4929 (N_4929,N_2954,N_2696);
nand U4930 (N_4930,N_2599,N_2937);
nor U4931 (N_4931,N_2605,N_2637);
xor U4932 (N_4932,N_2334,N_2234);
or U4933 (N_4933,N_2271,N_2247);
nor U4934 (N_4934,N_2131,N_2471);
and U4935 (N_4935,N_3932,N_3208);
nand U4936 (N_4936,N_3544,N_3091);
nor U4937 (N_4937,N_3276,N_2233);
and U4938 (N_4938,N_3102,N_3893);
nor U4939 (N_4939,N_2274,N_2815);
nand U4940 (N_4940,N_3297,N_2389);
and U4941 (N_4941,N_2348,N_2047);
and U4942 (N_4942,N_3353,N_3159);
nand U4943 (N_4943,N_3632,N_3642);
nand U4944 (N_4944,N_3079,N_2224);
nor U4945 (N_4945,N_2261,N_3926);
and U4946 (N_4946,N_3054,N_3255);
or U4947 (N_4947,N_3740,N_3440);
or U4948 (N_4948,N_2163,N_3837);
xor U4949 (N_4949,N_3389,N_3468);
and U4950 (N_4950,N_3594,N_2042);
nand U4951 (N_4951,N_2628,N_2790);
nor U4952 (N_4952,N_3348,N_2257);
nor U4953 (N_4953,N_2005,N_2473);
or U4954 (N_4954,N_2743,N_2456);
or U4955 (N_4955,N_3123,N_3442);
nor U4956 (N_4956,N_2313,N_2149);
nor U4957 (N_4957,N_3656,N_3343);
and U4958 (N_4958,N_2879,N_3792);
and U4959 (N_4959,N_3828,N_2544);
xor U4960 (N_4960,N_3170,N_2142);
xor U4961 (N_4961,N_2366,N_2651);
xor U4962 (N_4962,N_3711,N_2900);
nand U4963 (N_4963,N_3582,N_3980);
xnor U4964 (N_4964,N_2413,N_2086);
nor U4965 (N_4965,N_2252,N_3115);
and U4966 (N_4966,N_2330,N_2124);
nor U4967 (N_4967,N_2052,N_2107);
nor U4968 (N_4968,N_3347,N_2476);
nor U4969 (N_4969,N_3756,N_3630);
xnor U4970 (N_4970,N_2078,N_3766);
xor U4971 (N_4971,N_3537,N_2190);
nor U4972 (N_4972,N_2020,N_2376);
xor U4973 (N_4973,N_3401,N_2387);
xor U4974 (N_4974,N_3423,N_2759);
or U4975 (N_4975,N_3025,N_3886);
xor U4976 (N_4976,N_2518,N_2144);
nand U4977 (N_4977,N_3770,N_2081);
xnor U4978 (N_4978,N_2112,N_3919);
nor U4979 (N_4979,N_2251,N_3705);
and U4980 (N_4980,N_2527,N_2866);
and U4981 (N_4981,N_3368,N_3296);
nand U4982 (N_4982,N_3209,N_3829);
nor U4983 (N_4983,N_2661,N_3215);
nor U4984 (N_4984,N_2600,N_3161);
nand U4985 (N_4985,N_2160,N_3164);
or U4986 (N_4986,N_2849,N_2277);
nand U4987 (N_4987,N_2214,N_2926);
xor U4988 (N_4988,N_3817,N_3899);
xnor U4989 (N_4989,N_2774,N_3119);
nand U4990 (N_4990,N_2531,N_2742);
nor U4991 (N_4991,N_2699,N_3996);
or U4992 (N_4992,N_2750,N_2489);
or U4993 (N_4993,N_3262,N_2033);
and U4994 (N_4994,N_2517,N_2621);
xor U4995 (N_4995,N_2795,N_3217);
nor U4996 (N_4996,N_2796,N_2576);
and U4997 (N_4997,N_3654,N_2542);
xnor U4998 (N_4998,N_2152,N_2024);
nand U4999 (N_4999,N_2611,N_3636);
and U5000 (N_5000,N_2819,N_3085);
nand U5001 (N_5001,N_2402,N_2508);
and U5002 (N_5002,N_3686,N_2242);
and U5003 (N_5003,N_2858,N_3126);
and U5004 (N_5004,N_2670,N_3154);
or U5005 (N_5005,N_2362,N_3898);
nand U5006 (N_5006,N_2194,N_3996);
xnor U5007 (N_5007,N_2155,N_2847);
nand U5008 (N_5008,N_2412,N_2899);
xor U5009 (N_5009,N_2738,N_2426);
and U5010 (N_5010,N_3660,N_3450);
and U5011 (N_5011,N_2293,N_2201);
nand U5012 (N_5012,N_3271,N_3164);
nor U5013 (N_5013,N_3432,N_3005);
nand U5014 (N_5014,N_3791,N_2832);
or U5015 (N_5015,N_3109,N_3535);
xnor U5016 (N_5016,N_3227,N_3706);
xnor U5017 (N_5017,N_2212,N_3228);
and U5018 (N_5018,N_3478,N_3281);
xnor U5019 (N_5019,N_2734,N_3712);
nor U5020 (N_5020,N_2586,N_3738);
and U5021 (N_5021,N_2329,N_3221);
and U5022 (N_5022,N_3754,N_3208);
and U5023 (N_5023,N_3800,N_2155);
xor U5024 (N_5024,N_3584,N_3918);
and U5025 (N_5025,N_3813,N_3345);
xnor U5026 (N_5026,N_3971,N_2508);
nor U5027 (N_5027,N_2232,N_2705);
nand U5028 (N_5028,N_2704,N_2521);
or U5029 (N_5029,N_3575,N_3391);
and U5030 (N_5030,N_2386,N_3849);
and U5031 (N_5031,N_2233,N_3585);
or U5032 (N_5032,N_3211,N_3133);
and U5033 (N_5033,N_2516,N_2850);
xor U5034 (N_5034,N_2165,N_3134);
and U5035 (N_5035,N_2548,N_3067);
nor U5036 (N_5036,N_2969,N_2942);
and U5037 (N_5037,N_3369,N_2962);
xor U5038 (N_5038,N_2103,N_2224);
or U5039 (N_5039,N_2021,N_2507);
and U5040 (N_5040,N_2793,N_3888);
or U5041 (N_5041,N_2100,N_3938);
and U5042 (N_5042,N_3629,N_2348);
nand U5043 (N_5043,N_2541,N_2341);
or U5044 (N_5044,N_3652,N_2428);
and U5045 (N_5045,N_2902,N_2973);
nand U5046 (N_5046,N_2275,N_3413);
and U5047 (N_5047,N_2605,N_3154);
nand U5048 (N_5048,N_2794,N_3533);
xnor U5049 (N_5049,N_2888,N_2306);
nand U5050 (N_5050,N_2405,N_2851);
or U5051 (N_5051,N_3634,N_3366);
xnor U5052 (N_5052,N_2343,N_3028);
xnor U5053 (N_5053,N_3191,N_2972);
nand U5054 (N_5054,N_3741,N_3199);
xor U5055 (N_5055,N_2916,N_3152);
or U5056 (N_5056,N_2051,N_2940);
and U5057 (N_5057,N_2802,N_2338);
nand U5058 (N_5058,N_2505,N_3107);
nand U5059 (N_5059,N_3644,N_3649);
nand U5060 (N_5060,N_3388,N_3919);
and U5061 (N_5061,N_2597,N_3671);
nor U5062 (N_5062,N_2957,N_2096);
or U5063 (N_5063,N_2690,N_3943);
xor U5064 (N_5064,N_2290,N_2533);
or U5065 (N_5065,N_2938,N_2783);
nand U5066 (N_5066,N_3649,N_3533);
and U5067 (N_5067,N_3873,N_2518);
nor U5068 (N_5068,N_2760,N_3672);
xor U5069 (N_5069,N_3353,N_2640);
nand U5070 (N_5070,N_3635,N_3479);
or U5071 (N_5071,N_2736,N_2737);
xor U5072 (N_5072,N_3186,N_2117);
nand U5073 (N_5073,N_2266,N_3865);
or U5074 (N_5074,N_3672,N_3317);
xnor U5075 (N_5075,N_3222,N_2820);
and U5076 (N_5076,N_2248,N_2621);
nor U5077 (N_5077,N_2491,N_2604);
xor U5078 (N_5078,N_2692,N_2504);
or U5079 (N_5079,N_2615,N_2360);
nand U5080 (N_5080,N_3285,N_3048);
nand U5081 (N_5081,N_2039,N_2716);
or U5082 (N_5082,N_3946,N_3589);
nand U5083 (N_5083,N_3252,N_3638);
xor U5084 (N_5084,N_3384,N_2006);
or U5085 (N_5085,N_3475,N_2148);
and U5086 (N_5086,N_2031,N_2140);
or U5087 (N_5087,N_2609,N_2801);
and U5088 (N_5088,N_2328,N_3051);
xor U5089 (N_5089,N_3964,N_3663);
nand U5090 (N_5090,N_2421,N_3068);
and U5091 (N_5091,N_2299,N_3448);
nand U5092 (N_5092,N_2252,N_3274);
and U5093 (N_5093,N_2989,N_3898);
xnor U5094 (N_5094,N_2634,N_3980);
xor U5095 (N_5095,N_2978,N_3229);
and U5096 (N_5096,N_3383,N_3668);
xor U5097 (N_5097,N_3862,N_3350);
nand U5098 (N_5098,N_3149,N_2662);
nor U5099 (N_5099,N_3668,N_3976);
nor U5100 (N_5100,N_2109,N_2022);
and U5101 (N_5101,N_3398,N_3020);
nor U5102 (N_5102,N_2583,N_3333);
nand U5103 (N_5103,N_3129,N_2870);
or U5104 (N_5104,N_3335,N_3387);
and U5105 (N_5105,N_2841,N_3866);
nor U5106 (N_5106,N_2136,N_3973);
xnor U5107 (N_5107,N_2221,N_2152);
nor U5108 (N_5108,N_2991,N_2750);
and U5109 (N_5109,N_2743,N_2108);
and U5110 (N_5110,N_3185,N_2900);
xor U5111 (N_5111,N_2601,N_2937);
and U5112 (N_5112,N_2392,N_3892);
nand U5113 (N_5113,N_3389,N_2201);
or U5114 (N_5114,N_3910,N_3521);
nor U5115 (N_5115,N_2793,N_2105);
and U5116 (N_5116,N_3542,N_2463);
nor U5117 (N_5117,N_3297,N_3828);
and U5118 (N_5118,N_2530,N_2839);
nor U5119 (N_5119,N_3674,N_2817);
xnor U5120 (N_5120,N_2505,N_2945);
xnor U5121 (N_5121,N_3690,N_3741);
nor U5122 (N_5122,N_3668,N_2394);
or U5123 (N_5123,N_2381,N_2086);
nand U5124 (N_5124,N_3318,N_3569);
and U5125 (N_5125,N_2505,N_3724);
nor U5126 (N_5126,N_2113,N_3920);
or U5127 (N_5127,N_3918,N_2313);
xor U5128 (N_5128,N_3500,N_3228);
xor U5129 (N_5129,N_3834,N_3437);
nand U5130 (N_5130,N_2946,N_3383);
and U5131 (N_5131,N_2506,N_3666);
nor U5132 (N_5132,N_2682,N_2989);
xnor U5133 (N_5133,N_2622,N_2735);
nor U5134 (N_5134,N_3610,N_3291);
xor U5135 (N_5135,N_3814,N_2809);
or U5136 (N_5136,N_3943,N_3692);
and U5137 (N_5137,N_3755,N_3975);
and U5138 (N_5138,N_3936,N_2913);
or U5139 (N_5139,N_2788,N_2707);
xor U5140 (N_5140,N_2649,N_3262);
and U5141 (N_5141,N_3003,N_3350);
or U5142 (N_5142,N_3625,N_3033);
nor U5143 (N_5143,N_2526,N_2715);
nor U5144 (N_5144,N_2805,N_2178);
and U5145 (N_5145,N_2458,N_3999);
xnor U5146 (N_5146,N_3223,N_3183);
or U5147 (N_5147,N_2149,N_3238);
and U5148 (N_5148,N_2222,N_2299);
xor U5149 (N_5149,N_3615,N_3412);
and U5150 (N_5150,N_2717,N_3599);
and U5151 (N_5151,N_2011,N_2907);
xor U5152 (N_5152,N_2597,N_3208);
xor U5153 (N_5153,N_3931,N_2557);
nor U5154 (N_5154,N_2903,N_3973);
xor U5155 (N_5155,N_2849,N_3452);
and U5156 (N_5156,N_2998,N_3095);
nand U5157 (N_5157,N_3994,N_2735);
nand U5158 (N_5158,N_3725,N_3037);
or U5159 (N_5159,N_3457,N_2764);
and U5160 (N_5160,N_3336,N_2722);
nand U5161 (N_5161,N_3965,N_2811);
xnor U5162 (N_5162,N_2834,N_2138);
nor U5163 (N_5163,N_3270,N_2003);
xnor U5164 (N_5164,N_2282,N_3887);
xor U5165 (N_5165,N_3394,N_2013);
nand U5166 (N_5166,N_3169,N_2738);
nand U5167 (N_5167,N_2426,N_3732);
or U5168 (N_5168,N_2827,N_3727);
nor U5169 (N_5169,N_2331,N_3114);
nand U5170 (N_5170,N_3804,N_2762);
nor U5171 (N_5171,N_2211,N_2982);
and U5172 (N_5172,N_3346,N_2202);
nor U5173 (N_5173,N_3686,N_3990);
nor U5174 (N_5174,N_3419,N_2108);
xnor U5175 (N_5175,N_3712,N_2816);
nor U5176 (N_5176,N_2832,N_3446);
and U5177 (N_5177,N_3720,N_3257);
or U5178 (N_5178,N_3658,N_2786);
or U5179 (N_5179,N_3863,N_2694);
nor U5180 (N_5180,N_2730,N_2073);
and U5181 (N_5181,N_2580,N_2817);
nand U5182 (N_5182,N_2166,N_2735);
and U5183 (N_5183,N_3270,N_2992);
or U5184 (N_5184,N_2457,N_2080);
xnor U5185 (N_5185,N_2970,N_2651);
nand U5186 (N_5186,N_2945,N_2338);
nand U5187 (N_5187,N_2002,N_2412);
or U5188 (N_5188,N_3536,N_2596);
or U5189 (N_5189,N_2714,N_2264);
nand U5190 (N_5190,N_2635,N_3871);
xnor U5191 (N_5191,N_3317,N_3559);
and U5192 (N_5192,N_3235,N_2202);
nor U5193 (N_5193,N_3790,N_3409);
xor U5194 (N_5194,N_2409,N_2335);
and U5195 (N_5195,N_3033,N_3523);
xnor U5196 (N_5196,N_3771,N_3522);
xor U5197 (N_5197,N_3948,N_3588);
xnor U5198 (N_5198,N_2842,N_2599);
xor U5199 (N_5199,N_3427,N_3444);
and U5200 (N_5200,N_3793,N_2068);
nand U5201 (N_5201,N_2371,N_2637);
or U5202 (N_5202,N_3716,N_2320);
and U5203 (N_5203,N_3035,N_3085);
or U5204 (N_5204,N_3552,N_3153);
xnor U5205 (N_5205,N_3176,N_2350);
or U5206 (N_5206,N_3271,N_2234);
nand U5207 (N_5207,N_3200,N_2012);
xnor U5208 (N_5208,N_2178,N_2515);
or U5209 (N_5209,N_2209,N_2283);
nor U5210 (N_5210,N_2008,N_3620);
nor U5211 (N_5211,N_3085,N_2134);
nand U5212 (N_5212,N_2001,N_3533);
xnor U5213 (N_5213,N_3962,N_3039);
and U5214 (N_5214,N_3704,N_3224);
or U5215 (N_5215,N_2576,N_3299);
nand U5216 (N_5216,N_3394,N_2076);
nand U5217 (N_5217,N_2737,N_3281);
and U5218 (N_5218,N_3746,N_3409);
and U5219 (N_5219,N_2631,N_3874);
nor U5220 (N_5220,N_2850,N_3407);
nor U5221 (N_5221,N_3383,N_3667);
nor U5222 (N_5222,N_2883,N_2294);
nor U5223 (N_5223,N_2031,N_3497);
nand U5224 (N_5224,N_2625,N_3058);
and U5225 (N_5225,N_3722,N_2925);
and U5226 (N_5226,N_2887,N_3362);
or U5227 (N_5227,N_2518,N_3397);
and U5228 (N_5228,N_2900,N_3960);
xnor U5229 (N_5229,N_3386,N_3670);
nand U5230 (N_5230,N_3440,N_2204);
xor U5231 (N_5231,N_3151,N_2639);
nand U5232 (N_5232,N_2918,N_2058);
nor U5233 (N_5233,N_3342,N_3810);
or U5234 (N_5234,N_2461,N_3102);
and U5235 (N_5235,N_2870,N_3291);
xnor U5236 (N_5236,N_3238,N_2703);
nor U5237 (N_5237,N_2056,N_3042);
and U5238 (N_5238,N_2567,N_2083);
nand U5239 (N_5239,N_2552,N_3740);
nor U5240 (N_5240,N_3425,N_2924);
and U5241 (N_5241,N_3627,N_2960);
nor U5242 (N_5242,N_3655,N_2759);
and U5243 (N_5243,N_3356,N_2586);
nor U5244 (N_5244,N_2420,N_3506);
nand U5245 (N_5245,N_3955,N_3128);
xnor U5246 (N_5246,N_3978,N_3053);
or U5247 (N_5247,N_2869,N_2955);
xor U5248 (N_5248,N_3002,N_3069);
or U5249 (N_5249,N_2349,N_3839);
or U5250 (N_5250,N_2430,N_2406);
xor U5251 (N_5251,N_2229,N_3779);
nand U5252 (N_5252,N_2942,N_3650);
xor U5253 (N_5253,N_3162,N_2650);
and U5254 (N_5254,N_3817,N_2837);
xnor U5255 (N_5255,N_2213,N_2685);
nand U5256 (N_5256,N_2681,N_3640);
and U5257 (N_5257,N_2064,N_2337);
and U5258 (N_5258,N_3017,N_3324);
nand U5259 (N_5259,N_2175,N_3469);
and U5260 (N_5260,N_2475,N_3479);
or U5261 (N_5261,N_3669,N_2689);
and U5262 (N_5262,N_3939,N_2968);
nor U5263 (N_5263,N_2828,N_2221);
nand U5264 (N_5264,N_3709,N_3463);
nor U5265 (N_5265,N_2606,N_2297);
nor U5266 (N_5266,N_3696,N_2324);
or U5267 (N_5267,N_2045,N_2760);
xnor U5268 (N_5268,N_2519,N_2997);
nand U5269 (N_5269,N_2755,N_3904);
nor U5270 (N_5270,N_2928,N_3875);
xor U5271 (N_5271,N_2934,N_2025);
or U5272 (N_5272,N_3135,N_2558);
nor U5273 (N_5273,N_3428,N_3139);
xor U5274 (N_5274,N_3743,N_2891);
nor U5275 (N_5275,N_2737,N_3257);
and U5276 (N_5276,N_2504,N_3232);
or U5277 (N_5277,N_3403,N_3130);
xor U5278 (N_5278,N_3418,N_2731);
xnor U5279 (N_5279,N_3190,N_2937);
or U5280 (N_5280,N_2394,N_3125);
nor U5281 (N_5281,N_2941,N_3390);
xor U5282 (N_5282,N_3184,N_2240);
xor U5283 (N_5283,N_3918,N_2354);
xnor U5284 (N_5284,N_2179,N_3699);
nor U5285 (N_5285,N_3898,N_3049);
nand U5286 (N_5286,N_3072,N_2179);
or U5287 (N_5287,N_3639,N_3095);
nand U5288 (N_5288,N_3707,N_3744);
xor U5289 (N_5289,N_3034,N_2131);
nand U5290 (N_5290,N_2692,N_3529);
and U5291 (N_5291,N_3206,N_3155);
xnor U5292 (N_5292,N_2362,N_3529);
nand U5293 (N_5293,N_3397,N_2166);
and U5294 (N_5294,N_3693,N_3694);
or U5295 (N_5295,N_2948,N_2720);
or U5296 (N_5296,N_3089,N_3738);
nand U5297 (N_5297,N_3087,N_3673);
nor U5298 (N_5298,N_2917,N_3609);
xnor U5299 (N_5299,N_3213,N_2588);
nor U5300 (N_5300,N_3042,N_3456);
nand U5301 (N_5301,N_3069,N_3544);
nand U5302 (N_5302,N_2176,N_3190);
nand U5303 (N_5303,N_3876,N_2841);
xor U5304 (N_5304,N_2552,N_2233);
or U5305 (N_5305,N_2743,N_3681);
nor U5306 (N_5306,N_3065,N_3191);
or U5307 (N_5307,N_2609,N_2014);
and U5308 (N_5308,N_2407,N_3412);
nor U5309 (N_5309,N_3687,N_2789);
or U5310 (N_5310,N_2755,N_2100);
xor U5311 (N_5311,N_2046,N_2827);
nand U5312 (N_5312,N_3624,N_3139);
and U5313 (N_5313,N_3561,N_2706);
and U5314 (N_5314,N_3943,N_3463);
or U5315 (N_5315,N_3058,N_3377);
nor U5316 (N_5316,N_2697,N_3607);
nand U5317 (N_5317,N_3838,N_2696);
nor U5318 (N_5318,N_2210,N_2425);
or U5319 (N_5319,N_2408,N_3867);
nor U5320 (N_5320,N_3539,N_2732);
xor U5321 (N_5321,N_2930,N_3929);
or U5322 (N_5322,N_2891,N_2554);
xnor U5323 (N_5323,N_2935,N_2655);
or U5324 (N_5324,N_2330,N_2502);
nand U5325 (N_5325,N_3735,N_2375);
nor U5326 (N_5326,N_2245,N_2171);
nor U5327 (N_5327,N_3335,N_2151);
and U5328 (N_5328,N_3991,N_3859);
xnor U5329 (N_5329,N_3626,N_3045);
and U5330 (N_5330,N_3661,N_3148);
or U5331 (N_5331,N_2459,N_3397);
nor U5332 (N_5332,N_2668,N_3388);
xnor U5333 (N_5333,N_3982,N_3763);
or U5334 (N_5334,N_3235,N_2020);
xnor U5335 (N_5335,N_3347,N_2799);
and U5336 (N_5336,N_2463,N_3452);
nand U5337 (N_5337,N_2765,N_3413);
nor U5338 (N_5338,N_3164,N_3064);
and U5339 (N_5339,N_2599,N_3646);
and U5340 (N_5340,N_2674,N_2560);
nor U5341 (N_5341,N_3116,N_2537);
xor U5342 (N_5342,N_3560,N_2401);
xnor U5343 (N_5343,N_3677,N_3054);
or U5344 (N_5344,N_3186,N_3190);
nor U5345 (N_5345,N_2561,N_2919);
nand U5346 (N_5346,N_2984,N_3819);
xor U5347 (N_5347,N_3713,N_2582);
and U5348 (N_5348,N_2643,N_3123);
or U5349 (N_5349,N_2588,N_2698);
nor U5350 (N_5350,N_2875,N_3224);
nand U5351 (N_5351,N_2543,N_2547);
nand U5352 (N_5352,N_3195,N_3797);
xor U5353 (N_5353,N_3822,N_2327);
or U5354 (N_5354,N_2725,N_2994);
nand U5355 (N_5355,N_2459,N_2512);
nand U5356 (N_5356,N_2471,N_2623);
or U5357 (N_5357,N_3359,N_2293);
or U5358 (N_5358,N_2706,N_3584);
or U5359 (N_5359,N_3515,N_3386);
and U5360 (N_5360,N_2257,N_2551);
and U5361 (N_5361,N_3108,N_2140);
and U5362 (N_5362,N_3704,N_2080);
or U5363 (N_5363,N_2972,N_2832);
or U5364 (N_5364,N_2822,N_3706);
nand U5365 (N_5365,N_3580,N_2995);
xnor U5366 (N_5366,N_3622,N_3065);
or U5367 (N_5367,N_3470,N_2521);
and U5368 (N_5368,N_3595,N_3123);
nand U5369 (N_5369,N_2164,N_2440);
nor U5370 (N_5370,N_3015,N_3621);
and U5371 (N_5371,N_2730,N_3065);
xor U5372 (N_5372,N_2423,N_2507);
nor U5373 (N_5373,N_2268,N_2850);
or U5374 (N_5374,N_3388,N_2645);
or U5375 (N_5375,N_3779,N_3875);
nor U5376 (N_5376,N_3457,N_3589);
and U5377 (N_5377,N_3494,N_2013);
and U5378 (N_5378,N_2583,N_2483);
nand U5379 (N_5379,N_2252,N_3677);
xnor U5380 (N_5380,N_2395,N_2320);
nand U5381 (N_5381,N_2314,N_3934);
or U5382 (N_5382,N_2354,N_2133);
nor U5383 (N_5383,N_3174,N_3912);
nand U5384 (N_5384,N_2456,N_2527);
and U5385 (N_5385,N_2917,N_3412);
and U5386 (N_5386,N_2005,N_3087);
xnor U5387 (N_5387,N_3592,N_2967);
or U5388 (N_5388,N_2686,N_3630);
and U5389 (N_5389,N_3108,N_3151);
nand U5390 (N_5390,N_3400,N_3221);
or U5391 (N_5391,N_2053,N_2964);
and U5392 (N_5392,N_2506,N_2308);
nor U5393 (N_5393,N_3338,N_2814);
nand U5394 (N_5394,N_3342,N_2309);
and U5395 (N_5395,N_3640,N_2137);
nand U5396 (N_5396,N_3852,N_2525);
or U5397 (N_5397,N_2820,N_2815);
xor U5398 (N_5398,N_2124,N_2266);
xor U5399 (N_5399,N_2632,N_2243);
xnor U5400 (N_5400,N_3627,N_3908);
nor U5401 (N_5401,N_2980,N_2073);
nor U5402 (N_5402,N_2502,N_2483);
nand U5403 (N_5403,N_3414,N_2359);
xor U5404 (N_5404,N_2539,N_3483);
xnor U5405 (N_5405,N_3879,N_2830);
and U5406 (N_5406,N_3378,N_3904);
xor U5407 (N_5407,N_3685,N_2483);
nand U5408 (N_5408,N_3781,N_3065);
xnor U5409 (N_5409,N_2857,N_3267);
or U5410 (N_5410,N_3862,N_2853);
nand U5411 (N_5411,N_2440,N_3757);
xnor U5412 (N_5412,N_3783,N_2229);
nand U5413 (N_5413,N_3949,N_3634);
nor U5414 (N_5414,N_3072,N_2794);
nand U5415 (N_5415,N_3476,N_3413);
nand U5416 (N_5416,N_2159,N_2952);
nor U5417 (N_5417,N_2268,N_3033);
nand U5418 (N_5418,N_2376,N_3487);
nor U5419 (N_5419,N_3178,N_3200);
nand U5420 (N_5420,N_3722,N_2119);
and U5421 (N_5421,N_2599,N_2756);
or U5422 (N_5422,N_2711,N_3592);
nand U5423 (N_5423,N_2978,N_2875);
nor U5424 (N_5424,N_3764,N_2121);
and U5425 (N_5425,N_3906,N_3105);
nor U5426 (N_5426,N_3447,N_3446);
nand U5427 (N_5427,N_3755,N_2896);
xnor U5428 (N_5428,N_3100,N_3008);
nor U5429 (N_5429,N_2340,N_3619);
or U5430 (N_5430,N_3808,N_3313);
nand U5431 (N_5431,N_2500,N_3226);
and U5432 (N_5432,N_3182,N_2457);
nor U5433 (N_5433,N_3780,N_2612);
or U5434 (N_5434,N_2622,N_3523);
and U5435 (N_5435,N_3195,N_2244);
and U5436 (N_5436,N_3756,N_3547);
xnor U5437 (N_5437,N_2531,N_3171);
nand U5438 (N_5438,N_2422,N_2713);
and U5439 (N_5439,N_2848,N_3720);
nor U5440 (N_5440,N_3818,N_3514);
or U5441 (N_5441,N_3291,N_3289);
nand U5442 (N_5442,N_3155,N_2127);
and U5443 (N_5443,N_3751,N_3929);
xnor U5444 (N_5444,N_2759,N_2049);
nand U5445 (N_5445,N_3501,N_2036);
or U5446 (N_5446,N_3638,N_2314);
nand U5447 (N_5447,N_3024,N_3298);
nand U5448 (N_5448,N_3939,N_2547);
nand U5449 (N_5449,N_2079,N_2593);
or U5450 (N_5450,N_3226,N_3559);
and U5451 (N_5451,N_2034,N_3777);
nor U5452 (N_5452,N_3718,N_3703);
nand U5453 (N_5453,N_2194,N_2708);
or U5454 (N_5454,N_3076,N_3452);
nor U5455 (N_5455,N_3650,N_3448);
nand U5456 (N_5456,N_2911,N_3149);
xnor U5457 (N_5457,N_2903,N_2518);
nor U5458 (N_5458,N_3545,N_2625);
and U5459 (N_5459,N_2172,N_2674);
nor U5460 (N_5460,N_2990,N_3277);
or U5461 (N_5461,N_3849,N_3728);
nand U5462 (N_5462,N_2528,N_2514);
xor U5463 (N_5463,N_3878,N_2506);
and U5464 (N_5464,N_2180,N_2633);
and U5465 (N_5465,N_2510,N_3747);
and U5466 (N_5466,N_3042,N_2167);
nand U5467 (N_5467,N_2283,N_2500);
xor U5468 (N_5468,N_2302,N_3589);
nand U5469 (N_5469,N_3089,N_2186);
or U5470 (N_5470,N_2743,N_3060);
xor U5471 (N_5471,N_3618,N_3586);
nor U5472 (N_5472,N_3067,N_3926);
or U5473 (N_5473,N_2549,N_2867);
nand U5474 (N_5474,N_2788,N_3256);
xnor U5475 (N_5475,N_3158,N_2813);
or U5476 (N_5476,N_3793,N_3373);
nor U5477 (N_5477,N_2888,N_3004);
or U5478 (N_5478,N_2440,N_3701);
nand U5479 (N_5479,N_3262,N_3763);
or U5480 (N_5480,N_2656,N_2904);
or U5481 (N_5481,N_2554,N_2284);
nand U5482 (N_5482,N_3682,N_3948);
and U5483 (N_5483,N_2392,N_3497);
nand U5484 (N_5484,N_3848,N_2019);
xor U5485 (N_5485,N_2460,N_3706);
nand U5486 (N_5486,N_3407,N_3670);
and U5487 (N_5487,N_2744,N_3675);
and U5488 (N_5488,N_3059,N_2968);
xor U5489 (N_5489,N_2286,N_3559);
nor U5490 (N_5490,N_3529,N_2682);
nand U5491 (N_5491,N_3819,N_2853);
and U5492 (N_5492,N_2647,N_2940);
nor U5493 (N_5493,N_3067,N_3252);
nor U5494 (N_5494,N_3816,N_3185);
nand U5495 (N_5495,N_3785,N_2333);
xnor U5496 (N_5496,N_2924,N_2485);
or U5497 (N_5497,N_3946,N_2083);
nor U5498 (N_5498,N_3058,N_2052);
or U5499 (N_5499,N_2186,N_2281);
xnor U5500 (N_5500,N_2687,N_2482);
nor U5501 (N_5501,N_3760,N_3808);
and U5502 (N_5502,N_3069,N_2625);
nand U5503 (N_5503,N_3278,N_3486);
nand U5504 (N_5504,N_3093,N_2803);
or U5505 (N_5505,N_2238,N_2276);
nor U5506 (N_5506,N_3798,N_3347);
nor U5507 (N_5507,N_3589,N_3690);
and U5508 (N_5508,N_3744,N_3448);
or U5509 (N_5509,N_2059,N_2037);
or U5510 (N_5510,N_2755,N_2025);
nor U5511 (N_5511,N_2337,N_2916);
xnor U5512 (N_5512,N_3085,N_2440);
nand U5513 (N_5513,N_2343,N_3561);
and U5514 (N_5514,N_3722,N_2332);
or U5515 (N_5515,N_3061,N_3389);
nor U5516 (N_5516,N_2865,N_2109);
xnor U5517 (N_5517,N_2228,N_3150);
xor U5518 (N_5518,N_2138,N_3303);
nor U5519 (N_5519,N_3363,N_2238);
or U5520 (N_5520,N_3108,N_2037);
xor U5521 (N_5521,N_2317,N_2147);
nor U5522 (N_5522,N_3531,N_3070);
nand U5523 (N_5523,N_3537,N_2865);
and U5524 (N_5524,N_3590,N_3311);
nand U5525 (N_5525,N_3531,N_3123);
nand U5526 (N_5526,N_3553,N_3199);
and U5527 (N_5527,N_3562,N_3748);
nand U5528 (N_5528,N_3751,N_2272);
nor U5529 (N_5529,N_3631,N_2780);
and U5530 (N_5530,N_2687,N_3824);
or U5531 (N_5531,N_2710,N_2034);
nand U5532 (N_5532,N_2500,N_3253);
nor U5533 (N_5533,N_3521,N_3894);
xnor U5534 (N_5534,N_3808,N_2527);
nand U5535 (N_5535,N_2870,N_3124);
or U5536 (N_5536,N_2964,N_2680);
nand U5537 (N_5537,N_2561,N_2168);
xnor U5538 (N_5538,N_3982,N_2539);
xor U5539 (N_5539,N_3818,N_2082);
or U5540 (N_5540,N_2161,N_2953);
xor U5541 (N_5541,N_3948,N_2875);
nor U5542 (N_5542,N_3864,N_2453);
nor U5543 (N_5543,N_3123,N_3176);
xor U5544 (N_5544,N_2349,N_2296);
nor U5545 (N_5545,N_3616,N_3217);
or U5546 (N_5546,N_3791,N_3449);
nand U5547 (N_5547,N_2564,N_2201);
or U5548 (N_5548,N_3662,N_2045);
and U5549 (N_5549,N_2349,N_3166);
and U5550 (N_5550,N_2006,N_3536);
nand U5551 (N_5551,N_2815,N_3922);
nand U5552 (N_5552,N_2503,N_2096);
and U5553 (N_5553,N_3068,N_3367);
or U5554 (N_5554,N_2227,N_3982);
xor U5555 (N_5555,N_2495,N_3438);
nor U5556 (N_5556,N_2334,N_2675);
nor U5557 (N_5557,N_2102,N_2946);
nand U5558 (N_5558,N_3605,N_2389);
and U5559 (N_5559,N_3748,N_2798);
and U5560 (N_5560,N_3475,N_3670);
or U5561 (N_5561,N_3528,N_3571);
and U5562 (N_5562,N_2355,N_2308);
nand U5563 (N_5563,N_2656,N_3952);
xor U5564 (N_5564,N_2361,N_2868);
nor U5565 (N_5565,N_2743,N_3476);
xor U5566 (N_5566,N_3821,N_2194);
nor U5567 (N_5567,N_2824,N_3242);
xnor U5568 (N_5568,N_3818,N_3819);
nor U5569 (N_5569,N_3599,N_2963);
and U5570 (N_5570,N_3338,N_3754);
nand U5571 (N_5571,N_2547,N_3677);
or U5572 (N_5572,N_3143,N_3867);
or U5573 (N_5573,N_2430,N_2923);
xnor U5574 (N_5574,N_2185,N_3717);
nand U5575 (N_5575,N_3755,N_2839);
and U5576 (N_5576,N_3944,N_3456);
or U5577 (N_5577,N_2614,N_2435);
and U5578 (N_5578,N_3668,N_2576);
or U5579 (N_5579,N_2967,N_3862);
nand U5580 (N_5580,N_3476,N_3997);
xor U5581 (N_5581,N_2351,N_2851);
xor U5582 (N_5582,N_3999,N_2799);
or U5583 (N_5583,N_2664,N_3774);
nor U5584 (N_5584,N_2353,N_3312);
nor U5585 (N_5585,N_3694,N_3279);
nor U5586 (N_5586,N_2465,N_3729);
and U5587 (N_5587,N_2282,N_3572);
nor U5588 (N_5588,N_3607,N_3352);
or U5589 (N_5589,N_3332,N_2271);
or U5590 (N_5590,N_3170,N_3956);
nand U5591 (N_5591,N_2728,N_3244);
or U5592 (N_5592,N_3612,N_2892);
and U5593 (N_5593,N_2940,N_2869);
nand U5594 (N_5594,N_2358,N_3684);
xnor U5595 (N_5595,N_2599,N_2168);
xnor U5596 (N_5596,N_3641,N_2394);
nand U5597 (N_5597,N_2510,N_3578);
or U5598 (N_5598,N_3312,N_2485);
nor U5599 (N_5599,N_2296,N_3059);
nor U5600 (N_5600,N_2209,N_2680);
nor U5601 (N_5601,N_2188,N_3831);
nor U5602 (N_5602,N_2189,N_2030);
nand U5603 (N_5603,N_3466,N_2269);
nand U5604 (N_5604,N_2025,N_2843);
or U5605 (N_5605,N_2739,N_3936);
nand U5606 (N_5606,N_2897,N_3301);
nor U5607 (N_5607,N_2555,N_2139);
nand U5608 (N_5608,N_2455,N_3480);
and U5609 (N_5609,N_2259,N_2723);
or U5610 (N_5610,N_2870,N_3940);
xor U5611 (N_5611,N_3580,N_3776);
nand U5612 (N_5612,N_2119,N_2542);
xnor U5613 (N_5613,N_2816,N_3069);
xnor U5614 (N_5614,N_3740,N_3385);
xnor U5615 (N_5615,N_3041,N_3204);
nor U5616 (N_5616,N_3341,N_3153);
xnor U5617 (N_5617,N_3098,N_2430);
nor U5618 (N_5618,N_3814,N_2177);
xnor U5619 (N_5619,N_2358,N_3700);
nand U5620 (N_5620,N_3857,N_3163);
or U5621 (N_5621,N_2604,N_3198);
nand U5622 (N_5622,N_2458,N_3314);
nand U5623 (N_5623,N_3848,N_3709);
xnor U5624 (N_5624,N_2386,N_3062);
nor U5625 (N_5625,N_2663,N_2654);
and U5626 (N_5626,N_3951,N_3585);
or U5627 (N_5627,N_3976,N_3194);
and U5628 (N_5628,N_3340,N_2338);
nor U5629 (N_5629,N_2351,N_2520);
nand U5630 (N_5630,N_3541,N_2528);
and U5631 (N_5631,N_3310,N_2952);
xor U5632 (N_5632,N_3768,N_2164);
xor U5633 (N_5633,N_2865,N_2062);
nor U5634 (N_5634,N_2506,N_3614);
xnor U5635 (N_5635,N_3245,N_2018);
xnor U5636 (N_5636,N_3482,N_3124);
or U5637 (N_5637,N_3118,N_2582);
nand U5638 (N_5638,N_2373,N_3981);
nand U5639 (N_5639,N_3629,N_3294);
or U5640 (N_5640,N_3653,N_3422);
or U5641 (N_5641,N_3913,N_2855);
and U5642 (N_5642,N_2805,N_3135);
xor U5643 (N_5643,N_3970,N_3977);
or U5644 (N_5644,N_3537,N_3195);
nor U5645 (N_5645,N_2035,N_3941);
xnor U5646 (N_5646,N_2091,N_3151);
and U5647 (N_5647,N_3623,N_2598);
xor U5648 (N_5648,N_3648,N_2318);
xor U5649 (N_5649,N_3705,N_2878);
or U5650 (N_5650,N_3931,N_3986);
nor U5651 (N_5651,N_3641,N_3403);
or U5652 (N_5652,N_3996,N_2353);
or U5653 (N_5653,N_2517,N_2926);
nand U5654 (N_5654,N_3833,N_3585);
nand U5655 (N_5655,N_2153,N_3465);
xnor U5656 (N_5656,N_3618,N_2611);
nand U5657 (N_5657,N_2156,N_3278);
nand U5658 (N_5658,N_2405,N_2025);
or U5659 (N_5659,N_3884,N_3705);
nor U5660 (N_5660,N_3058,N_3466);
nor U5661 (N_5661,N_3666,N_3879);
and U5662 (N_5662,N_2534,N_3795);
xor U5663 (N_5663,N_2043,N_3934);
nand U5664 (N_5664,N_2180,N_3292);
or U5665 (N_5665,N_2497,N_2637);
nor U5666 (N_5666,N_2233,N_3769);
nand U5667 (N_5667,N_2047,N_2421);
nor U5668 (N_5668,N_3719,N_3769);
and U5669 (N_5669,N_3598,N_2004);
nor U5670 (N_5670,N_2334,N_3816);
and U5671 (N_5671,N_3549,N_3070);
xor U5672 (N_5672,N_2067,N_3481);
nand U5673 (N_5673,N_3242,N_3771);
or U5674 (N_5674,N_2804,N_2994);
xnor U5675 (N_5675,N_2491,N_2326);
nand U5676 (N_5676,N_2775,N_3298);
nand U5677 (N_5677,N_3459,N_2559);
xnor U5678 (N_5678,N_3894,N_2515);
nor U5679 (N_5679,N_3922,N_3666);
nor U5680 (N_5680,N_3672,N_2947);
and U5681 (N_5681,N_3691,N_3018);
nand U5682 (N_5682,N_2500,N_2134);
nor U5683 (N_5683,N_3854,N_2289);
nor U5684 (N_5684,N_3242,N_2456);
and U5685 (N_5685,N_2941,N_3419);
nand U5686 (N_5686,N_2727,N_2617);
or U5687 (N_5687,N_2945,N_2518);
nand U5688 (N_5688,N_3930,N_2012);
or U5689 (N_5689,N_3748,N_3194);
xnor U5690 (N_5690,N_3444,N_2848);
and U5691 (N_5691,N_3000,N_3559);
xor U5692 (N_5692,N_2053,N_2311);
nand U5693 (N_5693,N_2229,N_3709);
xor U5694 (N_5694,N_3563,N_2880);
nor U5695 (N_5695,N_3889,N_2813);
and U5696 (N_5696,N_3931,N_2548);
nand U5697 (N_5697,N_2422,N_3660);
nor U5698 (N_5698,N_3219,N_2751);
and U5699 (N_5699,N_3525,N_3810);
and U5700 (N_5700,N_3374,N_2085);
xnor U5701 (N_5701,N_3008,N_3459);
nor U5702 (N_5702,N_3368,N_3722);
and U5703 (N_5703,N_3445,N_3646);
and U5704 (N_5704,N_2174,N_3406);
nand U5705 (N_5705,N_2699,N_3900);
and U5706 (N_5706,N_2615,N_2364);
and U5707 (N_5707,N_3509,N_2765);
and U5708 (N_5708,N_3921,N_2545);
and U5709 (N_5709,N_2675,N_3359);
xor U5710 (N_5710,N_2625,N_2963);
and U5711 (N_5711,N_2540,N_2013);
xnor U5712 (N_5712,N_3936,N_3606);
or U5713 (N_5713,N_2215,N_3530);
nand U5714 (N_5714,N_3584,N_3953);
nand U5715 (N_5715,N_2111,N_2132);
nor U5716 (N_5716,N_2234,N_3460);
xor U5717 (N_5717,N_3909,N_2839);
nor U5718 (N_5718,N_3590,N_3125);
nand U5719 (N_5719,N_3352,N_3740);
or U5720 (N_5720,N_3702,N_3093);
nand U5721 (N_5721,N_3955,N_3343);
and U5722 (N_5722,N_3965,N_3842);
xnor U5723 (N_5723,N_2204,N_3448);
xor U5724 (N_5724,N_3632,N_2061);
or U5725 (N_5725,N_3280,N_2258);
nor U5726 (N_5726,N_3106,N_2604);
nand U5727 (N_5727,N_2909,N_2726);
nor U5728 (N_5728,N_3239,N_2668);
nand U5729 (N_5729,N_2896,N_3426);
nand U5730 (N_5730,N_2225,N_2506);
or U5731 (N_5731,N_3237,N_3941);
nand U5732 (N_5732,N_2104,N_3232);
nand U5733 (N_5733,N_2466,N_2012);
xor U5734 (N_5734,N_2285,N_3690);
and U5735 (N_5735,N_2034,N_2443);
or U5736 (N_5736,N_2903,N_2928);
nor U5737 (N_5737,N_2557,N_2388);
xor U5738 (N_5738,N_2498,N_3913);
nand U5739 (N_5739,N_3899,N_3364);
and U5740 (N_5740,N_2450,N_2518);
nand U5741 (N_5741,N_2174,N_2591);
and U5742 (N_5742,N_3289,N_2789);
nor U5743 (N_5743,N_2757,N_2639);
and U5744 (N_5744,N_2331,N_3977);
and U5745 (N_5745,N_2666,N_3957);
nor U5746 (N_5746,N_2777,N_3687);
xnor U5747 (N_5747,N_3605,N_2206);
nor U5748 (N_5748,N_2843,N_3411);
and U5749 (N_5749,N_3517,N_3919);
and U5750 (N_5750,N_3768,N_3475);
nor U5751 (N_5751,N_3132,N_3399);
and U5752 (N_5752,N_3242,N_2842);
xnor U5753 (N_5753,N_2347,N_2967);
or U5754 (N_5754,N_2069,N_3457);
nand U5755 (N_5755,N_2010,N_3533);
nand U5756 (N_5756,N_2871,N_3016);
xnor U5757 (N_5757,N_3803,N_2128);
and U5758 (N_5758,N_3836,N_3024);
nand U5759 (N_5759,N_2910,N_3731);
nor U5760 (N_5760,N_2195,N_2615);
nand U5761 (N_5761,N_3126,N_3849);
and U5762 (N_5762,N_2104,N_2469);
or U5763 (N_5763,N_2036,N_3932);
nand U5764 (N_5764,N_3766,N_3520);
and U5765 (N_5765,N_2642,N_3627);
and U5766 (N_5766,N_2841,N_2571);
nor U5767 (N_5767,N_2564,N_3720);
nand U5768 (N_5768,N_2479,N_3828);
nand U5769 (N_5769,N_2614,N_3347);
xnor U5770 (N_5770,N_2653,N_3067);
nor U5771 (N_5771,N_3482,N_3681);
xor U5772 (N_5772,N_3832,N_2496);
nand U5773 (N_5773,N_3577,N_3874);
xor U5774 (N_5774,N_2301,N_3797);
xor U5775 (N_5775,N_3484,N_2710);
xnor U5776 (N_5776,N_2583,N_2342);
and U5777 (N_5777,N_2348,N_3915);
nor U5778 (N_5778,N_3599,N_2419);
and U5779 (N_5779,N_2817,N_2322);
xnor U5780 (N_5780,N_3497,N_2925);
nor U5781 (N_5781,N_3309,N_3947);
xnor U5782 (N_5782,N_2043,N_2800);
nor U5783 (N_5783,N_2394,N_3846);
xor U5784 (N_5784,N_3359,N_3846);
nand U5785 (N_5785,N_3172,N_3787);
or U5786 (N_5786,N_2855,N_3571);
or U5787 (N_5787,N_2111,N_2956);
and U5788 (N_5788,N_2325,N_3676);
nand U5789 (N_5789,N_2123,N_3291);
or U5790 (N_5790,N_2402,N_3371);
nand U5791 (N_5791,N_2492,N_2446);
nor U5792 (N_5792,N_3186,N_3689);
nand U5793 (N_5793,N_3397,N_2825);
xor U5794 (N_5794,N_3567,N_3791);
or U5795 (N_5795,N_2327,N_2293);
nor U5796 (N_5796,N_3140,N_2749);
and U5797 (N_5797,N_2699,N_3088);
nand U5798 (N_5798,N_2762,N_2307);
nand U5799 (N_5799,N_2332,N_2152);
nand U5800 (N_5800,N_2586,N_3593);
nand U5801 (N_5801,N_3057,N_3032);
and U5802 (N_5802,N_2117,N_2340);
and U5803 (N_5803,N_3516,N_3786);
nand U5804 (N_5804,N_2054,N_3433);
nand U5805 (N_5805,N_2120,N_3323);
nand U5806 (N_5806,N_3936,N_3643);
nor U5807 (N_5807,N_2299,N_2803);
xnor U5808 (N_5808,N_2035,N_3617);
or U5809 (N_5809,N_2561,N_3240);
xnor U5810 (N_5810,N_2785,N_2935);
and U5811 (N_5811,N_2755,N_2122);
and U5812 (N_5812,N_2442,N_2896);
xor U5813 (N_5813,N_2575,N_2646);
nand U5814 (N_5814,N_2683,N_3044);
or U5815 (N_5815,N_2182,N_2890);
and U5816 (N_5816,N_2611,N_3264);
xnor U5817 (N_5817,N_2165,N_2390);
nand U5818 (N_5818,N_3691,N_3326);
nor U5819 (N_5819,N_2529,N_2123);
or U5820 (N_5820,N_2746,N_2908);
and U5821 (N_5821,N_2038,N_2443);
or U5822 (N_5822,N_3776,N_3459);
and U5823 (N_5823,N_2526,N_3754);
nor U5824 (N_5824,N_2607,N_2853);
nor U5825 (N_5825,N_2133,N_3047);
or U5826 (N_5826,N_3702,N_3349);
and U5827 (N_5827,N_2605,N_2747);
nand U5828 (N_5828,N_3676,N_2215);
and U5829 (N_5829,N_3577,N_2598);
nor U5830 (N_5830,N_3580,N_2371);
or U5831 (N_5831,N_2962,N_2031);
nand U5832 (N_5832,N_2937,N_2508);
nand U5833 (N_5833,N_3564,N_3949);
and U5834 (N_5834,N_3940,N_2909);
xnor U5835 (N_5835,N_2435,N_3684);
and U5836 (N_5836,N_2623,N_2089);
or U5837 (N_5837,N_2969,N_2348);
or U5838 (N_5838,N_3774,N_2677);
and U5839 (N_5839,N_2045,N_3798);
nand U5840 (N_5840,N_2294,N_3489);
and U5841 (N_5841,N_2515,N_3855);
xnor U5842 (N_5842,N_2253,N_2159);
or U5843 (N_5843,N_2444,N_2858);
nor U5844 (N_5844,N_2826,N_3163);
nand U5845 (N_5845,N_2942,N_2043);
xor U5846 (N_5846,N_2282,N_3307);
nand U5847 (N_5847,N_2413,N_3026);
xnor U5848 (N_5848,N_3462,N_3668);
nand U5849 (N_5849,N_2352,N_3795);
and U5850 (N_5850,N_2092,N_3660);
nor U5851 (N_5851,N_3316,N_2047);
or U5852 (N_5852,N_2441,N_2443);
nand U5853 (N_5853,N_2474,N_3642);
nor U5854 (N_5854,N_2489,N_3458);
or U5855 (N_5855,N_3384,N_2642);
nand U5856 (N_5856,N_3735,N_3859);
nor U5857 (N_5857,N_3024,N_3831);
nand U5858 (N_5858,N_3643,N_3294);
or U5859 (N_5859,N_2164,N_2101);
nor U5860 (N_5860,N_3456,N_2588);
or U5861 (N_5861,N_3591,N_2194);
or U5862 (N_5862,N_2505,N_2877);
and U5863 (N_5863,N_3334,N_3399);
nor U5864 (N_5864,N_3015,N_3363);
xor U5865 (N_5865,N_2068,N_3962);
nand U5866 (N_5866,N_3276,N_3922);
nor U5867 (N_5867,N_2396,N_2507);
xnor U5868 (N_5868,N_3534,N_2702);
xor U5869 (N_5869,N_2788,N_2305);
or U5870 (N_5870,N_2002,N_3491);
nor U5871 (N_5871,N_3450,N_3970);
xor U5872 (N_5872,N_2006,N_3310);
nor U5873 (N_5873,N_2696,N_2876);
and U5874 (N_5874,N_3843,N_2712);
and U5875 (N_5875,N_2957,N_3581);
nand U5876 (N_5876,N_3206,N_3185);
and U5877 (N_5877,N_2412,N_3817);
or U5878 (N_5878,N_2715,N_2153);
and U5879 (N_5879,N_3981,N_2912);
nor U5880 (N_5880,N_2940,N_2872);
xor U5881 (N_5881,N_2308,N_3523);
and U5882 (N_5882,N_3325,N_3665);
nand U5883 (N_5883,N_2936,N_3167);
nand U5884 (N_5884,N_2478,N_2441);
nor U5885 (N_5885,N_2683,N_2681);
xor U5886 (N_5886,N_2736,N_3137);
nand U5887 (N_5887,N_3493,N_2923);
nand U5888 (N_5888,N_2458,N_2298);
or U5889 (N_5889,N_3389,N_3208);
or U5890 (N_5890,N_3818,N_3281);
and U5891 (N_5891,N_3036,N_3756);
nor U5892 (N_5892,N_2376,N_3709);
or U5893 (N_5893,N_2182,N_3170);
nor U5894 (N_5894,N_3614,N_2461);
nand U5895 (N_5895,N_3957,N_3999);
xor U5896 (N_5896,N_3756,N_2253);
and U5897 (N_5897,N_3663,N_2928);
and U5898 (N_5898,N_3380,N_3720);
and U5899 (N_5899,N_2369,N_2581);
and U5900 (N_5900,N_2996,N_2463);
and U5901 (N_5901,N_3603,N_3476);
or U5902 (N_5902,N_3754,N_2303);
and U5903 (N_5903,N_2853,N_3598);
xor U5904 (N_5904,N_3921,N_2567);
nor U5905 (N_5905,N_2912,N_2750);
nand U5906 (N_5906,N_2468,N_2764);
xor U5907 (N_5907,N_2842,N_2147);
or U5908 (N_5908,N_2339,N_3789);
or U5909 (N_5909,N_3528,N_2177);
nor U5910 (N_5910,N_3118,N_3662);
nand U5911 (N_5911,N_2557,N_2491);
nand U5912 (N_5912,N_3171,N_3713);
and U5913 (N_5913,N_3242,N_2835);
nand U5914 (N_5914,N_2419,N_2358);
nand U5915 (N_5915,N_3936,N_2166);
xor U5916 (N_5916,N_3910,N_3192);
and U5917 (N_5917,N_3558,N_3498);
and U5918 (N_5918,N_2386,N_3842);
xnor U5919 (N_5919,N_2689,N_2902);
nand U5920 (N_5920,N_2707,N_3651);
or U5921 (N_5921,N_2773,N_3307);
nand U5922 (N_5922,N_2381,N_3012);
xor U5923 (N_5923,N_3160,N_2185);
or U5924 (N_5924,N_3825,N_2489);
nor U5925 (N_5925,N_2961,N_3040);
nand U5926 (N_5926,N_2254,N_3697);
or U5927 (N_5927,N_2724,N_3730);
xor U5928 (N_5928,N_2227,N_2236);
and U5929 (N_5929,N_3441,N_2376);
nand U5930 (N_5930,N_3229,N_3681);
and U5931 (N_5931,N_3748,N_3056);
and U5932 (N_5932,N_2799,N_2305);
nor U5933 (N_5933,N_2723,N_2999);
nor U5934 (N_5934,N_3260,N_3614);
nand U5935 (N_5935,N_2592,N_3751);
nor U5936 (N_5936,N_3454,N_3954);
xor U5937 (N_5937,N_3548,N_2404);
nand U5938 (N_5938,N_2746,N_3641);
and U5939 (N_5939,N_2919,N_2278);
nor U5940 (N_5940,N_3215,N_3922);
or U5941 (N_5941,N_2962,N_2647);
xnor U5942 (N_5942,N_2351,N_3541);
or U5943 (N_5943,N_2698,N_3766);
xnor U5944 (N_5944,N_3084,N_2456);
nor U5945 (N_5945,N_3368,N_2867);
and U5946 (N_5946,N_2460,N_2407);
or U5947 (N_5947,N_2897,N_3681);
and U5948 (N_5948,N_2640,N_3952);
nand U5949 (N_5949,N_3851,N_3675);
nor U5950 (N_5950,N_3216,N_2987);
and U5951 (N_5951,N_3998,N_3652);
and U5952 (N_5952,N_2701,N_2808);
xor U5953 (N_5953,N_2878,N_3206);
nand U5954 (N_5954,N_3935,N_3345);
or U5955 (N_5955,N_2872,N_2471);
nand U5956 (N_5956,N_2145,N_2462);
nor U5957 (N_5957,N_3355,N_2782);
and U5958 (N_5958,N_3345,N_3471);
xnor U5959 (N_5959,N_2832,N_3305);
nand U5960 (N_5960,N_2051,N_3569);
nor U5961 (N_5961,N_3600,N_2808);
or U5962 (N_5962,N_2697,N_2304);
or U5963 (N_5963,N_3166,N_2867);
and U5964 (N_5964,N_3633,N_3853);
xor U5965 (N_5965,N_3830,N_2489);
and U5966 (N_5966,N_2215,N_2587);
and U5967 (N_5967,N_3844,N_2370);
and U5968 (N_5968,N_2321,N_2426);
xor U5969 (N_5969,N_2263,N_2500);
nand U5970 (N_5970,N_2748,N_3164);
nand U5971 (N_5971,N_3299,N_2932);
and U5972 (N_5972,N_2360,N_3455);
or U5973 (N_5973,N_3040,N_3898);
or U5974 (N_5974,N_3165,N_3624);
or U5975 (N_5975,N_3741,N_2255);
and U5976 (N_5976,N_3969,N_2972);
xnor U5977 (N_5977,N_3284,N_2604);
and U5978 (N_5978,N_2117,N_3989);
or U5979 (N_5979,N_3489,N_3972);
xnor U5980 (N_5980,N_2589,N_3129);
xnor U5981 (N_5981,N_3533,N_2528);
nand U5982 (N_5982,N_3888,N_2319);
nand U5983 (N_5983,N_3035,N_2128);
nand U5984 (N_5984,N_2406,N_2380);
and U5985 (N_5985,N_2262,N_2427);
xor U5986 (N_5986,N_3496,N_3695);
and U5987 (N_5987,N_3019,N_2476);
xnor U5988 (N_5988,N_3507,N_3224);
xor U5989 (N_5989,N_2387,N_3732);
and U5990 (N_5990,N_3912,N_3837);
or U5991 (N_5991,N_3003,N_3075);
and U5992 (N_5992,N_2398,N_2708);
nor U5993 (N_5993,N_2923,N_2006);
or U5994 (N_5994,N_2347,N_3416);
and U5995 (N_5995,N_3347,N_2202);
and U5996 (N_5996,N_3663,N_3725);
or U5997 (N_5997,N_2791,N_3174);
nand U5998 (N_5998,N_3244,N_3759);
and U5999 (N_5999,N_3930,N_2945);
nand U6000 (N_6000,N_5296,N_4869);
or U6001 (N_6001,N_4667,N_5090);
nor U6002 (N_6002,N_4463,N_5882);
xnor U6003 (N_6003,N_5747,N_5202);
xor U6004 (N_6004,N_4118,N_5052);
or U6005 (N_6005,N_5042,N_4474);
and U6006 (N_6006,N_5932,N_5158);
xor U6007 (N_6007,N_5150,N_4498);
xnor U6008 (N_6008,N_4351,N_4984);
and U6009 (N_6009,N_5390,N_5737);
nand U6010 (N_6010,N_5652,N_5573);
nand U6011 (N_6011,N_5071,N_4049);
xnor U6012 (N_6012,N_4072,N_5358);
nor U6013 (N_6013,N_4142,N_4662);
nor U6014 (N_6014,N_4507,N_4535);
or U6015 (N_6015,N_4178,N_4727);
and U6016 (N_6016,N_4942,N_5783);
nor U6017 (N_6017,N_5845,N_4516);
or U6018 (N_6018,N_4374,N_5587);
xor U6019 (N_6019,N_4785,N_5899);
or U6020 (N_6020,N_4966,N_5876);
and U6021 (N_6021,N_5036,N_5033);
xnor U6022 (N_6022,N_4290,N_4429);
nand U6023 (N_6023,N_4513,N_4488);
nor U6024 (N_6024,N_4581,N_5471);
or U6025 (N_6025,N_5588,N_5641);
xor U6026 (N_6026,N_4519,N_5104);
nor U6027 (N_6027,N_5890,N_5482);
nand U6028 (N_6028,N_5487,N_4553);
nor U6029 (N_6029,N_4313,N_5211);
or U6030 (N_6030,N_5132,N_5732);
or U6031 (N_6031,N_4578,N_4679);
nor U6032 (N_6032,N_5782,N_5653);
and U6033 (N_6033,N_4393,N_5142);
nand U6034 (N_6034,N_4524,N_4823);
nand U6035 (N_6035,N_4509,N_5752);
nor U6036 (N_6036,N_5962,N_4273);
and U6037 (N_6037,N_5107,N_4872);
and U6038 (N_6038,N_5921,N_5183);
nand U6039 (N_6039,N_5746,N_4166);
xnor U6040 (N_6040,N_4717,N_5222);
nand U6041 (N_6041,N_5669,N_4639);
nand U6042 (N_6042,N_4892,N_4494);
or U6043 (N_6043,N_5209,N_5383);
and U6044 (N_6044,N_4218,N_4078);
nand U6045 (N_6045,N_5713,N_4226);
nand U6046 (N_6046,N_4833,N_5688);
or U6047 (N_6047,N_4499,N_4962);
and U6048 (N_6048,N_4480,N_5235);
and U6049 (N_6049,N_4903,N_5902);
xor U6050 (N_6050,N_4796,N_4481);
nor U6051 (N_6051,N_4599,N_5738);
or U6052 (N_6052,N_5528,N_4769);
or U6053 (N_6053,N_5494,N_5371);
and U6054 (N_6054,N_5024,N_4885);
and U6055 (N_6055,N_4155,N_5099);
nand U6056 (N_6056,N_4681,N_4501);
nand U6057 (N_6057,N_5015,N_4134);
or U6058 (N_6058,N_5268,N_4771);
and U6059 (N_6059,N_5165,N_4666);
or U6060 (N_6060,N_5595,N_4337);
nand U6061 (N_6061,N_4468,N_4238);
nor U6062 (N_6062,N_4661,N_4839);
xor U6063 (N_6063,N_5361,N_4087);
nor U6064 (N_6064,N_5365,N_5013);
xnor U6065 (N_6065,N_5097,N_5056);
nand U6066 (N_6066,N_5629,N_5239);
nor U6067 (N_6067,N_4389,N_5378);
nand U6068 (N_6068,N_5335,N_5016);
nor U6069 (N_6069,N_5830,N_4412);
nor U6070 (N_6070,N_4598,N_5352);
xnor U6071 (N_6071,N_4728,N_4128);
nand U6072 (N_6072,N_4850,N_5523);
xnor U6073 (N_6073,N_4467,N_5149);
nor U6074 (N_6074,N_5906,N_4704);
nor U6075 (N_6075,N_5866,N_4930);
nand U6076 (N_6076,N_4622,N_4212);
and U6077 (N_6077,N_5460,N_4675);
xor U6078 (N_6078,N_5708,N_4164);
and U6079 (N_6079,N_5127,N_4398);
xnor U6080 (N_6080,N_5977,N_4815);
nor U6081 (N_6081,N_5578,N_5644);
nand U6082 (N_6082,N_4712,N_4986);
and U6083 (N_6083,N_4109,N_5778);
nor U6084 (N_6084,N_5497,N_5492);
nor U6085 (N_6085,N_5401,N_4009);
or U6086 (N_6086,N_4898,N_4431);
nor U6087 (N_6087,N_5615,N_5186);
and U6088 (N_6088,N_5008,N_5260);
nor U6089 (N_6089,N_5425,N_5468);
and U6090 (N_6090,N_5685,N_5740);
and U6091 (N_6091,N_5831,N_4517);
xor U6092 (N_6092,N_5112,N_4824);
nand U6093 (N_6093,N_5905,N_5813);
nor U6094 (N_6094,N_4749,N_4572);
nand U6095 (N_6095,N_4574,N_5323);
nand U6096 (N_6096,N_5463,N_5147);
and U6097 (N_6097,N_4641,N_5662);
nand U6098 (N_6098,N_5267,N_5873);
nor U6099 (N_6099,N_4455,N_5440);
xnor U6100 (N_6100,N_4248,N_4117);
xor U6101 (N_6101,N_4151,N_4423);
and U6102 (N_6102,N_5837,N_4171);
xnor U6103 (N_6103,N_4645,N_4223);
or U6104 (N_6104,N_4910,N_4353);
and U6105 (N_6105,N_5152,N_4185);
and U6106 (N_6106,N_4649,N_4141);
nor U6107 (N_6107,N_4841,N_4294);
xnor U6108 (N_6108,N_4705,N_5934);
nor U6109 (N_6109,N_4779,N_4853);
nor U6110 (N_6110,N_5647,N_4448);
xnor U6111 (N_6111,N_5780,N_5557);
xnor U6112 (N_6112,N_5797,N_4340);
or U6113 (N_6113,N_5464,N_5987);
or U6114 (N_6114,N_4865,N_4766);
and U6115 (N_6115,N_4752,N_5901);
or U6116 (N_6116,N_5314,N_4417);
and U6117 (N_6117,N_4133,N_5290);
and U6118 (N_6118,N_4349,N_5166);
and U6119 (N_6119,N_5860,N_4857);
and U6120 (N_6120,N_4274,N_5035);
and U6121 (N_6121,N_5495,N_4344);
or U6122 (N_6122,N_4320,N_4307);
nand U6123 (N_6123,N_4026,N_5223);
nor U6124 (N_6124,N_5069,N_4821);
nand U6125 (N_6125,N_4363,N_4253);
or U6126 (N_6126,N_4416,N_5203);
and U6127 (N_6127,N_5619,N_5331);
or U6128 (N_6128,N_5591,N_4612);
or U6129 (N_6129,N_4953,N_4086);
or U6130 (N_6130,N_4420,N_5439);
and U6131 (N_6131,N_4476,N_4225);
or U6132 (N_6132,N_5230,N_4372);
xnor U6133 (N_6133,N_5691,N_4446);
and U6134 (N_6134,N_4500,N_4456);
or U6135 (N_6135,N_5540,N_4658);
nor U6136 (N_6136,N_5978,N_5885);
nor U6137 (N_6137,N_4056,N_4773);
and U6138 (N_6138,N_5304,N_4647);
xnor U6139 (N_6139,N_4309,N_5661);
xor U6140 (N_6140,N_5415,N_4169);
nor U6141 (N_6141,N_5293,N_5635);
xnor U6142 (N_6142,N_4855,N_5274);
and U6143 (N_6143,N_5287,N_5648);
nor U6144 (N_6144,N_4458,N_4751);
nor U6145 (N_6145,N_4471,N_5169);
nor U6146 (N_6146,N_5410,N_5000);
nand U6147 (N_6147,N_5639,N_5535);
and U6148 (N_6148,N_5347,N_5187);
nor U6149 (N_6149,N_5050,N_5544);
nand U6150 (N_6150,N_5431,N_5745);
or U6151 (N_6151,N_4718,N_4484);
xnor U6152 (N_6152,N_5911,N_5021);
nand U6153 (N_6153,N_5840,N_4259);
nand U6154 (N_6154,N_5846,N_4590);
and U6155 (N_6155,N_4654,N_5402);
or U6156 (N_6156,N_4556,N_4737);
or U6157 (N_6157,N_5546,N_4917);
or U6158 (N_6158,N_5909,N_5295);
and U6159 (N_6159,N_5275,N_4160);
and U6160 (N_6160,N_5469,N_5272);
nand U6161 (N_6161,N_4366,N_4099);
nor U6162 (N_6162,N_4945,N_5594);
nand U6163 (N_6163,N_5847,N_5602);
or U6164 (N_6164,N_5940,N_4080);
and U6165 (N_6165,N_5306,N_4395);
xnor U6166 (N_6166,N_5153,N_4386);
nand U6167 (N_6167,N_5828,N_4544);
and U6168 (N_6168,N_5930,N_4034);
and U6169 (N_6169,N_5959,N_5125);
and U6170 (N_6170,N_5521,N_5170);
or U6171 (N_6171,N_4810,N_4084);
or U6172 (N_6172,N_4470,N_4346);
and U6173 (N_6173,N_5915,N_4411);
xor U6174 (N_6174,N_5763,N_5118);
and U6175 (N_6175,N_5108,N_4775);
and U6176 (N_6176,N_4886,N_4995);
nand U6177 (N_6177,N_5214,N_5140);
and U6178 (N_6178,N_4672,N_5188);
nor U6179 (N_6179,N_4188,N_5518);
xnor U6180 (N_6180,N_5570,N_4098);
nor U6181 (N_6181,N_5251,N_4870);
nand U6182 (N_6182,N_4721,N_5174);
nor U6183 (N_6183,N_5950,N_4659);
nor U6184 (N_6184,N_4332,N_5096);
or U6185 (N_6185,N_4597,N_4505);
nor U6186 (N_6186,N_5997,N_5478);
nand U6187 (N_6187,N_4715,N_4017);
nor U6188 (N_6188,N_4299,N_4090);
xor U6189 (N_6189,N_4726,N_5633);
nor U6190 (N_6190,N_5037,N_4204);
nand U6191 (N_6191,N_5806,N_5031);
nand U6192 (N_6192,N_4835,N_4110);
and U6193 (N_6193,N_4235,N_4430);
and U6194 (N_6194,N_4807,N_4758);
and U6195 (N_6195,N_4187,N_5951);
and U6196 (N_6196,N_4061,N_4121);
nor U6197 (N_6197,N_5181,N_5726);
or U6198 (N_6198,N_5771,N_5271);
nand U6199 (N_6199,N_4634,N_5400);
xor U6200 (N_6200,N_5193,N_4167);
and U6201 (N_6201,N_5130,N_5109);
or U6202 (N_6202,N_5690,N_4573);
or U6203 (N_6203,N_4605,N_5409);
xnor U6204 (N_6204,N_5265,N_5605);
nor U6205 (N_6205,N_4297,N_5386);
or U6206 (N_6206,N_5580,N_5196);
and U6207 (N_6207,N_5632,N_5363);
and U6208 (N_6208,N_4100,N_5949);
or U6209 (N_6209,N_4940,N_5220);
or U6210 (N_6210,N_4768,N_4811);
or U6211 (N_6211,N_4148,N_4483);
nand U6212 (N_6212,N_4439,N_5422);
and U6213 (N_6213,N_5083,N_4311);
nand U6214 (N_6214,N_4381,N_4293);
or U6215 (N_6215,N_5451,N_4486);
or U6216 (N_6216,N_5994,N_4889);
xor U6217 (N_6217,N_5329,N_4030);
nor U6218 (N_6218,N_5728,N_4284);
nor U6219 (N_6219,N_4345,N_5277);
or U6220 (N_6220,N_5427,N_5834);
or U6221 (N_6221,N_4781,N_4999);
or U6222 (N_6222,N_4533,N_4184);
nand U6223 (N_6223,N_4514,N_4482);
xor U6224 (N_6224,N_5916,N_5408);
nand U6225 (N_6225,N_5559,N_5561);
nor U6226 (N_6226,N_5403,N_5821);
nand U6227 (N_6227,N_4371,N_4861);
and U6228 (N_6228,N_4035,N_5844);
nor U6229 (N_6229,N_5566,N_5190);
nor U6230 (N_6230,N_4530,N_5693);
nand U6231 (N_6231,N_4719,N_5825);
or U6232 (N_6232,N_5665,N_4050);
or U6233 (N_6233,N_4450,N_5353);
nor U6234 (N_6234,N_4348,N_4531);
nand U6235 (N_6235,N_4863,N_4720);
nand U6236 (N_6236,N_5743,N_4859);
and U6237 (N_6237,N_4563,N_5088);
and U6238 (N_6238,N_5106,N_5446);
and U6239 (N_6239,N_4829,N_4047);
or U6240 (N_6240,N_4627,N_5143);
nor U6241 (N_6241,N_5739,N_4778);
and U6242 (N_6242,N_5457,N_5862);
and U6243 (N_6243,N_5689,N_5655);
and U6244 (N_6244,N_4998,N_4046);
nand U6245 (N_6245,N_4441,N_4459);
xnor U6246 (N_6246,N_5488,N_5172);
nand U6247 (N_6247,N_5565,N_5770);
and U6248 (N_6248,N_4322,N_5355);
nand U6249 (N_6249,N_4960,N_5568);
nand U6250 (N_6250,N_5030,N_4376);
nor U6251 (N_6251,N_5551,N_4019);
nor U6252 (N_6252,N_5227,N_4541);
and U6253 (N_6253,N_5758,N_5856);
nand U6254 (N_6254,N_5113,N_5449);
xnor U6255 (N_6255,N_4053,N_5044);
nor U6256 (N_6256,N_5373,N_5102);
xor U6257 (N_6257,N_5418,N_5973);
nor U6258 (N_6258,N_5286,N_4608);
nor U6259 (N_6259,N_4676,N_5232);
xnor U6260 (N_6260,N_5980,N_5849);
xor U6261 (N_6261,N_5167,N_5381);
and U6262 (N_6262,N_4321,N_5618);
nand U6263 (N_6263,N_4566,N_5466);
xnor U6264 (N_6264,N_4215,N_4923);
nor U6265 (N_6265,N_4268,N_4096);
nand U6266 (N_6266,N_5279,N_4963);
nand U6267 (N_6267,N_5351,N_5435);
or U6268 (N_6268,N_5157,N_4880);
or U6269 (N_6269,N_4228,N_5918);
nand U6270 (N_6270,N_4323,N_5894);
nand U6271 (N_6271,N_4415,N_5419);
nand U6272 (N_6272,N_4767,N_5706);
nand U6273 (N_6273,N_4196,N_4380);
nand U6274 (N_6274,N_5240,N_5336);
xnor U6275 (N_6275,N_4979,N_4252);
and U6276 (N_6276,N_5105,N_4214);
nor U6277 (N_6277,N_4736,N_4162);
nand U6278 (N_6278,N_4918,N_5462);
nor U6279 (N_6279,N_4258,N_4631);
xor U6280 (N_6280,N_4511,N_4714);
or U6281 (N_6281,N_5316,N_5789);
nand U6282 (N_6282,N_5054,N_4489);
or U6283 (N_6283,N_4334,N_5714);
xnor U6284 (N_6284,N_5204,N_5716);
nand U6285 (N_6285,N_5455,N_5765);
or U6286 (N_6286,N_4025,N_5554);
and U6287 (N_6287,N_4015,N_4968);
nand U6288 (N_6288,N_5946,N_4787);
nand U6289 (N_6289,N_4656,N_4980);
or U6290 (N_6290,N_5480,N_4437);
xnor U6291 (N_6291,N_4042,N_5053);
nor U6292 (N_6292,N_5156,N_4744);
or U6293 (N_6293,N_4147,N_4614);
xnor U6294 (N_6294,N_4911,N_5879);
and U6295 (N_6295,N_5576,N_5803);
xor U6296 (N_6296,N_5184,N_4404);
or U6297 (N_6297,N_4652,N_4818);
or U6298 (N_6298,N_5673,N_5958);
nor U6299 (N_6299,N_5774,N_5715);
xor U6300 (N_6300,N_4479,N_4230);
or U6301 (N_6301,N_4532,N_5245);
xor U6302 (N_6302,N_4291,N_4684);
or U6303 (N_6303,N_5490,N_4445);
xnor U6304 (N_6304,N_4012,N_4936);
xor U6305 (N_6305,N_5450,N_4759);
nor U6306 (N_6306,N_5182,N_5965);
nand U6307 (N_6307,N_4747,N_5168);
or U6308 (N_6308,N_4276,N_4229);
xor U6309 (N_6309,N_4189,N_5908);
xor U6310 (N_6310,N_5020,N_4272);
and U6311 (N_6311,N_5319,N_5433);
nor U6312 (N_6312,N_4808,N_5062);
nor U6313 (N_6313,N_4593,N_4625);
nor U6314 (N_6314,N_4817,N_4438);
nand U6315 (N_6315,N_4948,N_4819);
and U6316 (N_6316,N_5189,N_4161);
nor U6317 (N_6317,N_5812,N_4591);
xor U6318 (N_6318,N_4874,N_4314);
or U6319 (N_6319,N_5801,N_5912);
nor U6320 (N_6320,N_5984,N_5826);
nand U6321 (N_6321,N_5676,N_4925);
or U6322 (N_6322,N_4640,N_4365);
or U6323 (N_6323,N_5601,N_4698);
xor U6324 (N_6324,N_5672,N_5923);
nor U6325 (N_6325,N_4559,N_4198);
or U6326 (N_6326,N_4551,N_5775);
xor U6327 (N_6327,N_4449,N_4440);
and U6328 (N_6328,N_5627,N_4806);
xnor U6329 (N_6329,N_5327,N_5804);
xnor U6330 (N_6330,N_4812,N_5590);
and U6331 (N_6331,N_4242,N_4579);
or U6332 (N_6332,N_5005,N_5404);
xor U6333 (N_6333,N_5026,N_4887);
and U6334 (N_6334,N_4526,N_4725);
or U6335 (N_6335,N_4939,N_5858);
xnor U6336 (N_6336,N_4250,N_5658);
nand U6337 (N_6337,N_4091,N_5667);
nand U6338 (N_6338,N_5560,N_5332);
or U6339 (N_6339,N_4643,N_5796);
or U6340 (N_6340,N_5971,N_4803);
xor U6341 (N_6341,N_4292,N_5004);
xor U6342 (N_6342,N_5808,N_4982);
or U6343 (N_6343,N_5541,N_4234);
or U6344 (N_6344,N_5871,N_4710);
or U6345 (N_6345,N_4542,N_5974);
nand U6346 (N_6346,N_4677,N_4701);
nor U6347 (N_6347,N_4864,N_4743);
and U6348 (N_6348,N_4862,N_4237);
and U6349 (N_6349,N_4444,N_5231);
or U6350 (N_6350,N_5148,N_4407);
nand U6351 (N_6351,N_4687,N_5481);
and U6352 (N_6352,N_5931,N_4368);
nor U6353 (N_6353,N_4275,N_4723);
nand U6354 (N_6354,N_5628,N_4914);
xor U6355 (N_6355,N_5760,N_5281);
and U6356 (N_6356,N_4183,N_5028);
nand U6357 (N_6357,N_4805,N_4359);
or U6358 (N_6358,N_5164,N_4326);
xor U6359 (N_6359,N_5524,N_4915);
nor U6360 (N_6360,N_5699,N_5776);
nand U6361 (N_6361,N_5799,N_5434);
or U6362 (N_6362,N_4052,N_4890);
xor U6363 (N_6363,N_4453,N_5967);
nor U6364 (N_6364,N_5589,N_4062);
or U6365 (N_6365,N_4010,N_4895);
and U6366 (N_6366,N_4739,N_4539);
and U6367 (N_6367,N_5459,N_5519);
or U6368 (N_6368,N_4665,N_5756);
and U6369 (N_6369,N_5357,N_5848);
nor U6370 (N_6370,N_4137,N_4152);
xor U6371 (N_6371,N_4973,N_4589);
nor U6372 (N_6372,N_4433,N_4338);
xor U6373 (N_6373,N_5791,N_5354);
xor U6374 (N_6374,N_4619,N_5944);
nand U6375 (N_6375,N_5677,N_4562);
or U6376 (N_6376,N_4944,N_5201);
or U6377 (N_6377,N_5620,N_5339);
and U6378 (N_6378,N_5646,N_4858);
nor U6379 (N_6379,N_4875,N_5228);
nor U6380 (N_6380,N_5836,N_4107);
or U6381 (N_6381,N_5160,N_5705);
or U6382 (N_6382,N_5094,N_5155);
nand U6383 (N_6383,N_4690,N_4904);
nor U6384 (N_6384,N_5309,N_5503);
xnor U6385 (N_6385,N_4660,N_5437);
nor U6386 (N_6386,N_4460,N_4174);
nand U6387 (N_6387,N_5116,N_4094);
and U6388 (N_6388,N_4079,N_4628);
and U6389 (N_6389,N_4452,N_4399);
nand U6390 (N_6390,N_5320,N_4985);
or U6391 (N_6391,N_4286,N_5388);
and U6392 (N_6392,N_5176,N_5511);
and U6393 (N_6393,N_4336,N_4713);
or U6394 (N_6394,N_4629,N_4126);
nand U6395 (N_6395,N_5423,N_5372);
and U6396 (N_6396,N_5454,N_4642);
and U6397 (N_6397,N_5522,N_5683);
nor U6398 (N_6398,N_5537,N_4776);
or U6399 (N_6399,N_5759,N_5315);
xor U6400 (N_6400,N_4600,N_4068);
and U6401 (N_6401,N_4131,N_4924);
xnor U6402 (N_6402,N_4277,N_5477);
nand U6403 (N_6403,N_5744,N_5330);
nor U6404 (N_6404,N_5426,N_4280);
or U6405 (N_6405,N_5872,N_4101);
or U6406 (N_6406,N_5269,N_5630);
and U6407 (N_6407,N_5406,N_5066);
nor U6408 (N_6408,N_4607,N_5680);
xnor U6409 (N_6409,N_4922,N_5089);
nand U6410 (N_6410,N_5798,N_4881);
nor U6411 (N_6411,N_5913,N_4285);
nand U6412 (N_6412,N_5970,N_4554);
nor U6413 (N_6413,N_4240,N_5273);
xor U6414 (N_6414,N_4088,N_5276);
nand U6415 (N_6415,N_4256,N_5659);
nor U6416 (N_6416,N_4860,N_5029);
and U6417 (N_6417,N_4011,N_5823);
and U6418 (N_6418,N_4996,N_5080);
or U6419 (N_6419,N_4495,N_4564);
or U6420 (N_6420,N_4342,N_5470);
and U6421 (N_6421,N_4442,N_5349);
nand U6422 (N_6422,N_4397,N_5047);
and U6423 (N_6423,N_4784,N_5059);
and U6424 (N_6424,N_5051,N_4388);
nor U6425 (N_6425,N_5623,N_5956);
and U6426 (N_6426,N_5489,N_5666);
and U6427 (N_6427,N_5943,N_4615);
nand U6428 (N_6428,N_5945,N_4269);
nor U6429 (N_6429,N_4632,N_4075);
and U6430 (N_6430,N_5698,N_4888);
and U6431 (N_6431,N_4617,N_4447);
xnor U6432 (N_6432,N_4765,N_4261);
nor U6433 (N_6433,N_5038,N_4798);
xnor U6434 (N_6434,N_4156,N_5542);
xor U6435 (N_6435,N_5195,N_5501);
nand U6436 (N_6436,N_5248,N_4753);
xor U6437 (N_6437,N_5072,N_5321);
xor U6438 (N_6438,N_5098,N_5505);
or U6439 (N_6439,N_5509,N_5121);
or U6440 (N_6440,N_5177,N_4648);
nor U6441 (N_6441,N_4064,N_4040);
nand U6442 (N_6442,N_5514,N_4493);
xnor U6443 (N_6443,N_4843,N_5988);
or U6444 (N_6444,N_4851,N_4876);
nor U6445 (N_6445,N_4135,N_5254);
xnor U6446 (N_6446,N_4920,N_5547);
xor U6447 (N_6447,N_4004,N_4538);
or U6448 (N_6448,N_5927,N_4067);
or U6449 (N_6449,N_4106,N_5843);
nand U6450 (N_6450,N_4221,N_4697);
nor U6451 (N_6451,N_5717,N_5709);
or U6452 (N_6452,N_5614,N_5622);
and U6453 (N_6453,N_5668,N_4023);
xnor U6454 (N_6454,N_5532,N_4319);
nor U6455 (N_6455,N_5888,N_5199);
and U6456 (N_6456,N_4896,N_4220);
xor U6457 (N_6457,N_5922,N_4303);
and U6458 (N_6458,N_4180,N_4587);
or U6459 (N_6459,N_4716,N_4491);
or U6460 (N_6460,N_4129,N_4473);
and U6461 (N_6461,N_5456,N_4085);
and U6462 (N_6462,N_5811,N_4754);
nor U6463 (N_6463,N_5857,N_5074);
and U6464 (N_6464,N_4621,N_4021);
and U6465 (N_6465,N_4550,N_4316);
and U6466 (N_6466,N_4018,N_5312);
xor U6467 (N_6467,N_5242,N_4197);
and U6468 (N_6468,N_5049,N_5407);
nor U6469 (N_6469,N_4971,N_5328);
xor U6470 (N_6470,N_5014,N_4847);
and U6471 (N_6471,N_4475,N_5374);
and U6472 (N_6472,N_4685,N_5835);
xor U6473 (N_6473,N_4310,N_4900);
nor U6474 (N_6474,N_4177,N_4424);
or U6475 (N_6475,N_4981,N_4831);
nand U6476 (N_6476,N_5237,N_5393);
nor U6477 (N_6477,N_4176,N_4504);
nor U6478 (N_6478,N_4244,N_4246);
xor U6479 (N_6479,N_5880,N_4469);
nand U6480 (N_6480,N_5527,N_4144);
and U6481 (N_6481,N_5225,N_4741);
nand U6482 (N_6482,N_4149,N_4111);
or U6483 (N_6483,N_5141,N_4199);
xor U6484 (N_6484,N_4873,N_4170);
xor U6485 (N_6485,N_5679,N_5784);
nand U6486 (N_6486,N_4680,N_5822);
nand U6487 (N_6487,N_4426,N_5144);
or U6488 (N_6488,N_4521,N_5731);
xnor U6489 (N_6489,N_4792,N_4655);
and U6490 (N_6490,N_4891,N_4419);
and U6491 (N_6491,N_5213,N_5636);
xnor U6492 (N_6492,N_5465,N_5907);
and U6493 (N_6493,N_4825,N_5886);
and U6494 (N_6494,N_4443,N_4799);
nand U6495 (N_6495,N_4425,N_5942);
and U6496 (N_6496,N_4795,N_4464);
xnor U6497 (N_6497,N_4906,N_4822);
and U6498 (N_6498,N_4492,N_4883);
xor U6499 (N_6499,N_5972,N_5534);
or U6500 (N_6500,N_4602,N_4478);
nand U6501 (N_6501,N_4699,N_5609);
or U6502 (N_6502,N_5078,N_4195);
and U6503 (N_6503,N_4988,N_5395);
or U6504 (N_6504,N_5583,N_5981);
nor U6505 (N_6505,N_5842,N_4793);
nand U6506 (N_6506,N_5138,N_4626);
and U6507 (N_6507,N_4827,N_5864);
nor U6508 (N_6508,N_5311,N_5058);
xor U6509 (N_6509,N_5100,N_5517);
nor U6510 (N_6510,N_4165,N_4558);
nand U6511 (N_6511,N_5350,N_5217);
xnor U6512 (N_6512,N_5173,N_5720);
nor U6513 (N_6513,N_4060,N_5095);
and U6514 (N_6514,N_4039,N_4897);
and U6515 (N_6515,N_5520,N_4696);
and U6516 (N_6516,N_5725,N_5345);
and U6517 (N_6517,N_5710,N_4636);
or U6518 (N_6518,N_4877,N_4379);
nand U6519 (N_6519,N_4912,N_4312);
nor U6520 (N_6520,N_4674,N_5244);
xor U6521 (N_6521,N_4606,N_5063);
xnor U6522 (N_6522,N_4987,N_4339);
and U6523 (N_6523,N_4330,N_5569);
and U6524 (N_6524,N_5671,N_5491);
nor U6525 (N_6525,N_5452,N_5179);
xor U6526 (N_6526,N_5226,N_5119);
or U6527 (N_6527,N_5417,N_4295);
nand U6528 (N_6528,N_5575,N_4071);
or U6529 (N_6529,N_4219,N_4919);
and U6530 (N_6530,N_4105,N_4213);
nor U6531 (N_6531,N_5421,N_4975);
nand U6532 (N_6532,N_5307,N_4066);
or U6533 (N_6533,N_5262,N_4194);
xnor U6534 (N_6534,N_5263,N_5389);
xnor U6535 (N_6535,N_4324,N_4159);
xor U6536 (N_6536,N_5079,N_5064);
xor U6537 (N_6537,N_5645,N_5762);
xnor U6538 (N_6538,N_4826,N_5530);
xnor U6539 (N_6539,N_5258,N_4757);
and U6540 (N_6540,N_5805,N_4964);
and U6541 (N_6541,N_4770,N_4582);
nand U6542 (N_6542,N_5914,N_4181);
xor U6543 (N_6543,N_4163,N_4421);
or U6544 (N_6544,N_5616,N_5682);
nand U6545 (N_6545,N_5384,N_4961);
xor U6546 (N_6546,N_5761,N_5289);
nor U6547 (N_6547,N_4731,N_4576);
and U6548 (N_6548,N_5815,N_5297);
xnor U6549 (N_6549,N_4378,N_4588);
nor U6550 (N_6550,N_4265,N_5800);
and U6551 (N_6551,N_5073,N_4568);
or U6552 (N_6552,N_4969,N_4179);
nand U6553 (N_6553,N_4462,N_5687);
xor U6554 (N_6554,N_4125,N_5076);
or U6555 (N_6555,N_4108,N_4938);
and U6556 (N_6556,N_5585,N_5584);
or U6557 (N_6557,N_5998,N_5122);
and U6558 (N_6558,N_5929,N_4298);
nand U6559 (N_6559,N_5742,N_5851);
or U6560 (N_6560,N_5294,N_5572);
nand U6561 (N_6561,N_4552,N_4270);
or U6562 (N_6562,N_5563,N_4729);
xnor U6563 (N_6563,N_4991,N_5443);
nand U6564 (N_6564,N_5827,N_4671);
xor U6565 (N_6565,N_4190,N_4529);
and U6566 (N_6566,N_5192,N_5249);
or U6567 (N_6567,N_5833,N_5868);
and U6568 (N_6568,N_5453,N_4510);
and U6569 (N_6569,N_5611,N_5055);
nor U6570 (N_6570,N_5712,N_5895);
or U6571 (N_6571,N_4217,N_5261);
and U6572 (N_6572,N_5983,N_5773);
nor U6573 (N_6573,N_5785,N_5824);
nor U6574 (N_6574,N_4029,N_5162);
nand U6575 (N_6575,N_5727,N_4092);
nor U6576 (N_6576,N_5545,N_5111);
nor U6577 (N_6577,N_4173,N_5617);
nand U6578 (N_6578,N_4364,N_5057);
and U6579 (N_6579,N_5502,N_4842);
or U6580 (N_6580,N_5485,N_5506);
xor U6581 (N_6581,N_5387,N_5077);
and U6582 (N_6582,N_4383,N_4761);
nor U6583 (N_6583,N_5234,N_5484);
and U6584 (N_6584,N_4852,N_5881);
and U6585 (N_6585,N_4227,N_4401);
or U6586 (N_6586,N_4175,N_4260);
xnor U6587 (N_6587,N_5577,N_5684);
nand U6588 (N_6588,N_4191,N_4014);
nand U6589 (N_6589,N_5458,N_5476);
xnor U6590 (N_6590,N_5702,N_5338);
or U6591 (N_6591,N_5625,N_4193);
or U6592 (N_6592,N_4267,N_4854);
and U6593 (N_6593,N_5087,N_4974);
xnor U6594 (N_6594,N_4089,N_5884);
or U6595 (N_6595,N_4816,N_4300);
nand U6596 (N_6596,N_4620,N_5865);
nor U6597 (N_6597,N_5543,N_5206);
nor U6598 (N_6598,N_4304,N_5009);
nand U6599 (N_6599,N_4651,N_5526);
xor U6600 (N_6600,N_5734,N_5654);
nor U6601 (N_6601,N_5936,N_4136);
or U6602 (N_6602,N_4027,N_5084);
nand U6603 (N_6603,N_5574,N_5810);
nor U6604 (N_6604,N_5198,N_4856);
or U6605 (N_6605,N_4764,N_5475);
and U6606 (N_6606,N_5975,N_5963);
nand U6607 (N_6607,N_4400,N_4878);
or U6608 (N_6608,N_5586,N_5781);
nor U6609 (N_6609,N_5396,N_5224);
nor U6610 (N_6610,N_4362,N_4802);
xor U6611 (N_6611,N_4609,N_5674);
or U6612 (N_6612,N_4051,N_5022);
or U6613 (N_6613,N_4132,N_5246);
xnor U6614 (N_6614,N_5010,N_4730);
nand U6615 (N_6615,N_5889,N_4350);
xnor U6616 (N_6616,N_4547,N_5562);
and U6617 (N_6617,N_4994,N_4518);
nand U6618 (N_6618,N_4536,N_4921);
and U6619 (N_6619,N_5788,N_4989);
nor U6620 (N_6620,N_5233,N_5070);
or U6621 (N_6621,N_5753,N_5718);
nand U6622 (N_6622,N_5555,N_4689);
or U6623 (N_6623,N_4251,N_5536);
nor U6624 (N_6624,N_4112,N_4522);
and U6625 (N_6625,N_4933,N_4373);
or U6626 (N_6626,N_4327,N_4503);
nand U6627 (N_6627,N_4746,N_5444);
and U6628 (N_6628,N_4992,N_5467);
xor U6629 (N_6629,N_4095,N_4664);
and U6630 (N_6630,N_5986,N_4772);
or U6631 (N_6631,N_4076,N_4560);
nor U6632 (N_6632,N_4624,N_4732);
nand U6633 (N_6633,N_5696,N_5748);
nor U6634 (N_6634,N_5838,N_4369);
nand U6635 (N_6635,N_5892,N_5136);
or U6636 (N_6636,N_5766,N_5208);
nand U6637 (N_6637,N_5292,N_5832);
and U6638 (N_6638,N_5250,N_4673);
nor U6639 (N_6639,N_5448,N_4585);
xnor U6640 (N_6640,N_5878,N_4678);
and U6641 (N_6641,N_4123,N_5510);
nor U6642 (N_6642,N_5960,N_4281);
xnor U6643 (N_6643,N_5678,N_4786);
nand U6644 (N_6644,N_4700,N_4143);
nor U6645 (N_6645,N_5606,N_5445);
or U6646 (N_6646,N_5893,N_5067);
nor U6647 (N_6647,N_5324,N_5085);
nand U6648 (N_6648,N_5953,N_5411);
or U6649 (N_6649,N_4436,N_5159);
or U6650 (N_6650,N_5700,N_4577);
nand U6651 (N_6651,N_4057,N_5976);
xnor U6652 (N_6652,N_5933,N_5928);
or U6653 (N_6653,N_4153,N_5032);
xnor U6654 (N_6654,N_4003,N_5852);
nor U6655 (N_6655,N_5308,N_4209);
nand U6656 (N_6656,N_4243,N_5473);
nand U6657 (N_6657,N_5252,N_5414);
nor U6658 (N_6658,N_4601,N_4352);
and U6659 (N_6659,N_4247,N_5769);
xor U6660 (N_6660,N_5829,N_5513);
or U6661 (N_6661,N_5681,N_4032);
nand U6662 (N_6662,N_4683,N_5604);
nand U6663 (N_6663,N_5379,N_5216);
xnor U6664 (N_6664,N_4977,N_4820);
nand U6665 (N_6665,N_5787,N_4392);
nor U6666 (N_6666,N_4804,N_4296);
or U6667 (N_6667,N_4611,N_5802);
xnor U6668 (N_6668,N_5145,N_4202);
nand U6669 (N_6669,N_5642,N_5081);
nand U6670 (N_6670,N_4055,N_5999);
nor U6671 (N_6671,N_4929,N_4210);
and U6672 (N_6672,N_5135,N_5795);
or U6673 (N_6673,N_4943,N_5043);
nand U6674 (N_6674,N_5356,N_5218);
nand U6675 (N_6675,N_5579,N_4748);
xor U6676 (N_6676,N_4257,N_4138);
nor U6677 (N_6677,N_4130,N_5180);
and U6678 (N_6678,N_5793,N_5424);
nand U6679 (N_6679,N_5461,N_4801);
and U6680 (N_6680,N_4168,N_4686);
and U6681 (N_6681,N_5134,N_4360);
nand U6682 (N_6682,N_4527,N_4990);
and U6683 (N_6683,N_4934,N_4435);
or U6684 (N_6684,N_5496,N_5723);
nand U6685 (N_6685,N_5229,N_4020);
nor U6686 (N_6686,N_5305,N_4158);
nor U6687 (N_6687,N_5952,N_5082);
nor U6688 (N_6688,N_4211,N_5075);
and U6689 (N_6689,N_5221,N_5367);
or U6690 (N_6690,N_5256,N_4633);
nor U6691 (N_6691,N_5650,N_5855);
or U6692 (N_6692,N_5567,N_4957);
or U6693 (N_6693,N_4846,N_5436);
nor U6694 (N_6694,N_5937,N_5398);
or U6695 (N_6695,N_4894,N_5300);
and U6696 (N_6696,N_5877,N_5091);
nor U6697 (N_6697,N_4670,N_5474);
and U6698 (N_6698,N_4931,N_5649);
and U6699 (N_6699,N_5549,N_4800);
xnor U6700 (N_6700,N_4201,N_4356);
and U6701 (N_6701,N_4472,N_5025);
nor U6702 (N_6702,N_4958,N_4735);
or U6703 (N_6703,N_4932,N_5814);
xnor U6704 (N_6704,N_4791,N_5129);
or U6705 (N_6705,N_4394,N_5935);
and U6706 (N_6706,N_5442,N_4537);
and U6707 (N_6707,N_4722,N_5638);
and U6708 (N_6708,N_4361,N_4384);
nor U6709 (N_6709,N_4007,N_5596);
or U6710 (N_6710,N_4882,N_4613);
and U6711 (N_6711,N_4899,N_4150);
or U6712 (N_6712,N_5048,N_5061);
and U6713 (N_6713,N_5185,N_5767);
nor U6714 (N_6714,N_5413,N_4318);
and U6715 (N_6715,N_5171,N_4301);
xor U6716 (N_6716,N_4789,N_4951);
nand U6717 (N_6717,N_4575,N_5663);
and U6718 (N_6718,N_5920,N_5807);
or U6719 (N_6719,N_5288,N_4005);
xnor U6720 (N_6720,N_5317,N_5366);
nor U6721 (N_6721,N_4837,N_4809);
and U6722 (N_6722,N_5412,N_4490);
nand U6723 (N_6723,N_4663,N_5750);
nand U6724 (N_6724,N_4580,N_5370);
and U6725 (N_6725,N_5344,N_4070);
nor U6726 (N_6726,N_4264,N_4341);
and U6727 (N_6727,N_5285,N_5253);
xor U6728 (N_6728,N_5957,N_4630);
and U6729 (N_6729,N_4236,N_4409);
nor U6730 (N_6730,N_5027,N_4565);
and U6731 (N_6731,N_4618,N_5298);
xnor U6732 (N_6732,N_4355,N_4054);
nor U6733 (N_6733,N_4797,N_5018);
and U6734 (N_6734,N_5007,N_5660);
and U6735 (N_6735,N_5777,N_4077);
or U6736 (N_6736,N_4434,N_4200);
xnor U6737 (N_6737,N_5969,N_5792);
xnor U6738 (N_6738,N_5139,N_5041);
nand U6739 (N_6739,N_4487,N_4774);
xor U6740 (N_6740,N_4422,N_4208);
nor U6741 (N_6741,N_5117,N_4413);
xnor U6742 (N_6742,N_4594,N_5735);
nand U6743 (N_6743,N_5515,N_4543);
nand U6744 (N_6744,N_5093,N_5280);
or U6745 (N_6745,N_5947,N_4755);
xnor U6746 (N_6746,N_4006,N_5954);
xor U6747 (N_6747,N_5303,N_5103);
nor U6748 (N_6748,N_5816,N_5626);
nor U6749 (N_6749,N_5302,N_4073);
or U6750 (N_6750,N_4909,N_5841);
and U6751 (N_6751,N_4465,N_5516);
or U6752 (N_6752,N_4466,N_4871);
or U6753 (N_6753,N_4840,N_4935);
or U6754 (N_6754,N_5247,N_4616);
or U6755 (N_6755,N_4884,N_5003);
nand U6756 (N_6756,N_4555,N_5123);
or U6757 (N_6757,N_4367,N_5961);
nor U6758 (N_6758,N_5755,N_5420);
xnor U6759 (N_6759,N_4044,N_4008);
and U6760 (N_6760,N_5525,N_5092);
xnor U6761 (N_6761,N_5023,N_4497);
nor U6762 (N_6762,N_4065,N_5867);
and U6763 (N_6763,N_5359,N_4952);
and U6764 (N_6764,N_5034,N_5416);
nand U6765 (N_6765,N_4287,N_4283);
xor U6766 (N_6766,N_4222,N_5019);
or U6767 (N_6767,N_5599,N_4879);
and U6768 (N_6768,N_4418,N_4734);
and U6769 (N_6769,N_4506,N_4120);
and U6770 (N_6770,N_4650,N_4867);
and U6771 (N_6771,N_4637,N_4549);
nand U6772 (N_6772,N_4534,N_5238);
or U6773 (N_6773,N_5236,N_4428);
and U6774 (N_6774,N_5794,N_5205);
xnor U6775 (N_6775,N_5995,N_5259);
nor U6776 (N_6776,N_4041,N_4926);
xnor U6777 (N_6777,N_5966,N_4031);
and U6778 (N_6778,N_4278,N_5613);
nand U6779 (N_6779,N_4644,N_4838);
nand U6780 (N_6780,N_5612,N_5854);
and U6781 (N_6781,N_4241,N_4059);
xnor U6782 (N_6782,N_4370,N_5657);
nor U6783 (N_6783,N_4097,N_4083);
nand U6784 (N_6784,N_4239,N_4127);
and U6785 (N_6785,N_4461,N_4738);
nor U6786 (N_6786,N_5175,N_4669);
nand U6787 (N_6787,N_5498,N_5380);
and U6788 (N_6788,N_5212,N_5751);
and U6789 (N_6789,N_5533,N_5210);
and U6790 (N_6790,N_4224,N_5243);
nand U6791 (N_6791,N_4058,N_4688);
nand U6792 (N_6792,N_4093,N_5741);
or U6793 (N_6793,N_5979,N_5017);
or U6794 (N_6794,N_4358,N_5863);
xor U6795 (N_6795,N_4950,N_5869);
or U6796 (N_6796,N_4115,N_5692);
and U6797 (N_6797,N_4646,N_4508);
nor U6798 (N_6798,N_4124,N_5817);
xnor U6799 (N_6799,N_4000,N_5124);
and U6800 (N_6800,N_4477,N_4354);
nor U6801 (N_6801,N_5340,N_4692);
nor U6802 (N_6802,N_4623,N_5610);
nand U6803 (N_6803,N_4103,N_4232);
nand U6804 (N_6804,N_5313,N_5006);
xor U6805 (N_6805,N_5656,N_4512);
nand U6806 (N_6806,N_5779,N_4830);
nand U6807 (N_6807,N_4834,N_5850);
and U6808 (N_6808,N_4231,N_5874);
xor U6809 (N_6809,N_4668,N_4289);
nor U6810 (N_6810,N_4742,N_4308);
xnor U6811 (N_6811,N_4082,N_5163);
nor U6812 (N_6812,N_5405,N_5120);
or U6813 (N_6813,N_5333,N_4203);
xor U6814 (N_6814,N_4907,N_5592);
nand U6815 (N_6815,N_5341,N_5640);
and U6816 (N_6816,N_5002,N_4288);
and U6817 (N_6817,N_5110,N_5137);
xor U6818 (N_6818,N_5115,N_4377);
and U6819 (N_6819,N_4548,N_5729);
nand U6820 (N_6820,N_4790,N_5197);
nor U6821 (N_6821,N_4913,N_4603);
xnor U6822 (N_6822,N_4694,N_4788);
and U6823 (N_6823,N_4836,N_5326);
and U6824 (N_6824,N_5040,N_4959);
nand U6825 (N_6825,N_5012,N_4396);
nand U6826 (N_6826,N_5200,N_5992);
nand U6827 (N_6827,N_5133,N_4596);
xnor U6828 (N_6828,N_4905,N_4357);
and U6829 (N_6829,N_5500,N_5675);
nor U6830 (N_6830,N_4970,N_4033);
xor U6831 (N_6831,N_4691,N_4610);
and U6832 (N_6832,N_5360,N_5207);
and U6833 (N_6833,N_4432,N_4782);
and U6834 (N_6834,N_5704,N_4653);
xor U6835 (N_6835,N_5701,N_5581);
or U6836 (N_6836,N_5508,N_4604);
and U6837 (N_6837,N_5664,N_5991);
nand U6838 (N_6838,N_5178,N_5839);
and U6839 (N_6839,N_4186,N_5891);
nor U6840 (N_6840,N_4385,N_5859);
and U6841 (N_6841,N_4707,N_5512);
xor U6842 (N_6842,N_4967,N_4406);
nor U6843 (N_6843,N_5399,N_4703);
nor U6844 (N_6844,N_5101,N_5870);
xor U6845 (N_6845,N_4266,N_4207);
xor U6846 (N_6846,N_4206,N_4740);
or U6847 (N_6847,N_4708,N_5342);
or U6848 (N_6848,N_5571,N_5046);
xor U6849 (N_6849,N_5917,N_4382);
nand U6850 (N_6850,N_5719,N_5131);
or U6851 (N_6851,N_4451,N_5948);
nand U6852 (N_6852,N_5924,N_5432);
nor U6853 (N_6853,N_4262,N_4457);
or U6854 (N_6854,N_4306,N_4941);
and U6855 (N_6855,N_5564,N_4557);
nand U6856 (N_6856,N_4595,N_4540);
nand U6857 (N_6857,N_4182,N_5809);
or U6858 (N_6858,N_5086,N_5697);
nor U6859 (N_6859,N_5897,N_4119);
nand U6860 (N_6860,N_4375,N_4122);
or U6861 (N_6861,N_4868,N_4502);
and U6862 (N_6862,N_5896,N_5493);
or U6863 (N_6863,N_4245,N_5903);
xor U6864 (N_6864,N_4045,N_5430);
nand U6865 (N_6865,N_4845,N_4331);
xnor U6866 (N_6866,N_5241,N_4733);
xnor U6867 (N_6867,N_4390,N_5376);
and U6868 (N_6868,N_5919,N_5257);
nor U6869 (N_6869,N_5900,N_4901);
or U6870 (N_6870,N_5368,N_4037);
and U6871 (N_6871,N_5558,N_5703);
nor U6872 (N_6872,N_4763,N_5472);
nand U6873 (N_6873,N_4104,N_4335);
nand U6874 (N_6874,N_5507,N_4525);
and U6875 (N_6875,N_5548,N_4794);
xor U6876 (N_6876,N_5556,N_4592);
nor U6877 (N_6877,N_4022,N_5910);
xnor U6878 (N_6878,N_4569,N_5154);
and U6879 (N_6879,N_4693,N_5722);
or U6880 (N_6880,N_5730,N_4546);
and U6881 (N_6881,N_4496,N_5550);
nor U6882 (N_6882,N_5875,N_4570);
nand U6883 (N_6883,N_5686,N_4523);
or U6884 (N_6884,N_5364,N_5539);
xnor U6885 (N_6885,N_4965,N_4978);
nor U6886 (N_6886,N_5045,N_5853);
and U6887 (N_6887,N_4016,N_5278);
or U6888 (N_6888,N_4638,N_4028);
or U6889 (N_6889,N_4972,N_5707);
and U6890 (N_6890,N_4949,N_4711);
nor U6891 (N_6891,N_5926,N_5441);
or U6892 (N_6892,N_4139,N_4709);
or U6893 (N_6893,N_5146,N_4571);
and U6894 (N_6894,N_5904,N_5597);
nor U6895 (N_6895,N_4993,N_4403);
xnor U6896 (N_6896,N_4402,N_4928);
and U6897 (N_6897,N_4024,N_4724);
xor U6898 (N_6898,N_5215,N_5318);
xor U6899 (N_6899,N_4997,N_4528);
or U6900 (N_6900,N_4848,N_4063);
and U6901 (N_6901,N_4205,N_5219);
and U6902 (N_6902,N_5711,N_5282);
nand U6903 (N_6903,N_5651,N_4983);
xnor U6904 (N_6904,N_5993,N_5499);
nand U6905 (N_6905,N_4192,N_4081);
and U6906 (N_6906,N_4140,N_5982);
xor U6907 (N_6907,N_5291,N_5757);
nand U6908 (N_6908,N_4956,N_5428);
xnor U6909 (N_6909,N_5382,N_5429);
and U6910 (N_6910,N_5887,N_5191);
and U6911 (N_6911,N_4955,N_4391);
nand U6912 (N_6912,N_4866,N_5325);
nand U6913 (N_6913,N_4410,N_4263);
and U6914 (N_6914,N_4271,N_5608);
nor U6915 (N_6915,N_5266,N_4414);
and U6916 (N_6916,N_5486,N_4254);
and U6917 (N_6917,N_5938,N_4255);
xnor U6918 (N_6918,N_5392,N_4584);
or U6919 (N_6919,N_5996,N_5039);
nor U6920 (N_6920,N_5637,N_5754);
and U6921 (N_6921,N_4515,N_4216);
and U6922 (N_6922,N_5299,N_4902);
xnor U6923 (N_6923,N_5264,N_5001);
nor U6924 (N_6924,N_5068,N_5786);
xor U6925 (N_6925,N_5736,N_5898);
or U6926 (N_6926,N_4893,N_5348);
nand U6927 (N_6927,N_4954,N_4760);
or U6928 (N_6928,N_5694,N_5531);
nor U6929 (N_6929,N_5447,N_5670);
xnor U6930 (N_6930,N_4702,N_5011);
nand U6931 (N_6931,N_4405,N_4908);
or U6932 (N_6932,N_4249,N_4333);
or U6933 (N_6933,N_4927,N_4780);
nand U6934 (N_6934,N_5861,N_5964);
xnor U6935 (N_6935,N_5819,N_5397);
and U6936 (N_6936,N_4317,N_4813);
nand U6937 (N_6937,N_5322,N_4113);
nand U6938 (N_6938,N_5818,N_5377);
or U6939 (N_6939,N_4583,N_5939);
and U6940 (N_6940,N_5284,N_5194);
and U6941 (N_6941,N_4157,N_5394);
and U6942 (N_6942,N_4657,N_5634);
xnor U6943 (N_6943,N_4561,N_4408);
nand U6944 (N_6944,N_5985,N_5151);
or U6945 (N_6945,N_4567,N_4328);
and U6946 (N_6946,N_4302,N_5643);
nand U6947 (N_6947,N_4844,N_5391);
nor U6948 (N_6948,N_4329,N_5438);
nor U6949 (N_6949,N_4116,N_5270);
xor U6950 (N_6950,N_5504,N_5695);
or U6951 (N_6951,N_5310,N_4946);
nand U6952 (N_6952,N_5883,N_4485);
and U6953 (N_6953,N_5334,N_5375);
xnor U6954 (N_6954,N_4427,N_5624);
or U6955 (N_6955,N_5126,N_5631);
or U6956 (N_6956,N_4013,N_4325);
nand U6957 (N_6957,N_5553,N_5343);
nand U6958 (N_6958,N_5369,N_4916);
and U6959 (N_6959,N_5749,N_5724);
and U6960 (N_6960,N_5733,N_5593);
or U6961 (N_6961,N_5065,N_5925);
and U6962 (N_6962,N_4315,N_4762);
nand U6963 (N_6963,N_5772,N_4154);
nand U6964 (N_6964,N_5621,N_5790);
and U6965 (N_6965,N_5362,N_4282);
and U6966 (N_6966,N_5114,N_4545);
nor U6967 (N_6967,N_4347,N_4145);
xor U6968 (N_6968,N_5603,N_4937);
and U6969 (N_6969,N_4832,N_4387);
xnor U6970 (N_6970,N_5721,N_4706);
nor U6971 (N_6971,N_4074,N_5582);
nand U6972 (N_6972,N_5255,N_4454);
and U6973 (N_6973,N_4586,N_4114);
and U6974 (N_6974,N_4038,N_5346);
xor U6975 (N_6975,N_4279,N_5479);
nand U6976 (N_6976,N_4745,N_5820);
nand U6977 (N_6977,N_4036,N_4783);
or U6978 (N_6978,N_4750,N_5060);
xor U6979 (N_6979,N_4001,N_5128);
and U6980 (N_6980,N_5301,N_5552);
nand U6981 (N_6981,N_5385,N_4102);
nor U6982 (N_6982,N_5990,N_5768);
xnor U6983 (N_6983,N_4849,N_4233);
or U6984 (N_6984,N_4002,N_4828);
and U6985 (N_6985,N_4172,N_5161);
nor U6986 (N_6986,N_5955,N_4146);
or U6987 (N_6987,N_5337,N_4305);
or U6988 (N_6988,N_4682,N_5283);
nand U6989 (N_6989,N_4695,N_4976);
xor U6990 (N_6990,N_4048,N_5989);
nand U6991 (N_6991,N_5607,N_4756);
xnor U6992 (N_6992,N_4069,N_5598);
and U6993 (N_6993,N_4343,N_5764);
nand U6994 (N_6994,N_5600,N_4043);
nor U6995 (N_6995,N_4777,N_5941);
and U6996 (N_6996,N_4814,N_5538);
xor U6997 (N_6997,N_5529,N_5483);
nand U6998 (N_6998,N_4635,N_4947);
nor U6999 (N_6999,N_4520,N_5968);
or U7000 (N_7000,N_5421,N_4042);
and U7001 (N_7001,N_4531,N_4061);
nor U7002 (N_7002,N_4620,N_4911);
nor U7003 (N_7003,N_4112,N_5358);
nand U7004 (N_7004,N_5376,N_4665);
and U7005 (N_7005,N_5483,N_5681);
or U7006 (N_7006,N_5107,N_5935);
nand U7007 (N_7007,N_5892,N_4079);
xnor U7008 (N_7008,N_5180,N_4520);
xnor U7009 (N_7009,N_4993,N_4794);
nor U7010 (N_7010,N_4849,N_4777);
xnor U7011 (N_7011,N_4745,N_5200);
and U7012 (N_7012,N_5281,N_4295);
nand U7013 (N_7013,N_5248,N_5261);
nand U7014 (N_7014,N_5774,N_4418);
or U7015 (N_7015,N_5515,N_5417);
or U7016 (N_7016,N_4044,N_4735);
nand U7017 (N_7017,N_5462,N_5724);
and U7018 (N_7018,N_5198,N_5730);
nand U7019 (N_7019,N_5226,N_4243);
and U7020 (N_7020,N_4886,N_4880);
and U7021 (N_7021,N_5965,N_4484);
or U7022 (N_7022,N_4516,N_5718);
xnor U7023 (N_7023,N_4559,N_5886);
or U7024 (N_7024,N_5091,N_4855);
and U7025 (N_7025,N_4924,N_5640);
xnor U7026 (N_7026,N_5893,N_4168);
xnor U7027 (N_7027,N_4894,N_4309);
nor U7028 (N_7028,N_4974,N_5877);
or U7029 (N_7029,N_4635,N_4289);
or U7030 (N_7030,N_4006,N_5767);
or U7031 (N_7031,N_5959,N_5057);
or U7032 (N_7032,N_4038,N_5303);
xor U7033 (N_7033,N_4754,N_4802);
nor U7034 (N_7034,N_4164,N_5731);
or U7035 (N_7035,N_4898,N_5576);
and U7036 (N_7036,N_5741,N_5950);
or U7037 (N_7037,N_4228,N_4998);
nand U7038 (N_7038,N_5638,N_4918);
nand U7039 (N_7039,N_4634,N_5691);
nor U7040 (N_7040,N_4372,N_5943);
or U7041 (N_7041,N_4810,N_5888);
xnor U7042 (N_7042,N_4061,N_4268);
nor U7043 (N_7043,N_5298,N_5997);
or U7044 (N_7044,N_4327,N_4029);
xnor U7045 (N_7045,N_5119,N_4714);
nand U7046 (N_7046,N_4094,N_5213);
nor U7047 (N_7047,N_4648,N_4944);
or U7048 (N_7048,N_4432,N_4064);
nand U7049 (N_7049,N_4959,N_4138);
xor U7050 (N_7050,N_5127,N_5785);
nor U7051 (N_7051,N_5852,N_4500);
nor U7052 (N_7052,N_4588,N_4129);
nand U7053 (N_7053,N_4525,N_4380);
xnor U7054 (N_7054,N_5486,N_4686);
nor U7055 (N_7055,N_5038,N_4482);
nor U7056 (N_7056,N_5544,N_5034);
or U7057 (N_7057,N_4935,N_4674);
or U7058 (N_7058,N_4656,N_4636);
and U7059 (N_7059,N_4069,N_4870);
nor U7060 (N_7060,N_4737,N_4574);
or U7061 (N_7061,N_4442,N_4607);
nand U7062 (N_7062,N_4260,N_5034);
nand U7063 (N_7063,N_5865,N_4795);
and U7064 (N_7064,N_4996,N_4765);
xnor U7065 (N_7065,N_5970,N_4418);
xor U7066 (N_7066,N_4930,N_5441);
and U7067 (N_7067,N_4003,N_4354);
nor U7068 (N_7068,N_4409,N_4800);
and U7069 (N_7069,N_5075,N_5129);
or U7070 (N_7070,N_4952,N_5175);
xnor U7071 (N_7071,N_5904,N_4535);
or U7072 (N_7072,N_5042,N_5086);
and U7073 (N_7073,N_4370,N_5403);
or U7074 (N_7074,N_4234,N_5407);
xnor U7075 (N_7075,N_4338,N_5820);
xor U7076 (N_7076,N_4904,N_4088);
and U7077 (N_7077,N_5034,N_5367);
or U7078 (N_7078,N_4619,N_5255);
xor U7079 (N_7079,N_5513,N_5973);
or U7080 (N_7080,N_4452,N_4660);
nor U7081 (N_7081,N_4757,N_5390);
nor U7082 (N_7082,N_5067,N_5750);
or U7083 (N_7083,N_5935,N_4822);
and U7084 (N_7084,N_4568,N_5048);
xnor U7085 (N_7085,N_5350,N_5649);
nand U7086 (N_7086,N_5090,N_4952);
or U7087 (N_7087,N_5001,N_5614);
nand U7088 (N_7088,N_5422,N_5514);
or U7089 (N_7089,N_5500,N_4980);
or U7090 (N_7090,N_4077,N_5627);
or U7091 (N_7091,N_5688,N_4194);
nand U7092 (N_7092,N_4420,N_5014);
xor U7093 (N_7093,N_5501,N_4258);
xnor U7094 (N_7094,N_5257,N_5029);
xnor U7095 (N_7095,N_5133,N_5219);
and U7096 (N_7096,N_5628,N_4645);
xor U7097 (N_7097,N_4057,N_5632);
nor U7098 (N_7098,N_5012,N_5840);
nand U7099 (N_7099,N_4267,N_4194);
nor U7100 (N_7100,N_4085,N_5407);
xor U7101 (N_7101,N_4457,N_5297);
or U7102 (N_7102,N_4211,N_5680);
and U7103 (N_7103,N_4086,N_4878);
xor U7104 (N_7104,N_4129,N_4424);
and U7105 (N_7105,N_5876,N_4748);
and U7106 (N_7106,N_4320,N_4834);
and U7107 (N_7107,N_5215,N_5685);
nor U7108 (N_7108,N_5079,N_5671);
nor U7109 (N_7109,N_5126,N_4334);
nand U7110 (N_7110,N_5421,N_5471);
or U7111 (N_7111,N_4799,N_4260);
nor U7112 (N_7112,N_4311,N_5988);
or U7113 (N_7113,N_4549,N_5373);
xor U7114 (N_7114,N_5399,N_4527);
xor U7115 (N_7115,N_4434,N_5786);
xnor U7116 (N_7116,N_4909,N_4988);
and U7117 (N_7117,N_4159,N_5877);
and U7118 (N_7118,N_5221,N_5198);
nor U7119 (N_7119,N_5174,N_4257);
and U7120 (N_7120,N_4019,N_5784);
and U7121 (N_7121,N_5728,N_4340);
nand U7122 (N_7122,N_5478,N_5635);
and U7123 (N_7123,N_4433,N_4537);
nor U7124 (N_7124,N_5480,N_4108);
nor U7125 (N_7125,N_4046,N_4394);
or U7126 (N_7126,N_5624,N_5207);
or U7127 (N_7127,N_5456,N_5196);
nand U7128 (N_7128,N_4200,N_5726);
nor U7129 (N_7129,N_4548,N_4814);
nand U7130 (N_7130,N_5539,N_4735);
nor U7131 (N_7131,N_5273,N_4614);
nor U7132 (N_7132,N_5205,N_5071);
nand U7133 (N_7133,N_4254,N_5239);
or U7134 (N_7134,N_4435,N_5634);
and U7135 (N_7135,N_4743,N_5639);
or U7136 (N_7136,N_5907,N_4607);
nand U7137 (N_7137,N_5329,N_5566);
nor U7138 (N_7138,N_4917,N_4458);
xor U7139 (N_7139,N_5435,N_5881);
nor U7140 (N_7140,N_4717,N_4364);
or U7141 (N_7141,N_5034,N_4217);
nor U7142 (N_7142,N_5027,N_4036);
or U7143 (N_7143,N_4864,N_4230);
or U7144 (N_7144,N_5705,N_4072);
or U7145 (N_7145,N_5843,N_5930);
xnor U7146 (N_7146,N_4010,N_5470);
and U7147 (N_7147,N_5718,N_5546);
nor U7148 (N_7148,N_5459,N_4243);
xnor U7149 (N_7149,N_4942,N_5892);
nor U7150 (N_7150,N_4307,N_4847);
and U7151 (N_7151,N_5836,N_5538);
nand U7152 (N_7152,N_5163,N_5691);
xnor U7153 (N_7153,N_4069,N_5491);
or U7154 (N_7154,N_5201,N_5024);
or U7155 (N_7155,N_4599,N_4359);
and U7156 (N_7156,N_4326,N_5736);
xnor U7157 (N_7157,N_5462,N_4357);
nand U7158 (N_7158,N_4765,N_4887);
xor U7159 (N_7159,N_5941,N_5642);
nand U7160 (N_7160,N_4660,N_5029);
nand U7161 (N_7161,N_4921,N_5551);
xor U7162 (N_7162,N_4045,N_5050);
or U7163 (N_7163,N_4435,N_5166);
nor U7164 (N_7164,N_4272,N_5704);
or U7165 (N_7165,N_5592,N_4355);
or U7166 (N_7166,N_4052,N_4559);
and U7167 (N_7167,N_4250,N_5721);
xnor U7168 (N_7168,N_5428,N_4979);
or U7169 (N_7169,N_5733,N_4096);
nor U7170 (N_7170,N_4145,N_5377);
xor U7171 (N_7171,N_5873,N_4362);
nand U7172 (N_7172,N_5912,N_5006);
or U7173 (N_7173,N_5780,N_4035);
or U7174 (N_7174,N_5514,N_4521);
and U7175 (N_7175,N_4582,N_4272);
or U7176 (N_7176,N_4186,N_5939);
or U7177 (N_7177,N_4150,N_5929);
or U7178 (N_7178,N_5300,N_5297);
nor U7179 (N_7179,N_4124,N_4843);
and U7180 (N_7180,N_5498,N_4576);
or U7181 (N_7181,N_5728,N_5173);
nor U7182 (N_7182,N_5585,N_4175);
xor U7183 (N_7183,N_4586,N_4623);
or U7184 (N_7184,N_5966,N_4332);
or U7185 (N_7185,N_5233,N_4179);
and U7186 (N_7186,N_4672,N_4631);
or U7187 (N_7187,N_4585,N_5464);
and U7188 (N_7188,N_5083,N_4767);
nor U7189 (N_7189,N_5888,N_4987);
or U7190 (N_7190,N_5944,N_4571);
xor U7191 (N_7191,N_4383,N_4831);
xnor U7192 (N_7192,N_4658,N_4197);
or U7193 (N_7193,N_4738,N_4255);
nor U7194 (N_7194,N_4563,N_4929);
xor U7195 (N_7195,N_5216,N_5775);
or U7196 (N_7196,N_4691,N_5653);
nand U7197 (N_7197,N_5113,N_5308);
or U7198 (N_7198,N_4996,N_4994);
and U7199 (N_7199,N_5168,N_5534);
nand U7200 (N_7200,N_4267,N_5904);
or U7201 (N_7201,N_4147,N_4573);
and U7202 (N_7202,N_5487,N_5736);
nand U7203 (N_7203,N_4647,N_5285);
nor U7204 (N_7204,N_4737,N_5822);
nand U7205 (N_7205,N_5418,N_4749);
or U7206 (N_7206,N_4654,N_4898);
and U7207 (N_7207,N_4085,N_4723);
and U7208 (N_7208,N_4583,N_5441);
and U7209 (N_7209,N_4329,N_5081);
xnor U7210 (N_7210,N_4744,N_4225);
nor U7211 (N_7211,N_4024,N_4551);
nor U7212 (N_7212,N_4827,N_5728);
and U7213 (N_7213,N_5324,N_4313);
or U7214 (N_7214,N_5096,N_4076);
and U7215 (N_7215,N_5617,N_4260);
or U7216 (N_7216,N_4141,N_5650);
and U7217 (N_7217,N_5894,N_5051);
nand U7218 (N_7218,N_5882,N_4458);
and U7219 (N_7219,N_5026,N_5728);
or U7220 (N_7220,N_4153,N_5439);
nor U7221 (N_7221,N_4397,N_5039);
xor U7222 (N_7222,N_5372,N_5928);
or U7223 (N_7223,N_4050,N_4118);
nor U7224 (N_7224,N_5782,N_4399);
xnor U7225 (N_7225,N_5130,N_5823);
xor U7226 (N_7226,N_5142,N_5809);
and U7227 (N_7227,N_5968,N_4380);
xnor U7228 (N_7228,N_4526,N_4399);
nand U7229 (N_7229,N_4441,N_4785);
xor U7230 (N_7230,N_5845,N_5671);
or U7231 (N_7231,N_5712,N_5598);
or U7232 (N_7232,N_5288,N_5592);
nor U7233 (N_7233,N_5374,N_4326);
or U7234 (N_7234,N_5131,N_4414);
nor U7235 (N_7235,N_5150,N_4946);
nand U7236 (N_7236,N_5479,N_5288);
nand U7237 (N_7237,N_5135,N_5489);
nand U7238 (N_7238,N_5105,N_4755);
and U7239 (N_7239,N_4074,N_4586);
nor U7240 (N_7240,N_5862,N_5135);
nor U7241 (N_7241,N_5498,N_4524);
xor U7242 (N_7242,N_4817,N_5033);
or U7243 (N_7243,N_5391,N_5129);
nor U7244 (N_7244,N_5458,N_5641);
and U7245 (N_7245,N_5716,N_4631);
xnor U7246 (N_7246,N_4150,N_5541);
xor U7247 (N_7247,N_4238,N_5360);
or U7248 (N_7248,N_5315,N_5517);
and U7249 (N_7249,N_5305,N_4551);
and U7250 (N_7250,N_5391,N_4183);
nor U7251 (N_7251,N_5749,N_5114);
nand U7252 (N_7252,N_5476,N_4897);
or U7253 (N_7253,N_4756,N_4358);
xor U7254 (N_7254,N_5760,N_5351);
or U7255 (N_7255,N_5427,N_4760);
xnor U7256 (N_7256,N_4451,N_5438);
or U7257 (N_7257,N_4704,N_4568);
and U7258 (N_7258,N_5734,N_5579);
or U7259 (N_7259,N_5745,N_4012);
and U7260 (N_7260,N_4769,N_4321);
nand U7261 (N_7261,N_4516,N_5811);
nor U7262 (N_7262,N_4806,N_4224);
or U7263 (N_7263,N_5526,N_5137);
or U7264 (N_7264,N_4609,N_4459);
nor U7265 (N_7265,N_4878,N_5333);
or U7266 (N_7266,N_4091,N_4128);
nor U7267 (N_7267,N_4802,N_4011);
xnor U7268 (N_7268,N_4226,N_4317);
xor U7269 (N_7269,N_4208,N_5934);
nor U7270 (N_7270,N_5190,N_4113);
xnor U7271 (N_7271,N_4426,N_5322);
and U7272 (N_7272,N_5981,N_4938);
nor U7273 (N_7273,N_5043,N_5129);
xnor U7274 (N_7274,N_5603,N_4571);
and U7275 (N_7275,N_4260,N_4952);
nand U7276 (N_7276,N_4627,N_4820);
nand U7277 (N_7277,N_4898,N_5832);
xnor U7278 (N_7278,N_4172,N_4750);
nand U7279 (N_7279,N_4473,N_4254);
and U7280 (N_7280,N_5030,N_5655);
and U7281 (N_7281,N_5134,N_4794);
and U7282 (N_7282,N_4594,N_5611);
xor U7283 (N_7283,N_5682,N_4250);
nand U7284 (N_7284,N_4915,N_4033);
and U7285 (N_7285,N_4111,N_4248);
and U7286 (N_7286,N_4093,N_4937);
xnor U7287 (N_7287,N_4964,N_5810);
or U7288 (N_7288,N_5631,N_5796);
and U7289 (N_7289,N_4731,N_4101);
and U7290 (N_7290,N_5618,N_5181);
nand U7291 (N_7291,N_5082,N_5894);
xnor U7292 (N_7292,N_5261,N_5463);
nor U7293 (N_7293,N_5524,N_5011);
nor U7294 (N_7294,N_5543,N_5182);
nand U7295 (N_7295,N_4926,N_5171);
or U7296 (N_7296,N_5811,N_4751);
and U7297 (N_7297,N_4243,N_5703);
and U7298 (N_7298,N_4998,N_5485);
xor U7299 (N_7299,N_4643,N_5785);
and U7300 (N_7300,N_5436,N_4077);
nand U7301 (N_7301,N_4862,N_4967);
nand U7302 (N_7302,N_4495,N_4776);
nor U7303 (N_7303,N_5637,N_4700);
or U7304 (N_7304,N_4665,N_4668);
nor U7305 (N_7305,N_4902,N_5922);
or U7306 (N_7306,N_5976,N_5258);
nor U7307 (N_7307,N_5250,N_4534);
nand U7308 (N_7308,N_5359,N_4605);
and U7309 (N_7309,N_5631,N_5719);
or U7310 (N_7310,N_5956,N_5412);
nor U7311 (N_7311,N_5381,N_5923);
nand U7312 (N_7312,N_5253,N_4210);
and U7313 (N_7313,N_5341,N_4103);
or U7314 (N_7314,N_4225,N_4585);
xor U7315 (N_7315,N_4297,N_5168);
nand U7316 (N_7316,N_4313,N_5016);
nand U7317 (N_7317,N_4156,N_4578);
and U7318 (N_7318,N_5459,N_5457);
and U7319 (N_7319,N_4694,N_5819);
and U7320 (N_7320,N_4212,N_5283);
and U7321 (N_7321,N_4097,N_5519);
xnor U7322 (N_7322,N_5174,N_4464);
or U7323 (N_7323,N_4726,N_5090);
xor U7324 (N_7324,N_5006,N_5072);
xor U7325 (N_7325,N_4188,N_5424);
nand U7326 (N_7326,N_4616,N_4843);
nand U7327 (N_7327,N_4554,N_4485);
and U7328 (N_7328,N_4150,N_4512);
nand U7329 (N_7329,N_5886,N_4776);
nand U7330 (N_7330,N_5632,N_4547);
nor U7331 (N_7331,N_4461,N_5189);
nor U7332 (N_7332,N_5186,N_4556);
and U7333 (N_7333,N_4836,N_4037);
xnor U7334 (N_7334,N_5353,N_5671);
and U7335 (N_7335,N_4596,N_5461);
xor U7336 (N_7336,N_5536,N_5353);
and U7337 (N_7337,N_4638,N_5024);
nor U7338 (N_7338,N_4796,N_5879);
xor U7339 (N_7339,N_4845,N_4590);
or U7340 (N_7340,N_5659,N_4299);
or U7341 (N_7341,N_4558,N_4928);
xor U7342 (N_7342,N_4899,N_4000);
or U7343 (N_7343,N_4794,N_5776);
or U7344 (N_7344,N_4620,N_5175);
xnor U7345 (N_7345,N_4540,N_5396);
or U7346 (N_7346,N_4436,N_4851);
xnor U7347 (N_7347,N_4782,N_4522);
and U7348 (N_7348,N_4930,N_5056);
nand U7349 (N_7349,N_5688,N_4081);
nor U7350 (N_7350,N_5743,N_5203);
or U7351 (N_7351,N_5058,N_4444);
or U7352 (N_7352,N_5356,N_5438);
nor U7353 (N_7353,N_4818,N_4076);
xnor U7354 (N_7354,N_5972,N_5731);
or U7355 (N_7355,N_5131,N_5752);
xor U7356 (N_7356,N_4627,N_4659);
nor U7357 (N_7357,N_4323,N_5655);
or U7358 (N_7358,N_5350,N_5670);
xor U7359 (N_7359,N_4123,N_4394);
or U7360 (N_7360,N_4606,N_5145);
or U7361 (N_7361,N_4601,N_4899);
nand U7362 (N_7362,N_4749,N_4299);
and U7363 (N_7363,N_5373,N_5128);
xor U7364 (N_7364,N_4834,N_4237);
or U7365 (N_7365,N_4732,N_5656);
nand U7366 (N_7366,N_5149,N_5104);
nor U7367 (N_7367,N_4956,N_5270);
and U7368 (N_7368,N_5358,N_5511);
and U7369 (N_7369,N_4872,N_5009);
or U7370 (N_7370,N_5319,N_4700);
and U7371 (N_7371,N_5694,N_5963);
and U7372 (N_7372,N_4400,N_5206);
nand U7373 (N_7373,N_5626,N_5025);
and U7374 (N_7374,N_4026,N_5035);
nand U7375 (N_7375,N_5201,N_5739);
nand U7376 (N_7376,N_5692,N_5746);
nor U7377 (N_7377,N_5799,N_5046);
nor U7378 (N_7378,N_5580,N_5965);
nor U7379 (N_7379,N_5485,N_4662);
and U7380 (N_7380,N_5040,N_5411);
and U7381 (N_7381,N_4001,N_5399);
or U7382 (N_7382,N_5845,N_5168);
or U7383 (N_7383,N_4114,N_4920);
or U7384 (N_7384,N_5889,N_5816);
xor U7385 (N_7385,N_5593,N_5912);
nor U7386 (N_7386,N_4964,N_5660);
and U7387 (N_7387,N_4412,N_5232);
nor U7388 (N_7388,N_4173,N_4023);
or U7389 (N_7389,N_5341,N_5768);
xor U7390 (N_7390,N_4019,N_4564);
or U7391 (N_7391,N_5225,N_4250);
nor U7392 (N_7392,N_5335,N_4329);
nor U7393 (N_7393,N_4554,N_4746);
and U7394 (N_7394,N_4577,N_4907);
and U7395 (N_7395,N_5835,N_4309);
xor U7396 (N_7396,N_4090,N_5456);
or U7397 (N_7397,N_5224,N_4153);
xnor U7398 (N_7398,N_5207,N_5552);
xnor U7399 (N_7399,N_5751,N_4731);
or U7400 (N_7400,N_4887,N_4640);
and U7401 (N_7401,N_4624,N_5172);
and U7402 (N_7402,N_4364,N_4623);
xor U7403 (N_7403,N_5909,N_4434);
or U7404 (N_7404,N_4166,N_5573);
nand U7405 (N_7405,N_5141,N_5906);
and U7406 (N_7406,N_4602,N_5878);
nor U7407 (N_7407,N_5842,N_4037);
or U7408 (N_7408,N_5880,N_5514);
xnor U7409 (N_7409,N_4818,N_4096);
and U7410 (N_7410,N_5908,N_4260);
nand U7411 (N_7411,N_5983,N_4825);
or U7412 (N_7412,N_4188,N_4160);
nor U7413 (N_7413,N_4504,N_5336);
nand U7414 (N_7414,N_4183,N_5961);
xor U7415 (N_7415,N_4329,N_5070);
nand U7416 (N_7416,N_4610,N_4361);
nand U7417 (N_7417,N_5239,N_4468);
nand U7418 (N_7418,N_5177,N_5275);
nor U7419 (N_7419,N_5305,N_4966);
nand U7420 (N_7420,N_4300,N_5963);
nand U7421 (N_7421,N_4322,N_5301);
xnor U7422 (N_7422,N_5682,N_5477);
nand U7423 (N_7423,N_4354,N_4671);
and U7424 (N_7424,N_5706,N_4956);
xnor U7425 (N_7425,N_5415,N_5234);
nor U7426 (N_7426,N_4631,N_5019);
nand U7427 (N_7427,N_5853,N_5518);
nand U7428 (N_7428,N_5554,N_4004);
or U7429 (N_7429,N_5195,N_5469);
xnor U7430 (N_7430,N_5892,N_5997);
and U7431 (N_7431,N_5514,N_5683);
and U7432 (N_7432,N_5475,N_5463);
xor U7433 (N_7433,N_4901,N_4956);
or U7434 (N_7434,N_5915,N_5433);
xor U7435 (N_7435,N_5190,N_4063);
or U7436 (N_7436,N_4470,N_5846);
or U7437 (N_7437,N_5753,N_5794);
or U7438 (N_7438,N_4151,N_4326);
nor U7439 (N_7439,N_5797,N_5137);
or U7440 (N_7440,N_5077,N_4170);
and U7441 (N_7441,N_5605,N_4252);
nand U7442 (N_7442,N_4744,N_5219);
and U7443 (N_7443,N_4047,N_5772);
or U7444 (N_7444,N_5007,N_4368);
and U7445 (N_7445,N_5827,N_4490);
or U7446 (N_7446,N_5197,N_4209);
or U7447 (N_7447,N_5204,N_4252);
xnor U7448 (N_7448,N_5154,N_4835);
nor U7449 (N_7449,N_4901,N_5815);
or U7450 (N_7450,N_5117,N_4366);
nor U7451 (N_7451,N_4450,N_5260);
nor U7452 (N_7452,N_5872,N_4864);
nand U7453 (N_7453,N_5236,N_5807);
nand U7454 (N_7454,N_4208,N_5722);
nor U7455 (N_7455,N_5591,N_5787);
and U7456 (N_7456,N_5062,N_5953);
and U7457 (N_7457,N_4701,N_4638);
or U7458 (N_7458,N_4469,N_4224);
or U7459 (N_7459,N_5328,N_5027);
nand U7460 (N_7460,N_4200,N_4276);
and U7461 (N_7461,N_5096,N_4003);
nand U7462 (N_7462,N_4940,N_5705);
xor U7463 (N_7463,N_5948,N_4753);
nor U7464 (N_7464,N_4984,N_4700);
or U7465 (N_7465,N_4921,N_4637);
nor U7466 (N_7466,N_4104,N_5773);
or U7467 (N_7467,N_4773,N_5807);
or U7468 (N_7468,N_4518,N_4066);
or U7469 (N_7469,N_4209,N_5599);
and U7470 (N_7470,N_5426,N_5919);
and U7471 (N_7471,N_4203,N_4807);
nand U7472 (N_7472,N_5222,N_5255);
xor U7473 (N_7473,N_4682,N_4625);
nor U7474 (N_7474,N_4265,N_5015);
or U7475 (N_7475,N_5252,N_5796);
or U7476 (N_7476,N_4026,N_4751);
nor U7477 (N_7477,N_4879,N_5097);
xor U7478 (N_7478,N_4018,N_4226);
or U7479 (N_7479,N_5296,N_5392);
nand U7480 (N_7480,N_5966,N_5191);
nand U7481 (N_7481,N_4493,N_5974);
and U7482 (N_7482,N_4265,N_4560);
and U7483 (N_7483,N_4841,N_4081);
or U7484 (N_7484,N_5571,N_5637);
nor U7485 (N_7485,N_5971,N_4069);
nor U7486 (N_7486,N_4582,N_5248);
nand U7487 (N_7487,N_5205,N_5366);
or U7488 (N_7488,N_4559,N_4648);
xor U7489 (N_7489,N_4235,N_5610);
and U7490 (N_7490,N_5317,N_4187);
and U7491 (N_7491,N_5965,N_4849);
nor U7492 (N_7492,N_5252,N_4275);
nand U7493 (N_7493,N_4246,N_5157);
nand U7494 (N_7494,N_4656,N_4674);
or U7495 (N_7495,N_5644,N_5972);
xnor U7496 (N_7496,N_5158,N_4693);
xor U7497 (N_7497,N_4547,N_4520);
and U7498 (N_7498,N_5239,N_4623);
and U7499 (N_7499,N_4394,N_4957);
nor U7500 (N_7500,N_4090,N_5328);
nor U7501 (N_7501,N_5338,N_5325);
xor U7502 (N_7502,N_5910,N_5413);
xor U7503 (N_7503,N_5789,N_4826);
or U7504 (N_7504,N_4922,N_4491);
or U7505 (N_7505,N_4045,N_4218);
nand U7506 (N_7506,N_5323,N_5826);
nor U7507 (N_7507,N_5956,N_5751);
and U7508 (N_7508,N_5293,N_4141);
nand U7509 (N_7509,N_5797,N_5574);
nand U7510 (N_7510,N_5005,N_5386);
and U7511 (N_7511,N_5294,N_4346);
and U7512 (N_7512,N_4958,N_4792);
nor U7513 (N_7513,N_4690,N_5226);
nand U7514 (N_7514,N_4998,N_4955);
nand U7515 (N_7515,N_4293,N_5104);
nor U7516 (N_7516,N_5457,N_5386);
and U7517 (N_7517,N_4612,N_5149);
nor U7518 (N_7518,N_5215,N_5285);
nand U7519 (N_7519,N_4227,N_5815);
nor U7520 (N_7520,N_5893,N_5022);
nand U7521 (N_7521,N_5662,N_5501);
nor U7522 (N_7522,N_5272,N_5003);
or U7523 (N_7523,N_5250,N_4439);
or U7524 (N_7524,N_4947,N_4908);
nor U7525 (N_7525,N_4523,N_5183);
or U7526 (N_7526,N_4341,N_5152);
or U7527 (N_7527,N_4316,N_5672);
and U7528 (N_7528,N_4584,N_4211);
nor U7529 (N_7529,N_4787,N_4180);
and U7530 (N_7530,N_5132,N_5574);
nand U7531 (N_7531,N_5479,N_4862);
nor U7532 (N_7532,N_4444,N_5107);
nand U7533 (N_7533,N_5049,N_4453);
or U7534 (N_7534,N_5718,N_5464);
nand U7535 (N_7535,N_4839,N_5830);
xor U7536 (N_7536,N_4758,N_5588);
or U7537 (N_7537,N_5282,N_4514);
xnor U7538 (N_7538,N_4804,N_4679);
nor U7539 (N_7539,N_5791,N_4208);
and U7540 (N_7540,N_5778,N_4254);
or U7541 (N_7541,N_4966,N_5416);
or U7542 (N_7542,N_4601,N_5218);
nor U7543 (N_7543,N_5582,N_5164);
and U7544 (N_7544,N_5952,N_4452);
nor U7545 (N_7545,N_4875,N_5147);
and U7546 (N_7546,N_5145,N_4503);
and U7547 (N_7547,N_4358,N_5251);
xor U7548 (N_7548,N_4275,N_5274);
or U7549 (N_7549,N_5322,N_4758);
xor U7550 (N_7550,N_4592,N_4494);
xnor U7551 (N_7551,N_5571,N_4534);
nor U7552 (N_7552,N_5110,N_4511);
nand U7553 (N_7553,N_4227,N_4566);
xor U7554 (N_7554,N_4263,N_5199);
or U7555 (N_7555,N_5532,N_4570);
xor U7556 (N_7556,N_4011,N_5743);
or U7557 (N_7557,N_4339,N_4875);
and U7558 (N_7558,N_5496,N_5309);
and U7559 (N_7559,N_5516,N_4235);
nor U7560 (N_7560,N_5957,N_5221);
and U7561 (N_7561,N_5688,N_5257);
and U7562 (N_7562,N_5577,N_5371);
and U7563 (N_7563,N_4598,N_4302);
and U7564 (N_7564,N_5189,N_4473);
xnor U7565 (N_7565,N_4592,N_4186);
xor U7566 (N_7566,N_4331,N_5699);
nand U7567 (N_7567,N_5837,N_5343);
and U7568 (N_7568,N_4549,N_4862);
nor U7569 (N_7569,N_4617,N_4655);
nand U7570 (N_7570,N_5206,N_4214);
xor U7571 (N_7571,N_4722,N_5291);
nand U7572 (N_7572,N_5020,N_4032);
nand U7573 (N_7573,N_4552,N_5490);
nand U7574 (N_7574,N_4313,N_4773);
or U7575 (N_7575,N_5413,N_4716);
and U7576 (N_7576,N_5752,N_4647);
and U7577 (N_7577,N_4377,N_5068);
or U7578 (N_7578,N_4892,N_5368);
nor U7579 (N_7579,N_5402,N_5383);
and U7580 (N_7580,N_4148,N_5332);
xnor U7581 (N_7581,N_4630,N_4260);
nand U7582 (N_7582,N_4920,N_4550);
or U7583 (N_7583,N_4892,N_4961);
xor U7584 (N_7584,N_5337,N_4318);
or U7585 (N_7585,N_4960,N_4415);
xor U7586 (N_7586,N_4093,N_5147);
xnor U7587 (N_7587,N_5185,N_4563);
or U7588 (N_7588,N_5661,N_5187);
nand U7589 (N_7589,N_5272,N_5972);
and U7590 (N_7590,N_4378,N_4543);
and U7591 (N_7591,N_4170,N_4887);
nor U7592 (N_7592,N_5284,N_5438);
nor U7593 (N_7593,N_4809,N_4896);
nand U7594 (N_7594,N_5096,N_4380);
nand U7595 (N_7595,N_4500,N_4288);
xor U7596 (N_7596,N_5702,N_5558);
or U7597 (N_7597,N_4611,N_5466);
xnor U7598 (N_7598,N_4364,N_5651);
and U7599 (N_7599,N_4656,N_5780);
and U7600 (N_7600,N_4007,N_5031);
xnor U7601 (N_7601,N_5439,N_4763);
or U7602 (N_7602,N_4677,N_4471);
and U7603 (N_7603,N_5874,N_5215);
or U7604 (N_7604,N_5541,N_5005);
xnor U7605 (N_7605,N_5182,N_5135);
and U7606 (N_7606,N_4297,N_5894);
xnor U7607 (N_7607,N_5523,N_4563);
or U7608 (N_7608,N_4602,N_5986);
and U7609 (N_7609,N_5990,N_5685);
or U7610 (N_7610,N_4634,N_4988);
and U7611 (N_7611,N_4116,N_4425);
nand U7612 (N_7612,N_5755,N_5967);
nand U7613 (N_7613,N_5765,N_5946);
or U7614 (N_7614,N_5568,N_4318);
or U7615 (N_7615,N_4486,N_4767);
nand U7616 (N_7616,N_4962,N_5232);
nand U7617 (N_7617,N_5693,N_4306);
nand U7618 (N_7618,N_4043,N_5191);
xnor U7619 (N_7619,N_4140,N_5083);
and U7620 (N_7620,N_5925,N_5124);
and U7621 (N_7621,N_4827,N_4561);
xnor U7622 (N_7622,N_4754,N_5133);
xnor U7623 (N_7623,N_5109,N_5092);
xnor U7624 (N_7624,N_5816,N_5741);
nor U7625 (N_7625,N_5142,N_4702);
or U7626 (N_7626,N_4044,N_5934);
xnor U7627 (N_7627,N_4573,N_5462);
or U7628 (N_7628,N_4461,N_4839);
nor U7629 (N_7629,N_4213,N_5618);
nand U7630 (N_7630,N_4202,N_5444);
xnor U7631 (N_7631,N_5572,N_5320);
or U7632 (N_7632,N_4602,N_5887);
nor U7633 (N_7633,N_4074,N_5350);
xor U7634 (N_7634,N_4283,N_5897);
nor U7635 (N_7635,N_5492,N_4953);
nand U7636 (N_7636,N_5184,N_4174);
xor U7637 (N_7637,N_4652,N_5260);
xor U7638 (N_7638,N_5210,N_4153);
nor U7639 (N_7639,N_4751,N_4373);
and U7640 (N_7640,N_4989,N_5507);
nor U7641 (N_7641,N_5172,N_5006);
xor U7642 (N_7642,N_4771,N_4669);
nand U7643 (N_7643,N_5397,N_5991);
nor U7644 (N_7644,N_5177,N_5658);
and U7645 (N_7645,N_4991,N_5308);
xor U7646 (N_7646,N_4107,N_5623);
or U7647 (N_7647,N_4368,N_5486);
xnor U7648 (N_7648,N_5034,N_5140);
xor U7649 (N_7649,N_5947,N_4083);
or U7650 (N_7650,N_5073,N_5742);
nand U7651 (N_7651,N_5317,N_4784);
or U7652 (N_7652,N_4856,N_5880);
and U7653 (N_7653,N_5680,N_5135);
and U7654 (N_7654,N_4747,N_5631);
xnor U7655 (N_7655,N_4309,N_5834);
xor U7656 (N_7656,N_5378,N_5163);
nand U7657 (N_7657,N_4501,N_4250);
nand U7658 (N_7658,N_5912,N_4911);
xor U7659 (N_7659,N_4350,N_5081);
or U7660 (N_7660,N_4315,N_5328);
or U7661 (N_7661,N_4696,N_4105);
xor U7662 (N_7662,N_5416,N_4750);
nand U7663 (N_7663,N_5366,N_5902);
and U7664 (N_7664,N_4009,N_4604);
nor U7665 (N_7665,N_4071,N_4805);
and U7666 (N_7666,N_5405,N_4826);
or U7667 (N_7667,N_5415,N_5525);
nor U7668 (N_7668,N_4764,N_5811);
nand U7669 (N_7669,N_5552,N_5098);
nor U7670 (N_7670,N_4191,N_5780);
nor U7671 (N_7671,N_4046,N_5366);
and U7672 (N_7672,N_5158,N_5768);
and U7673 (N_7673,N_4874,N_5665);
and U7674 (N_7674,N_5567,N_5831);
nor U7675 (N_7675,N_5041,N_5305);
nor U7676 (N_7676,N_5428,N_5224);
nand U7677 (N_7677,N_5746,N_5728);
nor U7678 (N_7678,N_4542,N_4590);
nor U7679 (N_7679,N_4314,N_4033);
and U7680 (N_7680,N_4346,N_4772);
and U7681 (N_7681,N_4677,N_5212);
or U7682 (N_7682,N_5935,N_4750);
nor U7683 (N_7683,N_5023,N_4355);
or U7684 (N_7684,N_4655,N_5722);
xor U7685 (N_7685,N_5145,N_5967);
xnor U7686 (N_7686,N_4836,N_4888);
nand U7687 (N_7687,N_4279,N_5214);
and U7688 (N_7688,N_4225,N_5263);
nor U7689 (N_7689,N_5749,N_4087);
xnor U7690 (N_7690,N_4310,N_5492);
or U7691 (N_7691,N_4661,N_5974);
xor U7692 (N_7692,N_4671,N_4058);
nor U7693 (N_7693,N_4148,N_5561);
nor U7694 (N_7694,N_5154,N_5439);
nand U7695 (N_7695,N_5634,N_5406);
xor U7696 (N_7696,N_4226,N_5140);
nor U7697 (N_7697,N_4373,N_5888);
nand U7698 (N_7698,N_4579,N_4282);
xor U7699 (N_7699,N_5814,N_4285);
or U7700 (N_7700,N_5753,N_4787);
or U7701 (N_7701,N_5644,N_5159);
nand U7702 (N_7702,N_5764,N_5645);
nor U7703 (N_7703,N_5300,N_4711);
nor U7704 (N_7704,N_5303,N_4969);
nor U7705 (N_7705,N_5426,N_5718);
and U7706 (N_7706,N_5347,N_4790);
or U7707 (N_7707,N_5820,N_5517);
nor U7708 (N_7708,N_4837,N_4480);
xor U7709 (N_7709,N_4383,N_4690);
nor U7710 (N_7710,N_5048,N_4523);
or U7711 (N_7711,N_4565,N_4209);
xor U7712 (N_7712,N_5420,N_5176);
and U7713 (N_7713,N_5835,N_5076);
and U7714 (N_7714,N_5696,N_5272);
nand U7715 (N_7715,N_5307,N_5112);
nand U7716 (N_7716,N_5496,N_5958);
and U7717 (N_7717,N_4458,N_5431);
nand U7718 (N_7718,N_5816,N_4107);
nor U7719 (N_7719,N_4562,N_4427);
and U7720 (N_7720,N_4723,N_4845);
and U7721 (N_7721,N_4219,N_5069);
nand U7722 (N_7722,N_4371,N_4607);
nor U7723 (N_7723,N_4328,N_4274);
or U7724 (N_7724,N_5996,N_5303);
and U7725 (N_7725,N_4446,N_4409);
nor U7726 (N_7726,N_5163,N_5476);
xor U7727 (N_7727,N_5890,N_4135);
nor U7728 (N_7728,N_5084,N_4978);
xnor U7729 (N_7729,N_4878,N_5619);
nand U7730 (N_7730,N_4106,N_5064);
nor U7731 (N_7731,N_5606,N_4209);
and U7732 (N_7732,N_5601,N_4397);
and U7733 (N_7733,N_5987,N_4005);
nand U7734 (N_7734,N_4406,N_4278);
xnor U7735 (N_7735,N_5000,N_4727);
and U7736 (N_7736,N_5227,N_4700);
and U7737 (N_7737,N_5949,N_5337);
and U7738 (N_7738,N_4049,N_5920);
nor U7739 (N_7739,N_4115,N_4958);
and U7740 (N_7740,N_5288,N_4547);
nor U7741 (N_7741,N_4692,N_5967);
xor U7742 (N_7742,N_5894,N_4977);
xor U7743 (N_7743,N_5596,N_5540);
and U7744 (N_7744,N_5318,N_4696);
nand U7745 (N_7745,N_5395,N_5223);
nor U7746 (N_7746,N_4322,N_4541);
nor U7747 (N_7747,N_5210,N_4329);
and U7748 (N_7748,N_4826,N_4410);
nand U7749 (N_7749,N_4792,N_5937);
nand U7750 (N_7750,N_4462,N_4381);
nor U7751 (N_7751,N_5080,N_5723);
nor U7752 (N_7752,N_4807,N_4416);
nor U7753 (N_7753,N_4995,N_4454);
nor U7754 (N_7754,N_4742,N_4939);
or U7755 (N_7755,N_5853,N_5064);
and U7756 (N_7756,N_4172,N_4895);
nor U7757 (N_7757,N_5884,N_5833);
nor U7758 (N_7758,N_4143,N_5262);
and U7759 (N_7759,N_5360,N_4086);
nand U7760 (N_7760,N_5689,N_5669);
xnor U7761 (N_7761,N_4417,N_5218);
or U7762 (N_7762,N_4465,N_4044);
or U7763 (N_7763,N_5941,N_4404);
and U7764 (N_7764,N_5005,N_5736);
nand U7765 (N_7765,N_4096,N_4200);
nand U7766 (N_7766,N_5371,N_5916);
nand U7767 (N_7767,N_5712,N_4138);
xnor U7768 (N_7768,N_4639,N_5114);
nand U7769 (N_7769,N_5372,N_4262);
nor U7770 (N_7770,N_5051,N_4174);
nand U7771 (N_7771,N_4960,N_4241);
nand U7772 (N_7772,N_5937,N_4940);
xor U7773 (N_7773,N_4744,N_5323);
and U7774 (N_7774,N_4528,N_4507);
nor U7775 (N_7775,N_5686,N_5648);
and U7776 (N_7776,N_5121,N_4666);
nand U7777 (N_7777,N_4644,N_5654);
nand U7778 (N_7778,N_5187,N_4515);
xor U7779 (N_7779,N_5450,N_5650);
or U7780 (N_7780,N_5211,N_5113);
xor U7781 (N_7781,N_5650,N_4859);
and U7782 (N_7782,N_5308,N_5852);
nand U7783 (N_7783,N_5398,N_4565);
or U7784 (N_7784,N_5587,N_5787);
and U7785 (N_7785,N_5509,N_5662);
nor U7786 (N_7786,N_4132,N_5261);
or U7787 (N_7787,N_4231,N_5052);
or U7788 (N_7788,N_4274,N_4907);
xor U7789 (N_7789,N_5127,N_5753);
nor U7790 (N_7790,N_4747,N_4283);
or U7791 (N_7791,N_5389,N_4327);
nand U7792 (N_7792,N_5785,N_5643);
or U7793 (N_7793,N_5596,N_4229);
nor U7794 (N_7794,N_4493,N_4921);
nor U7795 (N_7795,N_5446,N_5368);
xor U7796 (N_7796,N_5709,N_4168);
xnor U7797 (N_7797,N_4928,N_5309);
nand U7798 (N_7798,N_5807,N_5392);
nor U7799 (N_7799,N_5185,N_4692);
xnor U7800 (N_7800,N_4886,N_5848);
nand U7801 (N_7801,N_5171,N_4766);
nand U7802 (N_7802,N_5743,N_4907);
nor U7803 (N_7803,N_4712,N_4575);
nand U7804 (N_7804,N_4943,N_5121);
nand U7805 (N_7805,N_4229,N_5709);
and U7806 (N_7806,N_4044,N_5208);
or U7807 (N_7807,N_5025,N_4446);
or U7808 (N_7808,N_4541,N_4511);
and U7809 (N_7809,N_4776,N_4494);
nand U7810 (N_7810,N_4877,N_5322);
nor U7811 (N_7811,N_4376,N_5397);
xnor U7812 (N_7812,N_5741,N_4105);
xnor U7813 (N_7813,N_5008,N_4520);
nor U7814 (N_7814,N_5514,N_5110);
and U7815 (N_7815,N_5689,N_4410);
nor U7816 (N_7816,N_5721,N_4894);
nand U7817 (N_7817,N_4477,N_5961);
nand U7818 (N_7818,N_4534,N_5265);
and U7819 (N_7819,N_4270,N_4057);
nor U7820 (N_7820,N_5525,N_4563);
or U7821 (N_7821,N_5716,N_5925);
nand U7822 (N_7822,N_5699,N_5448);
xnor U7823 (N_7823,N_4917,N_4018);
xnor U7824 (N_7824,N_5665,N_5235);
nand U7825 (N_7825,N_4954,N_4318);
nand U7826 (N_7826,N_5883,N_4312);
nor U7827 (N_7827,N_4090,N_4801);
and U7828 (N_7828,N_5104,N_5143);
and U7829 (N_7829,N_5904,N_5331);
or U7830 (N_7830,N_4168,N_5641);
or U7831 (N_7831,N_4198,N_4798);
or U7832 (N_7832,N_4826,N_4560);
nand U7833 (N_7833,N_5305,N_4707);
xor U7834 (N_7834,N_5360,N_5180);
xor U7835 (N_7835,N_4972,N_5221);
or U7836 (N_7836,N_4269,N_5391);
nand U7837 (N_7837,N_4534,N_5425);
nand U7838 (N_7838,N_4652,N_5089);
nor U7839 (N_7839,N_4391,N_5802);
nor U7840 (N_7840,N_5847,N_4199);
nand U7841 (N_7841,N_5910,N_5780);
xnor U7842 (N_7842,N_4726,N_5122);
xnor U7843 (N_7843,N_4025,N_5410);
xor U7844 (N_7844,N_5178,N_4319);
nand U7845 (N_7845,N_5417,N_4504);
or U7846 (N_7846,N_4953,N_5455);
or U7847 (N_7847,N_5206,N_4157);
xor U7848 (N_7848,N_4679,N_4382);
and U7849 (N_7849,N_5054,N_4784);
and U7850 (N_7850,N_5324,N_4231);
xnor U7851 (N_7851,N_5309,N_4221);
and U7852 (N_7852,N_4051,N_5553);
nand U7853 (N_7853,N_4053,N_5128);
xor U7854 (N_7854,N_5785,N_5260);
or U7855 (N_7855,N_5659,N_5726);
nand U7856 (N_7856,N_5170,N_4923);
and U7857 (N_7857,N_4637,N_4135);
nand U7858 (N_7858,N_4988,N_4836);
nor U7859 (N_7859,N_5424,N_5329);
or U7860 (N_7860,N_4168,N_4809);
and U7861 (N_7861,N_4917,N_4709);
xnor U7862 (N_7862,N_4705,N_5017);
nand U7863 (N_7863,N_4843,N_5815);
nor U7864 (N_7864,N_4516,N_5828);
or U7865 (N_7865,N_4090,N_4120);
nand U7866 (N_7866,N_5021,N_5942);
xnor U7867 (N_7867,N_4082,N_5864);
nor U7868 (N_7868,N_4135,N_5763);
nand U7869 (N_7869,N_5037,N_4918);
nand U7870 (N_7870,N_5485,N_4846);
nand U7871 (N_7871,N_5903,N_5300);
nor U7872 (N_7872,N_5980,N_4570);
and U7873 (N_7873,N_4661,N_4467);
xnor U7874 (N_7874,N_4262,N_4271);
xor U7875 (N_7875,N_4884,N_5846);
or U7876 (N_7876,N_5562,N_5871);
xor U7877 (N_7877,N_4389,N_4395);
and U7878 (N_7878,N_4903,N_4651);
or U7879 (N_7879,N_5888,N_5412);
nor U7880 (N_7880,N_4561,N_4880);
xor U7881 (N_7881,N_5551,N_4491);
or U7882 (N_7882,N_4242,N_5963);
nor U7883 (N_7883,N_5034,N_4471);
or U7884 (N_7884,N_4085,N_4116);
nor U7885 (N_7885,N_4429,N_5832);
nor U7886 (N_7886,N_5194,N_4709);
xor U7887 (N_7887,N_5673,N_4018);
xnor U7888 (N_7888,N_5680,N_4695);
xor U7889 (N_7889,N_5807,N_4398);
or U7890 (N_7890,N_5062,N_5978);
xnor U7891 (N_7891,N_4273,N_5363);
xor U7892 (N_7892,N_5573,N_5856);
or U7893 (N_7893,N_5718,N_5134);
xnor U7894 (N_7894,N_5228,N_4043);
and U7895 (N_7895,N_5441,N_5014);
nand U7896 (N_7896,N_4802,N_5645);
and U7897 (N_7897,N_5995,N_5291);
and U7898 (N_7898,N_5734,N_5139);
or U7899 (N_7899,N_5581,N_4929);
or U7900 (N_7900,N_5698,N_5730);
xnor U7901 (N_7901,N_5220,N_4281);
nand U7902 (N_7902,N_5970,N_5942);
nor U7903 (N_7903,N_5150,N_5820);
nor U7904 (N_7904,N_5166,N_4207);
xnor U7905 (N_7905,N_5917,N_4520);
nand U7906 (N_7906,N_4982,N_5472);
or U7907 (N_7907,N_4295,N_5092);
and U7908 (N_7908,N_5671,N_5586);
or U7909 (N_7909,N_5578,N_4180);
xnor U7910 (N_7910,N_4006,N_4558);
or U7911 (N_7911,N_4662,N_4710);
xor U7912 (N_7912,N_4388,N_5770);
nor U7913 (N_7913,N_4465,N_5054);
or U7914 (N_7914,N_5042,N_5892);
xor U7915 (N_7915,N_5400,N_5712);
and U7916 (N_7916,N_4888,N_5351);
xnor U7917 (N_7917,N_5586,N_4182);
and U7918 (N_7918,N_4916,N_5665);
nor U7919 (N_7919,N_5135,N_5751);
xor U7920 (N_7920,N_5470,N_4577);
nor U7921 (N_7921,N_4045,N_5950);
nor U7922 (N_7922,N_5706,N_5191);
nand U7923 (N_7923,N_4664,N_4471);
nor U7924 (N_7924,N_5151,N_4692);
and U7925 (N_7925,N_5090,N_4134);
and U7926 (N_7926,N_4206,N_4958);
and U7927 (N_7927,N_4247,N_5963);
xnor U7928 (N_7928,N_5961,N_5191);
nand U7929 (N_7929,N_4793,N_5681);
and U7930 (N_7930,N_4336,N_5226);
nand U7931 (N_7931,N_4390,N_5582);
and U7932 (N_7932,N_5379,N_5117);
xnor U7933 (N_7933,N_5357,N_5111);
nand U7934 (N_7934,N_5527,N_4036);
xnor U7935 (N_7935,N_5600,N_5405);
nor U7936 (N_7936,N_4746,N_4081);
nand U7937 (N_7937,N_5808,N_5864);
and U7938 (N_7938,N_5279,N_4456);
nor U7939 (N_7939,N_5609,N_4032);
or U7940 (N_7940,N_4442,N_5604);
or U7941 (N_7941,N_5768,N_4753);
nor U7942 (N_7942,N_4787,N_5117);
xor U7943 (N_7943,N_5827,N_4609);
or U7944 (N_7944,N_4311,N_5156);
nand U7945 (N_7945,N_4050,N_4651);
and U7946 (N_7946,N_4033,N_5101);
xnor U7947 (N_7947,N_5430,N_4440);
and U7948 (N_7948,N_5478,N_4775);
nor U7949 (N_7949,N_5873,N_5969);
nand U7950 (N_7950,N_5910,N_4912);
and U7951 (N_7951,N_5836,N_5694);
or U7952 (N_7952,N_5427,N_4630);
or U7953 (N_7953,N_4404,N_4263);
nor U7954 (N_7954,N_4196,N_5965);
and U7955 (N_7955,N_4005,N_5606);
nor U7956 (N_7956,N_5634,N_4265);
nand U7957 (N_7957,N_5297,N_5229);
nand U7958 (N_7958,N_4982,N_5681);
and U7959 (N_7959,N_4557,N_4830);
xnor U7960 (N_7960,N_4192,N_5492);
or U7961 (N_7961,N_4279,N_4359);
and U7962 (N_7962,N_4467,N_5430);
xnor U7963 (N_7963,N_5066,N_5909);
nor U7964 (N_7964,N_4652,N_5667);
nand U7965 (N_7965,N_5305,N_5768);
nand U7966 (N_7966,N_4264,N_4265);
nand U7967 (N_7967,N_5280,N_5419);
nand U7968 (N_7968,N_5699,N_4069);
xor U7969 (N_7969,N_5758,N_5688);
nand U7970 (N_7970,N_5935,N_4988);
xor U7971 (N_7971,N_4130,N_4124);
xor U7972 (N_7972,N_5753,N_5186);
xor U7973 (N_7973,N_5116,N_4481);
xor U7974 (N_7974,N_5877,N_5197);
or U7975 (N_7975,N_5965,N_4417);
and U7976 (N_7976,N_4184,N_4002);
and U7977 (N_7977,N_5280,N_5071);
and U7978 (N_7978,N_5911,N_4821);
nand U7979 (N_7979,N_4204,N_5184);
xor U7980 (N_7980,N_5975,N_4973);
and U7981 (N_7981,N_4624,N_5214);
and U7982 (N_7982,N_4384,N_4460);
or U7983 (N_7983,N_5188,N_4535);
and U7984 (N_7984,N_5356,N_4695);
and U7985 (N_7985,N_5213,N_4980);
and U7986 (N_7986,N_4155,N_4682);
and U7987 (N_7987,N_5421,N_4781);
or U7988 (N_7988,N_5054,N_5805);
nand U7989 (N_7989,N_4573,N_4631);
nor U7990 (N_7990,N_5365,N_5930);
and U7991 (N_7991,N_4076,N_4936);
or U7992 (N_7992,N_4574,N_5877);
nor U7993 (N_7993,N_4877,N_5228);
xnor U7994 (N_7994,N_5375,N_4556);
and U7995 (N_7995,N_5600,N_4286);
or U7996 (N_7996,N_4526,N_5078);
nor U7997 (N_7997,N_5075,N_4158);
nor U7998 (N_7998,N_4386,N_5312);
and U7999 (N_7999,N_4965,N_5782);
or U8000 (N_8000,N_7118,N_6405);
nand U8001 (N_8001,N_6656,N_6657);
nor U8002 (N_8002,N_7822,N_7471);
nand U8003 (N_8003,N_7314,N_6203);
or U8004 (N_8004,N_6160,N_6000);
and U8005 (N_8005,N_6157,N_6618);
or U8006 (N_8006,N_7240,N_6635);
nor U8007 (N_8007,N_7417,N_6577);
xor U8008 (N_8008,N_6295,N_7920);
xnor U8009 (N_8009,N_6254,N_7651);
nand U8010 (N_8010,N_7156,N_7371);
or U8011 (N_8011,N_7015,N_7835);
and U8012 (N_8012,N_6463,N_7029);
or U8013 (N_8013,N_7621,N_7506);
or U8014 (N_8014,N_7923,N_6630);
or U8015 (N_8015,N_6015,N_6290);
and U8016 (N_8016,N_6883,N_7250);
xor U8017 (N_8017,N_6511,N_6029);
or U8018 (N_8018,N_7768,N_6143);
nor U8019 (N_8019,N_6934,N_6425);
nor U8020 (N_8020,N_7065,N_7262);
xor U8021 (N_8021,N_6276,N_7280);
nand U8022 (N_8022,N_7163,N_7007);
nand U8023 (N_8023,N_6146,N_7339);
or U8024 (N_8024,N_7806,N_6447);
and U8025 (N_8025,N_7890,N_6600);
xnor U8026 (N_8026,N_6858,N_6815);
xnor U8027 (N_8027,N_6662,N_6011);
and U8028 (N_8028,N_6754,N_6768);
or U8029 (N_8029,N_6285,N_7529);
or U8030 (N_8030,N_6536,N_6046);
nor U8031 (N_8031,N_7041,N_6386);
or U8032 (N_8032,N_6054,N_6204);
or U8033 (N_8033,N_7964,N_6082);
nand U8034 (N_8034,N_7660,N_7642);
or U8035 (N_8035,N_6636,N_7242);
nor U8036 (N_8036,N_6987,N_7000);
and U8037 (N_8037,N_7198,N_6352);
xnor U8038 (N_8038,N_7539,N_6264);
nor U8039 (N_8039,N_6691,N_6003);
nor U8040 (N_8040,N_6225,N_7188);
and U8041 (N_8041,N_7721,N_6593);
nand U8042 (N_8042,N_7450,N_7828);
and U8043 (N_8043,N_7808,N_6108);
or U8044 (N_8044,N_6701,N_6296);
or U8045 (N_8045,N_6414,N_7243);
nor U8046 (N_8046,N_6823,N_7310);
nand U8047 (N_8047,N_7357,N_6240);
and U8048 (N_8048,N_7291,N_6783);
or U8049 (N_8049,N_7845,N_6497);
xor U8050 (N_8050,N_6266,N_6098);
and U8051 (N_8051,N_6931,N_7916);
nand U8052 (N_8052,N_6149,N_7825);
nor U8053 (N_8053,N_6210,N_6507);
nor U8054 (N_8054,N_6299,N_7360);
nor U8055 (N_8055,N_7930,N_6742);
nand U8056 (N_8056,N_6661,N_6592);
or U8057 (N_8057,N_6455,N_7879);
or U8058 (N_8058,N_7810,N_7018);
nand U8059 (N_8059,N_7998,N_7337);
or U8060 (N_8060,N_6229,N_6523);
or U8061 (N_8061,N_7988,N_6840);
nand U8062 (N_8062,N_6698,N_6695);
or U8063 (N_8063,N_7862,N_7716);
and U8064 (N_8064,N_7790,N_6867);
nand U8065 (N_8065,N_6647,N_6492);
nand U8066 (N_8066,N_6154,N_7286);
or U8067 (N_8067,N_7372,N_6104);
xnor U8068 (N_8068,N_6936,N_7281);
nor U8069 (N_8069,N_6216,N_6699);
xor U8070 (N_8070,N_7535,N_6394);
nor U8071 (N_8071,N_7048,N_6306);
xor U8072 (N_8072,N_7678,N_6268);
xnor U8073 (N_8073,N_6800,N_7134);
nor U8074 (N_8074,N_7781,N_7246);
and U8075 (N_8075,N_6803,N_7207);
and U8076 (N_8076,N_6179,N_7638);
xnor U8077 (N_8077,N_6366,N_7206);
and U8078 (N_8078,N_6688,N_7072);
nor U8079 (N_8079,N_7389,N_6059);
and U8080 (N_8080,N_6186,N_6498);
nand U8081 (N_8081,N_7510,N_6176);
xor U8082 (N_8082,N_6850,N_7724);
or U8083 (N_8083,N_7353,N_6704);
nor U8084 (N_8084,N_7616,N_7555);
or U8085 (N_8085,N_6966,N_7715);
xnor U8086 (N_8086,N_7472,N_7871);
xnor U8087 (N_8087,N_6779,N_6416);
and U8088 (N_8088,N_6709,N_7123);
and U8089 (N_8089,N_6866,N_7269);
nor U8090 (N_8090,N_6017,N_7965);
xor U8091 (N_8091,N_7222,N_7384);
nor U8092 (N_8092,N_7053,N_6617);
nor U8093 (N_8093,N_6300,N_7159);
xnor U8094 (N_8094,N_6232,N_7830);
xor U8095 (N_8095,N_6193,N_7312);
nand U8096 (N_8096,N_7729,N_7838);
or U8097 (N_8097,N_7549,N_7869);
and U8098 (N_8098,N_6608,N_7829);
nand U8099 (N_8099,N_6342,N_6144);
xnor U8100 (N_8100,N_7058,N_7500);
or U8101 (N_8101,N_7001,N_6245);
or U8102 (N_8102,N_7152,N_6317);
xor U8103 (N_8103,N_7338,N_6753);
xnor U8104 (N_8104,N_6215,N_7727);
xor U8105 (N_8105,N_6616,N_7753);
nor U8106 (N_8106,N_7073,N_7897);
and U8107 (N_8107,N_6458,N_6786);
or U8108 (N_8108,N_7725,N_6591);
nor U8109 (N_8109,N_7199,N_7573);
nor U8110 (N_8110,N_7287,N_7665);
nor U8111 (N_8111,N_6838,N_7276);
nor U8112 (N_8112,N_6814,N_6465);
xor U8113 (N_8113,N_7027,N_6664);
xor U8114 (N_8114,N_6148,N_6621);
nor U8115 (N_8115,N_7074,N_7764);
nand U8116 (N_8116,N_7225,N_6963);
nand U8117 (N_8117,N_6911,N_7478);
xor U8118 (N_8118,N_6622,N_6192);
nor U8119 (N_8119,N_7900,N_6286);
nand U8120 (N_8120,N_6520,N_6065);
and U8121 (N_8121,N_7083,N_6354);
nor U8122 (N_8122,N_7905,N_6989);
nand U8123 (N_8123,N_7311,N_6727);
nor U8124 (N_8124,N_6522,N_7590);
or U8125 (N_8125,N_7346,N_7003);
and U8126 (N_8126,N_7087,N_6234);
xnor U8127 (N_8127,N_7336,N_7610);
xor U8128 (N_8128,N_7615,N_6693);
or U8129 (N_8129,N_7982,N_6977);
and U8130 (N_8130,N_7775,N_7130);
or U8131 (N_8131,N_7558,N_7398);
and U8132 (N_8132,N_6561,N_7426);
nand U8133 (N_8133,N_7100,N_7416);
nor U8134 (N_8134,N_6620,N_6150);
xor U8135 (N_8135,N_6272,N_6574);
nor U8136 (N_8136,N_6292,N_6023);
and U8137 (N_8137,N_6832,N_6315);
nand U8138 (N_8138,N_6820,N_7388);
and U8139 (N_8139,N_7076,N_6161);
nor U8140 (N_8140,N_7889,N_6269);
and U8141 (N_8141,N_6393,N_6928);
nand U8142 (N_8142,N_6220,N_7435);
nand U8143 (N_8143,N_6380,N_6588);
and U8144 (N_8144,N_6095,N_6728);
or U8145 (N_8145,N_7801,N_7523);
nand U8146 (N_8146,N_6787,N_7846);
nor U8147 (N_8147,N_7881,N_6532);
xor U8148 (N_8148,N_7304,N_6951);
nand U8149 (N_8149,N_6848,N_7141);
nand U8150 (N_8150,N_6710,N_7180);
and U8151 (N_8151,N_6667,N_6093);
or U8152 (N_8152,N_7369,N_6795);
nor U8153 (N_8153,N_6159,N_6646);
and U8154 (N_8154,N_7874,N_6469);
xor U8155 (N_8155,N_6898,N_7238);
and U8156 (N_8156,N_6674,N_7751);
nor U8157 (N_8157,N_7170,N_7814);
and U8158 (N_8158,N_7819,N_6696);
nand U8159 (N_8159,N_6196,N_7972);
nor U8160 (N_8160,N_6938,N_7359);
nand U8161 (N_8161,N_6756,N_7200);
or U8162 (N_8162,N_6995,N_7750);
nor U8163 (N_8163,N_7030,N_7902);
nand U8164 (N_8164,N_6810,N_7096);
or U8165 (N_8165,N_6175,N_6164);
xor U8166 (N_8166,N_6933,N_7386);
nor U8167 (N_8167,N_7383,N_6700);
xor U8168 (N_8168,N_7974,N_6340);
xnor U8169 (N_8169,N_7899,N_6547);
nand U8170 (N_8170,N_6861,N_7533);
nand U8171 (N_8171,N_6399,N_6729);
or U8172 (N_8172,N_7632,N_7832);
xnor U8173 (N_8173,N_6505,N_6530);
xnor U8174 (N_8174,N_6835,N_7347);
xnor U8175 (N_8175,N_6055,N_6542);
xnor U8176 (N_8176,N_7016,N_6859);
and U8177 (N_8177,N_7758,N_7301);
xnor U8178 (N_8178,N_6402,N_7955);
nand U8179 (N_8179,N_6822,N_6604);
nor U8180 (N_8180,N_7315,N_6002);
xnor U8181 (N_8181,N_7184,N_7161);
or U8182 (N_8182,N_7348,N_7462);
xor U8183 (N_8183,N_6706,N_7952);
xor U8184 (N_8184,N_7335,N_7865);
nand U8185 (N_8185,N_6279,N_6680);
xor U8186 (N_8186,N_7979,N_6641);
nand U8187 (N_8187,N_7052,N_6271);
nor U8188 (N_8188,N_7668,N_7517);
or U8189 (N_8189,N_7316,N_6723);
xnor U8190 (N_8190,N_6298,N_6854);
nor U8191 (N_8191,N_7444,N_6576);
xnor U8192 (N_8192,N_7425,N_7913);
nor U8193 (N_8193,N_6156,N_7547);
nor U8194 (N_8194,N_7989,N_6813);
nand U8195 (N_8195,N_6006,N_6589);
or U8196 (N_8196,N_7625,N_6287);
nor U8197 (N_8197,N_6501,N_7367);
and U8198 (N_8198,N_7319,N_7994);
or U8199 (N_8199,N_7142,N_7635);
nor U8200 (N_8200,N_6255,N_7609);
or U8201 (N_8201,N_7875,N_6111);
nor U8202 (N_8202,N_7449,N_7205);
nand U8203 (N_8203,N_6844,N_6797);
and U8204 (N_8204,N_6304,N_6560);
nand U8205 (N_8205,N_6128,N_7396);
nand U8206 (N_8206,N_7581,N_7707);
and U8207 (N_8207,N_7543,N_6294);
nor U8208 (N_8208,N_6750,N_7731);
nand U8209 (N_8209,N_6929,N_7737);
nand U8210 (N_8210,N_6598,N_7231);
nor U8211 (N_8211,N_7672,N_7299);
and U8212 (N_8212,N_6716,N_7748);
nand U8213 (N_8213,N_6894,N_6913);
nand U8214 (N_8214,N_6022,N_7309);
and U8215 (N_8215,N_6714,N_7933);
nor U8216 (N_8216,N_7230,N_6889);
or U8217 (N_8217,N_6058,N_6243);
nor U8218 (N_8218,N_6280,N_7241);
and U8219 (N_8219,N_6430,N_6955);
and U8220 (N_8220,N_6774,N_6817);
and U8221 (N_8221,N_7631,N_6660);
nor U8222 (N_8222,N_7483,N_6169);
nor U8223 (N_8223,N_7976,N_6663);
and U8224 (N_8224,N_7894,N_7585);
or U8225 (N_8225,N_7352,N_7203);
and U8226 (N_8226,N_6615,N_7214);
xnor U8227 (N_8227,N_6719,N_6401);
nand U8228 (N_8228,N_7518,N_7597);
nor U8229 (N_8229,N_6624,N_7308);
or U8230 (N_8230,N_6671,N_6816);
nor U8231 (N_8231,N_6921,N_7447);
nand U8232 (N_8232,N_7767,N_6993);
xor U8233 (N_8233,N_7834,N_6811);
and U8234 (N_8234,N_7612,N_7049);
and U8235 (N_8235,N_6796,N_6632);
nand U8236 (N_8236,N_7823,N_6431);
and U8237 (N_8237,N_6089,N_6760);
nand U8238 (N_8238,N_6724,N_7971);
or U8239 (N_8239,N_6348,N_6263);
xor U8240 (N_8240,N_7996,N_7436);
xor U8241 (N_8241,N_7811,N_7962);
xor U8242 (N_8242,N_7224,N_7582);
and U8243 (N_8243,N_7694,N_7826);
or U8244 (N_8244,N_6182,N_7006);
xnor U8245 (N_8245,N_7204,N_6311);
or U8246 (N_8246,N_6368,N_6676);
xnor U8247 (N_8247,N_7085,N_7605);
xor U8248 (N_8248,N_6557,N_6361);
nand U8249 (N_8249,N_6666,N_6759);
and U8250 (N_8250,N_6328,N_6551);
or U8251 (N_8251,N_7486,N_7508);
and U8252 (N_8252,N_7567,N_6445);
or U8253 (N_8253,N_6812,N_7749);
and U8254 (N_8254,N_6851,N_6106);
or U8255 (N_8255,N_7370,N_7321);
xor U8256 (N_8256,N_6923,N_7010);
or U8257 (N_8257,N_7968,N_7734);
or U8258 (N_8258,N_7057,N_6491);
and U8259 (N_8259,N_7192,N_6969);
nor U8260 (N_8260,N_6440,N_6241);
nor U8261 (N_8261,N_6071,N_6376);
or U8262 (N_8262,N_6162,N_6310);
and U8263 (N_8263,N_7466,N_6749);
xnor U8264 (N_8264,N_6541,N_7685);
nor U8265 (N_8265,N_7710,N_7218);
and U8266 (N_8266,N_6433,N_6504);
xnor U8267 (N_8267,N_6423,N_6490);
nor U8268 (N_8268,N_6101,N_6322);
or U8269 (N_8269,N_6238,N_6484);
nand U8270 (N_8270,N_7324,N_6262);
or U8271 (N_8271,N_7220,N_7233);
and U8272 (N_8272,N_6733,N_6439);
xnor U8273 (N_8273,N_7151,N_6201);
xnor U8274 (N_8274,N_6946,N_7634);
and U8275 (N_8275,N_7940,N_6045);
or U8276 (N_8276,N_6606,N_7528);
nor U8277 (N_8277,N_7780,N_6471);
and U8278 (N_8278,N_6183,N_6605);
and U8279 (N_8279,N_7591,N_7714);
and U8280 (N_8280,N_7244,N_7410);
xor U8281 (N_8281,N_6918,N_6222);
nand U8282 (N_8282,N_7643,N_6525);
nand U8283 (N_8283,N_7226,N_6109);
or U8284 (N_8284,N_7429,N_7223);
nor U8285 (N_8285,N_6968,N_6556);
nor U8286 (N_8286,N_6387,N_7211);
or U8287 (N_8287,N_7385,N_7494);
nor U8288 (N_8288,N_6078,N_6697);
nor U8289 (N_8289,N_6199,N_7300);
nand U8290 (N_8290,N_6195,N_6964);
nor U8291 (N_8291,N_7068,N_7927);
nor U8292 (N_8292,N_7926,N_7329);
and U8293 (N_8293,N_7005,N_6367);
xnor U8294 (N_8294,N_7813,N_7014);
nand U8295 (N_8295,N_6785,N_7358);
and U8296 (N_8296,N_7575,N_7511);
nand U8297 (N_8297,N_7031,N_7305);
or U8298 (N_8298,N_7055,N_6070);
nand U8299 (N_8299,N_6665,N_6242);
and U8300 (N_8300,N_6990,N_6527);
xnor U8301 (N_8301,N_7481,N_7559);
and U8302 (N_8302,N_6337,N_6777);
and U8303 (N_8303,N_7945,N_7081);
or U8304 (N_8304,N_6864,N_6138);
xor U8305 (N_8305,N_6669,N_7765);
nand U8306 (N_8306,N_7522,N_6611);
nand U8307 (N_8307,N_6332,N_6942);
nand U8308 (N_8308,N_6074,N_6345);
and U8309 (N_8309,N_7807,N_7644);
xor U8310 (N_8310,N_6247,N_6226);
or U8311 (N_8311,N_6550,N_6862);
nor U8312 (N_8312,N_6515,N_7062);
nor U8313 (N_8313,N_6601,N_6578);
nor U8314 (N_8314,N_6088,N_6853);
and U8315 (N_8315,N_7885,N_7661);
and U8316 (N_8316,N_7627,N_6218);
nor U8317 (N_8317,N_7190,N_6775);
xor U8318 (N_8318,N_6718,N_6683);
nor U8319 (N_8319,N_7824,N_6582);
or U8320 (N_8320,N_6948,N_7467);
or U8321 (N_8321,N_6407,N_7676);
or U8322 (N_8322,N_7611,N_6091);
or U8323 (N_8323,N_6424,N_6571);
nand U8324 (N_8324,N_7553,N_7176);
xor U8325 (N_8325,N_6922,N_6094);
and U8326 (N_8326,N_7659,N_7317);
nor U8327 (N_8327,N_7744,N_7080);
nand U8328 (N_8328,N_6763,N_7387);
nand U8329 (N_8329,N_7201,N_6427);
or U8330 (N_8330,N_6004,N_7669);
xor U8331 (N_8331,N_6284,N_7424);
nor U8332 (N_8332,N_7195,N_7354);
and U8333 (N_8333,N_6645,N_6908);
xor U8334 (N_8334,N_6583,N_7787);
and U8335 (N_8335,N_6979,N_7999);
xor U8336 (N_8336,N_7606,N_6897);
and U8337 (N_8337,N_7095,N_7400);
nor U8338 (N_8338,N_7756,N_7960);
nor U8339 (N_8339,N_7699,N_6950);
nand U8340 (N_8340,N_7479,N_6917);
nand U8341 (N_8341,N_6566,N_6350);
nor U8342 (N_8342,N_6468,N_7932);
nor U8343 (N_8343,N_7969,N_6573);
nand U8344 (N_8344,N_6012,N_6267);
or U8345 (N_8345,N_7414,N_7437);
or U8346 (N_8346,N_7364,N_6442);
and U8347 (N_8347,N_7351,N_7380);
or U8348 (N_8348,N_7586,N_6119);
or U8349 (N_8349,N_6060,N_7056);
nand U8350 (N_8350,N_6562,N_7991);
and U8351 (N_8351,N_6944,N_6726);
nor U8352 (N_8352,N_7961,N_6535);
and U8353 (N_8353,N_6151,N_6528);
xor U8354 (N_8354,N_6147,N_7114);
nand U8355 (N_8355,N_7264,N_6049);
xor U8356 (N_8356,N_7043,N_7148);
nor U8357 (N_8357,N_6828,N_7812);
and U8358 (N_8358,N_6248,N_6301);
and U8359 (N_8359,N_7911,N_6681);
nand U8360 (N_8360,N_6249,N_7702);
xor U8361 (N_8361,N_6771,N_6791);
or U8362 (N_8362,N_7534,N_7135);
nand U8363 (N_8363,N_7645,N_7563);
nor U8364 (N_8364,N_7432,N_7139);
or U8365 (N_8365,N_6991,N_7548);
nor U8366 (N_8366,N_7235,N_7746);
nor U8367 (N_8367,N_6824,N_7022);
or U8368 (N_8368,N_7884,N_7265);
nand U8369 (N_8369,N_7763,N_7677);
and U8370 (N_8370,N_7173,N_7579);
xnor U8371 (N_8371,N_7033,N_6260);
nand U8372 (N_8372,N_6313,N_6901);
nor U8373 (N_8373,N_7588,N_6420);
xor U8374 (N_8374,N_7442,N_7088);
xnor U8375 (N_8375,N_7116,N_7598);
or U8376 (N_8376,N_6793,N_7782);
nor U8377 (N_8377,N_6025,N_6112);
nor U8378 (N_8378,N_7692,N_6035);
xnor U8379 (N_8379,N_7102,N_6524);
and U8380 (N_8380,N_7743,N_6805);
nor U8381 (N_8381,N_6110,N_6168);
and U8382 (N_8382,N_6397,N_6237);
nor U8383 (N_8383,N_6937,N_6529);
nand U8384 (N_8384,N_7596,N_6634);
xnor U8385 (N_8385,N_6010,N_6872);
nand U8386 (N_8386,N_6947,N_6075);
or U8387 (N_8387,N_6041,N_6596);
nor U8388 (N_8388,N_7121,N_7978);
nand U8389 (N_8389,N_6782,N_6752);
nor U8390 (N_8390,N_6852,N_7892);
nand U8391 (N_8391,N_7208,N_7182);
nor U8392 (N_8392,N_6021,N_7490);
xnor U8393 (N_8393,N_6435,N_6347);
nand U8394 (N_8394,N_6548,N_6945);
nand U8395 (N_8395,N_6741,N_6005);
and U8396 (N_8396,N_6554,N_6409);
nor U8397 (N_8397,N_6998,N_6213);
xnor U8398 (N_8398,N_7907,N_7788);
xnor U8399 (N_8399,N_7906,N_7652);
xor U8400 (N_8400,N_7883,N_6178);
nor U8401 (N_8401,N_7938,N_7816);
nor U8402 (N_8402,N_6357,N_6673);
nand U8403 (N_8403,N_6682,N_6533);
or U8404 (N_8404,N_6545,N_7171);
and U8405 (N_8405,N_7382,N_7904);
nand U8406 (N_8406,N_6235,N_7452);
nor U8407 (N_8407,N_7390,N_7392);
nor U8408 (N_8408,N_6976,N_7026);
nor U8409 (N_8409,N_7740,N_6765);
and U8410 (N_8410,N_6312,N_6390);
and U8411 (N_8411,N_6564,N_6694);
nand U8412 (N_8412,N_7629,N_7708);
nor U8413 (N_8413,N_6865,N_6980);
nand U8414 (N_8414,N_6735,N_7602);
and U8415 (N_8415,N_6125,N_6818);
xor U8416 (N_8416,N_6239,N_7791);
or U8417 (N_8417,N_6289,N_7012);
or U8418 (N_8418,N_6961,N_6102);
nor U8419 (N_8419,N_7290,N_7556);
nor U8420 (N_8420,N_6739,N_6308);
nor U8421 (N_8421,N_7446,N_6932);
and U8422 (N_8422,N_6016,N_6751);
xor U8423 (N_8423,N_6770,N_6473);
and U8424 (N_8424,N_7657,N_6227);
xnor U8425 (N_8425,N_7229,N_6489);
nor U8426 (N_8426,N_6481,N_7106);
nand U8427 (N_8427,N_7255,N_7109);
and U8428 (N_8428,N_6132,N_7272);
or U8429 (N_8429,N_6597,N_7381);
xnor U8430 (N_8430,N_7178,N_7115);
nor U8431 (N_8431,N_7040,N_7851);
or U8432 (N_8432,N_7079,N_6236);
xnor U8433 (N_8433,N_7306,N_7008);
or U8434 (N_8434,N_7720,N_6485);
nor U8435 (N_8435,N_7491,N_7592);
nand U8436 (N_8436,N_6493,N_7860);
nor U8437 (N_8437,N_6909,N_6069);
xnor U8438 (N_8438,N_7407,N_7655);
and U8439 (N_8439,N_6107,N_7408);
nand U8440 (N_8440,N_6685,N_7423);
xnor U8441 (N_8441,N_6062,N_7108);
or U8442 (N_8442,N_7039,N_7175);
nor U8443 (N_8443,N_6336,N_6957);
nor U8444 (N_8444,N_7909,N_6382);
xnor U8445 (N_8445,N_6999,N_7473);
or U8446 (N_8446,N_7530,N_7430);
nor U8447 (N_8447,N_6303,N_6130);
nand U8448 (N_8448,N_7993,N_6612);
and U8449 (N_8449,N_7837,N_7818);
nand U8450 (N_8450,N_6849,N_6517);
or U8451 (N_8451,N_6398,N_7562);
or U8452 (N_8452,N_6880,N_7421);
nor U8453 (N_8453,N_6039,N_7261);
xnor U8454 (N_8454,N_6040,N_7997);
nor U8455 (N_8455,N_7090,N_6194);
or U8456 (N_8456,N_7608,N_7460);
or U8457 (N_8457,N_7735,N_7804);
nand U8458 (N_8458,N_7448,N_6653);
or U8459 (N_8459,N_7754,N_7850);
nor U8460 (N_8460,N_7071,N_6637);
or U8461 (N_8461,N_7326,N_6712);
xor U8462 (N_8462,N_7613,N_6586);
nor U8463 (N_8463,N_6136,N_7594);
nand U8464 (N_8464,N_7480,N_6044);
nor U8465 (N_8465,N_7967,N_7798);
and U8466 (N_8466,N_6329,N_6282);
or U8467 (N_8467,N_7908,N_7474);
and U8468 (N_8468,N_7546,N_6028);
or U8469 (N_8469,N_6396,N_6326);
or U8470 (N_8470,N_6857,N_6799);
xor U8471 (N_8471,N_6821,N_6819);
xnor U8472 (N_8472,N_6212,N_6537);
or U8473 (N_8473,N_6997,N_6170);
or U8474 (N_8474,N_7428,N_6640);
and U8475 (N_8475,N_7844,N_7705);
and U8476 (N_8476,N_7453,N_7641);
or U8477 (N_8477,N_6064,N_7896);
nor U8478 (N_8478,N_7847,N_6068);
nand U8479 (N_8479,N_6808,N_7463);
xor U8480 (N_8480,N_6057,N_6037);
nor U8481 (N_8481,N_7021,N_7046);
xor U8482 (N_8482,N_7193,N_7696);
and U8483 (N_8483,N_7542,N_6043);
or U8484 (N_8484,N_6356,N_7540);
nor U8485 (N_8485,N_7797,N_6140);
xor U8486 (N_8486,N_6474,N_6483);
xor U8487 (N_8487,N_7733,N_6827);
nor U8488 (N_8488,N_7137,N_6277);
xor U8489 (N_8489,N_6459,N_6869);
or U8490 (N_8490,N_7375,N_6900);
or U8491 (N_8491,N_7514,N_6429);
xor U8492 (N_8492,N_7949,N_7516);
and U8493 (N_8493,N_6549,N_7455);
xor U8494 (N_8494,N_6377,N_6806);
xor U8495 (N_8495,N_7568,N_6422);
and U8496 (N_8496,N_6434,N_7915);
nor U8497 (N_8497,N_6885,N_6346);
and U8498 (N_8498,N_6772,N_7526);
nor U8499 (N_8499,N_6141,N_6625);
or U8500 (N_8500,N_6383,N_7674);
or U8501 (N_8501,N_6072,N_7561);
xnor U8502 (N_8502,N_6686,N_6887);
nor U8503 (N_8503,N_6659,N_6167);
or U8504 (N_8504,N_6644,N_7683);
nor U8505 (N_8505,N_6926,N_7795);
or U8506 (N_8506,N_6392,N_7160);
xnor U8507 (N_8507,N_6940,N_6137);
nand U8508 (N_8508,N_6842,N_6142);
or U8509 (N_8509,N_7289,N_7537);
or U8510 (N_8510,N_6538,N_6677);
nor U8511 (N_8511,N_6978,N_6516);
nor U8512 (N_8512,N_6500,N_7939);
and U8513 (N_8513,N_7356,N_7587);
nand U8514 (N_8514,N_7623,N_6834);
nand U8515 (N_8515,N_6411,N_6081);
nor U8516 (N_8516,N_6134,N_7693);
xnor U8517 (N_8517,N_6339,N_6323);
nand U8518 (N_8518,N_7209,N_7215);
nor U8519 (N_8519,N_7378,N_7794);
xor U8520 (N_8520,N_7792,N_6281);
and U8521 (N_8521,N_7482,N_7957);
nor U8522 (N_8522,N_7082,N_6954);
and U8523 (N_8523,N_7237,N_7332);
or U8524 (N_8524,N_7009,N_6103);
nand U8525 (N_8525,N_6708,N_7785);
and U8526 (N_8526,N_7273,N_7987);
nand U8527 (N_8527,N_6353,N_6224);
or U8528 (N_8528,N_6825,N_7420);
or U8529 (N_8529,N_6893,N_6184);
or U8530 (N_8530,N_6231,N_6001);
and U8531 (N_8531,N_6324,N_6873);
or U8532 (N_8532,N_6745,N_6090);
and U8533 (N_8533,N_6257,N_7910);
or U8534 (N_8534,N_7980,N_7017);
nand U8535 (N_8535,N_6767,N_7566);
nand U8536 (N_8536,N_6400,N_7155);
or U8537 (N_8537,N_7903,N_6766);
or U8538 (N_8538,N_7020,N_6984);
and U8539 (N_8539,N_7002,N_6623);
nand U8540 (N_8540,N_6121,N_7888);
nor U8541 (N_8541,N_7532,N_7355);
and U8542 (N_8542,N_6454,N_7512);
nand U8543 (N_8543,N_6096,N_6837);
and U8544 (N_8544,N_7666,N_6609);
nor U8545 (N_8545,N_7941,N_6967);
and U8546 (N_8546,N_6185,N_6344);
nand U8547 (N_8547,N_6325,N_7270);
xnor U8548 (N_8548,N_7284,N_7164);
nand U8549 (N_8549,N_7963,N_7105);
nor U8550 (N_8550,N_6907,N_7443);
or U8551 (N_8551,N_7942,N_7334);
xor U8552 (N_8552,N_6715,N_7493);
and U8553 (N_8553,N_7126,N_7799);
and U8554 (N_8554,N_7762,N_6047);
nand U8555 (N_8555,N_6365,N_6030);
xor U8556 (N_8556,N_7583,N_7552);
xor U8557 (N_8557,N_7232,N_6654);
and U8558 (N_8558,N_6341,N_6668);
nor U8559 (N_8559,N_7662,N_7285);
or U8560 (N_8560,N_6910,N_6316);
nand U8561 (N_8561,N_7653,N_7919);
or U8562 (N_8562,N_7140,N_7525);
and U8563 (N_8563,N_7527,N_7433);
and U8564 (N_8564,N_6935,N_7469);
or U8565 (N_8565,N_6924,N_6919);
or U8566 (N_8566,N_6448,N_7647);
and U8567 (N_8567,N_6443,N_6076);
xnor U8568 (N_8568,N_7034,N_6629);
xnor U8569 (N_8569,N_7394,N_7409);
xor U8570 (N_8570,N_6233,N_7368);
and U8571 (N_8571,N_7411,N_6568);
nor U8572 (N_8572,N_6165,N_6158);
xor U8573 (N_8573,N_7113,N_7187);
xor U8574 (N_8574,N_7047,N_7259);
nand U8575 (N_8575,N_7165,N_7817);
nor U8576 (N_8576,N_7701,N_7495);
xor U8577 (N_8577,N_7709,N_7504);
or U8578 (N_8578,N_7044,N_7554);
xnor U8579 (N_8579,N_6270,N_7228);
or U8580 (N_8580,N_6958,N_7872);
or U8581 (N_8581,N_6736,N_6126);
and U8582 (N_8582,N_6648,N_6208);
or U8583 (N_8583,N_6116,N_6747);
or U8584 (N_8584,N_6338,N_6903);
and U8585 (N_8585,N_7477,N_7691);
and U8586 (N_8586,N_7127,N_6860);
and U8587 (N_8587,N_6855,N_6692);
or U8588 (N_8588,N_7028,N_7350);
nor U8589 (N_8589,N_7279,N_6521);
xor U8590 (N_8590,N_6221,N_7803);
and U8591 (N_8591,N_6711,N_7564);
nor U8592 (N_8592,N_7344,N_6180);
nor U8593 (N_8593,N_6385,N_7248);
xor U8594 (N_8594,N_6902,N_6467);
xnor U8595 (N_8595,N_6187,N_6962);
or U8596 (N_8596,N_7684,N_7268);
nor U8597 (N_8597,N_7107,N_6334);
or U8598 (N_8598,N_7427,N_6077);
nand U8599 (N_8599,N_7831,N_7893);
and U8600 (N_8600,N_6705,N_7931);
nand U8601 (N_8601,N_6746,N_7595);
nor U8602 (N_8602,N_6584,N_6559);
and U8603 (N_8603,N_6495,N_7624);
xor U8604 (N_8604,N_7227,N_6839);
nand U8605 (N_8605,N_7841,N_7886);
nand U8606 (N_8606,N_6020,N_7626);
nor U8607 (N_8607,N_6707,N_6305);
nor U8608 (N_8608,N_7718,N_6163);
xnor U8609 (N_8609,N_6475,N_6690);
and U8610 (N_8610,N_7956,N_6956);
or U8611 (N_8611,N_6446,N_7404);
xnor U8612 (N_8612,N_7091,N_7440);
and U8613 (N_8613,N_6478,N_6080);
xnor U8614 (N_8614,N_7133,N_7536);
nand U8615 (N_8615,N_6152,N_7687);
and U8616 (N_8616,N_7833,N_6449);
xor U8617 (N_8617,N_7499,N_7944);
and U8618 (N_8618,N_7771,N_7019);
nand U8619 (N_8619,N_7042,N_7412);
and U8620 (N_8620,N_7550,N_7675);
nor U8621 (N_8621,N_7294,N_6063);
or U8622 (N_8622,N_6722,N_6223);
and U8623 (N_8623,N_6905,N_6720);
nand U8624 (N_8624,N_6730,N_7258);
nand U8625 (N_8625,N_6960,N_6914);
nand U8626 (N_8626,N_6802,N_6503);
nor U8627 (N_8627,N_7458,N_6689);
nor U8628 (N_8628,N_6114,N_7217);
xnor U8629 (N_8629,N_7954,N_7600);
nor U8630 (N_8630,N_6563,N_6544);
or U8631 (N_8631,N_6079,N_7174);
xor U8632 (N_8632,N_6655,N_6274);
nand U8633 (N_8633,N_6876,N_6992);
and U8634 (N_8634,N_6036,N_6293);
xor U8635 (N_8635,N_7601,N_6265);
nand U8636 (N_8636,N_6450,N_7593);
xnor U8637 (N_8637,N_7747,N_7565);
or U8638 (N_8638,N_6371,N_7663);
xnor U8639 (N_8639,N_7323,N_7322);
nor U8640 (N_8640,N_6488,N_7092);
or U8641 (N_8641,N_7342,N_6027);
xor U8642 (N_8642,N_6097,N_6477);
or U8643 (N_8643,N_7580,N_6895);
nand U8644 (N_8644,N_7330,N_7509);
nor U8645 (N_8645,N_7636,N_6975);
nor U8646 (N_8646,N_6731,N_6155);
and U8647 (N_8647,N_7366,N_7796);
nand U8648 (N_8648,N_6291,N_7617);
and U8649 (N_8649,N_7650,N_6567);
or U8650 (N_8650,N_7599,N_7895);
nand U8651 (N_8651,N_7431,N_7604);
nor U8652 (N_8652,N_7465,N_7487);
nand U8653 (N_8653,N_7531,N_7779);
and U8654 (N_8654,N_7327,N_7093);
and U8655 (N_8655,N_7111,N_6758);
or U8656 (N_8656,N_6331,N_7880);
and U8657 (N_8657,N_7395,N_6129);
nor U8658 (N_8658,N_7545,N_7158);
and U8659 (N_8659,N_7809,N_7736);
and U8660 (N_8660,N_7025,N_6879);
xnor U8661 (N_8661,N_6757,N_6438);
xor U8662 (N_8662,N_6061,N_7891);
nor U8663 (N_8663,N_7973,N_6649);
nand U8664 (N_8664,N_7439,N_6413);
xnor U8665 (N_8665,N_6217,N_7492);
or U8666 (N_8666,N_7786,N_7325);
or U8667 (N_8667,N_6762,N_6798);
and U8668 (N_8668,N_7901,N_6575);
xnor U8669 (N_8669,N_7419,N_7569);
xnor U8670 (N_8670,N_7345,N_7037);
xor U8671 (N_8671,N_7524,N_7059);
nand U8672 (N_8672,N_7827,N_7898);
nand U8673 (N_8673,N_6570,N_6558);
nand U8674 (N_8674,N_7391,N_7147);
nand U8675 (N_8675,N_6881,N_7066);
nand U8676 (N_8676,N_7853,N_6139);
xor U8677 (N_8677,N_6379,N_7700);
nand U8678 (N_8678,N_6008,N_7800);
or U8679 (N_8679,N_6679,N_6166);
xnor U8680 (N_8680,N_7067,N_7153);
nand U8681 (N_8681,N_7098,N_6092);
and U8682 (N_8682,N_7766,N_7985);
or U8683 (N_8683,N_7373,N_7282);
and U8684 (N_8684,N_6457,N_6886);
and U8685 (N_8685,N_6228,N_6408);
xnor U8686 (N_8686,N_6122,N_6451);
nand U8687 (N_8687,N_7497,N_6920);
nor U8688 (N_8688,N_6513,N_6572);
nor U8689 (N_8689,N_7275,N_7741);
and U8690 (N_8690,N_6014,N_6871);
nand U8691 (N_8691,N_7144,N_7713);
and U8692 (N_8692,N_7202,N_6744);
xnor U8693 (N_8693,N_7870,N_6870);
or U8694 (N_8694,N_7630,N_7303);
or U8695 (N_8695,N_6836,N_7719);
or U8696 (N_8696,N_6594,N_6496);
or U8697 (N_8697,N_6190,N_6042);
nor U8698 (N_8698,N_6743,N_7622);
and U8699 (N_8699,N_6256,N_7664);
or U8700 (N_8700,N_7513,N_6512);
xor U8701 (N_8701,N_7397,N_7607);
and U8702 (N_8702,N_6807,N_7413);
or U8703 (N_8703,N_7489,N_7256);
xnor U8704 (N_8704,N_6675,N_6988);
xnor U8705 (N_8705,N_7959,N_6482);
xnor U8706 (N_8706,N_6487,N_6780);
and U8707 (N_8707,N_7866,N_7247);
and U8708 (N_8708,N_7488,N_7278);
nand U8709 (N_8709,N_7815,N_7726);
nand U8710 (N_8710,N_6388,N_6619);
nand U8711 (N_8711,N_6153,N_6804);
nand U8712 (N_8712,N_7464,N_7947);
or U8713 (N_8713,N_6764,N_6965);
and U8714 (N_8714,N_6453,N_6684);
nand U8715 (N_8715,N_7679,N_7362);
xor U8716 (N_8716,N_6581,N_6891);
nor U8717 (N_8717,N_7341,N_7732);
and U8718 (N_8718,N_6330,N_7966);
xnor U8719 (N_8719,N_7363,N_6246);
or U8720 (N_8720,N_6539,N_7169);
xor U8721 (N_8721,N_7377,N_7149);
nand U8722 (N_8722,N_6333,N_6437);
nor U8723 (N_8723,N_6788,N_6355);
nor U8724 (N_8724,N_6856,N_7730);
nand U8725 (N_8725,N_7288,N_6105);
or U8726 (N_8726,N_7496,N_6320);
or U8727 (N_8727,N_6275,N_7162);
and U8728 (N_8728,N_7112,N_6971);
xor U8729 (N_8729,N_6373,N_7221);
xor U8730 (N_8730,N_6627,N_7867);
xnor U8731 (N_8731,N_6177,N_6552);
nor U8732 (N_8732,N_6278,N_6610);
xnor U8733 (N_8733,N_7711,N_6048);
or U8734 (N_8734,N_7934,N_6941);
or U8735 (N_8735,N_7103,N_6826);
xnor U8736 (N_8736,N_6358,N_7097);
nor U8737 (N_8737,N_6406,N_6461);
nor U8738 (N_8738,N_7254,N_7928);
nor U8739 (N_8739,N_6725,N_6925);
nand U8740 (N_8740,N_6884,N_6127);
nor U8741 (N_8741,N_6738,N_7628);
nor U8742 (N_8742,N_7946,N_6363);
nor U8743 (N_8743,N_6996,N_7197);
nor U8744 (N_8744,N_7541,N_6748);
nor U8745 (N_8745,N_7249,N_7618);
nor U8746 (N_8746,N_6877,N_7614);
nor U8747 (N_8747,N_7054,N_6959);
nor U8748 (N_8748,N_6056,N_7219);
or U8749 (N_8749,N_6890,N_6801);
and U8750 (N_8750,N_7124,N_6436);
xor U8751 (N_8751,N_6013,N_6173);
nor U8752 (N_8752,N_7656,N_6024);
xnor U8753 (N_8753,N_6587,N_7984);
nor U8754 (N_8754,N_6643,N_6702);
nor U8755 (N_8755,N_7456,N_6018);
xnor U8756 (N_8756,N_7951,N_7406);
nor U8757 (N_8757,N_6784,N_7475);
nand U8758 (N_8758,N_7131,N_6642);
and U8759 (N_8759,N_7292,N_6174);
and U8760 (N_8760,N_7637,N_6509);
or U8761 (N_8761,N_7917,N_6607);
xnor U8762 (N_8762,N_6372,N_6638);
nor U8763 (N_8763,N_6009,N_6651);
or U8764 (N_8764,N_7854,N_6335);
nor U8765 (N_8765,N_6983,N_7584);
nor U8766 (N_8766,N_6085,N_6565);
or U8767 (N_8767,N_6831,N_7445);
and U8768 (N_8768,N_7328,N_7061);
xnor U8769 (N_8769,N_6419,N_6982);
or U8770 (N_8770,N_6362,N_6868);
xnor U8771 (N_8771,N_6480,N_7723);
or U8772 (N_8772,N_7935,N_7051);
xor U8773 (N_8773,N_6410,N_7544);
and U8774 (N_8774,N_7520,N_7212);
nor U8775 (N_8775,N_6906,N_7864);
nor U8776 (N_8776,N_7013,N_6740);
xnor U8777 (N_8777,N_7277,N_6230);
and U8778 (N_8778,N_7302,N_6833);
and U8779 (N_8779,N_7557,N_7857);
nor U8780 (N_8780,N_7745,N_6073);
nand U8781 (N_8781,N_7878,N_6863);
nor U8782 (N_8782,N_6628,N_7077);
xor U8783 (N_8783,N_6343,N_7402);
nand U8784 (N_8784,N_6543,N_7189);
xnor U8785 (N_8785,N_7977,N_6052);
xor U8786 (N_8786,N_6404,N_6713);
and U8787 (N_8787,N_7181,N_6253);
and U8788 (N_8788,N_6829,N_6579);
xnor U8789 (N_8789,N_7589,N_6084);
nor U8790 (N_8790,N_7914,N_6845);
or U8791 (N_8791,N_6633,N_6776);
and U8792 (N_8792,N_7990,N_7101);
or U8793 (N_8793,N_7104,N_6441);
and U8794 (N_8794,N_7760,N_7924);
nand U8795 (N_8795,N_7717,N_6384);
xnor U8796 (N_8796,N_6214,N_6734);
or U8797 (N_8797,N_7856,N_6321);
xnor U8798 (N_8798,N_6830,N_7138);
nand U8799 (N_8799,N_7297,N_6841);
nand U8800 (N_8800,N_6672,N_6370);
or U8801 (N_8801,N_6972,N_6172);
and U8802 (N_8802,N_6670,N_7929);
and U8803 (N_8803,N_6452,N_6145);
nand U8804 (N_8804,N_7770,N_7922);
xnor U8805 (N_8805,N_7742,N_6502);
nor U8806 (N_8806,N_7873,N_6007);
nand U8807 (N_8807,N_6781,N_7136);
xor U8808 (N_8808,N_6479,N_7283);
and U8809 (N_8809,N_7441,N_7658);
or U8810 (N_8810,N_6508,N_7502);
and U8811 (N_8811,N_6066,N_7454);
and U8812 (N_8812,N_6930,N_6171);
nand U8813 (N_8813,N_7777,N_7120);
nor U8814 (N_8814,N_7697,N_7680);
nand U8815 (N_8815,N_6703,N_7125);
nand U8816 (N_8816,N_7078,N_7157);
and U8817 (N_8817,N_7146,N_7122);
nand U8818 (N_8818,N_6518,N_6789);
nor U8819 (N_8819,N_7937,N_7172);
nor U8820 (N_8820,N_7925,N_6252);
nor U8821 (N_8821,N_7063,N_6421);
nor U8822 (N_8822,N_6994,N_7434);
nor U8823 (N_8823,N_7263,N_7343);
xor U8824 (N_8824,N_7099,N_6067);
nor U8825 (N_8825,N_7476,N_7468);
nand U8826 (N_8826,N_6117,N_7802);
nand U8827 (N_8827,N_6083,N_6389);
or U8828 (N_8828,N_6019,N_7374);
nand U8829 (N_8829,N_6211,N_6878);
nor U8830 (N_8830,N_7451,N_7789);
nor U8831 (N_8831,N_6974,N_7086);
nor U8832 (N_8832,N_6050,N_6953);
and U8833 (N_8833,N_6133,N_6639);
and U8834 (N_8834,N_7185,N_6113);
and U8835 (N_8835,N_6952,N_6099);
nor U8836 (N_8836,N_7236,N_6534);
or U8837 (N_8837,N_6882,N_6658);
and U8838 (N_8838,N_7399,N_6318);
nor U8839 (N_8839,N_6973,N_7686);
nand U8840 (N_8840,N_6273,N_7752);
and U8841 (N_8841,N_6364,N_6205);
xor U8842 (N_8842,N_7117,N_6131);
nand U8843 (N_8843,N_6519,N_7855);
nand U8844 (N_8844,N_7577,N_7143);
nand U8845 (N_8845,N_7576,N_6580);
or U8846 (N_8846,N_7045,N_7843);
nand U8847 (N_8847,N_6374,N_6319);
and U8848 (N_8848,N_6732,N_7050);
xor U8849 (N_8849,N_6755,N_7757);
nand U8850 (N_8850,N_7578,N_7868);
xor U8851 (N_8851,N_6051,N_7877);
nand U8852 (N_8852,N_6790,N_7772);
nand U8853 (N_8853,N_6939,N_6031);
and U8854 (N_8854,N_7438,N_6916);
nor U8855 (N_8855,N_6896,N_6631);
nand U8856 (N_8856,N_7572,N_7267);
xnor U8857 (N_8857,N_6288,N_7950);
nand U8858 (N_8858,N_7035,N_7461);
xor U8859 (N_8859,N_7293,N_7690);
nand U8860 (N_8860,N_6378,N_7179);
xnor U8861 (N_8861,N_7110,N_7671);
or U8862 (N_8862,N_7739,N_7603);
nand U8863 (N_8863,N_7761,N_7863);
and U8864 (N_8864,N_6188,N_6444);
and U8865 (N_8865,N_6470,N_7769);
nor U8866 (N_8866,N_7738,N_7689);
nor U8867 (N_8867,N_7667,N_7084);
nand U8868 (N_8868,N_6599,N_7129);
and U8869 (N_8869,N_6456,N_7257);
and U8870 (N_8870,N_6053,N_7986);
nor U8871 (N_8871,N_6678,N_7571);
xor U8872 (N_8872,N_7075,N_6874);
nor U8873 (N_8873,N_7953,N_6360);
nand U8874 (N_8874,N_7501,N_6569);
xor U8875 (N_8875,N_7070,N_7698);
or U8876 (N_8876,N_7970,N_7975);
nand U8877 (N_8877,N_7239,N_6297);
and U8878 (N_8878,N_6135,N_6847);
nand U8879 (N_8879,N_6412,N_6846);
nand U8880 (N_8880,N_6809,N_7861);
nor U8881 (N_8881,N_6904,N_6375);
xor U8882 (N_8882,N_6553,N_7194);
xnor U8883 (N_8883,N_6189,N_7712);
nor U8884 (N_8884,N_6915,N_6395);
xor U8885 (N_8885,N_6981,N_7981);
nand U8886 (N_8886,N_7820,N_7704);
xnor U8887 (N_8887,N_7849,N_6595);
nor U8888 (N_8888,N_6927,N_7340);
nand U8889 (N_8889,N_7183,N_7648);
nand U8890 (N_8890,N_6514,N_6369);
nor U8891 (N_8891,N_7253,N_6875);
or U8892 (N_8892,N_7484,N_6403);
or U8893 (N_8893,N_6261,N_7470);
nand U8894 (N_8894,N_6259,N_7361);
or U8895 (N_8895,N_7839,N_7936);
nor U8896 (N_8896,N_6843,N_7405);
nand U8897 (N_8897,N_7295,N_7252);
and U8898 (N_8898,N_7186,N_7912);
nor U8899 (N_8899,N_7393,N_7640);
or U8900 (N_8900,N_7415,N_6087);
and U8901 (N_8901,N_7485,N_7505);
and U8902 (N_8902,N_7654,N_6086);
xor U8903 (N_8903,N_7234,N_7836);
nand U8904 (N_8904,N_7154,N_7992);
and U8905 (N_8905,N_7274,N_6462);
nand U8906 (N_8906,N_7089,N_7943);
nand U8907 (N_8907,N_6526,N_7728);
nor U8908 (N_8908,N_6349,N_6033);
or U8909 (N_8909,N_7271,N_6912);
xnor U8910 (N_8910,N_6207,N_6197);
xnor U8911 (N_8911,N_7682,N_6200);
xnor U8912 (N_8912,N_6769,N_7876);
or U8913 (N_8913,N_7307,N_6026);
and U8914 (N_8914,N_6773,N_6191);
or U8915 (N_8915,N_7245,N_7150);
xor U8916 (N_8916,N_7521,N_6250);
or U8917 (N_8917,N_6432,N_7032);
or U8918 (N_8918,N_6100,N_7848);
and U8919 (N_8919,N_7784,N_6460);
or U8920 (N_8920,N_7210,N_6590);
xor U8921 (N_8921,N_7503,N_7570);
or U8922 (N_8922,N_6499,N_6283);
or U8923 (N_8923,N_7459,N_7023);
nand U8924 (N_8924,N_6943,N_7773);
and U8925 (N_8925,N_7064,N_6494);
nor U8926 (N_8926,N_6721,N_6555);
xnor U8927 (N_8927,N_6181,N_7376);
or U8928 (N_8928,N_6038,N_6687);
or U8929 (N_8929,N_7574,N_7216);
or U8930 (N_8930,N_7649,N_7793);
nor U8931 (N_8931,N_7958,N_7060);
nand U8932 (N_8932,N_7706,N_7094);
nor U8933 (N_8933,N_6466,N_7776);
xor U8934 (N_8934,N_7859,N_7703);
xor U8935 (N_8935,N_7639,N_7403);
nor U8936 (N_8936,N_7296,N_7515);
or U8937 (N_8937,N_7858,N_7457);
nand U8938 (N_8938,N_7365,N_7755);
nand U8939 (N_8939,N_6985,N_6206);
xor U8940 (N_8940,N_7498,N_7852);
nand U8941 (N_8941,N_7298,N_6464);
nor U8942 (N_8942,N_6794,N_6540);
or U8943 (N_8943,N_7921,N_7145);
nand U8944 (N_8944,N_7011,N_7805);
nor U8945 (N_8945,N_7313,N_7213);
and U8946 (N_8946,N_7995,N_6351);
xnor U8947 (N_8947,N_7024,N_7783);
nand U8948 (N_8948,N_6202,N_7688);
nand U8949 (N_8949,N_7918,N_6602);
and U8950 (N_8950,N_7507,N_6034);
nand U8951 (N_8951,N_6209,N_6124);
nor U8952 (N_8952,N_6585,N_6613);
nand U8953 (N_8953,N_7695,N_7842);
nor U8954 (N_8954,N_6472,N_6381);
xnor U8955 (N_8955,N_7177,N_6652);
nand U8956 (N_8956,N_7722,N_7004);
xnor U8957 (N_8957,N_6761,N_7778);
nand U8958 (N_8958,N_6892,N_6486);
xor U8959 (N_8959,N_7260,N_7560);
nand U8960 (N_8960,N_6510,N_6359);
nor U8961 (N_8961,N_7538,N_6219);
or U8962 (N_8962,N_6614,N_6888);
nand U8963 (N_8963,N_6118,N_7620);
nor U8964 (N_8964,N_7681,N_6426);
or U8965 (N_8965,N_7196,N_7132);
and U8966 (N_8966,N_7774,N_6778);
or U8967 (N_8967,N_6531,N_6970);
xor U8968 (N_8968,N_6327,N_6251);
or U8969 (N_8969,N_6792,N_7670);
nor U8970 (N_8970,N_7887,N_6417);
and U8971 (N_8971,N_6123,N_7251);
xnor U8972 (N_8972,N_7821,N_7519);
xnor U8973 (N_8973,N_7401,N_6476);
and U8974 (N_8974,N_6949,N_7418);
nand U8975 (N_8975,N_7166,N_6115);
nor U8976 (N_8976,N_7167,N_7882);
nand U8977 (N_8977,N_6626,N_6717);
and U8978 (N_8978,N_6899,N_6120);
nor U8979 (N_8979,N_7266,N_6198);
or U8980 (N_8980,N_7036,N_6986);
or U8981 (N_8981,N_7331,N_6428);
nor U8982 (N_8982,N_6506,N_7038);
xor U8983 (N_8983,N_7349,N_7191);
xnor U8984 (N_8984,N_6418,N_7646);
xnor U8985 (N_8985,N_7983,N_7069);
nand U8986 (N_8986,N_6546,N_6391);
or U8987 (N_8987,N_6314,N_6603);
nor U8988 (N_8988,N_6258,N_7551);
or U8989 (N_8989,N_7168,N_7673);
or U8990 (N_8990,N_7759,N_7333);
and U8991 (N_8991,N_6309,N_6302);
nor U8992 (N_8992,N_7318,N_7619);
nand U8993 (N_8993,N_7633,N_7128);
nor U8994 (N_8994,N_7422,N_7948);
and U8995 (N_8995,N_6032,N_7379);
nand U8996 (N_8996,N_7840,N_7119);
or U8997 (N_8997,N_6415,N_7320);
and U8998 (N_8998,N_6737,N_6650);
nor U8999 (N_8999,N_6307,N_6244);
nor U9000 (N_9000,N_7848,N_6021);
and U9001 (N_9001,N_7028,N_7747);
xnor U9002 (N_9002,N_7038,N_6346);
nor U9003 (N_9003,N_7941,N_7349);
xor U9004 (N_9004,N_6982,N_6407);
or U9005 (N_9005,N_7082,N_6267);
xnor U9006 (N_9006,N_7510,N_6852);
nand U9007 (N_9007,N_7642,N_6525);
xor U9008 (N_9008,N_6312,N_7357);
nor U9009 (N_9009,N_7211,N_7846);
nor U9010 (N_9010,N_7864,N_6577);
or U9011 (N_9011,N_6083,N_6383);
xnor U9012 (N_9012,N_6928,N_7391);
and U9013 (N_9013,N_7197,N_6296);
or U9014 (N_9014,N_6743,N_6123);
nand U9015 (N_9015,N_6434,N_7700);
or U9016 (N_9016,N_6037,N_7191);
xnor U9017 (N_9017,N_7238,N_7972);
nand U9018 (N_9018,N_7065,N_6927);
xor U9019 (N_9019,N_7205,N_6113);
and U9020 (N_9020,N_7752,N_6859);
xor U9021 (N_9021,N_6615,N_7567);
or U9022 (N_9022,N_6305,N_7989);
nor U9023 (N_9023,N_6385,N_7857);
or U9024 (N_9024,N_6675,N_6503);
and U9025 (N_9025,N_7476,N_7206);
and U9026 (N_9026,N_7350,N_7463);
and U9027 (N_9027,N_6450,N_6371);
nand U9028 (N_9028,N_6515,N_6818);
and U9029 (N_9029,N_6083,N_7967);
nand U9030 (N_9030,N_7178,N_6643);
and U9031 (N_9031,N_7381,N_7348);
nor U9032 (N_9032,N_6839,N_7352);
and U9033 (N_9033,N_6163,N_7933);
nor U9034 (N_9034,N_7240,N_6165);
xor U9035 (N_9035,N_7628,N_7470);
or U9036 (N_9036,N_7884,N_7429);
xnor U9037 (N_9037,N_6266,N_7593);
nand U9038 (N_9038,N_7690,N_7541);
xor U9039 (N_9039,N_7404,N_6173);
nand U9040 (N_9040,N_7588,N_7873);
or U9041 (N_9041,N_6039,N_6077);
nor U9042 (N_9042,N_6426,N_7801);
xor U9043 (N_9043,N_6893,N_6174);
or U9044 (N_9044,N_7391,N_6334);
and U9045 (N_9045,N_6416,N_6289);
xnor U9046 (N_9046,N_7104,N_7941);
nor U9047 (N_9047,N_7914,N_6239);
nor U9048 (N_9048,N_7670,N_6420);
and U9049 (N_9049,N_6812,N_7540);
nand U9050 (N_9050,N_7295,N_6775);
nand U9051 (N_9051,N_7669,N_7211);
or U9052 (N_9052,N_6138,N_6884);
and U9053 (N_9053,N_6813,N_6744);
and U9054 (N_9054,N_6298,N_6594);
nor U9055 (N_9055,N_7902,N_6694);
xor U9056 (N_9056,N_6511,N_7607);
nor U9057 (N_9057,N_7475,N_7419);
xnor U9058 (N_9058,N_7376,N_7354);
nor U9059 (N_9059,N_7263,N_7758);
nand U9060 (N_9060,N_7271,N_6997);
xor U9061 (N_9061,N_6307,N_7600);
nor U9062 (N_9062,N_7051,N_7082);
nand U9063 (N_9063,N_7793,N_6582);
and U9064 (N_9064,N_6643,N_6737);
xnor U9065 (N_9065,N_7143,N_7738);
nand U9066 (N_9066,N_7251,N_7526);
nand U9067 (N_9067,N_7999,N_7386);
or U9068 (N_9068,N_6877,N_7039);
or U9069 (N_9069,N_6147,N_7551);
or U9070 (N_9070,N_6317,N_6816);
and U9071 (N_9071,N_7119,N_6115);
and U9072 (N_9072,N_6915,N_7028);
xor U9073 (N_9073,N_7366,N_6689);
xor U9074 (N_9074,N_6330,N_6298);
or U9075 (N_9075,N_7966,N_7880);
nor U9076 (N_9076,N_6088,N_6810);
nand U9077 (N_9077,N_7591,N_6374);
and U9078 (N_9078,N_7190,N_7266);
or U9079 (N_9079,N_6366,N_6587);
xnor U9080 (N_9080,N_6469,N_7165);
or U9081 (N_9081,N_6958,N_6252);
nor U9082 (N_9082,N_6673,N_6100);
nand U9083 (N_9083,N_7601,N_6123);
nor U9084 (N_9084,N_7770,N_7777);
nand U9085 (N_9085,N_6430,N_6989);
and U9086 (N_9086,N_7172,N_6417);
xnor U9087 (N_9087,N_6735,N_7764);
nand U9088 (N_9088,N_7128,N_6851);
nand U9089 (N_9089,N_6644,N_6546);
xor U9090 (N_9090,N_7351,N_7814);
xnor U9091 (N_9091,N_6188,N_6977);
nand U9092 (N_9092,N_6092,N_7937);
or U9093 (N_9093,N_6109,N_6302);
nor U9094 (N_9094,N_6337,N_6050);
and U9095 (N_9095,N_7001,N_6028);
or U9096 (N_9096,N_6996,N_7070);
and U9097 (N_9097,N_7655,N_6562);
or U9098 (N_9098,N_7338,N_6618);
nand U9099 (N_9099,N_7588,N_7178);
and U9100 (N_9100,N_6512,N_6517);
nor U9101 (N_9101,N_7354,N_6808);
nand U9102 (N_9102,N_7851,N_7714);
xnor U9103 (N_9103,N_7978,N_7557);
nor U9104 (N_9104,N_6409,N_7870);
nand U9105 (N_9105,N_7041,N_6257);
nor U9106 (N_9106,N_6719,N_7769);
xor U9107 (N_9107,N_6863,N_6693);
xnor U9108 (N_9108,N_7190,N_7340);
nor U9109 (N_9109,N_7493,N_7941);
and U9110 (N_9110,N_7678,N_6314);
or U9111 (N_9111,N_7085,N_6503);
and U9112 (N_9112,N_6060,N_6003);
or U9113 (N_9113,N_7355,N_6320);
nor U9114 (N_9114,N_6966,N_7758);
and U9115 (N_9115,N_6572,N_6315);
or U9116 (N_9116,N_7197,N_6006);
nor U9117 (N_9117,N_7128,N_7046);
and U9118 (N_9118,N_7272,N_6190);
xor U9119 (N_9119,N_7153,N_6789);
xor U9120 (N_9120,N_6558,N_6702);
nand U9121 (N_9121,N_6633,N_6658);
xor U9122 (N_9122,N_7649,N_7023);
and U9123 (N_9123,N_7273,N_6011);
nand U9124 (N_9124,N_6891,N_6148);
nor U9125 (N_9125,N_6618,N_6827);
or U9126 (N_9126,N_7114,N_7499);
xnor U9127 (N_9127,N_6087,N_6763);
nand U9128 (N_9128,N_7315,N_6062);
nor U9129 (N_9129,N_6306,N_7772);
xor U9130 (N_9130,N_6050,N_6493);
and U9131 (N_9131,N_7141,N_6700);
nor U9132 (N_9132,N_7155,N_6713);
or U9133 (N_9133,N_7514,N_6570);
xor U9134 (N_9134,N_7784,N_6578);
nand U9135 (N_9135,N_6073,N_6674);
or U9136 (N_9136,N_6905,N_7762);
nand U9137 (N_9137,N_6743,N_6018);
nor U9138 (N_9138,N_6875,N_6498);
and U9139 (N_9139,N_6097,N_6653);
xor U9140 (N_9140,N_7004,N_6534);
or U9141 (N_9141,N_6946,N_6408);
or U9142 (N_9142,N_7358,N_7279);
nor U9143 (N_9143,N_7711,N_6278);
nand U9144 (N_9144,N_6728,N_7062);
and U9145 (N_9145,N_7407,N_6136);
and U9146 (N_9146,N_6468,N_6226);
nand U9147 (N_9147,N_7999,N_7677);
nor U9148 (N_9148,N_6791,N_7310);
xor U9149 (N_9149,N_6291,N_7037);
nand U9150 (N_9150,N_7348,N_7200);
or U9151 (N_9151,N_6074,N_7471);
nor U9152 (N_9152,N_6389,N_7991);
or U9153 (N_9153,N_7639,N_7415);
xnor U9154 (N_9154,N_6574,N_6896);
xor U9155 (N_9155,N_7826,N_6729);
nand U9156 (N_9156,N_7978,N_6437);
nor U9157 (N_9157,N_6559,N_6090);
nand U9158 (N_9158,N_7770,N_7821);
xnor U9159 (N_9159,N_6414,N_6690);
nand U9160 (N_9160,N_6724,N_6379);
nor U9161 (N_9161,N_7618,N_6702);
nand U9162 (N_9162,N_7745,N_6201);
nand U9163 (N_9163,N_6967,N_7059);
and U9164 (N_9164,N_6513,N_6746);
nand U9165 (N_9165,N_6871,N_6547);
or U9166 (N_9166,N_7811,N_6832);
nor U9167 (N_9167,N_6532,N_7132);
and U9168 (N_9168,N_7818,N_7852);
xnor U9169 (N_9169,N_7105,N_7967);
nand U9170 (N_9170,N_6044,N_7083);
nand U9171 (N_9171,N_6410,N_6883);
xor U9172 (N_9172,N_6148,N_7449);
or U9173 (N_9173,N_7156,N_7498);
nand U9174 (N_9174,N_7506,N_6265);
nor U9175 (N_9175,N_6598,N_6450);
nor U9176 (N_9176,N_7444,N_7092);
nand U9177 (N_9177,N_7366,N_7092);
or U9178 (N_9178,N_7870,N_6620);
and U9179 (N_9179,N_6942,N_6617);
and U9180 (N_9180,N_7849,N_6899);
nand U9181 (N_9181,N_6412,N_7484);
and U9182 (N_9182,N_6580,N_6172);
nor U9183 (N_9183,N_6876,N_7583);
nand U9184 (N_9184,N_6002,N_6957);
nand U9185 (N_9185,N_7805,N_7866);
nand U9186 (N_9186,N_7389,N_7457);
xnor U9187 (N_9187,N_7095,N_6035);
xnor U9188 (N_9188,N_6341,N_6412);
or U9189 (N_9189,N_7426,N_6967);
or U9190 (N_9190,N_7550,N_6916);
xor U9191 (N_9191,N_7564,N_6174);
nor U9192 (N_9192,N_7405,N_6835);
and U9193 (N_9193,N_6323,N_7102);
or U9194 (N_9194,N_7401,N_7205);
nand U9195 (N_9195,N_6034,N_7048);
or U9196 (N_9196,N_7390,N_6883);
nor U9197 (N_9197,N_7786,N_6624);
nor U9198 (N_9198,N_6391,N_6632);
nor U9199 (N_9199,N_7919,N_6840);
nand U9200 (N_9200,N_7351,N_7261);
or U9201 (N_9201,N_7094,N_7765);
nor U9202 (N_9202,N_7894,N_6929);
xnor U9203 (N_9203,N_7691,N_6591);
nor U9204 (N_9204,N_6908,N_7117);
xnor U9205 (N_9205,N_6658,N_6506);
nand U9206 (N_9206,N_7535,N_6599);
nand U9207 (N_9207,N_6622,N_6750);
nand U9208 (N_9208,N_6573,N_7545);
and U9209 (N_9209,N_7600,N_7702);
xor U9210 (N_9210,N_7813,N_6475);
nor U9211 (N_9211,N_6340,N_6317);
and U9212 (N_9212,N_7221,N_7402);
or U9213 (N_9213,N_6269,N_6102);
and U9214 (N_9214,N_7720,N_6331);
or U9215 (N_9215,N_6256,N_7522);
and U9216 (N_9216,N_7964,N_7155);
or U9217 (N_9217,N_7913,N_7463);
nand U9218 (N_9218,N_7338,N_6509);
nor U9219 (N_9219,N_6078,N_7175);
nor U9220 (N_9220,N_7753,N_6721);
or U9221 (N_9221,N_6166,N_6646);
or U9222 (N_9222,N_7374,N_6508);
xnor U9223 (N_9223,N_7691,N_6057);
or U9224 (N_9224,N_7381,N_6259);
nor U9225 (N_9225,N_6765,N_6949);
or U9226 (N_9226,N_6990,N_7421);
xnor U9227 (N_9227,N_6884,N_6663);
xnor U9228 (N_9228,N_7471,N_7605);
nand U9229 (N_9229,N_7497,N_6121);
nor U9230 (N_9230,N_7698,N_6523);
xor U9231 (N_9231,N_6125,N_6351);
nor U9232 (N_9232,N_7205,N_6293);
nand U9233 (N_9233,N_7651,N_6629);
nor U9234 (N_9234,N_7958,N_7109);
nor U9235 (N_9235,N_7016,N_7250);
or U9236 (N_9236,N_7845,N_7905);
nand U9237 (N_9237,N_7067,N_6603);
nand U9238 (N_9238,N_7957,N_7549);
nor U9239 (N_9239,N_6070,N_7201);
xnor U9240 (N_9240,N_7548,N_6046);
nor U9241 (N_9241,N_6208,N_7888);
nand U9242 (N_9242,N_6597,N_7267);
xor U9243 (N_9243,N_7991,N_7941);
nand U9244 (N_9244,N_6275,N_7745);
and U9245 (N_9245,N_6241,N_7474);
and U9246 (N_9246,N_6012,N_6128);
nand U9247 (N_9247,N_7090,N_6095);
and U9248 (N_9248,N_6983,N_7723);
and U9249 (N_9249,N_6800,N_7607);
nor U9250 (N_9250,N_6824,N_6153);
xnor U9251 (N_9251,N_6979,N_7437);
xnor U9252 (N_9252,N_6708,N_6131);
xnor U9253 (N_9253,N_7921,N_7331);
nand U9254 (N_9254,N_7428,N_7461);
and U9255 (N_9255,N_7154,N_7231);
xor U9256 (N_9256,N_7724,N_7738);
nand U9257 (N_9257,N_6450,N_6955);
nand U9258 (N_9258,N_7546,N_6290);
xnor U9259 (N_9259,N_7332,N_6878);
and U9260 (N_9260,N_7309,N_6127);
or U9261 (N_9261,N_6293,N_7246);
nand U9262 (N_9262,N_6751,N_7140);
xor U9263 (N_9263,N_7976,N_7320);
nor U9264 (N_9264,N_6812,N_6507);
xor U9265 (N_9265,N_7831,N_7626);
or U9266 (N_9266,N_6488,N_6119);
nand U9267 (N_9267,N_6173,N_6352);
and U9268 (N_9268,N_7334,N_7660);
nand U9269 (N_9269,N_6598,N_6734);
nor U9270 (N_9270,N_7683,N_7709);
nor U9271 (N_9271,N_6229,N_7414);
or U9272 (N_9272,N_6800,N_6706);
or U9273 (N_9273,N_6981,N_7217);
or U9274 (N_9274,N_6076,N_6444);
and U9275 (N_9275,N_6069,N_7293);
or U9276 (N_9276,N_7058,N_6287);
or U9277 (N_9277,N_6388,N_7112);
or U9278 (N_9278,N_6820,N_7475);
or U9279 (N_9279,N_6131,N_7416);
nand U9280 (N_9280,N_7695,N_6352);
nand U9281 (N_9281,N_6686,N_7154);
and U9282 (N_9282,N_6903,N_6459);
nor U9283 (N_9283,N_7735,N_7465);
nand U9284 (N_9284,N_7978,N_6313);
nor U9285 (N_9285,N_6411,N_7910);
xnor U9286 (N_9286,N_7596,N_6357);
xnor U9287 (N_9287,N_7625,N_7724);
or U9288 (N_9288,N_7836,N_7891);
xnor U9289 (N_9289,N_7101,N_6749);
nor U9290 (N_9290,N_6434,N_6064);
nor U9291 (N_9291,N_6868,N_7079);
nand U9292 (N_9292,N_6028,N_6479);
nand U9293 (N_9293,N_7196,N_6912);
or U9294 (N_9294,N_7751,N_7081);
and U9295 (N_9295,N_6767,N_6656);
nand U9296 (N_9296,N_6218,N_6546);
xor U9297 (N_9297,N_7885,N_7665);
or U9298 (N_9298,N_7791,N_7260);
nor U9299 (N_9299,N_6348,N_7461);
xor U9300 (N_9300,N_7238,N_6496);
xor U9301 (N_9301,N_7629,N_6318);
or U9302 (N_9302,N_6028,N_7218);
nor U9303 (N_9303,N_7374,N_7175);
xor U9304 (N_9304,N_6702,N_6790);
nand U9305 (N_9305,N_7230,N_6013);
and U9306 (N_9306,N_6660,N_7699);
and U9307 (N_9307,N_6537,N_6766);
xnor U9308 (N_9308,N_7424,N_7461);
nand U9309 (N_9309,N_7481,N_6347);
and U9310 (N_9310,N_7617,N_7411);
or U9311 (N_9311,N_6200,N_7951);
nand U9312 (N_9312,N_6351,N_6539);
and U9313 (N_9313,N_7711,N_6649);
nor U9314 (N_9314,N_7273,N_7017);
nand U9315 (N_9315,N_7982,N_6895);
xor U9316 (N_9316,N_6074,N_6039);
nor U9317 (N_9317,N_6295,N_7602);
and U9318 (N_9318,N_6913,N_7055);
xor U9319 (N_9319,N_6909,N_7708);
nand U9320 (N_9320,N_6242,N_7215);
nor U9321 (N_9321,N_6660,N_7608);
nor U9322 (N_9322,N_7193,N_6758);
nand U9323 (N_9323,N_6501,N_7268);
and U9324 (N_9324,N_6891,N_6253);
nor U9325 (N_9325,N_6607,N_6639);
or U9326 (N_9326,N_7100,N_6825);
nor U9327 (N_9327,N_7969,N_6866);
xnor U9328 (N_9328,N_6719,N_6648);
and U9329 (N_9329,N_7533,N_7516);
or U9330 (N_9330,N_7287,N_7468);
nand U9331 (N_9331,N_6767,N_6117);
nor U9332 (N_9332,N_7722,N_6179);
nor U9333 (N_9333,N_7741,N_7022);
and U9334 (N_9334,N_6936,N_7432);
nor U9335 (N_9335,N_6284,N_7612);
nor U9336 (N_9336,N_7635,N_6737);
and U9337 (N_9337,N_6224,N_6027);
or U9338 (N_9338,N_6186,N_7474);
or U9339 (N_9339,N_7252,N_6861);
or U9340 (N_9340,N_7800,N_7147);
or U9341 (N_9341,N_7845,N_6681);
or U9342 (N_9342,N_7230,N_6954);
nor U9343 (N_9343,N_7776,N_7609);
or U9344 (N_9344,N_6040,N_6813);
and U9345 (N_9345,N_6756,N_7194);
xor U9346 (N_9346,N_6876,N_7637);
nor U9347 (N_9347,N_7659,N_6482);
nor U9348 (N_9348,N_7490,N_6313);
or U9349 (N_9349,N_7073,N_7220);
and U9350 (N_9350,N_6556,N_7282);
nor U9351 (N_9351,N_7891,N_7054);
nand U9352 (N_9352,N_7303,N_7878);
or U9353 (N_9353,N_6608,N_6639);
and U9354 (N_9354,N_6986,N_7394);
nand U9355 (N_9355,N_6512,N_7763);
or U9356 (N_9356,N_6859,N_6868);
or U9357 (N_9357,N_7769,N_7692);
xor U9358 (N_9358,N_6318,N_7298);
nor U9359 (N_9359,N_6566,N_7043);
nor U9360 (N_9360,N_6946,N_7291);
nor U9361 (N_9361,N_7232,N_6642);
nor U9362 (N_9362,N_7963,N_6759);
or U9363 (N_9363,N_6102,N_6576);
nor U9364 (N_9364,N_6961,N_7278);
nand U9365 (N_9365,N_6796,N_6104);
or U9366 (N_9366,N_7974,N_7300);
and U9367 (N_9367,N_7382,N_7755);
nand U9368 (N_9368,N_6589,N_7817);
nor U9369 (N_9369,N_6750,N_6496);
xor U9370 (N_9370,N_7358,N_7355);
or U9371 (N_9371,N_7020,N_6334);
or U9372 (N_9372,N_7462,N_7708);
nor U9373 (N_9373,N_7248,N_6595);
nor U9374 (N_9374,N_7231,N_6937);
or U9375 (N_9375,N_6321,N_6119);
nand U9376 (N_9376,N_7586,N_6268);
and U9377 (N_9377,N_6913,N_6575);
nand U9378 (N_9378,N_6053,N_6181);
or U9379 (N_9379,N_7899,N_7310);
nor U9380 (N_9380,N_7578,N_6331);
or U9381 (N_9381,N_7869,N_7688);
nor U9382 (N_9382,N_6464,N_7562);
nand U9383 (N_9383,N_7804,N_6529);
xnor U9384 (N_9384,N_7569,N_6306);
and U9385 (N_9385,N_6602,N_7645);
or U9386 (N_9386,N_6488,N_7145);
nor U9387 (N_9387,N_6499,N_6007);
xor U9388 (N_9388,N_6935,N_6739);
nand U9389 (N_9389,N_6206,N_6931);
nand U9390 (N_9390,N_7603,N_6895);
nor U9391 (N_9391,N_6872,N_6852);
nand U9392 (N_9392,N_7508,N_7614);
nor U9393 (N_9393,N_6060,N_6477);
and U9394 (N_9394,N_6929,N_6390);
and U9395 (N_9395,N_6346,N_6090);
nand U9396 (N_9396,N_7420,N_6360);
nor U9397 (N_9397,N_6653,N_6453);
nand U9398 (N_9398,N_7786,N_6256);
nor U9399 (N_9399,N_7726,N_6959);
xor U9400 (N_9400,N_6210,N_6075);
or U9401 (N_9401,N_6234,N_7230);
and U9402 (N_9402,N_7811,N_7464);
or U9403 (N_9403,N_7724,N_7735);
nor U9404 (N_9404,N_7731,N_7347);
xnor U9405 (N_9405,N_7158,N_6797);
nand U9406 (N_9406,N_6906,N_6368);
nand U9407 (N_9407,N_7512,N_6324);
or U9408 (N_9408,N_6698,N_6516);
and U9409 (N_9409,N_7383,N_6362);
or U9410 (N_9410,N_6735,N_6121);
nor U9411 (N_9411,N_7866,N_7385);
nor U9412 (N_9412,N_7854,N_6571);
nand U9413 (N_9413,N_7673,N_7861);
nor U9414 (N_9414,N_6509,N_6564);
nand U9415 (N_9415,N_7295,N_6725);
xnor U9416 (N_9416,N_6679,N_7231);
nor U9417 (N_9417,N_6893,N_7916);
and U9418 (N_9418,N_6727,N_7271);
and U9419 (N_9419,N_7582,N_7340);
xor U9420 (N_9420,N_7363,N_7400);
and U9421 (N_9421,N_7669,N_7467);
nand U9422 (N_9422,N_6430,N_6581);
or U9423 (N_9423,N_6204,N_7716);
and U9424 (N_9424,N_7168,N_6200);
or U9425 (N_9425,N_6113,N_6097);
xor U9426 (N_9426,N_6266,N_6965);
and U9427 (N_9427,N_7545,N_7212);
nor U9428 (N_9428,N_7477,N_6707);
nor U9429 (N_9429,N_6849,N_7445);
and U9430 (N_9430,N_6259,N_7279);
xnor U9431 (N_9431,N_7076,N_6894);
xnor U9432 (N_9432,N_6490,N_7892);
xor U9433 (N_9433,N_6102,N_7246);
or U9434 (N_9434,N_6173,N_6917);
or U9435 (N_9435,N_7738,N_7500);
nor U9436 (N_9436,N_7585,N_7344);
or U9437 (N_9437,N_6692,N_7921);
nand U9438 (N_9438,N_7709,N_6953);
xnor U9439 (N_9439,N_7160,N_6860);
nand U9440 (N_9440,N_6026,N_7026);
or U9441 (N_9441,N_7021,N_6670);
xor U9442 (N_9442,N_7218,N_6549);
and U9443 (N_9443,N_7184,N_7403);
nor U9444 (N_9444,N_6905,N_6088);
xnor U9445 (N_9445,N_7785,N_7871);
or U9446 (N_9446,N_6121,N_7646);
nand U9447 (N_9447,N_7788,N_6237);
or U9448 (N_9448,N_7530,N_6340);
and U9449 (N_9449,N_6083,N_6598);
or U9450 (N_9450,N_7934,N_7086);
and U9451 (N_9451,N_6315,N_7515);
xnor U9452 (N_9452,N_6715,N_7437);
nand U9453 (N_9453,N_6777,N_7999);
xnor U9454 (N_9454,N_7785,N_7907);
or U9455 (N_9455,N_6618,N_6684);
nand U9456 (N_9456,N_7797,N_7850);
nor U9457 (N_9457,N_6064,N_6310);
or U9458 (N_9458,N_6111,N_7475);
or U9459 (N_9459,N_6993,N_6726);
or U9460 (N_9460,N_6121,N_6663);
nor U9461 (N_9461,N_7967,N_7175);
and U9462 (N_9462,N_7874,N_6739);
nor U9463 (N_9463,N_7777,N_7727);
nor U9464 (N_9464,N_7344,N_6870);
nor U9465 (N_9465,N_6673,N_7054);
or U9466 (N_9466,N_7414,N_7792);
nand U9467 (N_9467,N_7260,N_6393);
and U9468 (N_9468,N_6086,N_7894);
nand U9469 (N_9469,N_6181,N_6692);
and U9470 (N_9470,N_6689,N_6723);
or U9471 (N_9471,N_6740,N_6630);
or U9472 (N_9472,N_6621,N_6560);
nand U9473 (N_9473,N_6268,N_6573);
and U9474 (N_9474,N_7593,N_6417);
nand U9475 (N_9475,N_7901,N_6312);
or U9476 (N_9476,N_7114,N_7027);
or U9477 (N_9477,N_7426,N_6422);
or U9478 (N_9478,N_7164,N_7142);
and U9479 (N_9479,N_6597,N_7213);
nor U9480 (N_9480,N_7148,N_7628);
or U9481 (N_9481,N_7240,N_7742);
or U9482 (N_9482,N_7053,N_6741);
or U9483 (N_9483,N_6538,N_6748);
xnor U9484 (N_9484,N_7078,N_6250);
xor U9485 (N_9485,N_6631,N_6985);
and U9486 (N_9486,N_7085,N_7121);
nor U9487 (N_9487,N_6288,N_7069);
xor U9488 (N_9488,N_6212,N_6187);
nand U9489 (N_9489,N_7042,N_7850);
nand U9490 (N_9490,N_6749,N_6937);
and U9491 (N_9491,N_6325,N_7956);
and U9492 (N_9492,N_6777,N_7360);
nor U9493 (N_9493,N_6566,N_7847);
and U9494 (N_9494,N_7186,N_6213);
and U9495 (N_9495,N_7159,N_6473);
nor U9496 (N_9496,N_6683,N_7929);
xor U9497 (N_9497,N_6054,N_7938);
and U9498 (N_9498,N_7783,N_7720);
xnor U9499 (N_9499,N_7124,N_6389);
xnor U9500 (N_9500,N_7650,N_6782);
and U9501 (N_9501,N_6939,N_7053);
or U9502 (N_9502,N_6471,N_7679);
or U9503 (N_9503,N_7022,N_7509);
xnor U9504 (N_9504,N_7517,N_7771);
nor U9505 (N_9505,N_6371,N_6719);
nor U9506 (N_9506,N_7365,N_7413);
xor U9507 (N_9507,N_7550,N_6934);
xnor U9508 (N_9508,N_7698,N_6107);
nor U9509 (N_9509,N_6170,N_7074);
or U9510 (N_9510,N_7071,N_7503);
or U9511 (N_9511,N_7901,N_7450);
or U9512 (N_9512,N_6263,N_7889);
and U9513 (N_9513,N_7088,N_6341);
or U9514 (N_9514,N_6065,N_6402);
or U9515 (N_9515,N_7257,N_7528);
nor U9516 (N_9516,N_7671,N_6692);
and U9517 (N_9517,N_6386,N_6739);
nor U9518 (N_9518,N_7006,N_7115);
or U9519 (N_9519,N_6175,N_6828);
nor U9520 (N_9520,N_6081,N_7913);
xnor U9521 (N_9521,N_7242,N_7745);
xnor U9522 (N_9522,N_7327,N_7056);
nor U9523 (N_9523,N_7766,N_6181);
or U9524 (N_9524,N_6595,N_7146);
and U9525 (N_9525,N_6184,N_7976);
xnor U9526 (N_9526,N_7834,N_6719);
and U9527 (N_9527,N_7804,N_6588);
or U9528 (N_9528,N_7850,N_7544);
or U9529 (N_9529,N_7730,N_7702);
nor U9530 (N_9530,N_7716,N_7267);
nand U9531 (N_9531,N_6698,N_7646);
and U9532 (N_9532,N_6937,N_6327);
and U9533 (N_9533,N_7162,N_7610);
or U9534 (N_9534,N_7795,N_6263);
nand U9535 (N_9535,N_6984,N_7777);
xnor U9536 (N_9536,N_7865,N_7517);
and U9537 (N_9537,N_6724,N_6188);
or U9538 (N_9538,N_7448,N_6291);
and U9539 (N_9539,N_7641,N_7081);
xor U9540 (N_9540,N_6779,N_6103);
nor U9541 (N_9541,N_6849,N_7171);
nor U9542 (N_9542,N_7784,N_6872);
nor U9543 (N_9543,N_7097,N_6733);
nor U9544 (N_9544,N_7293,N_7510);
nand U9545 (N_9545,N_6725,N_7080);
nor U9546 (N_9546,N_6887,N_7576);
and U9547 (N_9547,N_7830,N_7693);
nand U9548 (N_9548,N_7727,N_6502);
xor U9549 (N_9549,N_6780,N_6875);
or U9550 (N_9550,N_7074,N_7482);
or U9551 (N_9551,N_7936,N_7660);
nor U9552 (N_9552,N_6056,N_7968);
xor U9553 (N_9553,N_6338,N_6601);
and U9554 (N_9554,N_7160,N_6044);
nand U9555 (N_9555,N_6713,N_7611);
and U9556 (N_9556,N_7233,N_7839);
or U9557 (N_9557,N_7001,N_7827);
xnor U9558 (N_9558,N_7548,N_6303);
nand U9559 (N_9559,N_6508,N_6906);
or U9560 (N_9560,N_7460,N_6898);
nand U9561 (N_9561,N_7151,N_7100);
nand U9562 (N_9562,N_7400,N_7973);
nand U9563 (N_9563,N_6030,N_7202);
nand U9564 (N_9564,N_7971,N_6929);
or U9565 (N_9565,N_6145,N_7541);
or U9566 (N_9566,N_7699,N_6603);
and U9567 (N_9567,N_6477,N_7748);
or U9568 (N_9568,N_6456,N_6461);
or U9569 (N_9569,N_6757,N_7556);
nor U9570 (N_9570,N_6034,N_7006);
or U9571 (N_9571,N_7877,N_6492);
nand U9572 (N_9572,N_7684,N_7720);
or U9573 (N_9573,N_6518,N_7668);
nor U9574 (N_9574,N_6853,N_7470);
and U9575 (N_9575,N_6715,N_7188);
nand U9576 (N_9576,N_7553,N_7555);
nand U9577 (N_9577,N_7458,N_7947);
nand U9578 (N_9578,N_6661,N_6353);
xor U9579 (N_9579,N_7064,N_6549);
or U9580 (N_9580,N_6153,N_7771);
and U9581 (N_9581,N_7309,N_6149);
nor U9582 (N_9582,N_7379,N_6781);
nand U9583 (N_9583,N_7743,N_7801);
nor U9584 (N_9584,N_6713,N_6750);
or U9585 (N_9585,N_7519,N_7990);
and U9586 (N_9586,N_6033,N_6166);
and U9587 (N_9587,N_6395,N_7805);
and U9588 (N_9588,N_7014,N_6995);
nor U9589 (N_9589,N_6854,N_7296);
nor U9590 (N_9590,N_7657,N_6545);
nand U9591 (N_9591,N_6539,N_7376);
and U9592 (N_9592,N_6589,N_6795);
nor U9593 (N_9593,N_6188,N_7664);
nand U9594 (N_9594,N_6433,N_7199);
and U9595 (N_9595,N_7119,N_6684);
nand U9596 (N_9596,N_6059,N_6065);
and U9597 (N_9597,N_7089,N_7677);
xnor U9598 (N_9598,N_7911,N_6110);
and U9599 (N_9599,N_7437,N_6997);
xnor U9600 (N_9600,N_7875,N_7756);
nor U9601 (N_9601,N_7302,N_7350);
or U9602 (N_9602,N_6283,N_6877);
nand U9603 (N_9603,N_6117,N_7658);
nor U9604 (N_9604,N_7083,N_7851);
nand U9605 (N_9605,N_6931,N_7058);
nor U9606 (N_9606,N_7799,N_7018);
xor U9607 (N_9607,N_7505,N_7384);
and U9608 (N_9608,N_6568,N_7126);
or U9609 (N_9609,N_6955,N_6178);
nand U9610 (N_9610,N_6633,N_7431);
nand U9611 (N_9611,N_7203,N_7156);
nor U9612 (N_9612,N_6027,N_6052);
and U9613 (N_9613,N_6125,N_6155);
nor U9614 (N_9614,N_6311,N_7861);
xnor U9615 (N_9615,N_6009,N_7630);
xor U9616 (N_9616,N_7782,N_7567);
xor U9617 (N_9617,N_6904,N_7897);
or U9618 (N_9618,N_7804,N_7516);
nand U9619 (N_9619,N_6742,N_7305);
xor U9620 (N_9620,N_6998,N_7509);
or U9621 (N_9621,N_7978,N_7822);
and U9622 (N_9622,N_7868,N_6963);
or U9623 (N_9623,N_7334,N_7994);
nand U9624 (N_9624,N_7249,N_7712);
nor U9625 (N_9625,N_6755,N_7307);
nor U9626 (N_9626,N_6672,N_7688);
xnor U9627 (N_9627,N_7195,N_6755);
or U9628 (N_9628,N_6555,N_7329);
nor U9629 (N_9629,N_6306,N_7502);
xnor U9630 (N_9630,N_7291,N_6318);
nand U9631 (N_9631,N_7411,N_7979);
nor U9632 (N_9632,N_6860,N_7613);
and U9633 (N_9633,N_7382,N_7076);
xnor U9634 (N_9634,N_7743,N_6037);
nand U9635 (N_9635,N_6426,N_6941);
nor U9636 (N_9636,N_7297,N_6119);
or U9637 (N_9637,N_7907,N_6404);
nand U9638 (N_9638,N_7128,N_6524);
and U9639 (N_9639,N_6675,N_6365);
and U9640 (N_9640,N_7949,N_7523);
nor U9641 (N_9641,N_7943,N_6514);
nand U9642 (N_9642,N_7831,N_7442);
nor U9643 (N_9643,N_6225,N_6666);
xnor U9644 (N_9644,N_7016,N_7165);
nand U9645 (N_9645,N_7746,N_6530);
and U9646 (N_9646,N_7044,N_7954);
nor U9647 (N_9647,N_6462,N_7648);
nand U9648 (N_9648,N_7072,N_7219);
nand U9649 (N_9649,N_7344,N_6642);
or U9650 (N_9650,N_7406,N_6509);
xor U9651 (N_9651,N_7639,N_7628);
or U9652 (N_9652,N_6735,N_6378);
nor U9653 (N_9653,N_6398,N_7252);
xnor U9654 (N_9654,N_6812,N_7139);
and U9655 (N_9655,N_7964,N_7685);
or U9656 (N_9656,N_7787,N_6561);
xor U9657 (N_9657,N_6439,N_6070);
nand U9658 (N_9658,N_7444,N_7562);
nor U9659 (N_9659,N_7966,N_7406);
xnor U9660 (N_9660,N_6910,N_6265);
xnor U9661 (N_9661,N_6029,N_6085);
nor U9662 (N_9662,N_6743,N_6733);
nor U9663 (N_9663,N_7023,N_7673);
xor U9664 (N_9664,N_7215,N_7274);
nor U9665 (N_9665,N_6521,N_6464);
nor U9666 (N_9666,N_6010,N_6296);
nand U9667 (N_9667,N_6684,N_7354);
nand U9668 (N_9668,N_7808,N_6689);
nor U9669 (N_9669,N_6476,N_6979);
nor U9670 (N_9670,N_6303,N_7778);
xor U9671 (N_9671,N_7711,N_6002);
or U9672 (N_9672,N_6249,N_6270);
xor U9673 (N_9673,N_7409,N_7357);
xnor U9674 (N_9674,N_7865,N_6561);
or U9675 (N_9675,N_7952,N_6579);
nor U9676 (N_9676,N_7720,N_6403);
or U9677 (N_9677,N_6429,N_6160);
xor U9678 (N_9678,N_7301,N_7855);
xor U9679 (N_9679,N_6454,N_6719);
xnor U9680 (N_9680,N_7226,N_7628);
or U9681 (N_9681,N_6095,N_7332);
nor U9682 (N_9682,N_6789,N_6470);
or U9683 (N_9683,N_6777,N_6560);
xor U9684 (N_9684,N_6773,N_6709);
nand U9685 (N_9685,N_6158,N_6308);
or U9686 (N_9686,N_7761,N_6862);
and U9687 (N_9687,N_6053,N_7644);
or U9688 (N_9688,N_6945,N_6070);
or U9689 (N_9689,N_7780,N_7925);
nand U9690 (N_9690,N_6884,N_7704);
or U9691 (N_9691,N_7433,N_7996);
and U9692 (N_9692,N_7321,N_7644);
nand U9693 (N_9693,N_6228,N_6420);
or U9694 (N_9694,N_6617,N_7276);
nor U9695 (N_9695,N_7852,N_6818);
nand U9696 (N_9696,N_7572,N_7731);
and U9697 (N_9697,N_6958,N_6401);
and U9698 (N_9698,N_6472,N_6253);
or U9699 (N_9699,N_7474,N_7694);
or U9700 (N_9700,N_7074,N_6847);
xnor U9701 (N_9701,N_7491,N_7070);
nand U9702 (N_9702,N_7997,N_7832);
and U9703 (N_9703,N_7705,N_7714);
nor U9704 (N_9704,N_6220,N_7993);
nor U9705 (N_9705,N_6949,N_7226);
xor U9706 (N_9706,N_6560,N_7023);
and U9707 (N_9707,N_6625,N_7925);
or U9708 (N_9708,N_6542,N_7655);
nand U9709 (N_9709,N_6109,N_6116);
or U9710 (N_9710,N_7565,N_6269);
or U9711 (N_9711,N_7927,N_6536);
nor U9712 (N_9712,N_6071,N_6070);
nand U9713 (N_9713,N_7624,N_6254);
xnor U9714 (N_9714,N_7010,N_7119);
and U9715 (N_9715,N_7904,N_6608);
nand U9716 (N_9716,N_7652,N_6054);
and U9717 (N_9717,N_6007,N_7207);
and U9718 (N_9718,N_7912,N_6833);
nand U9719 (N_9719,N_7598,N_7183);
nor U9720 (N_9720,N_7602,N_7724);
nand U9721 (N_9721,N_7327,N_7571);
and U9722 (N_9722,N_6758,N_6550);
or U9723 (N_9723,N_6190,N_7864);
nor U9724 (N_9724,N_6444,N_7571);
and U9725 (N_9725,N_6314,N_7453);
and U9726 (N_9726,N_6383,N_7598);
and U9727 (N_9727,N_6016,N_7711);
xor U9728 (N_9728,N_7759,N_7426);
nand U9729 (N_9729,N_6793,N_6756);
nor U9730 (N_9730,N_7227,N_7427);
or U9731 (N_9731,N_6831,N_6200);
xor U9732 (N_9732,N_7663,N_7014);
xor U9733 (N_9733,N_6969,N_6543);
nor U9734 (N_9734,N_6421,N_6101);
nand U9735 (N_9735,N_6028,N_7307);
nor U9736 (N_9736,N_7194,N_6823);
xnor U9737 (N_9737,N_6969,N_7434);
and U9738 (N_9738,N_7719,N_7606);
nand U9739 (N_9739,N_6712,N_6390);
nand U9740 (N_9740,N_6713,N_7904);
xor U9741 (N_9741,N_6548,N_7988);
xnor U9742 (N_9742,N_7361,N_6292);
and U9743 (N_9743,N_6505,N_6727);
xor U9744 (N_9744,N_7771,N_6566);
and U9745 (N_9745,N_7949,N_6213);
nor U9746 (N_9746,N_7482,N_7587);
nand U9747 (N_9747,N_6182,N_7921);
and U9748 (N_9748,N_7089,N_6256);
xnor U9749 (N_9749,N_6756,N_7964);
xnor U9750 (N_9750,N_7571,N_6874);
nor U9751 (N_9751,N_6154,N_7703);
nand U9752 (N_9752,N_6249,N_7749);
nor U9753 (N_9753,N_6976,N_6865);
nand U9754 (N_9754,N_7979,N_6978);
nand U9755 (N_9755,N_6442,N_6380);
or U9756 (N_9756,N_7830,N_7236);
and U9757 (N_9757,N_6098,N_7757);
nor U9758 (N_9758,N_7483,N_6605);
or U9759 (N_9759,N_6455,N_7674);
nand U9760 (N_9760,N_6859,N_7620);
and U9761 (N_9761,N_6080,N_6040);
nand U9762 (N_9762,N_6639,N_7571);
nand U9763 (N_9763,N_7454,N_6241);
nand U9764 (N_9764,N_6323,N_7636);
or U9765 (N_9765,N_6867,N_6498);
or U9766 (N_9766,N_7662,N_7134);
xnor U9767 (N_9767,N_6573,N_7474);
and U9768 (N_9768,N_7545,N_6771);
nor U9769 (N_9769,N_7375,N_6572);
or U9770 (N_9770,N_7824,N_7984);
nor U9771 (N_9771,N_7118,N_7260);
xnor U9772 (N_9772,N_6629,N_7195);
xnor U9773 (N_9773,N_7782,N_7082);
xor U9774 (N_9774,N_7001,N_6408);
nor U9775 (N_9775,N_6021,N_6152);
nand U9776 (N_9776,N_7334,N_7474);
nor U9777 (N_9777,N_6479,N_6976);
or U9778 (N_9778,N_6425,N_6713);
and U9779 (N_9779,N_6355,N_6562);
nand U9780 (N_9780,N_7470,N_6274);
and U9781 (N_9781,N_7705,N_6311);
nor U9782 (N_9782,N_6357,N_7384);
nor U9783 (N_9783,N_6388,N_7674);
nor U9784 (N_9784,N_7327,N_7483);
or U9785 (N_9785,N_6587,N_6306);
nand U9786 (N_9786,N_6360,N_7130);
nor U9787 (N_9787,N_6436,N_6422);
and U9788 (N_9788,N_7318,N_6656);
or U9789 (N_9789,N_6028,N_6669);
xnor U9790 (N_9790,N_6612,N_6471);
xnor U9791 (N_9791,N_7253,N_6326);
nand U9792 (N_9792,N_7337,N_7784);
nor U9793 (N_9793,N_6574,N_6374);
nor U9794 (N_9794,N_6928,N_6361);
and U9795 (N_9795,N_6653,N_6445);
xor U9796 (N_9796,N_6145,N_6015);
and U9797 (N_9797,N_6247,N_7060);
or U9798 (N_9798,N_7271,N_7670);
nand U9799 (N_9799,N_7367,N_6875);
xor U9800 (N_9800,N_6131,N_7248);
nand U9801 (N_9801,N_6052,N_6945);
xnor U9802 (N_9802,N_7183,N_6915);
xnor U9803 (N_9803,N_7832,N_6745);
nor U9804 (N_9804,N_6249,N_7898);
nand U9805 (N_9805,N_7713,N_6488);
and U9806 (N_9806,N_7339,N_7522);
xor U9807 (N_9807,N_6999,N_7178);
xnor U9808 (N_9808,N_6211,N_7312);
xor U9809 (N_9809,N_7391,N_6344);
nand U9810 (N_9810,N_6777,N_7561);
xor U9811 (N_9811,N_6252,N_6669);
and U9812 (N_9812,N_7641,N_6449);
xor U9813 (N_9813,N_6125,N_6148);
and U9814 (N_9814,N_7939,N_7561);
and U9815 (N_9815,N_7361,N_7295);
or U9816 (N_9816,N_6706,N_6501);
and U9817 (N_9817,N_7530,N_6375);
nor U9818 (N_9818,N_6455,N_7596);
nand U9819 (N_9819,N_6076,N_7199);
xnor U9820 (N_9820,N_7328,N_7166);
xnor U9821 (N_9821,N_6431,N_6936);
or U9822 (N_9822,N_6989,N_6075);
nand U9823 (N_9823,N_6103,N_6338);
nor U9824 (N_9824,N_6295,N_7366);
nor U9825 (N_9825,N_7801,N_6121);
or U9826 (N_9826,N_7382,N_6081);
and U9827 (N_9827,N_6243,N_6727);
nor U9828 (N_9828,N_7915,N_6980);
nand U9829 (N_9829,N_7244,N_6135);
xnor U9830 (N_9830,N_6579,N_6595);
and U9831 (N_9831,N_7613,N_7970);
and U9832 (N_9832,N_6979,N_6609);
xor U9833 (N_9833,N_7545,N_7325);
or U9834 (N_9834,N_7351,N_6687);
or U9835 (N_9835,N_7528,N_6401);
nor U9836 (N_9836,N_6034,N_6799);
or U9837 (N_9837,N_6461,N_7831);
or U9838 (N_9838,N_6849,N_6017);
and U9839 (N_9839,N_6884,N_6673);
and U9840 (N_9840,N_7240,N_7613);
xnor U9841 (N_9841,N_7091,N_7975);
nor U9842 (N_9842,N_7217,N_7777);
or U9843 (N_9843,N_6822,N_6692);
or U9844 (N_9844,N_6353,N_6762);
nor U9845 (N_9845,N_6213,N_7375);
or U9846 (N_9846,N_7780,N_6743);
nand U9847 (N_9847,N_6452,N_6098);
nand U9848 (N_9848,N_7472,N_6245);
or U9849 (N_9849,N_6225,N_7543);
nand U9850 (N_9850,N_7419,N_7117);
and U9851 (N_9851,N_7821,N_6386);
xor U9852 (N_9852,N_6596,N_7408);
and U9853 (N_9853,N_6082,N_6007);
nor U9854 (N_9854,N_6962,N_6708);
xor U9855 (N_9855,N_6164,N_6555);
nor U9856 (N_9856,N_7367,N_7017);
xor U9857 (N_9857,N_7748,N_7830);
xnor U9858 (N_9858,N_7206,N_6517);
or U9859 (N_9859,N_6728,N_6748);
and U9860 (N_9860,N_6778,N_7478);
and U9861 (N_9861,N_7961,N_7099);
nor U9862 (N_9862,N_7004,N_6122);
nand U9863 (N_9863,N_7714,N_7465);
nor U9864 (N_9864,N_7616,N_7656);
or U9865 (N_9865,N_7051,N_7494);
xor U9866 (N_9866,N_7290,N_6653);
or U9867 (N_9867,N_7639,N_7660);
and U9868 (N_9868,N_7513,N_7127);
nand U9869 (N_9869,N_7286,N_7270);
nor U9870 (N_9870,N_7247,N_7293);
nor U9871 (N_9871,N_6591,N_6316);
or U9872 (N_9872,N_6164,N_6927);
and U9873 (N_9873,N_6260,N_6195);
xor U9874 (N_9874,N_6534,N_7260);
xnor U9875 (N_9875,N_7413,N_6430);
or U9876 (N_9876,N_7470,N_7008);
and U9877 (N_9877,N_7373,N_6253);
nand U9878 (N_9878,N_7257,N_6166);
nor U9879 (N_9879,N_6447,N_6142);
and U9880 (N_9880,N_7152,N_6638);
nand U9881 (N_9881,N_6786,N_7272);
or U9882 (N_9882,N_7051,N_7453);
nor U9883 (N_9883,N_7542,N_7726);
nand U9884 (N_9884,N_6932,N_7532);
xor U9885 (N_9885,N_7529,N_6379);
nand U9886 (N_9886,N_7564,N_7642);
nand U9887 (N_9887,N_7355,N_6107);
and U9888 (N_9888,N_7995,N_7578);
or U9889 (N_9889,N_7652,N_6226);
or U9890 (N_9890,N_7607,N_6340);
or U9891 (N_9891,N_7567,N_6564);
nand U9892 (N_9892,N_6025,N_7243);
xnor U9893 (N_9893,N_6625,N_6939);
nand U9894 (N_9894,N_7372,N_7359);
xnor U9895 (N_9895,N_6590,N_6351);
nor U9896 (N_9896,N_6245,N_6660);
xnor U9897 (N_9897,N_7277,N_7385);
or U9898 (N_9898,N_6946,N_7990);
or U9899 (N_9899,N_7170,N_7430);
or U9900 (N_9900,N_6128,N_7905);
or U9901 (N_9901,N_7678,N_6545);
and U9902 (N_9902,N_7092,N_7003);
xor U9903 (N_9903,N_7560,N_7451);
or U9904 (N_9904,N_6943,N_6435);
and U9905 (N_9905,N_6070,N_6155);
xnor U9906 (N_9906,N_7069,N_7353);
nor U9907 (N_9907,N_6891,N_7286);
xnor U9908 (N_9908,N_6558,N_7083);
nand U9909 (N_9909,N_7251,N_7792);
or U9910 (N_9910,N_7005,N_7923);
and U9911 (N_9911,N_6258,N_6743);
nor U9912 (N_9912,N_7377,N_6104);
nand U9913 (N_9913,N_6737,N_7286);
nand U9914 (N_9914,N_7848,N_6102);
nor U9915 (N_9915,N_6930,N_6505);
nor U9916 (N_9916,N_7401,N_6716);
nand U9917 (N_9917,N_6621,N_7375);
nand U9918 (N_9918,N_6168,N_7556);
nor U9919 (N_9919,N_6081,N_6338);
nand U9920 (N_9920,N_7342,N_7610);
and U9921 (N_9921,N_7414,N_7353);
nor U9922 (N_9922,N_7658,N_6254);
nor U9923 (N_9923,N_6639,N_6761);
or U9924 (N_9924,N_6996,N_6106);
nand U9925 (N_9925,N_7661,N_7130);
xor U9926 (N_9926,N_7994,N_6033);
or U9927 (N_9927,N_6640,N_6392);
xnor U9928 (N_9928,N_6855,N_7047);
nand U9929 (N_9929,N_6957,N_7274);
and U9930 (N_9930,N_6341,N_7643);
nor U9931 (N_9931,N_7012,N_7686);
xnor U9932 (N_9932,N_7103,N_7998);
nand U9933 (N_9933,N_6797,N_6344);
nand U9934 (N_9934,N_6384,N_6377);
xor U9935 (N_9935,N_7758,N_6263);
nand U9936 (N_9936,N_6828,N_6244);
and U9937 (N_9937,N_6009,N_7261);
and U9938 (N_9938,N_6705,N_6793);
and U9939 (N_9939,N_7432,N_7656);
nand U9940 (N_9940,N_6429,N_7897);
or U9941 (N_9941,N_7415,N_6991);
or U9942 (N_9942,N_7750,N_7771);
xor U9943 (N_9943,N_6549,N_6451);
xnor U9944 (N_9944,N_7020,N_7098);
xor U9945 (N_9945,N_6362,N_7270);
nand U9946 (N_9946,N_6191,N_7503);
or U9947 (N_9947,N_6342,N_7939);
or U9948 (N_9948,N_7652,N_6325);
and U9949 (N_9949,N_7118,N_7247);
xor U9950 (N_9950,N_7637,N_7541);
nand U9951 (N_9951,N_7914,N_6904);
nor U9952 (N_9952,N_6360,N_6262);
xnor U9953 (N_9953,N_7825,N_6104);
and U9954 (N_9954,N_7939,N_6490);
xor U9955 (N_9955,N_6826,N_7312);
xor U9956 (N_9956,N_6733,N_7303);
and U9957 (N_9957,N_7104,N_6746);
or U9958 (N_9958,N_6464,N_7406);
nor U9959 (N_9959,N_6029,N_7876);
nor U9960 (N_9960,N_7570,N_6090);
nand U9961 (N_9961,N_6860,N_7010);
nand U9962 (N_9962,N_6714,N_6369);
xor U9963 (N_9963,N_6512,N_6001);
and U9964 (N_9964,N_6741,N_7290);
nor U9965 (N_9965,N_7604,N_6841);
nor U9966 (N_9966,N_6056,N_6332);
nor U9967 (N_9967,N_7193,N_6613);
or U9968 (N_9968,N_6739,N_7637);
xor U9969 (N_9969,N_7224,N_6756);
or U9970 (N_9970,N_6698,N_6444);
and U9971 (N_9971,N_6392,N_6505);
xnor U9972 (N_9972,N_6972,N_6361);
nand U9973 (N_9973,N_7466,N_6810);
and U9974 (N_9974,N_7562,N_7536);
nand U9975 (N_9975,N_6774,N_7572);
nand U9976 (N_9976,N_6142,N_6286);
nor U9977 (N_9977,N_7685,N_6263);
nor U9978 (N_9978,N_7233,N_7353);
xnor U9979 (N_9979,N_7234,N_7115);
nor U9980 (N_9980,N_6533,N_7903);
nand U9981 (N_9981,N_6536,N_7100);
nor U9982 (N_9982,N_7975,N_6748);
or U9983 (N_9983,N_6853,N_7220);
or U9984 (N_9984,N_7557,N_7806);
nor U9985 (N_9985,N_7555,N_6941);
nand U9986 (N_9986,N_7057,N_6599);
or U9987 (N_9987,N_6543,N_6051);
or U9988 (N_9988,N_7857,N_6557);
nand U9989 (N_9989,N_6127,N_6413);
and U9990 (N_9990,N_6469,N_6307);
nor U9991 (N_9991,N_7205,N_6574);
xor U9992 (N_9992,N_6230,N_7876);
or U9993 (N_9993,N_7132,N_7365);
xnor U9994 (N_9994,N_7789,N_6659);
or U9995 (N_9995,N_6233,N_7322);
and U9996 (N_9996,N_7739,N_7573);
xor U9997 (N_9997,N_7325,N_6153);
or U9998 (N_9998,N_7160,N_6681);
nor U9999 (N_9999,N_7813,N_6299);
and U10000 (N_10000,N_8227,N_8661);
nand U10001 (N_10001,N_9230,N_8954);
and U10002 (N_10002,N_9714,N_9962);
nor U10003 (N_10003,N_8689,N_8885);
or U10004 (N_10004,N_9130,N_8075);
or U10005 (N_10005,N_9410,N_8360);
nor U10006 (N_10006,N_8042,N_9666);
nor U10007 (N_10007,N_9805,N_9196);
or U10008 (N_10008,N_9886,N_9832);
and U10009 (N_10009,N_8394,N_8573);
or U10010 (N_10010,N_8977,N_9577);
nor U10011 (N_10011,N_9680,N_9476);
and U10012 (N_10012,N_8780,N_9199);
or U10013 (N_10013,N_8072,N_9379);
nand U10014 (N_10014,N_8028,N_9665);
nor U10015 (N_10015,N_9361,N_8945);
xnor U10016 (N_10016,N_8578,N_9037);
nand U10017 (N_10017,N_9109,N_9801);
or U10018 (N_10018,N_8126,N_8402);
or U10019 (N_10019,N_9789,N_9466);
or U10020 (N_10020,N_9259,N_8836);
nand U10021 (N_10021,N_8988,N_9648);
xor U10022 (N_10022,N_9930,N_9946);
or U10023 (N_10023,N_9926,N_9482);
and U10024 (N_10024,N_9375,N_8163);
nor U10025 (N_10025,N_9343,N_8485);
xnor U10026 (N_10026,N_9991,N_8388);
and U10027 (N_10027,N_9241,N_8098);
or U10028 (N_10028,N_8446,N_8299);
nor U10029 (N_10029,N_8551,N_8572);
xnor U10030 (N_10030,N_8241,N_8681);
or U10031 (N_10031,N_9856,N_9568);
or U10032 (N_10032,N_9131,N_8957);
nand U10033 (N_10033,N_8368,N_9561);
or U10034 (N_10034,N_9253,N_8916);
nand U10035 (N_10035,N_9041,N_9516);
nand U10036 (N_10036,N_8853,N_8658);
nor U10037 (N_10037,N_9175,N_9281);
xnor U10038 (N_10038,N_9055,N_8191);
xnor U10039 (N_10039,N_8375,N_8674);
nand U10040 (N_10040,N_9256,N_8678);
or U10041 (N_10041,N_8708,N_9104);
and U10042 (N_10042,N_8750,N_9236);
xnor U10043 (N_10043,N_9618,N_8540);
nor U10044 (N_10044,N_8513,N_8563);
nand U10045 (N_10045,N_9066,N_9693);
nor U10046 (N_10046,N_9574,N_9077);
xor U10047 (N_10047,N_8285,N_9772);
and U10048 (N_10048,N_9933,N_9943);
or U10049 (N_10049,N_9505,N_8127);
xnor U10050 (N_10050,N_9018,N_9490);
xnor U10051 (N_10051,N_9397,N_9209);
or U10052 (N_10052,N_8065,N_9790);
or U10053 (N_10053,N_8183,N_9803);
and U10054 (N_10054,N_8649,N_9050);
or U10055 (N_10055,N_8997,N_8264);
and U10056 (N_10056,N_9558,N_8637);
nand U10057 (N_10057,N_8453,N_8574);
and U10058 (N_10058,N_9099,N_9146);
nand U10059 (N_10059,N_9826,N_9017);
nand U10060 (N_10060,N_8583,N_8426);
and U10061 (N_10061,N_8165,N_9860);
nor U10062 (N_10062,N_9087,N_9645);
and U10063 (N_10063,N_9903,N_9807);
and U10064 (N_10064,N_8137,N_9566);
and U10065 (N_10065,N_9800,N_9300);
and U10066 (N_10066,N_8892,N_8036);
nor U10067 (N_10067,N_9294,N_9553);
xnor U10068 (N_10068,N_9865,N_8272);
and U10069 (N_10069,N_8209,N_8000);
or U10070 (N_10070,N_8735,N_9634);
nor U10071 (N_10071,N_9474,N_8867);
nand U10072 (N_10072,N_9108,N_8917);
and U10073 (N_10073,N_8921,N_9782);
nand U10074 (N_10074,N_9312,N_9464);
or U10075 (N_10075,N_9461,N_9289);
nor U10076 (N_10076,N_8639,N_8123);
xor U10077 (N_10077,N_9609,N_9834);
or U10078 (N_10078,N_8675,N_9337);
and U10079 (N_10079,N_8015,N_9033);
nand U10080 (N_10080,N_9435,N_8890);
xnor U10081 (N_10081,N_8912,N_9870);
xor U10082 (N_10082,N_8259,N_8159);
or U10083 (N_10083,N_8587,N_9963);
nor U10084 (N_10084,N_9433,N_8952);
or U10085 (N_10085,N_8062,N_9625);
and U10086 (N_10086,N_9016,N_9941);
nand U10087 (N_10087,N_9092,N_9871);
or U10088 (N_10088,N_8422,N_8470);
or U10089 (N_10089,N_8635,N_9203);
or U10090 (N_10090,N_8815,N_8320);
or U10091 (N_10091,N_9023,N_8502);
xor U10092 (N_10092,N_8162,N_9849);
nor U10093 (N_10093,N_9355,N_9046);
and U10094 (N_10094,N_8330,N_8489);
and U10095 (N_10095,N_9164,N_9757);
or U10096 (N_10096,N_9346,N_8447);
and U10097 (N_10097,N_9382,N_9749);
nand U10098 (N_10098,N_9258,N_9595);
nor U10099 (N_10099,N_9949,N_9034);
nor U10100 (N_10100,N_9458,N_9310);
nand U10101 (N_10101,N_9833,N_8425);
nand U10102 (N_10102,N_8410,N_8145);
and U10103 (N_10103,N_8647,N_9938);
nand U10104 (N_10104,N_8791,N_8991);
nor U10105 (N_10105,N_8802,N_9770);
or U10106 (N_10106,N_8309,N_9855);
nand U10107 (N_10107,N_8588,N_9530);
nand U10108 (N_10108,N_9829,N_8501);
or U10109 (N_10109,N_8932,N_9897);
xnor U10110 (N_10110,N_8673,N_8367);
nor U10111 (N_10111,N_8499,N_9244);
or U10112 (N_10112,N_8033,N_8862);
nor U10113 (N_10113,N_8558,N_9389);
and U10114 (N_10114,N_8292,N_8886);
xor U10115 (N_10115,N_8773,N_9194);
nand U10116 (N_10116,N_8353,N_9787);
nand U10117 (N_10117,N_8395,N_8451);
nand U10118 (N_10118,N_8434,N_8949);
nor U10119 (N_10119,N_8757,N_8281);
nand U10120 (N_10120,N_8117,N_9811);
xnor U10121 (N_10121,N_8919,N_8129);
xor U10122 (N_10122,N_9298,N_8046);
nand U10123 (N_10123,N_8304,N_9998);
and U10124 (N_10124,N_8418,N_9740);
xnor U10125 (N_10125,N_8408,N_8414);
xnor U10126 (N_10126,N_8128,N_9135);
nand U10127 (N_10127,N_9057,N_9830);
nand U10128 (N_10128,N_9635,N_8203);
and U10129 (N_10129,N_8266,N_9073);
nand U10130 (N_10130,N_9126,N_9575);
and U10131 (N_10131,N_8239,N_9027);
nor U10132 (N_10132,N_9845,N_9081);
nor U10133 (N_10133,N_8296,N_8344);
xor U10134 (N_10134,N_8101,N_8358);
and U10135 (N_10135,N_9891,N_8920);
or U10136 (N_10136,N_8719,N_9485);
and U10137 (N_10137,N_8785,N_8595);
nor U10138 (N_10138,N_9923,N_9438);
and U10139 (N_10139,N_8923,N_9582);
or U10140 (N_10140,N_9139,N_9525);
xnor U10141 (N_10141,N_9799,N_9412);
xnor U10142 (N_10142,N_9842,N_8910);
or U10143 (N_10143,N_9548,N_9628);
nand U10144 (N_10144,N_9959,N_9650);
nand U10145 (N_10145,N_8519,N_9232);
nor U10146 (N_10146,N_8171,N_8454);
or U10147 (N_10147,N_9719,N_9419);
and U10148 (N_10148,N_8986,N_8269);
or U10149 (N_10149,N_9186,N_9174);
xnor U10150 (N_10150,N_9867,N_9528);
and U10151 (N_10151,N_9285,N_9942);
nand U10152 (N_10152,N_9824,N_9979);
nand U10153 (N_10153,N_9987,N_8534);
or U10154 (N_10154,N_9791,N_8751);
or U10155 (N_10155,N_9619,N_9908);
nor U10156 (N_10156,N_9904,N_8003);
and U10157 (N_10157,N_8354,N_8262);
xnor U10158 (N_10158,N_8657,N_8550);
and U10159 (N_10159,N_8797,N_9040);
xor U10160 (N_10160,N_9264,N_8893);
or U10161 (N_10161,N_8905,N_8077);
or U10162 (N_10162,N_9978,N_8250);
nor U10163 (N_10163,N_9712,N_9877);
nand U10164 (N_10164,N_8226,N_9899);
xnor U10165 (N_10165,N_9425,N_8745);
nor U10166 (N_10166,N_9497,N_8192);
and U10167 (N_10167,N_8788,N_9231);
nand U10168 (N_10168,N_9409,N_9990);
and U10169 (N_10169,N_8532,N_8172);
xnor U10170 (N_10170,N_8059,N_9301);
and U10171 (N_10171,N_9919,N_8160);
or U10172 (N_10172,N_8190,N_9754);
nor U10173 (N_10173,N_9658,N_9721);
or U10174 (N_10174,N_8896,N_9894);
xor U10175 (N_10175,N_9065,N_8373);
and U10176 (N_10176,N_8616,N_9111);
nand U10177 (N_10177,N_8312,N_8032);
nor U10178 (N_10178,N_9197,N_9031);
nor U10179 (N_10179,N_8477,N_9106);
nor U10180 (N_10180,N_8476,N_8242);
and U10181 (N_10181,N_9268,N_8514);
xnor U10182 (N_10182,N_9014,N_9818);
nand U10183 (N_10183,N_9171,N_9339);
nor U10184 (N_10184,N_9202,N_8288);
or U10185 (N_10185,N_9083,N_8260);
or U10186 (N_10186,N_8363,N_9150);
or U10187 (N_10187,N_8684,N_8517);
nand U10188 (N_10188,N_8467,N_9290);
nor U10189 (N_10189,N_8324,N_8630);
nor U10190 (N_10190,N_8473,N_8804);
or U10191 (N_10191,N_8733,N_9322);
and U10192 (N_10192,N_9837,N_9531);
nand U10193 (N_10193,N_9000,N_9159);
nor U10194 (N_10194,N_8759,N_8734);
and U10195 (N_10195,N_8598,N_8752);
nand U10196 (N_10196,N_8781,N_9598);
and U10197 (N_10197,N_8297,N_9205);
xnor U10198 (N_10198,N_8974,N_9667);
or U10199 (N_10199,N_8818,N_9551);
or U10200 (N_10200,N_8581,N_8186);
nor U10201 (N_10201,N_9121,N_9694);
xor U10202 (N_10202,N_9844,N_8268);
nand U10203 (N_10203,N_9659,N_9004);
nand U10204 (N_10204,N_8826,N_9679);
xnor U10205 (N_10205,N_9475,N_8557);
xnor U10206 (N_10206,N_8342,N_9736);
and U10207 (N_10207,N_8529,N_9567);
nor U10208 (N_10208,N_8727,N_8531);
and U10209 (N_10209,N_9612,N_9641);
nand U10210 (N_10210,N_8051,N_9536);
or U10211 (N_10211,N_9545,N_8010);
or U10212 (N_10212,N_9279,N_8860);
nor U10213 (N_10213,N_8692,N_9396);
nor U10214 (N_10214,N_8690,N_9304);
and U10215 (N_10215,N_9359,N_9644);
or U10216 (N_10216,N_8198,N_9215);
nand U10217 (N_10217,N_9102,N_8329);
and U10218 (N_10218,N_9292,N_8817);
xor U10219 (N_10219,N_9411,N_8984);
or U10220 (N_10220,N_8680,N_8440);
or U10221 (N_10221,N_8082,N_8141);
nand U10222 (N_10222,N_8108,N_8359);
or U10223 (N_10223,N_8486,N_8723);
and U10224 (N_10224,N_8528,N_9690);
xnor U10225 (N_10225,N_8287,N_9036);
xor U10226 (N_10226,N_9827,N_8810);
xnor U10227 (N_10227,N_8083,N_9399);
xnor U10228 (N_10228,N_9723,N_8482);
xnor U10229 (N_10229,N_8107,N_8048);
or U10230 (N_10230,N_8377,N_8475);
nand U10231 (N_10231,N_8355,N_9638);
and U10232 (N_10232,N_8423,N_9890);
or U10233 (N_10233,N_9299,N_9333);
nor U10234 (N_10234,N_8942,N_9165);
nand U10235 (N_10235,N_9936,N_8911);
nor U10236 (N_10236,N_8011,N_8922);
nor U10237 (N_10237,N_8442,N_9564);
nand U10238 (N_10238,N_8045,N_8516);
or U10239 (N_10239,N_8686,N_9413);
nor U10240 (N_10240,N_8717,N_8261);
nand U10241 (N_10241,N_8302,N_9363);
or U10242 (N_10242,N_8496,N_8877);
and U10243 (N_10243,N_8212,N_9085);
and U10244 (N_10244,N_9204,N_8668);
nor U10245 (N_10245,N_8074,N_9056);
nand U10246 (N_10246,N_8087,N_9808);
and U10247 (N_10247,N_8654,N_9585);
nor U10248 (N_10248,N_9424,N_8286);
and U10249 (N_10249,N_9738,N_8973);
nand U10250 (N_10250,N_9670,N_8390);
nor U10251 (N_10251,N_8234,N_8090);
or U10252 (N_10252,N_9030,N_8542);
nand U10253 (N_10253,N_9320,N_8953);
or U10254 (N_10254,N_9400,N_8113);
nor U10255 (N_10255,N_8216,N_8725);
nor U10256 (N_10256,N_9624,N_9814);
and U10257 (N_10257,N_9091,N_8566);
or U10258 (N_10258,N_9463,N_8707);
nor U10259 (N_10259,N_9506,N_8672);
or U10260 (N_10260,N_9900,N_9873);
and U10261 (N_10261,N_9816,N_9813);
nor U10262 (N_10262,N_9980,N_9045);
or U10263 (N_10263,N_8567,N_8962);
or U10264 (N_10264,N_8995,N_8115);
or U10265 (N_10265,N_9181,N_8197);
or U10266 (N_10266,N_8915,N_8020);
or U10267 (N_10267,N_8387,N_9927);
or U10268 (N_10268,N_9520,N_9220);
nand U10269 (N_10269,N_9539,N_8770);
nor U10270 (N_10270,N_8865,N_9513);
or U10271 (N_10271,N_9847,N_9662);
nand U10272 (N_10272,N_9348,N_8792);
nor U10273 (N_10273,N_8095,N_8136);
and U10274 (N_10274,N_8291,N_8899);
xnor U10275 (N_10275,N_8319,N_9144);
xnor U10276 (N_10276,N_9302,N_9200);
xnor U10277 (N_10277,N_8561,N_9840);
xnor U10278 (N_10278,N_9436,N_9151);
or U10279 (N_10279,N_9122,N_9010);
nand U10280 (N_10280,N_8705,N_8200);
or U10281 (N_10281,N_9327,N_9695);
or U10282 (N_10282,N_9243,N_9078);
xor U10283 (N_10283,N_8503,N_8295);
xnor U10284 (N_10284,N_9557,N_9597);
nand U10285 (N_10285,N_9542,N_9724);
or U10286 (N_10286,N_9604,N_8497);
nor U10287 (N_10287,N_9395,N_9062);
nand U10288 (N_10288,N_8432,N_8794);
and U10289 (N_10289,N_8168,N_8968);
xor U10290 (N_10290,N_9836,N_8610);
xnor U10291 (N_10291,N_9647,N_9058);
and U10292 (N_10292,N_9212,N_9535);
nand U10293 (N_10293,N_8385,N_8800);
nand U10294 (N_10294,N_9173,N_8199);
xor U10295 (N_10295,N_9495,N_8600);
xnor U10296 (N_10296,N_9885,N_8456);
xor U10297 (N_10297,N_8450,N_8498);
nand U10298 (N_10298,N_8455,N_9246);
or U10299 (N_10299,N_8652,N_8022);
nand U10300 (N_10300,N_8509,N_8691);
or U10301 (N_10301,N_8992,N_9878);
and U10302 (N_10302,N_8348,N_8131);
xnor U10303 (N_10303,N_9972,N_9201);
nor U10304 (N_10304,N_9141,N_9701);
nor U10305 (N_10305,N_8783,N_9707);
xnor U10306 (N_10306,N_8303,N_9291);
xnor U10307 (N_10307,N_8628,N_9371);
xor U10308 (N_10308,N_9123,N_9430);
nand U10309 (N_10309,N_8645,N_8118);
xnor U10310 (N_10310,N_8824,N_9858);
xnor U10311 (N_10311,N_9716,N_8270);
xnor U10312 (N_10312,N_9527,N_8060);
nor U10313 (N_10313,N_8774,N_9902);
nand U10314 (N_10314,N_8361,N_9771);
nand U10315 (N_10315,N_9912,N_8546);
nand U10316 (N_10316,N_8832,N_9169);
nand U10317 (N_10317,N_8080,N_9512);
nand U10318 (N_10318,N_9732,N_9214);
and U10319 (N_10319,N_9261,N_8933);
xor U10320 (N_10320,N_8946,N_9706);
xnor U10321 (N_10321,N_8007,N_8655);
and U10322 (N_10322,N_8006,N_9571);
nor U10323 (N_10323,N_9623,N_9052);
or U10324 (N_10324,N_9021,N_8554);
xor U10325 (N_10325,N_8530,N_9145);
xnor U10326 (N_10326,N_9937,N_9219);
xor U10327 (N_10327,N_8666,N_9893);
or U10328 (N_10328,N_8093,N_8805);
and U10329 (N_10329,N_8364,N_9002);
xor U10330 (N_10330,N_9611,N_9708);
nand U10331 (N_10331,N_9794,N_8710);
and U10332 (N_10332,N_8881,N_9443);
xor U10333 (N_10333,N_8960,N_8421);
nand U10334 (N_10334,N_8799,N_9517);
nor U10335 (N_10335,N_9183,N_8228);
xnor U10336 (N_10336,N_9850,N_8790);
xnor U10337 (N_10337,N_8584,N_8043);
and U10338 (N_10338,N_8855,N_9368);
nand U10339 (N_10339,N_8525,N_8372);
and U10340 (N_10340,N_8606,N_9705);
or U10341 (N_10341,N_9793,N_9970);
or U10342 (N_10342,N_8839,N_8591);
xor U10343 (N_10343,N_8008,N_9001);
nor U10344 (N_10344,N_8134,N_9781);
and U10345 (N_10345,N_8430,N_9133);
nand U10346 (N_10346,N_9742,N_8013);
or U10347 (N_10347,N_8976,N_9472);
xor U10348 (N_10348,N_8282,N_8850);
nor U10349 (N_10349,N_8740,N_9182);
xor U10350 (N_10350,N_9428,N_9103);
or U10351 (N_10351,N_9583,N_8934);
and U10352 (N_10352,N_9335,N_8187);
and U10353 (N_10353,N_9643,N_9616);
nand U10354 (N_10354,N_9717,N_8721);
nand U10355 (N_10355,N_8362,N_8906);
nand U10356 (N_10356,N_8184,N_8274);
nand U10357 (N_10357,N_8771,N_8100);
nand U10358 (N_10358,N_8125,N_8088);
xor U10359 (N_10359,N_8883,N_9272);
nand U10360 (N_10360,N_9263,N_8135);
and U10361 (N_10361,N_8903,N_8963);
xnor U10362 (N_10362,N_9600,N_8601);
nor U10363 (N_10363,N_9418,N_8222);
nor U10364 (N_10364,N_8267,N_9550);
or U10365 (N_10365,N_9935,N_9415);
and U10366 (N_10366,N_8146,N_9391);
or U10367 (N_10367,N_8869,N_8712);
xor U10368 (N_10368,N_9007,N_9688);
nand U10369 (N_10369,N_9627,N_9277);
or U10370 (N_10370,N_9009,N_8806);
xor U10371 (N_10371,N_8050,N_9589);
nor U10372 (N_10372,N_8596,N_9608);
and U10373 (N_10373,N_8902,N_8311);
nor U10374 (N_10374,N_9297,N_8170);
and U10375 (N_10375,N_9426,N_9768);
and U10376 (N_10376,N_9154,N_8218);
xnor U10377 (N_10377,N_8687,N_9168);
nand U10378 (N_10378,N_9269,N_8258);
nor U10379 (N_10379,N_8801,N_9500);
or U10380 (N_10380,N_9431,N_9654);
and U10381 (N_10381,N_8640,N_9223);
or U10382 (N_10382,N_8256,N_8114);
xor U10383 (N_10383,N_9163,N_8961);
nor U10384 (N_10384,N_9465,N_9462);
nor U10385 (N_10385,N_9118,N_8054);
and U10386 (N_10386,N_9629,N_9861);
or U10387 (N_10387,N_8586,N_8231);
and U10388 (N_10388,N_8615,N_9709);
nand U10389 (N_10389,N_9868,N_9866);
nand U10390 (N_10390,N_8769,N_9445);
and U10391 (N_10391,N_8180,N_9649);
xor U10392 (N_10392,N_9427,N_9778);
nor U10393 (N_10393,N_9317,N_8807);
and U10394 (N_10394,N_9821,N_8958);
or U10395 (N_10395,N_9915,N_8061);
xor U10396 (N_10396,N_9332,N_9839);
or U10397 (N_10397,N_8289,N_8702);
nand U10398 (N_10398,N_9284,N_9370);
or U10399 (N_10399,N_9934,N_8732);
xor U10400 (N_10400,N_9697,N_9115);
xnor U10401 (N_10401,N_9968,N_9404);
and U10402 (N_10402,N_9766,N_8219);
and U10403 (N_10403,N_9555,N_8429);
xnor U10404 (N_10404,N_8392,N_9112);
and U10405 (N_10405,N_8709,N_8111);
nor U10406 (N_10406,N_8398,N_9931);
xor U10407 (N_10407,N_8469,N_9082);
nand U10408 (N_10408,N_9526,N_8808);
or U10409 (N_10409,N_9470,N_9060);
nor U10410 (N_10410,N_8603,N_8841);
and U10411 (N_10411,N_9751,N_8458);
nor U10412 (N_10412,N_9592,N_8318);
xor U10413 (N_10413,N_8873,N_8547);
xor U10414 (N_10414,N_8279,N_8030);
nand U10415 (N_10415,N_8173,N_9964);
or U10416 (N_10416,N_9533,N_8230);
nand U10417 (N_10417,N_9384,N_8164);
or U10418 (N_10418,N_8122,N_9651);
or U10419 (N_10419,N_9313,N_9992);
xnor U10420 (N_10420,N_8938,N_9234);
nor U10421 (N_10421,N_8357,N_8156);
nor U10422 (N_10422,N_8576,N_8907);
and U10423 (N_10423,N_9765,N_9210);
nand U10424 (N_10424,N_9718,N_8564);
or U10425 (N_10425,N_8491,N_9601);
xnor U10426 (N_10426,N_9248,N_9660);
or U10427 (N_10427,N_9483,N_8848);
nor U10428 (N_10428,N_9161,N_8820);
nor U10429 (N_10429,N_9906,N_9067);
nand U10430 (N_10430,N_8474,N_9090);
nor U10431 (N_10431,N_8592,N_9344);
or U10432 (N_10432,N_8631,N_9510);
nor U10433 (N_10433,N_9563,N_8724);
nand U10434 (N_10434,N_8646,N_9167);
and U10435 (N_10435,N_8047,N_8851);
nand U10436 (N_10436,N_8021,N_8238);
nor U10437 (N_10437,N_9993,N_8811);
and U10438 (N_10438,N_8293,N_8328);
and U10439 (N_10439,N_8510,N_8849);
nor U10440 (N_10440,N_8055,N_9098);
and U10441 (N_10441,N_9823,N_8271);
nand U10442 (N_10442,N_8948,N_8351);
nor U10443 (N_10443,N_8908,N_9127);
or U10444 (N_10444,N_9459,N_9283);
xnor U10445 (N_10445,N_9704,N_8703);
or U10446 (N_10446,N_8374,N_9245);
nor U10447 (N_10447,N_9812,N_9769);
and U10448 (N_10448,N_9452,N_9072);
xnor U10449 (N_10449,N_8431,N_8436);
or U10450 (N_10450,N_9969,N_8753);
and U10451 (N_10451,N_8301,N_8210);
nor U10452 (N_10452,N_8859,N_9351);
and U10453 (N_10453,N_8428,N_8660);
and U10454 (N_10454,N_9522,N_9883);
nand U10455 (N_10455,N_8110,N_8812);
nand U10456 (N_10456,N_8931,N_8864);
and U10457 (N_10457,N_9255,N_9270);
xnor U10458 (N_10458,N_8840,N_8939);
and U10459 (N_10459,N_9663,N_8393);
and U10460 (N_10460,N_8955,N_9854);
xor U10461 (N_10461,N_9652,N_9869);
nand U10462 (N_10462,N_9828,N_9124);
xor U10463 (N_10463,N_9994,N_8167);
and U10464 (N_10464,N_9989,N_9080);
or U10465 (N_10465,N_8989,N_8221);
nor U10466 (N_10466,N_8625,N_9636);
xor U10467 (N_10467,N_9341,N_8380);
and U10468 (N_10468,N_8665,N_9190);
nand U10469 (N_10469,N_9703,N_8208);
nand U10470 (N_10470,N_9094,N_8755);
nor U10471 (N_10471,N_9921,N_9511);
or U10472 (N_10472,N_8166,N_9074);
or U10473 (N_10473,N_9982,N_8336);
nor U10474 (N_10474,N_9493,N_9362);
or U10475 (N_10475,N_8343,N_9044);
nor U10476 (N_10476,N_9398,N_8798);
nand U10477 (N_10477,N_8814,N_9773);
xnor U10478 (N_10478,N_9226,N_9977);
nor U10479 (N_10479,N_8760,N_8994);
nand U10480 (N_10480,N_9965,N_9119);
or U10481 (N_10481,N_9729,N_9653);
and U10482 (N_10482,N_9365,N_9378);
and U10483 (N_10483,N_8403,N_8768);
nor U10484 (N_10484,N_8452,N_9606);
nor U10485 (N_10485,N_9222,N_9184);
and U10486 (N_10486,N_9071,N_9988);
nor U10487 (N_10487,N_8073,N_8838);
or U10488 (N_10488,N_8878,N_9314);
and U10489 (N_10489,N_9621,N_9380);
nand U10490 (N_10490,N_8650,N_8555);
and U10491 (N_10491,N_9862,N_8697);
xnor U10492 (N_10492,N_8322,N_8070);
nor U10493 (N_10493,N_9013,N_9125);
or U10494 (N_10494,N_8831,N_8633);
nand U10495 (N_10495,N_9678,N_8682);
and U10496 (N_10496,N_8492,N_8144);
xor U10497 (N_10497,N_9468,N_8715);
nand U10498 (N_10498,N_9615,N_9939);
nand U10499 (N_10499,N_9831,N_9405);
nand U10500 (N_10500,N_8830,N_8305);
nand U10501 (N_10501,N_9213,N_9851);
and U10502 (N_10502,N_9274,N_8505);
and U10503 (N_10503,N_9967,N_8121);
nor U10504 (N_10504,N_8593,N_9806);
nor U10505 (N_10505,N_8809,N_9105);
or U10506 (N_10506,N_9143,N_8914);
nand U10507 (N_10507,N_9265,N_9003);
xor U10508 (N_10508,N_8462,N_9129);
xnor U10509 (N_10509,N_8659,N_8204);
nand U10510 (N_10510,N_8016,N_8928);
and U10511 (N_10511,N_9918,N_9664);
and U10512 (N_10512,N_8420,N_8834);
and U10513 (N_10513,N_9407,N_8941);
nor U10514 (N_10514,N_8313,N_8688);
xor U10515 (N_10515,N_9944,N_9315);
nor U10516 (N_10516,N_9096,N_9590);
or U10517 (N_10517,N_8323,N_8205);
and U10518 (N_10518,N_9329,N_9737);
nand U10519 (N_10519,N_9309,N_8193);
and U10520 (N_10520,N_8527,N_9100);
and U10521 (N_10521,N_9889,N_9120);
and U10522 (N_10522,N_8488,N_8972);
nand U10523 (N_10523,N_9477,N_8026);
xor U10524 (N_10524,N_8177,N_9841);
and U10525 (N_10525,N_8930,N_9288);
or U10526 (N_10526,N_8448,N_8762);
xnor U10527 (N_10527,N_8944,N_8176);
xnor U10528 (N_10528,N_8314,N_8504);
xor U10529 (N_10529,N_8823,N_9605);
nor U10530 (N_10530,N_8449,N_8148);
xor U10531 (N_10531,N_9024,N_8178);
xor U10532 (N_10532,N_9012,N_8718);
and U10533 (N_10533,N_9153,N_8340);
nand U10534 (N_10534,N_9776,N_8653);
nor U10535 (N_10535,N_8094,N_9881);
or U10536 (N_10536,N_8726,N_9086);
xor U10537 (N_10537,N_9626,N_8866);
and U10538 (N_10538,N_9392,N_9211);
and U10539 (N_10539,N_8552,N_9715);
and U10540 (N_10540,N_8404,N_9759);
nor U10541 (N_10541,N_9677,N_9049);
xnor U10542 (N_10542,N_8993,N_9432);
or U10543 (N_10543,N_8443,N_8133);
nor U10544 (N_10544,N_8844,N_8777);
nand U10545 (N_10545,N_8063,N_9913);
nor U10546 (N_10546,N_8679,N_9884);
nor U10547 (N_10547,N_9882,N_8396);
nand U10548 (N_10548,N_8700,N_9306);
nand U10549 (N_10549,N_9479,N_8220);
and U10550 (N_10550,N_8037,N_9579);
and U10551 (N_10551,N_8966,N_9303);
xnor U10552 (N_10552,N_9385,N_8427);
or U10553 (N_10553,N_9328,N_9570);
or U10554 (N_10554,N_8255,N_8294);
and U10555 (N_10555,N_8049,N_9838);
nand U10556 (N_10556,N_9743,N_9434);
xor U10557 (N_10557,N_9494,N_8959);
nor U10558 (N_10558,N_9491,N_9504);
and U10559 (N_10559,N_8276,N_9429);
nor U10560 (N_10560,N_8782,N_9307);
xor U10561 (N_10561,N_9975,N_9581);
and U10562 (N_10562,N_9673,N_8696);
or U10563 (N_10563,N_9916,N_8251);
nor U10564 (N_10564,N_8150,N_8109);
nand U10565 (N_10565,N_9971,N_8580);
nand U10566 (N_10566,N_9305,N_8597);
or U10567 (N_10567,N_8412,N_8904);
xor U10568 (N_10568,N_9521,N_8982);
nand U10569 (N_10569,N_8548,N_8341);
and U10570 (N_10570,N_9725,N_8787);
nand U10571 (N_10571,N_9901,N_9321);
xor U10572 (N_10572,N_9720,N_9880);
nand U10573 (N_10573,N_8099,N_9039);
or U10574 (N_10574,N_9020,N_8175);
or U10575 (N_10575,N_9614,N_8002);
xor U10576 (N_10576,N_9848,N_9981);
and U10577 (N_10577,N_8215,N_9417);
or U10578 (N_10578,N_9138,N_8536);
nor U10579 (N_10579,N_9997,N_9674);
nor U10580 (N_10580,N_9722,N_8089);
nor U10581 (N_10581,N_9110,N_9689);
and U10582 (N_10582,N_9602,N_8041);
nor U10583 (N_10583,N_8518,N_9480);
nor U10584 (N_10584,N_9691,N_9364);
and U10585 (N_10585,N_9532,N_9198);
and U10586 (N_10586,N_9353,N_9043);
nand U10587 (N_10587,N_8748,N_9961);
xor U10588 (N_10588,N_9180,N_9745);
and U10589 (N_10589,N_8460,N_8971);
and U10590 (N_10590,N_9454,N_9763);
nand U10591 (N_10591,N_9026,N_9661);
nor U10592 (N_10592,N_8409,N_9273);
or U10593 (N_10593,N_8439,N_8711);
nand U10594 (N_10594,N_8181,N_8280);
nor U10595 (N_10595,N_9107,N_8039);
or U10596 (N_10596,N_9656,N_9051);
xnor U10597 (N_10597,N_8024,N_9455);
or U10598 (N_10598,N_8034,N_8624);
and U10599 (N_10599,N_9240,N_8594);
nor U10600 (N_10600,N_9149,N_8506);
xor U10601 (N_10601,N_8669,N_9170);
nand U10602 (N_10602,N_9408,N_8213);
nand U10603 (N_10603,N_8943,N_9403);
nand U10604 (N_10604,N_9367,N_8520);
and U10605 (N_10605,N_8092,N_8901);
nor U10606 (N_10606,N_8875,N_8614);
xnor U10607 (N_10607,N_9179,N_9330);
xnor U10608 (N_10608,N_9529,N_8999);
xnor U10609 (N_10609,N_8233,N_9448);
and U10610 (N_10610,N_9334,N_8683);
or U10611 (N_10611,N_9728,N_9177);
nor U10612 (N_10612,N_8067,N_9336);
nand U10613 (N_10613,N_8940,N_8803);
xnor U10614 (N_10614,N_9888,N_8185);
xor U10615 (N_10615,N_8854,N_9857);
nor U10616 (N_10616,N_9762,N_8174);
nor U10617 (N_10617,N_9217,N_8217);
xor U10618 (N_10618,N_8613,N_9879);
xor U10619 (N_10619,N_9549,N_8334);
or U10620 (N_10620,N_9218,N_8626);
and U10621 (N_10621,N_8487,N_8868);
and U10622 (N_10622,N_8909,N_9233);
nand U10623 (N_10623,N_8521,N_8339);
nor U10624 (N_10624,N_8981,N_9733);
xnor U10625 (N_10625,N_9785,N_9756);
or U10626 (N_10626,N_9859,N_8085);
or U10627 (N_10627,N_9178,N_9457);
and U10628 (N_10628,N_8382,N_8035);
nor U10629 (N_10629,N_9132,N_8068);
or U10630 (N_10630,N_8979,N_9795);
nor U10631 (N_10631,N_9402,N_9358);
and U10632 (N_10632,N_9249,N_9376);
xor U10633 (N_10633,N_9158,N_8247);
nand U10634 (N_10634,N_8612,N_9280);
and U10635 (N_10635,N_8964,N_8772);
nand U10636 (N_10636,N_8017,N_9565);
or U10637 (N_10637,N_9922,N_8664);
xor U10638 (N_10638,N_9774,N_8913);
nand U10639 (N_10639,N_8196,N_8463);
or U10640 (N_10640,N_9503,N_8722);
and U10641 (N_10641,N_9239,N_9788);
and U10642 (N_10642,N_8438,N_9917);
nand U10643 (N_10643,N_9610,N_9669);
and U10644 (N_10644,N_8194,N_8562);
nand U10645 (N_10645,N_8369,N_8401);
or U10646 (N_10646,N_8605,N_9440);
nand U10647 (N_10647,N_8371,N_8257);
nor U10648 (N_10648,N_9140,N_8023);
and U10649 (N_10649,N_8819,N_8656);
nand U10650 (N_10650,N_9746,N_9655);
or U10651 (N_10651,N_9576,N_8816);
nor U10652 (N_10652,N_8927,N_9599);
or U10653 (N_10653,N_8179,N_8124);
or U10654 (N_10654,N_9887,N_9986);
and U10655 (N_10655,N_8967,N_9038);
or U10656 (N_10656,N_9646,N_8437);
or U10657 (N_10657,N_8478,N_8829);
nor U10658 (N_10658,N_8764,N_9925);
xor U10659 (N_10659,N_8161,N_9537);
and U10660 (N_10660,N_9955,N_8189);
or U10661 (N_10661,N_8766,N_8120);
xnor U10662 (N_10662,N_8157,N_8663);
or U10663 (N_10663,N_9456,N_8706);
nand U10664 (N_10664,N_9741,N_9898);
and U10665 (N_10665,N_9948,N_8779);
xnor U10666 (N_10666,N_9326,N_9488);
nor U10667 (N_10667,N_9632,N_8714);
xnor U10668 (N_10668,N_8796,N_9172);
and U10669 (N_10669,N_9254,N_9095);
and U10670 (N_10670,N_8424,N_9401);
or U10671 (N_10671,N_9687,N_8151);
or U10672 (N_10672,N_9137,N_9267);
nor U10673 (N_10673,N_8545,N_9995);
nand U10674 (N_10674,N_8698,N_9113);
nor U10675 (N_10675,N_9560,N_9872);
xor U10676 (N_10676,N_8263,N_8602);
and U10677 (N_10677,N_9069,N_8195);
nand U10678 (N_10678,N_8240,N_8879);
nor U10679 (N_10679,N_9029,N_9815);
nand U10680 (N_10680,N_9668,N_8352);
xnor U10681 (N_10681,N_8575,N_9508);
or U10682 (N_10682,N_8321,N_8347);
nand U10683 (N_10683,N_8604,N_8139);
and U10684 (N_10684,N_8880,N_8356);
nand U10685 (N_10685,N_9338,N_9206);
or U10686 (N_10686,N_8335,N_9097);
and U10687 (N_10687,N_8627,N_8538);
nand U10688 (N_10688,N_9414,N_8894);
xor U10689 (N_10689,N_8887,N_9620);
nand U10690 (N_10690,N_9640,N_9752);
nand U10691 (N_10691,N_9958,N_9686);
nand U10692 (N_10692,N_9999,N_9562);
or U10693 (N_10693,N_8490,N_9515);
nand U10694 (N_10694,N_9657,N_9863);
xnor U10695 (N_10695,N_8747,N_9798);
nand U10696 (N_10696,N_9032,N_8307);
nand U10697 (N_10697,N_8632,N_9775);
xnor U10698 (N_10698,N_9940,N_9698);
nor U10699 (N_10699,N_9155,N_8214);
xnor U10700 (N_10700,N_9156,N_9473);
and U10701 (N_10701,N_8235,N_9260);
xnor U10702 (N_10702,N_9498,N_9054);
or U10703 (N_10703,N_8524,N_9372);
xnor U10704 (N_10704,N_8852,N_9381);
nor U10705 (N_10705,N_9420,N_9366);
or U10706 (N_10706,N_8236,N_9726);
and U10707 (N_10707,N_9286,N_9323);
and U10708 (N_10708,N_8225,N_8756);
xor U10709 (N_10709,N_9932,N_8029);
nand U10710 (N_10710,N_8936,N_8622);
nand U10711 (N_10711,N_8599,N_8253);
xnor U10712 (N_10712,N_8076,N_9804);
or U10713 (N_10713,N_8778,N_8386);
xnor U10714 (N_10714,N_8104,N_9053);
nor U10715 (N_10715,N_8978,N_8677);
or U10716 (N_10716,N_8027,N_8623);
or U10717 (N_10717,N_8577,N_8246);
nand U10718 (N_10718,N_8201,N_8856);
nor U10719 (N_10719,N_9594,N_9262);
nor U10720 (N_10720,N_8248,N_9406);
and U10721 (N_10721,N_9817,N_8758);
or U10722 (N_10722,N_8419,N_8644);
and U10723 (N_10723,N_8445,N_8541);
or U10724 (N_10724,N_9896,N_8019);
xnor U10725 (N_10725,N_8537,N_8106);
and U10726 (N_10726,N_8071,N_9221);
and U10727 (N_10727,N_9633,N_8847);
and U10728 (N_10728,N_8483,N_8332);
nand U10729 (N_10729,N_8947,N_8565);
and U10730 (N_10730,N_8776,N_9193);
nor U10731 (N_10731,N_8091,N_9059);
nor U10732 (N_10732,N_9509,N_9192);
or U10733 (N_10733,N_9852,N_8956);
or U10734 (N_10734,N_9784,N_8457);
xnor U10735 (N_10735,N_9188,N_9252);
or U10736 (N_10736,N_9682,N_9622);
nor U10737 (N_10737,N_8998,N_8618);
and U10738 (N_10738,N_8784,N_9699);
and U10739 (N_10739,N_8699,N_8265);
nand U10740 (N_10740,N_9453,N_9064);
nand U10741 (N_10741,N_9907,N_8694);
and U10742 (N_10742,N_8370,N_9136);
xnor U10743 (N_10743,N_9352,N_9349);
xor U10744 (N_10744,N_9700,N_8500);
nand U10745 (N_10745,N_9481,N_9208);
or U10746 (N_10746,N_8872,N_8407);
xnor U10747 (N_10747,N_9157,N_9713);
nor U10748 (N_10748,N_9764,N_9547);
and U10749 (N_10749,N_8112,N_8619);
nor U10750 (N_10750,N_8132,N_8924);
or U10751 (N_10751,N_8290,N_9727);
nor U10752 (N_10752,N_9388,N_9390);
or U10753 (N_10753,N_9676,N_9166);
or U10754 (N_10754,N_9028,N_8481);
nor U10755 (N_10755,N_9631,N_9295);
and U10756 (N_10756,N_9681,N_8079);
nand U10757 (N_10757,N_8084,N_9584);
nor U10758 (N_10758,N_9683,N_9162);
xor U10759 (N_10759,N_9296,N_9238);
or U10760 (N_10760,N_9541,N_8950);
and U10761 (N_10761,N_9393,N_8786);
or U10762 (N_10762,N_9947,N_9487);
and U10763 (N_10763,N_8086,N_9325);
xor U10764 (N_10764,N_8479,N_8549);
nand U10765 (N_10765,N_9437,N_8105);
and U10766 (N_10766,N_9318,N_9731);
nand U10767 (N_10767,N_8767,N_9777);
or U10768 (N_10768,N_9853,N_9596);
nand U10769 (N_10769,N_8638,N_8040);
or U10770 (N_10770,N_9101,N_8582);
or U10771 (N_10771,N_8237,N_8158);
and U10772 (N_10772,N_9360,N_8965);
or U10773 (N_10773,N_8278,N_9518);
or U10774 (N_10774,N_8069,N_8254);
nand U10775 (N_10775,N_9760,N_8397);
or U10776 (N_10776,N_9331,N_8651);
nor U10777 (N_10777,N_8739,N_9696);
nand U10778 (N_10778,N_9451,N_8898);
nand U10779 (N_10779,N_9953,N_8742);
xnor U10780 (N_10780,N_8789,N_9282);
or U10781 (N_10781,N_9460,N_8140);
nor U10782 (N_10782,N_8466,N_8730);
nor U10783 (N_10783,N_9734,N_8444);
or U10784 (N_10784,N_9876,N_8746);
and U10785 (N_10785,N_9984,N_9523);
nand U10786 (N_10786,N_8232,N_9779);
nor U10787 (N_10787,N_8081,N_8900);
xor U10788 (N_10788,N_9735,N_9187);
nor U10789 (N_10789,N_8889,N_9819);
nand U10790 (N_10790,N_9496,N_8980);
nor U10791 (N_10791,N_8793,N_8471);
nor U10792 (N_10792,N_8389,N_8337);
or U10793 (N_10793,N_8837,N_9767);
and U10794 (N_10794,N_8495,N_8152);
or U10795 (N_10795,N_8147,N_9189);
nand U10796 (N_10796,N_8569,N_8493);
or U10797 (N_10797,N_8641,N_8737);
nand U10798 (N_10798,N_9357,N_9802);
or U10799 (N_10799,N_9637,N_8004);
and U10800 (N_10800,N_9761,N_8202);
or U10801 (N_10801,N_9786,N_8713);
and U10802 (N_10802,N_8349,N_9228);
nor U10803 (N_10803,N_9195,N_8350);
xnor U10804 (N_10804,N_9247,N_8685);
nor U10805 (N_10805,N_9809,N_8053);
xnor U10806 (N_10806,N_8828,N_8102);
nor U10807 (N_10807,N_9237,N_8097);
or U10808 (N_10808,N_9369,N_8507);
xor U10809 (N_10809,N_8138,N_9783);
or U10810 (N_10810,N_9711,N_9546);
nand U10811 (N_10811,N_9976,N_8842);
nand U10812 (N_10812,N_9895,N_9552);
nand U10813 (N_10813,N_8858,N_9758);
or U10814 (N_10814,N_9702,N_9910);
nand U10815 (N_10815,N_9499,N_8951);
and U10816 (N_10816,N_9928,N_8249);
nor U10817 (N_10817,N_8895,N_9954);
nor U10818 (N_10818,N_9951,N_8935);
nand U10819 (N_10819,N_9047,N_9797);
nand U10820 (N_10820,N_8560,N_8025);
or U10821 (N_10821,N_8720,N_8996);
xor U10822 (N_10822,N_8704,N_9920);
or U10823 (N_10823,N_9675,N_9242);
and U10824 (N_10824,N_8435,N_9063);
xor U10825 (N_10825,N_9471,N_9191);
and U10826 (N_10826,N_9739,N_9973);
and U10827 (N_10827,N_9974,N_9792);
and U10828 (N_10828,N_8399,N_9117);
xnor U10829 (N_10829,N_9005,N_9316);
nand U10830 (N_10830,N_9810,N_9588);
nand U10831 (N_10831,N_9914,N_9229);
nor U10832 (N_10832,N_9755,N_8897);
xor U10833 (N_10833,N_8001,N_8472);
xor U10834 (N_10834,N_8662,N_8512);
nor U10835 (N_10835,N_9075,N_8544);
and U10836 (N_10836,N_8012,N_9613);
nand U10837 (N_10837,N_9266,N_9324);
xor U10838 (N_10838,N_9492,N_8005);
or U10839 (N_10839,N_9985,N_9672);
xnor U10840 (N_10840,N_9484,N_8031);
and U10841 (N_10841,N_8857,N_9543);
and U10842 (N_10842,N_8511,N_8821);
nand U10843 (N_10843,N_9011,N_9275);
nor U10844 (N_10844,N_8273,N_9554);
and U10845 (N_10845,N_8738,N_9394);
nand U10846 (N_10846,N_8096,N_8835);
or U10847 (N_10847,N_8153,N_8813);
xnor U10848 (N_10848,N_8570,N_9084);
xor U10849 (N_10849,N_8741,N_8579);
nor U10850 (N_10850,N_9416,N_9572);
nand U10851 (N_10851,N_9386,N_9593);
nor U10852 (N_10852,N_9905,N_8515);
xor U10853 (N_10853,N_9287,N_8338);
or U10854 (N_10854,N_8775,N_8381);
or U10855 (N_10855,N_9607,N_9293);
nand U10856 (N_10856,N_8252,N_8494);
nor U10857 (N_10857,N_8882,N_9671);
or U10858 (N_10858,N_8667,N_9446);
xnor U10859 (N_10859,N_9070,N_8103);
or U10860 (N_10860,N_8441,N_8413);
or U10861 (N_10861,N_8155,N_9642);
or U10862 (N_10862,N_8078,N_8308);
nand U10863 (N_10863,N_9796,N_8317);
and U10864 (N_10864,N_8559,N_8018);
xnor U10865 (N_10865,N_9354,N_8316);
or U10866 (N_10866,N_8629,N_8188);
and U10867 (N_10867,N_8611,N_9825);
or U10868 (N_10868,N_9076,N_9983);
and U10869 (N_10869,N_9134,N_9311);
xor U10870 (N_10870,N_8621,N_8736);
nor U10871 (N_10871,N_9068,N_8609);
xnor U10872 (N_10872,N_8891,N_8607);
nand U10873 (N_10873,N_8553,N_8376);
or U10874 (N_10874,N_8244,N_9350);
nor U10875 (N_10875,N_9225,N_8416);
and U10876 (N_10876,N_9250,N_8384);
or U10877 (N_10877,N_8333,N_9586);
xor U10878 (N_10878,N_8636,N_9780);
nor U10879 (N_10879,N_8671,N_9128);
xor U10880 (N_10880,N_8417,N_9875);
or U10881 (N_10881,N_9227,N_8822);
nand U10882 (N_10882,N_8731,N_8038);
and U10883 (N_10883,N_9820,N_8585);
nand U10884 (N_10884,N_9556,N_9093);
nand U10885 (N_10885,N_9692,N_8009);
nand U10886 (N_10886,N_8224,N_8533);
nor U10887 (N_10887,N_8876,N_8014);
xor U10888 (N_10888,N_9630,N_8058);
nor U10889 (N_10889,N_9148,N_8643);
and U10890 (N_10890,N_8149,N_9540);
xor U10891 (N_10891,N_9501,N_9449);
nand U10892 (N_10892,N_9750,N_9079);
or U10893 (N_10893,N_8365,N_8245);
nor U10894 (N_10894,N_8464,N_8182);
nand U10895 (N_10895,N_9929,N_8535);
nor U10896 (N_10896,N_9224,N_9015);
xnor U10897 (N_10897,N_8116,N_9088);
and U10898 (N_10898,N_8484,N_9061);
and U10899 (N_10899,N_9048,N_9278);
or U10900 (N_10900,N_9603,N_8937);
nand U10901 (N_10901,N_8670,N_8845);
nor U10902 (N_10902,N_8379,N_8154);
nor U10903 (N_10903,N_8975,N_8743);
or U10904 (N_10904,N_9469,N_9373);
and U10905 (N_10905,N_9892,N_9639);
or U10906 (N_10906,N_8763,N_8056);
and U10907 (N_10907,N_8130,N_8676);
xnor U10908 (N_10908,N_9035,N_8143);
nand U10909 (N_10909,N_9347,N_8874);
and U10910 (N_10910,N_9569,N_9152);
nand U10911 (N_10911,N_9374,N_8985);
xnor U10912 (N_10912,N_9216,N_9960);
and U10913 (N_10913,N_9864,N_9843);
xnor U10914 (N_10914,N_8325,N_9846);
nand U10915 (N_10915,N_8729,N_8526);
xor U10916 (N_10916,N_8523,N_9423);
nand U10917 (N_10917,N_9514,N_9486);
and U10918 (N_10918,N_9956,N_8620);
and U10919 (N_10919,N_8391,N_8701);
and U10920 (N_10920,N_9019,N_9909);
xnor U10921 (N_10921,N_8648,N_8990);
or U10922 (N_10922,N_9685,N_9578);
or U10923 (N_10923,N_8211,N_8207);
or U10924 (N_10924,N_9489,N_9952);
or U10925 (N_10925,N_8617,N_9271);
and U10926 (N_10926,N_9251,N_8884);
and U10927 (N_10927,N_8761,N_8556);
xnor U10928 (N_10928,N_8433,N_8406);
and U10929 (N_10929,N_9753,N_9684);
or U10930 (N_10930,N_9022,N_8833);
nor U10931 (N_10931,N_8749,N_9116);
nor U10932 (N_10932,N_8508,N_8223);
nor U10933 (N_10933,N_8987,N_9276);
nand U10934 (N_10934,N_8983,N_9114);
or U10935 (N_10935,N_8795,N_9559);
xor U10936 (N_10936,N_8522,N_9441);
xnor U10937 (N_10937,N_9383,N_8044);
nand U10938 (N_10938,N_8843,N_9387);
nor U10939 (N_10939,N_8608,N_8589);
xor U10940 (N_10940,N_9008,N_9710);
nor U10941 (N_10941,N_8366,N_8693);
or U10942 (N_10942,N_8926,N_9006);
xnor U10943 (N_10943,N_9147,N_8744);
nor U10944 (N_10944,N_8052,N_9502);
nand U10945 (N_10945,N_8825,N_9207);
or U10946 (N_10946,N_9345,N_8411);
xor U10947 (N_10947,N_8465,N_9235);
xor U10948 (N_10948,N_8861,N_9340);
or U10949 (N_10949,N_8243,N_9911);
nor U10950 (N_10950,N_8765,N_8277);
and U10951 (N_10951,N_9748,N_9587);
nor U10952 (N_10952,N_9447,N_8066);
or U10953 (N_10953,N_9996,N_8306);
and U10954 (N_10954,N_8863,N_8400);
nand U10955 (N_10955,N_8754,N_9342);
nor U10956 (N_10956,N_8275,N_9730);
xor U10957 (N_10957,N_9747,N_9874);
xnor U10958 (N_10958,N_8480,N_8571);
or U10959 (N_10959,N_8539,N_9089);
nor U10960 (N_10960,N_9591,N_9308);
nor U10961 (N_10961,N_9444,N_8870);
or U10962 (N_10962,N_9319,N_8300);
nand U10963 (N_10963,N_9478,N_8716);
or U10964 (N_10964,N_8543,N_9534);
and U10965 (N_10965,N_8695,N_8728);
nor U10966 (N_10966,N_9025,N_9257);
or U10967 (N_10967,N_9467,N_8568);
and U10968 (N_10968,N_8827,N_8970);
or U10969 (N_10969,N_9356,N_8929);
or U10970 (N_10970,N_8415,N_9185);
xor U10971 (N_10971,N_8383,N_9945);
nor U10972 (N_10972,N_8590,N_9142);
xor U10973 (N_10973,N_9377,N_8064);
and U10974 (N_10974,N_9042,N_8345);
nor U10975 (N_10975,N_9957,N_8310);
or U10976 (N_10976,N_8326,N_8405);
or U10977 (N_10977,N_8298,N_8057);
and U10978 (N_10978,N_9422,N_9507);
or U10979 (N_10979,N_9519,N_8315);
xor U10980 (N_10980,N_8346,N_8119);
nand U10981 (N_10981,N_8229,N_8206);
xor U10982 (N_10982,N_8459,N_8283);
or U10983 (N_10983,N_9524,N_9160);
or U10984 (N_10984,N_9617,N_9835);
xor U10985 (N_10985,N_8327,N_9439);
nand U10986 (N_10986,N_8925,N_8331);
and U10987 (N_10987,N_8461,N_8888);
and U10988 (N_10988,N_8871,N_8846);
nor U10989 (N_10989,N_9950,N_8468);
nand U10990 (N_10990,N_9442,N_9544);
and U10991 (N_10991,N_9573,N_8642);
or U10992 (N_10992,N_9450,N_8634);
xnor U10993 (N_10993,N_9744,N_8918);
nand U10994 (N_10994,N_8969,N_9924);
and U10995 (N_10995,N_8378,N_8142);
nand U10996 (N_10996,N_8169,N_9538);
or U10997 (N_10997,N_9176,N_9421);
nor U10998 (N_10998,N_9966,N_9822);
and U10999 (N_10999,N_9580,N_8284);
and U11000 (N_11000,N_9396,N_9789);
or U11001 (N_11001,N_9443,N_9273);
or U11002 (N_11002,N_8738,N_8598);
or U11003 (N_11003,N_9884,N_9388);
nor U11004 (N_11004,N_9111,N_8072);
and U11005 (N_11005,N_8285,N_8364);
nand U11006 (N_11006,N_9753,N_9573);
xor U11007 (N_11007,N_8161,N_9143);
and U11008 (N_11008,N_9720,N_9798);
or U11009 (N_11009,N_8696,N_8752);
or U11010 (N_11010,N_9011,N_9186);
xor U11011 (N_11011,N_9781,N_9582);
and U11012 (N_11012,N_8927,N_9420);
nor U11013 (N_11013,N_9303,N_9667);
and U11014 (N_11014,N_9732,N_8424);
and U11015 (N_11015,N_9776,N_8683);
or U11016 (N_11016,N_9161,N_9250);
and U11017 (N_11017,N_9435,N_8041);
nand U11018 (N_11018,N_8916,N_9180);
and U11019 (N_11019,N_9318,N_8782);
and U11020 (N_11020,N_8031,N_8326);
nor U11021 (N_11021,N_9409,N_8879);
xnor U11022 (N_11022,N_8653,N_8964);
or U11023 (N_11023,N_8689,N_8800);
and U11024 (N_11024,N_9114,N_8810);
or U11025 (N_11025,N_9952,N_9327);
nand U11026 (N_11026,N_9973,N_8685);
or U11027 (N_11027,N_9551,N_9036);
or U11028 (N_11028,N_8733,N_9627);
nand U11029 (N_11029,N_9722,N_8944);
or U11030 (N_11030,N_9154,N_8103);
xor U11031 (N_11031,N_8414,N_8109);
and U11032 (N_11032,N_8679,N_9348);
or U11033 (N_11033,N_8982,N_8620);
xnor U11034 (N_11034,N_8867,N_8691);
or U11035 (N_11035,N_9230,N_9323);
nor U11036 (N_11036,N_9525,N_9129);
nand U11037 (N_11037,N_9403,N_9137);
nand U11038 (N_11038,N_9426,N_9956);
nor U11039 (N_11039,N_9683,N_8427);
or U11040 (N_11040,N_8420,N_9490);
xor U11041 (N_11041,N_9280,N_8445);
and U11042 (N_11042,N_8333,N_9805);
nand U11043 (N_11043,N_8614,N_8190);
xnor U11044 (N_11044,N_9544,N_8214);
nand U11045 (N_11045,N_9336,N_8950);
or U11046 (N_11046,N_9664,N_9747);
and U11047 (N_11047,N_8441,N_8448);
or U11048 (N_11048,N_9068,N_9050);
xor U11049 (N_11049,N_9732,N_8840);
xnor U11050 (N_11050,N_8336,N_9715);
xnor U11051 (N_11051,N_8871,N_9392);
and U11052 (N_11052,N_8238,N_8936);
nand U11053 (N_11053,N_9717,N_9777);
nand U11054 (N_11054,N_9620,N_9563);
nand U11055 (N_11055,N_8322,N_8955);
nand U11056 (N_11056,N_8206,N_8253);
and U11057 (N_11057,N_8455,N_8571);
or U11058 (N_11058,N_9044,N_9199);
nor U11059 (N_11059,N_8002,N_9867);
nor U11060 (N_11060,N_9875,N_8350);
xnor U11061 (N_11061,N_8865,N_9002);
nor U11062 (N_11062,N_8692,N_8800);
or U11063 (N_11063,N_9760,N_9199);
nor U11064 (N_11064,N_9487,N_8438);
or U11065 (N_11065,N_9433,N_8341);
nand U11066 (N_11066,N_9186,N_9989);
and U11067 (N_11067,N_8521,N_8519);
or U11068 (N_11068,N_9754,N_9560);
nand U11069 (N_11069,N_8205,N_9353);
nor U11070 (N_11070,N_9324,N_8923);
nand U11071 (N_11071,N_9971,N_8601);
nand U11072 (N_11072,N_9222,N_8668);
and U11073 (N_11073,N_9190,N_8329);
xnor U11074 (N_11074,N_8534,N_9276);
nand U11075 (N_11075,N_9625,N_9065);
xor U11076 (N_11076,N_9571,N_8043);
and U11077 (N_11077,N_8140,N_9502);
or U11078 (N_11078,N_9698,N_8923);
or U11079 (N_11079,N_8366,N_8531);
or U11080 (N_11080,N_9796,N_8347);
xnor U11081 (N_11081,N_8183,N_9975);
or U11082 (N_11082,N_8294,N_9536);
and U11083 (N_11083,N_9079,N_9252);
and U11084 (N_11084,N_9528,N_9110);
nor U11085 (N_11085,N_9770,N_9079);
nor U11086 (N_11086,N_8420,N_8223);
nand U11087 (N_11087,N_9193,N_9303);
nand U11088 (N_11088,N_8803,N_9647);
and U11089 (N_11089,N_9404,N_9858);
xor U11090 (N_11090,N_9387,N_8264);
nand U11091 (N_11091,N_8857,N_8443);
and U11092 (N_11092,N_9010,N_9102);
or U11093 (N_11093,N_8111,N_9104);
nor U11094 (N_11094,N_8011,N_9366);
and U11095 (N_11095,N_8586,N_8708);
nand U11096 (N_11096,N_9433,N_9159);
xor U11097 (N_11097,N_8761,N_8549);
xnor U11098 (N_11098,N_8976,N_9868);
or U11099 (N_11099,N_9478,N_9775);
nand U11100 (N_11100,N_9354,N_8383);
nand U11101 (N_11101,N_8586,N_8748);
and U11102 (N_11102,N_8201,N_8921);
or U11103 (N_11103,N_9961,N_9273);
or U11104 (N_11104,N_9091,N_9789);
nand U11105 (N_11105,N_8202,N_9738);
and U11106 (N_11106,N_8080,N_9510);
or U11107 (N_11107,N_9392,N_8534);
nor U11108 (N_11108,N_8696,N_9178);
nor U11109 (N_11109,N_8657,N_8415);
or U11110 (N_11110,N_9968,N_8701);
nor U11111 (N_11111,N_8655,N_9535);
or U11112 (N_11112,N_9156,N_9487);
and U11113 (N_11113,N_8148,N_8243);
nand U11114 (N_11114,N_8024,N_9494);
or U11115 (N_11115,N_8822,N_8587);
nand U11116 (N_11116,N_8670,N_9450);
nand U11117 (N_11117,N_9342,N_9535);
or U11118 (N_11118,N_9840,N_9193);
nor U11119 (N_11119,N_9724,N_9405);
xor U11120 (N_11120,N_9346,N_9777);
and U11121 (N_11121,N_9636,N_9425);
xnor U11122 (N_11122,N_8759,N_8753);
xor U11123 (N_11123,N_8020,N_9825);
and U11124 (N_11124,N_8803,N_8400);
or U11125 (N_11125,N_8045,N_8588);
nand U11126 (N_11126,N_8885,N_8671);
xnor U11127 (N_11127,N_8083,N_8748);
nor U11128 (N_11128,N_9164,N_8227);
xnor U11129 (N_11129,N_8763,N_9509);
or U11130 (N_11130,N_9030,N_9527);
xnor U11131 (N_11131,N_9657,N_9011);
and U11132 (N_11132,N_9231,N_9779);
and U11133 (N_11133,N_9000,N_9421);
or U11134 (N_11134,N_8886,N_8106);
nor U11135 (N_11135,N_9590,N_8335);
and U11136 (N_11136,N_9857,N_9971);
nor U11137 (N_11137,N_9430,N_8507);
or U11138 (N_11138,N_9057,N_9564);
nand U11139 (N_11139,N_9281,N_8385);
xor U11140 (N_11140,N_8279,N_8817);
nor U11141 (N_11141,N_8153,N_8981);
and U11142 (N_11142,N_8945,N_8356);
and U11143 (N_11143,N_9004,N_8760);
xnor U11144 (N_11144,N_8617,N_9312);
or U11145 (N_11145,N_9031,N_8274);
nand U11146 (N_11146,N_8368,N_9150);
nor U11147 (N_11147,N_8731,N_9437);
nand U11148 (N_11148,N_8352,N_9403);
nor U11149 (N_11149,N_9612,N_8567);
nand U11150 (N_11150,N_9182,N_8419);
nor U11151 (N_11151,N_9488,N_9907);
nand U11152 (N_11152,N_8371,N_8429);
nor U11153 (N_11153,N_8883,N_9713);
nor U11154 (N_11154,N_9204,N_8730);
xnor U11155 (N_11155,N_9423,N_9245);
nand U11156 (N_11156,N_9297,N_8074);
nor U11157 (N_11157,N_9946,N_8929);
and U11158 (N_11158,N_9525,N_8315);
or U11159 (N_11159,N_8613,N_8957);
xor U11160 (N_11160,N_9440,N_9241);
or U11161 (N_11161,N_8572,N_9479);
nor U11162 (N_11162,N_9675,N_8952);
and U11163 (N_11163,N_9870,N_9535);
nor U11164 (N_11164,N_9916,N_9561);
xor U11165 (N_11165,N_9545,N_8441);
nor U11166 (N_11166,N_8362,N_9146);
nand U11167 (N_11167,N_9760,N_8641);
nand U11168 (N_11168,N_9211,N_8754);
or U11169 (N_11169,N_8267,N_9557);
nand U11170 (N_11170,N_8481,N_9282);
nor U11171 (N_11171,N_9091,N_9208);
and U11172 (N_11172,N_9985,N_9831);
xnor U11173 (N_11173,N_9717,N_9162);
and U11174 (N_11174,N_9185,N_9986);
nor U11175 (N_11175,N_8976,N_8971);
nor U11176 (N_11176,N_9002,N_8094);
xor U11177 (N_11177,N_9646,N_8485);
or U11178 (N_11178,N_8505,N_9124);
nand U11179 (N_11179,N_9186,N_8644);
and U11180 (N_11180,N_9461,N_8357);
nor U11181 (N_11181,N_9048,N_9384);
nor U11182 (N_11182,N_8557,N_8967);
or U11183 (N_11183,N_8502,N_9000);
nor U11184 (N_11184,N_8388,N_9484);
nor U11185 (N_11185,N_9917,N_9996);
or U11186 (N_11186,N_8767,N_9541);
and U11187 (N_11187,N_8222,N_8469);
nand U11188 (N_11188,N_9241,N_8765);
xor U11189 (N_11189,N_9601,N_9674);
nand U11190 (N_11190,N_9583,N_9856);
and U11191 (N_11191,N_8387,N_8935);
nor U11192 (N_11192,N_8068,N_8291);
nor U11193 (N_11193,N_9305,N_9273);
xnor U11194 (N_11194,N_8139,N_9208);
xor U11195 (N_11195,N_8560,N_8688);
nand U11196 (N_11196,N_9634,N_9421);
nand U11197 (N_11197,N_8350,N_9315);
and U11198 (N_11198,N_8105,N_9098);
nand U11199 (N_11199,N_8692,N_8391);
or U11200 (N_11200,N_8974,N_9499);
xnor U11201 (N_11201,N_9881,N_8250);
or U11202 (N_11202,N_8955,N_9080);
xnor U11203 (N_11203,N_8562,N_9364);
and U11204 (N_11204,N_8459,N_8362);
nand U11205 (N_11205,N_9951,N_8464);
nand U11206 (N_11206,N_8567,N_8038);
or U11207 (N_11207,N_9598,N_9200);
or U11208 (N_11208,N_8771,N_9837);
xnor U11209 (N_11209,N_8796,N_9071);
nor U11210 (N_11210,N_9768,N_8707);
xnor U11211 (N_11211,N_9646,N_8638);
nor U11212 (N_11212,N_9953,N_8138);
nand U11213 (N_11213,N_9603,N_9580);
nand U11214 (N_11214,N_9337,N_9712);
nand U11215 (N_11215,N_9330,N_9103);
nand U11216 (N_11216,N_8901,N_9712);
or U11217 (N_11217,N_9153,N_8128);
and U11218 (N_11218,N_9571,N_8287);
xor U11219 (N_11219,N_9956,N_9319);
xnor U11220 (N_11220,N_8395,N_8825);
or U11221 (N_11221,N_9720,N_8587);
or U11222 (N_11222,N_8895,N_8471);
nand U11223 (N_11223,N_9161,N_9301);
nand U11224 (N_11224,N_8969,N_8931);
nor U11225 (N_11225,N_8991,N_9295);
nor U11226 (N_11226,N_8279,N_9621);
nand U11227 (N_11227,N_8058,N_8728);
xor U11228 (N_11228,N_9430,N_8786);
nor U11229 (N_11229,N_9594,N_8433);
nand U11230 (N_11230,N_9610,N_9856);
xnor U11231 (N_11231,N_9148,N_9155);
and U11232 (N_11232,N_8232,N_9667);
or U11233 (N_11233,N_8055,N_9013);
or U11234 (N_11234,N_9069,N_8888);
and U11235 (N_11235,N_8102,N_8729);
nand U11236 (N_11236,N_9072,N_8268);
or U11237 (N_11237,N_8341,N_8413);
or U11238 (N_11238,N_8721,N_9329);
nor U11239 (N_11239,N_8951,N_8721);
xor U11240 (N_11240,N_9612,N_9658);
and U11241 (N_11241,N_8556,N_8974);
or U11242 (N_11242,N_8891,N_9403);
nor U11243 (N_11243,N_9424,N_8631);
nor U11244 (N_11244,N_8773,N_9258);
and U11245 (N_11245,N_9220,N_9688);
or U11246 (N_11246,N_9778,N_9238);
nor U11247 (N_11247,N_8221,N_8862);
nand U11248 (N_11248,N_9301,N_9998);
nor U11249 (N_11249,N_9259,N_9058);
xor U11250 (N_11250,N_9273,N_9208);
and U11251 (N_11251,N_9015,N_9709);
xnor U11252 (N_11252,N_9893,N_8810);
nor U11253 (N_11253,N_8332,N_9911);
nand U11254 (N_11254,N_9671,N_8231);
or U11255 (N_11255,N_9392,N_9922);
nand U11256 (N_11256,N_8417,N_9347);
and U11257 (N_11257,N_8525,N_9148);
and U11258 (N_11258,N_9649,N_8635);
and U11259 (N_11259,N_9549,N_9938);
nor U11260 (N_11260,N_8710,N_9231);
nor U11261 (N_11261,N_9592,N_9867);
xnor U11262 (N_11262,N_8416,N_9434);
or U11263 (N_11263,N_9179,N_9191);
nand U11264 (N_11264,N_8419,N_9085);
or U11265 (N_11265,N_8985,N_8393);
and U11266 (N_11266,N_8152,N_8510);
nand U11267 (N_11267,N_9902,N_9900);
or U11268 (N_11268,N_8915,N_9050);
and U11269 (N_11269,N_8704,N_8245);
and U11270 (N_11270,N_9545,N_9482);
and U11271 (N_11271,N_8194,N_8365);
and U11272 (N_11272,N_8143,N_9771);
nor U11273 (N_11273,N_9671,N_9693);
xor U11274 (N_11274,N_9552,N_8950);
or U11275 (N_11275,N_9007,N_8097);
and U11276 (N_11276,N_9468,N_9510);
xnor U11277 (N_11277,N_8385,N_8162);
nand U11278 (N_11278,N_8369,N_8968);
or U11279 (N_11279,N_9654,N_9515);
xor U11280 (N_11280,N_8143,N_9143);
nand U11281 (N_11281,N_8188,N_9770);
xnor U11282 (N_11282,N_9525,N_8204);
xor U11283 (N_11283,N_8486,N_9952);
or U11284 (N_11284,N_9420,N_9101);
nor U11285 (N_11285,N_8645,N_9052);
and U11286 (N_11286,N_9883,N_8028);
or U11287 (N_11287,N_9846,N_8502);
or U11288 (N_11288,N_8499,N_9289);
and U11289 (N_11289,N_8057,N_9140);
xnor U11290 (N_11290,N_9013,N_9456);
xnor U11291 (N_11291,N_8277,N_9362);
nand U11292 (N_11292,N_9535,N_9586);
nor U11293 (N_11293,N_8709,N_8789);
nor U11294 (N_11294,N_9751,N_8930);
nor U11295 (N_11295,N_9697,N_8409);
nand U11296 (N_11296,N_9751,N_9282);
or U11297 (N_11297,N_8235,N_8033);
and U11298 (N_11298,N_8613,N_8831);
or U11299 (N_11299,N_9837,N_9571);
nor U11300 (N_11300,N_8651,N_9313);
xnor U11301 (N_11301,N_9528,N_8180);
nand U11302 (N_11302,N_9317,N_8762);
xnor U11303 (N_11303,N_8107,N_8795);
xor U11304 (N_11304,N_9518,N_8815);
and U11305 (N_11305,N_9611,N_8251);
nand U11306 (N_11306,N_8558,N_9566);
or U11307 (N_11307,N_8503,N_8937);
nor U11308 (N_11308,N_8684,N_8952);
nand U11309 (N_11309,N_9858,N_9278);
or U11310 (N_11310,N_8938,N_9647);
xor U11311 (N_11311,N_9441,N_8042);
xnor U11312 (N_11312,N_9449,N_9899);
or U11313 (N_11313,N_9455,N_8120);
nand U11314 (N_11314,N_9139,N_9517);
or U11315 (N_11315,N_9675,N_9322);
and U11316 (N_11316,N_8531,N_8105);
and U11317 (N_11317,N_8066,N_8275);
nor U11318 (N_11318,N_8926,N_9345);
and U11319 (N_11319,N_9207,N_9965);
xnor U11320 (N_11320,N_9274,N_8447);
xor U11321 (N_11321,N_8306,N_8811);
nor U11322 (N_11322,N_9331,N_8811);
nand U11323 (N_11323,N_8343,N_8924);
or U11324 (N_11324,N_8546,N_8958);
and U11325 (N_11325,N_8114,N_9308);
nor U11326 (N_11326,N_9769,N_8045);
xnor U11327 (N_11327,N_9528,N_8361);
and U11328 (N_11328,N_8212,N_8787);
or U11329 (N_11329,N_9417,N_8275);
nor U11330 (N_11330,N_9904,N_8726);
nor U11331 (N_11331,N_8527,N_9007);
nor U11332 (N_11332,N_9174,N_9339);
nand U11333 (N_11333,N_9698,N_9449);
and U11334 (N_11334,N_9288,N_9577);
or U11335 (N_11335,N_8817,N_8386);
nand U11336 (N_11336,N_8563,N_9097);
and U11337 (N_11337,N_9750,N_8627);
and U11338 (N_11338,N_9445,N_8492);
or U11339 (N_11339,N_8838,N_8543);
nor U11340 (N_11340,N_8084,N_9913);
xnor U11341 (N_11341,N_9427,N_8715);
and U11342 (N_11342,N_8339,N_9512);
and U11343 (N_11343,N_9741,N_9987);
xnor U11344 (N_11344,N_8147,N_8226);
nor U11345 (N_11345,N_9173,N_8638);
nor U11346 (N_11346,N_8430,N_8804);
or U11347 (N_11347,N_9865,N_8217);
and U11348 (N_11348,N_8575,N_9498);
nand U11349 (N_11349,N_8126,N_9459);
xnor U11350 (N_11350,N_9110,N_9052);
xor U11351 (N_11351,N_9871,N_9578);
xnor U11352 (N_11352,N_8717,N_9425);
and U11353 (N_11353,N_9332,N_9494);
nor U11354 (N_11354,N_8836,N_8418);
and U11355 (N_11355,N_9710,N_8770);
or U11356 (N_11356,N_8894,N_8462);
xor U11357 (N_11357,N_9334,N_9597);
nand U11358 (N_11358,N_8492,N_9720);
or U11359 (N_11359,N_8408,N_9394);
nand U11360 (N_11360,N_9790,N_9285);
or U11361 (N_11361,N_8403,N_9276);
nand U11362 (N_11362,N_9093,N_9813);
or U11363 (N_11363,N_9722,N_9516);
and U11364 (N_11364,N_9669,N_9552);
or U11365 (N_11365,N_9935,N_8701);
nand U11366 (N_11366,N_8566,N_9184);
and U11367 (N_11367,N_9490,N_9398);
xnor U11368 (N_11368,N_8092,N_8330);
xnor U11369 (N_11369,N_9112,N_9828);
and U11370 (N_11370,N_8010,N_9538);
and U11371 (N_11371,N_8409,N_8289);
or U11372 (N_11372,N_9960,N_9399);
xor U11373 (N_11373,N_8507,N_9885);
xnor U11374 (N_11374,N_8140,N_8136);
and U11375 (N_11375,N_9165,N_9820);
or U11376 (N_11376,N_9736,N_8774);
nand U11377 (N_11377,N_8642,N_8029);
nand U11378 (N_11378,N_8213,N_9632);
and U11379 (N_11379,N_9079,N_9546);
and U11380 (N_11380,N_8870,N_9162);
and U11381 (N_11381,N_9505,N_9203);
and U11382 (N_11382,N_8118,N_8181);
xor U11383 (N_11383,N_8256,N_8224);
and U11384 (N_11384,N_9227,N_8571);
nand U11385 (N_11385,N_9373,N_9423);
or U11386 (N_11386,N_8178,N_9385);
nand U11387 (N_11387,N_9639,N_9969);
and U11388 (N_11388,N_9331,N_9080);
or U11389 (N_11389,N_9875,N_9979);
nand U11390 (N_11390,N_8044,N_9269);
nor U11391 (N_11391,N_9748,N_9935);
and U11392 (N_11392,N_9534,N_9808);
or U11393 (N_11393,N_9098,N_8370);
nor U11394 (N_11394,N_8151,N_9693);
or U11395 (N_11395,N_9093,N_9213);
nand U11396 (N_11396,N_8430,N_8940);
nand U11397 (N_11397,N_8742,N_8643);
and U11398 (N_11398,N_9490,N_9654);
and U11399 (N_11399,N_8864,N_9229);
and U11400 (N_11400,N_9118,N_8231);
or U11401 (N_11401,N_8934,N_8244);
nand U11402 (N_11402,N_8696,N_8857);
nand U11403 (N_11403,N_8712,N_8713);
nand U11404 (N_11404,N_8342,N_8509);
xnor U11405 (N_11405,N_9426,N_8435);
nand U11406 (N_11406,N_9189,N_9539);
nand U11407 (N_11407,N_9025,N_8485);
nor U11408 (N_11408,N_8443,N_8525);
or U11409 (N_11409,N_8005,N_9078);
nand U11410 (N_11410,N_8606,N_8252);
and U11411 (N_11411,N_9441,N_8977);
xnor U11412 (N_11412,N_9931,N_9992);
or U11413 (N_11413,N_9236,N_8643);
nand U11414 (N_11414,N_9326,N_8743);
or U11415 (N_11415,N_8925,N_9648);
and U11416 (N_11416,N_8062,N_9564);
and U11417 (N_11417,N_9217,N_8532);
nor U11418 (N_11418,N_9531,N_9218);
or U11419 (N_11419,N_8325,N_9726);
nand U11420 (N_11420,N_9711,N_8038);
nor U11421 (N_11421,N_9541,N_8839);
or U11422 (N_11422,N_9856,N_9558);
and U11423 (N_11423,N_8088,N_9009);
nand U11424 (N_11424,N_9953,N_8351);
nand U11425 (N_11425,N_9027,N_8225);
and U11426 (N_11426,N_8701,N_9809);
and U11427 (N_11427,N_8806,N_9403);
and U11428 (N_11428,N_8411,N_9379);
or U11429 (N_11429,N_9946,N_9303);
xor U11430 (N_11430,N_8061,N_9144);
nor U11431 (N_11431,N_8360,N_9532);
xor U11432 (N_11432,N_9973,N_8180);
nand U11433 (N_11433,N_8169,N_8841);
nor U11434 (N_11434,N_8400,N_9742);
nor U11435 (N_11435,N_8521,N_9809);
nand U11436 (N_11436,N_8368,N_8656);
nand U11437 (N_11437,N_8388,N_8947);
xor U11438 (N_11438,N_8541,N_8759);
nor U11439 (N_11439,N_8257,N_8433);
or U11440 (N_11440,N_9158,N_8793);
and U11441 (N_11441,N_8524,N_8616);
xor U11442 (N_11442,N_9085,N_9079);
xor U11443 (N_11443,N_8000,N_9243);
nand U11444 (N_11444,N_8776,N_8432);
nor U11445 (N_11445,N_8915,N_9762);
or U11446 (N_11446,N_8001,N_9620);
nand U11447 (N_11447,N_9019,N_9471);
and U11448 (N_11448,N_9598,N_9279);
or U11449 (N_11449,N_8722,N_9061);
nor U11450 (N_11450,N_9111,N_8594);
nor U11451 (N_11451,N_9688,N_9516);
nand U11452 (N_11452,N_8692,N_8617);
or U11453 (N_11453,N_8929,N_9297);
or U11454 (N_11454,N_8433,N_9743);
xor U11455 (N_11455,N_8814,N_9665);
xor U11456 (N_11456,N_8510,N_8706);
or U11457 (N_11457,N_8001,N_8186);
xnor U11458 (N_11458,N_9491,N_8072);
nand U11459 (N_11459,N_8158,N_8038);
nor U11460 (N_11460,N_8736,N_8159);
nand U11461 (N_11461,N_8218,N_8049);
and U11462 (N_11462,N_9188,N_8020);
and U11463 (N_11463,N_8242,N_9487);
or U11464 (N_11464,N_8028,N_9930);
and U11465 (N_11465,N_8862,N_8276);
and U11466 (N_11466,N_8261,N_9845);
nor U11467 (N_11467,N_9363,N_9549);
nand U11468 (N_11468,N_8476,N_8367);
nand U11469 (N_11469,N_8528,N_8220);
xor U11470 (N_11470,N_9647,N_8535);
xor U11471 (N_11471,N_8968,N_8254);
xnor U11472 (N_11472,N_9842,N_9522);
xor U11473 (N_11473,N_9319,N_9499);
or U11474 (N_11474,N_9855,N_9688);
nor U11475 (N_11475,N_8096,N_8516);
and U11476 (N_11476,N_8411,N_8566);
xnor U11477 (N_11477,N_9990,N_8491);
nand U11478 (N_11478,N_9900,N_8320);
nor U11479 (N_11479,N_9715,N_9164);
and U11480 (N_11480,N_9032,N_8823);
nor U11481 (N_11481,N_9970,N_9418);
or U11482 (N_11482,N_8960,N_9173);
nand U11483 (N_11483,N_9658,N_9986);
nand U11484 (N_11484,N_8164,N_8586);
or U11485 (N_11485,N_8718,N_8157);
nor U11486 (N_11486,N_8941,N_8218);
xor U11487 (N_11487,N_8623,N_8924);
xnor U11488 (N_11488,N_8318,N_8077);
xnor U11489 (N_11489,N_8075,N_8510);
or U11490 (N_11490,N_9082,N_9706);
or U11491 (N_11491,N_9330,N_9328);
nor U11492 (N_11492,N_9879,N_8442);
or U11493 (N_11493,N_9430,N_8076);
nand U11494 (N_11494,N_8257,N_9885);
nand U11495 (N_11495,N_8906,N_9790);
and U11496 (N_11496,N_9870,N_9717);
and U11497 (N_11497,N_8181,N_8415);
nand U11498 (N_11498,N_9129,N_9483);
and U11499 (N_11499,N_8920,N_8541);
nor U11500 (N_11500,N_9798,N_8801);
nor U11501 (N_11501,N_9644,N_8576);
or U11502 (N_11502,N_9188,N_8967);
or U11503 (N_11503,N_8775,N_9536);
xor U11504 (N_11504,N_9797,N_9922);
xnor U11505 (N_11505,N_9862,N_9623);
xnor U11506 (N_11506,N_8893,N_8933);
nor U11507 (N_11507,N_8585,N_8776);
and U11508 (N_11508,N_8086,N_9953);
and U11509 (N_11509,N_9559,N_8830);
nand U11510 (N_11510,N_9409,N_9596);
nand U11511 (N_11511,N_8172,N_9638);
xor U11512 (N_11512,N_9312,N_9540);
nor U11513 (N_11513,N_8534,N_8112);
nor U11514 (N_11514,N_8671,N_8938);
or U11515 (N_11515,N_8537,N_9949);
xor U11516 (N_11516,N_9870,N_8574);
nor U11517 (N_11517,N_9370,N_8522);
xnor U11518 (N_11518,N_9660,N_8487);
nand U11519 (N_11519,N_9931,N_9892);
and U11520 (N_11520,N_9991,N_9774);
or U11521 (N_11521,N_8868,N_8556);
nand U11522 (N_11522,N_9542,N_8677);
xor U11523 (N_11523,N_9988,N_9922);
or U11524 (N_11524,N_9886,N_8770);
nand U11525 (N_11525,N_9535,N_8414);
xnor U11526 (N_11526,N_8302,N_9162);
or U11527 (N_11527,N_8989,N_8245);
and U11528 (N_11528,N_9478,N_8954);
xnor U11529 (N_11529,N_8487,N_8387);
nand U11530 (N_11530,N_9948,N_9793);
and U11531 (N_11531,N_8671,N_8633);
xor U11532 (N_11532,N_9233,N_8929);
nand U11533 (N_11533,N_9138,N_9529);
nand U11534 (N_11534,N_9751,N_9394);
or U11535 (N_11535,N_8808,N_9767);
nand U11536 (N_11536,N_8474,N_8608);
xnor U11537 (N_11537,N_8739,N_9296);
xnor U11538 (N_11538,N_8127,N_8792);
nor U11539 (N_11539,N_9876,N_9893);
or U11540 (N_11540,N_9445,N_8767);
nor U11541 (N_11541,N_8338,N_8884);
nor U11542 (N_11542,N_9222,N_9117);
or U11543 (N_11543,N_8644,N_9285);
nand U11544 (N_11544,N_8328,N_9116);
nand U11545 (N_11545,N_9288,N_9346);
nand U11546 (N_11546,N_8929,N_8367);
or U11547 (N_11547,N_9471,N_8161);
nor U11548 (N_11548,N_9513,N_9326);
xor U11549 (N_11549,N_8207,N_8682);
or U11550 (N_11550,N_8790,N_8752);
or U11551 (N_11551,N_9961,N_8579);
xnor U11552 (N_11552,N_9170,N_9072);
xor U11553 (N_11553,N_8014,N_9628);
and U11554 (N_11554,N_9031,N_8429);
nand U11555 (N_11555,N_8830,N_8643);
nor U11556 (N_11556,N_8678,N_8479);
xnor U11557 (N_11557,N_8816,N_9486);
and U11558 (N_11558,N_8519,N_8477);
nor U11559 (N_11559,N_9467,N_8158);
and U11560 (N_11560,N_9851,N_8639);
or U11561 (N_11561,N_8101,N_8348);
xor U11562 (N_11562,N_8467,N_9640);
or U11563 (N_11563,N_8050,N_8841);
nand U11564 (N_11564,N_9539,N_9609);
xnor U11565 (N_11565,N_8783,N_8409);
nor U11566 (N_11566,N_8942,N_8647);
or U11567 (N_11567,N_8908,N_9920);
and U11568 (N_11568,N_9524,N_8634);
or U11569 (N_11569,N_8836,N_9922);
and U11570 (N_11570,N_8626,N_8906);
xor U11571 (N_11571,N_8026,N_8905);
xor U11572 (N_11572,N_8753,N_9847);
and U11573 (N_11573,N_8585,N_9376);
and U11574 (N_11574,N_9379,N_9081);
or U11575 (N_11575,N_9260,N_9447);
nand U11576 (N_11576,N_9067,N_9056);
nand U11577 (N_11577,N_9085,N_9071);
nand U11578 (N_11578,N_9427,N_9873);
and U11579 (N_11579,N_8127,N_8013);
and U11580 (N_11580,N_9470,N_9600);
nand U11581 (N_11581,N_9423,N_9100);
xnor U11582 (N_11582,N_8101,N_9869);
xor U11583 (N_11583,N_8801,N_8605);
nand U11584 (N_11584,N_9847,N_8879);
nor U11585 (N_11585,N_8060,N_9270);
and U11586 (N_11586,N_9326,N_8642);
and U11587 (N_11587,N_9943,N_9301);
nor U11588 (N_11588,N_9483,N_8489);
nor U11589 (N_11589,N_8515,N_8914);
nor U11590 (N_11590,N_8363,N_9618);
nor U11591 (N_11591,N_9093,N_8751);
nand U11592 (N_11592,N_9737,N_9550);
xnor U11593 (N_11593,N_8594,N_9109);
nor U11594 (N_11594,N_8487,N_8075);
nand U11595 (N_11595,N_8293,N_9539);
nand U11596 (N_11596,N_8017,N_9344);
nand U11597 (N_11597,N_9324,N_8585);
xnor U11598 (N_11598,N_9292,N_8868);
or U11599 (N_11599,N_9867,N_9337);
or U11600 (N_11600,N_9462,N_8318);
nand U11601 (N_11601,N_8920,N_9549);
nand U11602 (N_11602,N_9443,N_9055);
xor U11603 (N_11603,N_8390,N_9639);
nor U11604 (N_11604,N_9622,N_8810);
or U11605 (N_11605,N_8019,N_8693);
nand U11606 (N_11606,N_9416,N_8267);
and U11607 (N_11607,N_8763,N_9436);
nor U11608 (N_11608,N_9242,N_8383);
and U11609 (N_11609,N_8501,N_8331);
or U11610 (N_11610,N_9100,N_8946);
nand U11611 (N_11611,N_9188,N_8258);
nand U11612 (N_11612,N_9388,N_8437);
nand U11613 (N_11613,N_9902,N_9735);
xor U11614 (N_11614,N_8254,N_9102);
and U11615 (N_11615,N_9247,N_9251);
nand U11616 (N_11616,N_8833,N_9137);
nand U11617 (N_11617,N_9437,N_8268);
xnor U11618 (N_11618,N_9382,N_9894);
nor U11619 (N_11619,N_9294,N_9229);
or U11620 (N_11620,N_9474,N_8598);
nor U11621 (N_11621,N_9304,N_8178);
nor U11622 (N_11622,N_8060,N_8240);
nor U11623 (N_11623,N_9201,N_9834);
nor U11624 (N_11624,N_8400,N_9922);
or U11625 (N_11625,N_9292,N_8343);
nand U11626 (N_11626,N_9621,N_9225);
nor U11627 (N_11627,N_9603,N_9813);
and U11628 (N_11628,N_9962,N_9936);
xnor U11629 (N_11629,N_8503,N_8123);
nand U11630 (N_11630,N_8011,N_9655);
nor U11631 (N_11631,N_9526,N_8203);
and U11632 (N_11632,N_9757,N_8868);
xor U11633 (N_11633,N_9319,N_8403);
and U11634 (N_11634,N_8919,N_8456);
nor U11635 (N_11635,N_9973,N_8476);
and U11636 (N_11636,N_8794,N_8219);
or U11637 (N_11637,N_9758,N_9358);
nand U11638 (N_11638,N_9990,N_8481);
xnor U11639 (N_11639,N_8222,N_8519);
or U11640 (N_11640,N_8558,N_9075);
or U11641 (N_11641,N_9739,N_9922);
nand U11642 (N_11642,N_9907,N_8011);
nand U11643 (N_11643,N_9114,N_8271);
xor U11644 (N_11644,N_8097,N_9078);
or U11645 (N_11645,N_8708,N_9437);
xnor U11646 (N_11646,N_8676,N_9262);
xnor U11647 (N_11647,N_9535,N_8366);
or U11648 (N_11648,N_9228,N_8274);
nand U11649 (N_11649,N_9826,N_8890);
nand U11650 (N_11650,N_8090,N_9165);
xnor U11651 (N_11651,N_8123,N_8238);
nand U11652 (N_11652,N_8918,N_9466);
nor U11653 (N_11653,N_9236,N_8045);
nand U11654 (N_11654,N_8293,N_8013);
and U11655 (N_11655,N_8287,N_9054);
or U11656 (N_11656,N_8113,N_9425);
nand U11657 (N_11657,N_8089,N_8183);
nand U11658 (N_11658,N_8969,N_8463);
nor U11659 (N_11659,N_9960,N_8548);
xnor U11660 (N_11660,N_8769,N_9163);
and U11661 (N_11661,N_8686,N_8751);
nor U11662 (N_11662,N_9410,N_8870);
nand U11663 (N_11663,N_8547,N_9856);
xnor U11664 (N_11664,N_8639,N_9937);
nand U11665 (N_11665,N_8528,N_8487);
nor U11666 (N_11666,N_8039,N_8421);
nor U11667 (N_11667,N_9186,N_9923);
or U11668 (N_11668,N_8615,N_9339);
and U11669 (N_11669,N_8563,N_9065);
xnor U11670 (N_11670,N_8850,N_9177);
xor U11671 (N_11671,N_8912,N_9858);
xnor U11672 (N_11672,N_8059,N_9025);
and U11673 (N_11673,N_9829,N_8384);
xnor U11674 (N_11674,N_8780,N_8731);
nand U11675 (N_11675,N_9387,N_9839);
or U11676 (N_11676,N_8169,N_8237);
xor U11677 (N_11677,N_8840,N_8459);
nand U11678 (N_11678,N_8209,N_9924);
nor U11679 (N_11679,N_8718,N_8800);
and U11680 (N_11680,N_9695,N_9789);
nor U11681 (N_11681,N_8026,N_8675);
nand U11682 (N_11682,N_8178,N_9584);
nand U11683 (N_11683,N_9413,N_9062);
or U11684 (N_11684,N_9380,N_9718);
and U11685 (N_11685,N_9663,N_9490);
and U11686 (N_11686,N_9598,N_8406);
nand U11687 (N_11687,N_9944,N_8956);
nor U11688 (N_11688,N_8828,N_9207);
nor U11689 (N_11689,N_9794,N_9483);
nor U11690 (N_11690,N_9543,N_8061);
nor U11691 (N_11691,N_9903,N_9661);
or U11692 (N_11692,N_9207,N_8190);
nand U11693 (N_11693,N_9865,N_9891);
nand U11694 (N_11694,N_9288,N_9304);
or U11695 (N_11695,N_9716,N_9022);
nand U11696 (N_11696,N_8596,N_8626);
nand U11697 (N_11697,N_9844,N_8764);
or U11698 (N_11698,N_9119,N_8574);
and U11699 (N_11699,N_8952,N_9207);
or U11700 (N_11700,N_9130,N_8377);
nor U11701 (N_11701,N_8195,N_8679);
nor U11702 (N_11702,N_9729,N_8465);
xor U11703 (N_11703,N_8723,N_9057);
nand U11704 (N_11704,N_9776,N_9957);
or U11705 (N_11705,N_8960,N_8447);
nand U11706 (N_11706,N_9433,N_8402);
or U11707 (N_11707,N_9919,N_8174);
nand U11708 (N_11708,N_8524,N_9171);
nor U11709 (N_11709,N_9906,N_9478);
or U11710 (N_11710,N_9773,N_9815);
nor U11711 (N_11711,N_9688,N_9037);
xor U11712 (N_11712,N_8893,N_9860);
xor U11713 (N_11713,N_9184,N_9697);
xor U11714 (N_11714,N_9380,N_9101);
and U11715 (N_11715,N_9767,N_8229);
xnor U11716 (N_11716,N_9473,N_9786);
xnor U11717 (N_11717,N_9287,N_8801);
or U11718 (N_11718,N_9899,N_8189);
nor U11719 (N_11719,N_9152,N_8608);
or U11720 (N_11720,N_8345,N_8811);
or U11721 (N_11721,N_9118,N_8969);
and U11722 (N_11722,N_9723,N_9712);
xnor U11723 (N_11723,N_9867,N_8150);
nor U11724 (N_11724,N_9429,N_8968);
nor U11725 (N_11725,N_8309,N_8740);
and U11726 (N_11726,N_8059,N_9936);
nor U11727 (N_11727,N_9193,N_8308);
or U11728 (N_11728,N_8502,N_8372);
xor U11729 (N_11729,N_9392,N_9980);
xnor U11730 (N_11730,N_8716,N_9526);
xnor U11731 (N_11731,N_8251,N_8974);
or U11732 (N_11732,N_9188,N_8511);
nor U11733 (N_11733,N_8340,N_9028);
nand U11734 (N_11734,N_9813,N_9744);
nand U11735 (N_11735,N_8470,N_8821);
nor U11736 (N_11736,N_9135,N_8022);
and U11737 (N_11737,N_9430,N_8114);
nand U11738 (N_11738,N_8182,N_8988);
nand U11739 (N_11739,N_9311,N_8642);
nand U11740 (N_11740,N_8765,N_8147);
and U11741 (N_11741,N_8058,N_8800);
or U11742 (N_11742,N_9989,N_8058);
xor U11743 (N_11743,N_9924,N_9677);
nor U11744 (N_11744,N_8293,N_9735);
xnor U11745 (N_11745,N_8208,N_8981);
and U11746 (N_11746,N_8672,N_9198);
nand U11747 (N_11747,N_8986,N_9422);
and U11748 (N_11748,N_8707,N_9083);
or U11749 (N_11749,N_9929,N_8037);
or U11750 (N_11750,N_8802,N_8981);
xor U11751 (N_11751,N_9687,N_9519);
xor U11752 (N_11752,N_8097,N_9556);
nor U11753 (N_11753,N_9093,N_9160);
or U11754 (N_11754,N_8969,N_8921);
nor U11755 (N_11755,N_9708,N_9100);
or U11756 (N_11756,N_9580,N_9850);
and U11757 (N_11757,N_8525,N_9425);
xor U11758 (N_11758,N_9008,N_9140);
nor U11759 (N_11759,N_8634,N_8002);
nand U11760 (N_11760,N_9288,N_8084);
xnor U11761 (N_11761,N_9603,N_8774);
xor U11762 (N_11762,N_9782,N_8316);
and U11763 (N_11763,N_8006,N_8583);
and U11764 (N_11764,N_8067,N_9022);
xnor U11765 (N_11765,N_9604,N_8705);
or U11766 (N_11766,N_9216,N_9134);
nand U11767 (N_11767,N_9860,N_9120);
nand U11768 (N_11768,N_8109,N_8708);
and U11769 (N_11769,N_9597,N_9638);
xor U11770 (N_11770,N_9774,N_8550);
xnor U11771 (N_11771,N_8779,N_8631);
or U11772 (N_11772,N_9373,N_8112);
nor U11773 (N_11773,N_9010,N_8672);
nor U11774 (N_11774,N_9603,N_9688);
xor U11775 (N_11775,N_8059,N_9776);
xnor U11776 (N_11776,N_9223,N_8765);
xnor U11777 (N_11777,N_9060,N_9362);
xor U11778 (N_11778,N_8710,N_8837);
or U11779 (N_11779,N_8944,N_9823);
and U11780 (N_11780,N_9594,N_9240);
or U11781 (N_11781,N_8926,N_9468);
xnor U11782 (N_11782,N_8557,N_9303);
nor U11783 (N_11783,N_8241,N_9792);
xnor U11784 (N_11784,N_8123,N_8195);
and U11785 (N_11785,N_8532,N_8043);
xnor U11786 (N_11786,N_9708,N_8994);
or U11787 (N_11787,N_8510,N_9633);
and U11788 (N_11788,N_8980,N_9260);
xor U11789 (N_11789,N_8646,N_9700);
xor U11790 (N_11790,N_8285,N_9619);
nor U11791 (N_11791,N_9577,N_9170);
nor U11792 (N_11792,N_9829,N_9465);
xor U11793 (N_11793,N_9876,N_9905);
nor U11794 (N_11794,N_8859,N_9418);
nor U11795 (N_11795,N_9356,N_9615);
nor U11796 (N_11796,N_9255,N_8729);
nand U11797 (N_11797,N_9744,N_8323);
nor U11798 (N_11798,N_9172,N_8418);
nand U11799 (N_11799,N_8336,N_9416);
or U11800 (N_11800,N_8505,N_9506);
or U11801 (N_11801,N_9299,N_8176);
and U11802 (N_11802,N_9560,N_8246);
and U11803 (N_11803,N_8243,N_8713);
xnor U11804 (N_11804,N_9354,N_8986);
nor U11805 (N_11805,N_8949,N_9921);
or U11806 (N_11806,N_8433,N_9688);
nand U11807 (N_11807,N_9459,N_8296);
xor U11808 (N_11808,N_9845,N_8747);
nand U11809 (N_11809,N_8150,N_8192);
and U11810 (N_11810,N_9467,N_8577);
nor U11811 (N_11811,N_9552,N_8850);
xor U11812 (N_11812,N_9731,N_8247);
xnor U11813 (N_11813,N_9391,N_8812);
and U11814 (N_11814,N_8178,N_9665);
or U11815 (N_11815,N_8537,N_8741);
and U11816 (N_11816,N_8371,N_9330);
nor U11817 (N_11817,N_9457,N_9682);
xor U11818 (N_11818,N_9492,N_9933);
xnor U11819 (N_11819,N_9558,N_9119);
nand U11820 (N_11820,N_8760,N_9727);
nand U11821 (N_11821,N_8790,N_9099);
and U11822 (N_11822,N_8234,N_8921);
nand U11823 (N_11823,N_8984,N_9601);
nand U11824 (N_11824,N_8439,N_9143);
and U11825 (N_11825,N_8185,N_8397);
and U11826 (N_11826,N_9079,N_8493);
nand U11827 (N_11827,N_9870,N_9979);
xor U11828 (N_11828,N_9396,N_9792);
or U11829 (N_11829,N_8464,N_9555);
or U11830 (N_11830,N_8867,N_9860);
xor U11831 (N_11831,N_8333,N_9437);
xor U11832 (N_11832,N_9876,N_8165);
xor U11833 (N_11833,N_8171,N_8140);
nor U11834 (N_11834,N_8931,N_9604);
xnor U11835 (N_11835,N_8090,N_8526);
nor U11836 (N_11836,N_8262,N_9080);
and U11837 (N_11837,N_9722,N_9732);
or U11838 (N_11838,N_8451,N_8748);
nand U11839 (N_11839,N_8668,N_9724);
nand U11840 (N_11840,N_8878,N_9272);
or U11841 (N_11841,N_8278,N_9711);
nor U11842 (N_11842,N_9013,N_9417);
xor U11843 (N_11843,N_8666,N_9581);
nand U11844 (N_11844,N_9421,N_8441);
and U11845 (N_11845,N_8527,N_9782);
nor U11846 (N_11846,N_9845,N_8558);
or U11847 (N_11847,N_8901,N_8622);
nand U11848 (N_11848,N_9649,N_9036);
and U11849 (N_11849,N_8434,N_8999);
nor U11850 (N_11850,N_9414,N_8349);
or U11851 (N_11851,N_9479,N_9363);
xnor U11852 (N_11852,N_9864,N_9023);
or U11853 (N_11853,N_9007,N_8065);
xnor U11854 (N_11854,N_8694,N_9283);
nand U11855 (N_11855,N_8996,N_9990);
and U11856 (N_11856,N_8144,N_9742);
xnor U11857 (N_11857,N_8637,N_8349);
nor U11858 (N_11858,N_8892,N_8831);
xor U11859 (N_11859,N_8441,N_9073);
xor U11860 (N_11860,N_9714,N_8534);
or U11861 (N_11861,N_9397,N_8333);
and U11862 (N_11862,N_8142,N_9324);
nand U11863 (N_11863,N_8088,N_8590);
nor U11864 (N_11864,N_8360,N_9318);
nand U11865 (N_11865,N_8423,N_9767);
nor U11866 (N_11866,N_8473,N_9627);
or U11867 (N_11867,N_9816,N_8847);
nor U11868 (N_11868,N_9113,N_9618);
nor U11869 (N_11869,N_8981,N_9145);
nand U11870 (N_11870,N_8287,N_9471);
nand U11871 (N_11871,N_9600,N_8047);
and U11872 (N_11872,N_8505,N_9790);
or U11873 (N_11873,N_8796,N_8656);
nand U11874 (N_11874,N_8340,N_9161);
nor U11875 (N_11875,N_9382,N_8185);
and U11876 (N_11876,N_9044,N_9272);
nand U11877 (N_11877,N_8194,N_8809);
and U11878 (N_11878,N_8993,N_8289);
nand U11879 (N_11879,N_8238,N_8280);
and U11880 (N_11880,N_8273,N_8665);
or U11881 (N_11881,N_9933,N_9920);
and U11882 (N_11882,N_9368,N_9870);
xor U11883 (N_11883,N_8808,N_9159);
nor U11884 (N_11884,N_8889,N_9029);
or U11885 (N_11885,N_9288,N_8538);
nand U11886 (N_11886,N_9707,N_9009);
and U11887 (N_11887,N_9788,N_9412);
nor U11888 (N_11888,N_9800,N_9147);
nor U11889 (N_11889,N_8297,N_9329);
and U11890 (N_11890,N_8416,N_8183);
or U11891 (N_11891,N_9018,N_8459);
xnor U11892 (N_11892,N_9232,N_8591);
and U11893 (N_11893,N_8810,N_8989);
and U11894 (N_11894,N_8457,N_8149);
nand U11895 (N_11895,N_9944,N_8252);
and U11896 (N_11896,N_9123,N_8100);
nand U11897 (N_11897,N_9720,N_9573);
and U11898 (N_11898,N_9371,N_9171);
nand U11899 (N_11899,N_9363,N_9087);
and U11900 (N_11900,N_8640,N_9604);
xnor U11901 (N_11901,N_8648,N_8280);
or U11902 (N_11902,N_9192,N_8162);
xor U11903 (N_11903,N_8549,N_8831);
or U11904 (N_11904,N_8189,N_8772);
and U11905 (N_11905,N_9596,N_8111);
or U11906 (N_11906,N_9403,N_8494);
xnor U11907 (N_11907,N_9276,N_9279);
xnor U11908 (N_11908,N_9827,N_8267);
xor U11909 (N_11909,N_8821,N_9114);
nor U11910 (N_11910,N_8411,N_8974);
nand U11911 (N_11911,N_8510,N_8107);
or U11912 (N_11912,N_9763,N_9570);
or U11913 (N_11913,N_8629,N_9271);
nand U11914 (N_11914,N_8966,N_8249);
nand U11915 (N_11915,N_8884,N_8125);
and U11916 (N_11916,N_9931,N_8199);
xnor U11917 (N_11917,N_8032,N_9468);
nor U11918 (N_11918,N_9700,N_8355);
or U11919 (N_11919,N_9052,N_9299);
and U11920 (N_11920,N_8810,N_9233);
nor U11921 (N_11921,N_8541,N_8818);
xor U11922 (N_11922,N_9688,N_8598);
xnor U11923 (N_11923,N_9604,N_9575);
xnor U11924 (N_11924,N_9998,N_8463);
nor U11925 (N_11925,N_9341,N_9737);
or U11926 (N_11926,N_9459,N_9749);
xor U11927 (N_11927,N_9892,N_9504);
xor U11928 (N_11928,N_9904,N_9508);
xor U11929 (N_11929,N_9121,N_9688);
or U11930 (N_11930,N_9102,N_8685);
xor U11931 (N_11931,N_9354,N_9443);
xnor U11932 (N_11932,N_8724,N_9370);
and U11933 (N_11933,N_9024,N_8209);
xnor U11934 (N_11934,N_8164,N_9293);
and U11935 (N_11935,N_8650,N_8554);
nand U11936 (N_11936,N_9642,N_8803);
and U11937 (N_11937,N_9606,N_8192);
nor U11938 (N_11938,N_9098,N_8874);
or U11939 (N_11939,N_9283,N_9040);
nor U11940 (N_11940,N_8060,N_9536);
or U11941 (N_11941,N_9095,N_9993);
xnor U11942 (N_11942,N_9861,N_9006);
and U11943 (N_11943,N_9481,N_8702);
nand U11944 (N_11944,N_9105,N_8625);
and U11945 (N_11945,N_8403,N_9239);
and U11946 (N_11946,N_9798,N_9883);
and U11947 (N_11947,N_8915,N_8666);
and U11948 (N_11948,N_8746,N_8484);
nand U11949 (N_11949,N_8683,N_8657);
nor U11950 (N_11950,N_9780,N_8117);
and U11951 (N_11951,N_8044,N_9280);
xnor U11952 (N_11952,N_9638,N_9649);
nand U11953 (N_11953,N_8595,N_8131);
nand U11954 (N_11954,N_8624,N_8413);
or U11955 (N_11955,N_8738,N_8008);
nand U11956 (N_11956,N_9295,N_8807);
xnor U11957 (N_11957,N_9286,N_9440);
or U11958 (N_11958,N_8337,N_9069);
nand U11959 (N_11959,N_8924,N_8181);
nand U11960 (N_11960,N_9457,N_9310);
nor U11961 (N_11961,N_9959,N_8920);
nor U11962 (N_11962,N_8594,N_9178);
or U11963 (N_11963,N_8535,N_8008);
nand U11964 (N_11964,N_8361,N_9020);
nor U11965 (N_11965,N_9146,N_9420);
nand U11966 (N_11966,N_9682,N_9811);
and U11967 (N_11967,N_8600,N_9380);
nand U11968 (N_11968,N_9708,N_9187);
or U11969 (N_11969,N_8159,N_8876);
xnor U11970 (N_11970,N_9909,N_9509);
nand U11971 (N_11971,N_9007,N_8465);
nand U11972 (N_11972,N_8746,N_9429);
nand U11973 (N_11973,N_9905,N_8227);
nor U11974 (N_11974,N_8934,N_8505);
xor U11975 (N_11975,N_8169,N_8890);
nand U11976 (N_11976,N_8096,N_8573);
nand U11977 (N_11977,N_8653,N_8745);
or U11978 (N_11978,N_9279,N_8101);
or U11979 (N_11979,N_8711,N_8921);
or U11980 (N_11980,N_8406,N_8304);
and U11981 (N_11981,N_9351,N_9681);
nand U11982 (N_11982,N_8935,N_9264);
and U11983 (N_11983,N_9592,N_8797);
or U11984 (N_11984,N_8180,N_8148);
or U11985 (N_11985,N_8807,N_8179);
xnor U11986 (N_11986,N_8275,N_9817);
nor U11987 (N_11987,N_8547,N_9411);
xor U11988 (N_11988,N_8732,N_9517);
xor U11989 (N_11989,N_8415,N_9435);
or U11990 (N_11990,N_9053,N_8336);
nor U11991 (N_11991,N_9234,N_9574);
and U11992 (N_11992,N_8844,N_9099);
or U11993 (N_11993,N_8309,N_8088);
xor U11994 (N_11994,N_8867,N_9715);
and U11995 (N_11995,N_9739,N_8633);
or U11996 (N_11996,N_8617,N_9072);
xor U11997 (N_11997,N_9818,N_8159);
or U11998 (N_11998,N_8507,N_8570);
or U11999 (N_11999,N_8788,N_9668);
and U12000 (N_12000,N_11014,N_11092);
or U12001 (N_12001,N_11737,N_11394);
or U12002 (N_12002,N_11911,N_10586);
nand U12003 (N_12003,N_10004,N_11081);
and U12004 (N_12004,N_11691,N_11122);
nor U12005 (N_12005,N_10332,N_10320);
or U12006 (N_12006,N_10317,N_10327);
nor U12007 (N_12007,N_11304,N_11258);
nor U12008 (N_12008,N_11802,N_11758);
or U12009 (N_12009,N_10633,N_10905);
xnor U12010 (N_12010,N_11809,N_10909);
xor U12011 (N_12011,N_11896,N_10189);
nor U12012 (N_12012,N_11702,N_10597);
xnor U12013 (N_12013,N_11769,N_11409);
nor U12014 (N_12014,N_11217,N_10802);
nand U12015 (N_12015,N_11167,N_11635);
xor U12016 (N_12016,N_11271,N_10057);
and U12017 (N_12017,N_10995,N_10834);
xnor U12018 (N_12018,N_11999,N_11786);
and U12019 (N_12019,N_11124,N_10810);
nor U12020 (N_12020,N_10750,N_10977);
or U12021 (N_12021,N_10770,N_10484);
nor U12022 (N_12022,N_11406,N_10165);
xor U12023 (N_12023,N_10291,N_10140);
nor U12024 (N_12024,N_11593,N_11608);
nand U12025 (N_12025,N_10061,N_11178);
or U12026 (N_12026,N_11004,N_11823);
nand U12027 (N_12027,N_11865,N_10574);
nor U12028 (N_12028,N_11622,N_10869);
nor U12029 (N_12029,N_10578,N_10263);
and U12030 (N_12030,N_10322,N_11936);
and U12031 (N_12031,N_10210,N_10573);
or U12032 (N_12032,N_10981,N_10715);
nand U12033 (N_12033,N_10756,N_11528);
nand U12034 (N_12034,N_10654,N_10224);
and U12035 (N_12035,N_10042,N_10379);
nand U12036 (N_12036,N_10174,N_10538);
nor U12037 (N_12037,N_11246,N_11041);
nor U12038 (N_12038,N_11472,N_10676);
nand U12039 (N_12039,N_10141,N_10817);
nand U12040 (N_12040,N_11760,N_11424);
nor U12041 (N_12041,N_10704,N_11642);
nor U12042 (N_12042,N_11662,N_10473);
nand U12043 (N_12043,N_10645,N_10562);
xnor U12044 (N_12044,N_10114,N_11425);
or U12045 (N_12045,N_10634,N_10130);
nor U12046 (N_12046,N_11940,N_11159);
xor U12047 (N_12047,N_10585,N_11334);
and U12048 (N_12048,N_11360,N_10326);
nand U12049 (N_12049,N_11188,N_11184);
xor U12050 (N_12050,N_10438,N_11356);
and U12051 (N_12051,N_10912,N_11413);
nor U12052 (N_12052,N_10465,N_10630);
xnor U12053 (N_12053,N_11020,N_11794);
or U12054 (N_12054,N_10010,N_10844);
and U12055 (N_12055,N_10423,N_11108);
or U12056 (N_12056,N_11981,N_11992);
nor U12057 (N_12057,N_11000,N_10591);
nor U12058 (N_12058,N_11066,N_11759);
nor U12059 (N_12059,N_11820,N_10413);
nand U12060 (N_12060,N_11187,N_10510);
nand U12061 (N_12061,N_11799,N_11433);
xor U12062 (N_12062,N_10662,N_11652);
nor U12063 (N_12063,N_11288,N_11135);
nand U12064 (N_12064,N_11777,N_11856);
xnor U12065 (N_12065,N_11620,N_10858);
or U12066 (N_12066,N_10713,N_10250);
nor U12067 (N_12067,N_10726,N_10493);
and U12068 (N_12068,N_10962,N_11416);
nand U12069 (N_12069,N_11491,N_10358);
nor U12070 (N_12070,N_10648,N_11382);
xor U12071 (N_12071,N_11971,N_11705);
and U12072 (N_12072,N_10580,N_11561);
or U12073 (N_12073,N_11723,N_11682);
or U12074 (N_12074,N_11945,N_11090);
and U12075 (N_12075,N_11895,N_10357);
nand U12076 (N_12076,N_11436,N_11350);
nor U12077 (N_12077,N_11630,N_11480);
xnor U12078 (N_12078,N_10786,N_11136);
nand U12079 (N_12079,N_10078,N_10093);
xor U12080 (N_12080,N_11263,N_10319);
nor U12081 (N_12081,N_10097,N_10699);
xor U12082 (N_12082,N_10897,N_11882);
nor U12083 (N_12083,N_10702,N_11358);
or U12084 (N_12084,N_10370,N_10103);
nor U12085 (N_12085,N_10246,N_11997);
nor U12086 (N_12086,N_10583,N_10553);
nand U12087 (N_12087,N_10677,N_10318);
or U12088 (N_12088,N_11907,N_10062);
xor U12089 (N_12089,N_11881,N_10352);
nand U12090 (N_12090,N_11496,N_10498);
and U12091 (N_12091,N_11452,N_11570);
nand U12092 (N_12092,N_11191,N_11072);
xnor U12093 (N_12093,N_10711,N_10231);
and U12094 (N_12094,N_10254,N_11193);
or U12095 (N_12095,N_11498,N_10641);
xor U12096 (N_12096,N_11114,N_10748);
and U12097 (N_12097,N_10839,N_11559);
and U12098 (N_12098,N_10712,N_10054);
xor U12099 (N_12099,N_11380,N_10164);
and U12100 (N_12100,N_11657,N_10549);
or U12101 (N_12101,N_10482,N_10669);
nand U12102 (N_12102,N_10674,N_10226);
or U12103 (N_12103,N_10282,N_11176);
xnor U12104 (N_12104,N_10667,N_11289);
and U12105 (N_12105,N_10403,N_11505);
and U12106 (N_12106,N_11840,N_10518);
and U12107 (N_12107,N_11242,N_11353);
or U12108 (N_12108,N_11422,N_10952);
xnor U12109 (N_12109,N_10592,N_11924);
nor U12110 (N_12110,N_11497,N_10273);
xnor U12111 (N_12111,N_10421,N_10094);
nand U12112 (N_12112,N_11901,N_11477);
xor U12113 (N_12113,N_11451,N_11859);
and U12114 (N_12114,N_11224,N_10168);
nor U12115 (N_12115,N_11339,N_10980);
or U12116 (N_12116,N_11698,N_11488);
xnor U12117 (N_12117,N_11716,N_10611);
or U12118 (N_12118,N_10735,N_10820);
and U12119 (N_12119,N_10038,N_10560);
or U12120 (N_12120,N_11316,N_11269);
nand U12121 (N_12121,N_11457,N_11509);
nor U12122 (N_12122,N_11419,N_10896);
or U12123 (N_12123,N_10460,N_10960);
and U12124 (N_12124,N_10074,N_10201);
nand U12125 (N_12125,N_11764,N_10229);
nor U12126 (N_12126,N_11367,N_11625);
or U12127 (N_12127,N_11085,N_11851);
nand U12128 (N_12128,N_11552,N_10171);
or U12129 (N_12129,N_11955,N_10668);
nor U12130 (N_12130,N_11717,N_11673);
and U12131 (N_12131,N_10664,N_10529);
nand U12132 (N_12132,N_11137,N_10339);
xor U12133 (N_12133,N_11321,N_10619);
or U12134 (N_12134,N_11916,N_10182);
or U12135 (N_12135,N_10218,N_11162);
or U12136 (N_12136,N_10800,N_10945);
nand U12137 (N_12137,N_10132,N_10060);
and U12138 (N_12138,N_11629,N_10657);
nand U12139 (N_12139,N_10405,N_10558);
and U12140 (N_12140,N_11686,N_11525);
and U12141 (N_12141,N_10887,N_10431);
nand U12142 (N_12142,N_10342,N_11152);
nand U12143 (N_12143,N_11910,N_10033);
nand U12144 (N_12144,N_10565,N_11349);
nor U12145 (N_12145,N_10581,N_11161);
or U12146 (N_12146,N_10507,N_10516);
or U12147 (N_12147,N_10148,N_11526);
or U12148 (N_12148,N_11780,N_10050);
or U12149 (N_12149,N_11318,N_10566);
nor U12150 (N_12150,N_11059,N_11954);
nand U12151 (N_12151,N_11824,N_10972);
nor U12152 (N_12152,N_11511,N_10416);
nand U12153 (N_12153,N_10515,N_10249);
xnor U12154 (N_12154,N_11689,N_10838);
nor U12155 (N_12155,N_11011,N_10749);
nor U12156 (N_12156,N_11942,N_10823);
and U12157 (N_12157,N_11833,N_10769);
xor U12158 (N_12158,N_10512,N_11886);
xor U12159 (N_12159,N_11984,N_10939);
nand U12160 (N_12160,N_10106,N_10391);
and U12161 (N_12161,N_10655,N_10197);
or U12162 (N_12162,N_11565,N_10175);
nor U12163 (N_12163,N_10979,N_10154);
and U12164 (N_12164,N_11903,N_11140);
nor U12165 (N_12165,N_11335,N_10483);
or U12166 (N_12166,N_10430,N_10771);
xnor U12167 (N_12167,N_11364,N_11993);
and U12168 (N_12168,N_10624,N_11157);
xor U12169 (N_12169,N_11079,N_10364);
nor U12170 (N_12170,N_11442,N_11766);
xor U12171 (N_12171,N_11839,N_10703);
nor U12172 (N_12172,N_10819,N_11355);
and U12173 (N_12173,N_10865,N_10190);
and U12174 (N_12174,N_10524,N_10765);
or U12175 (N_12175,N_11572,N_11266);
or U12176 (N_12176,N_10485,N_11342);
and U12177 (N_12177,N_10248,N_10888);
xnor U12178 (N_12178,N_11305,N_11329);
or U12179 (N_12179,N_11170,N_11675);
and U12180 (N_12180,N_11431,N_11236);
nor U12181 (N_12181,N_11607,N_10388);
nor U12182 (N_12182,N_11646,N_10324);
xor U12183 (N_12183,N_11478,N_11727);
nand U12184 (N_12184,N_11724,N_11423);
nor U12185 (N_12185,N_10118,N_10880);
nand U12186 (N_12186,N_11308,N_11659);
or U12187 (N_12187,N_11492,N_10564);
nor U12188 (N_12188,N_11384,N_11194);
nand U12189 (N_12189,N_11641,N_11273);
nand U12190 (N_12190,N_11848,N_10768);
nand U12191 (N_12191,N_10505,N_10588);
nor U12192 (N_12192,N_11206,N_10757);
or U12193 (N_12193,N_10395,N_10974);
nor U12194 (N_12194,N_11420,N_10292);
or U12195 (N_12195,N_11715,N_10862);
nand U12196 (N_12196,N_11805,N_10690);
and U12197 (N_12197,N_10293,N_10520);
xnor U12198 (N_12198,N_10763,N_10067);
nor U12199 (N_12199,N_11133,N_11665);
nor U12200 (N_12200,N_11791,N_11991);
and U12201 (N_12201,N_10257,N_11551);
xor U12202 (N_12202,N_10933,N_10990);
and U12203 (N_12203,N_11026,N_11567);
or U12204 (N_12204,N_11776,N_10700);
xor U12205 (N_12205,N_10812,N_10453);
nand U12206 (N_12206,N_11919,N_10491);
nor U12207 (N_12207,N_11482,N_11668);
nor U12208 (N_12208,N_11746,N_11393);
or U12209 (N_12209,N_10968,N_11199);
nor U12210 (N_12210,N_11411,N_11464);
nand U12211 (N_12211,N_11044,N_10283);
nor U12212 (N_12212,N_10816,N_11040);
and U12213 (N_12213,N_11510,N_11696);
or U12214 (N_12214,N_10546,N_11333);
or U12215 (N_12215,N_11885,N_10077);
xor U12216 (N_12216,N_10501,N_10940);
nand U12217 (N_12217,N_10809,N_10036);
xor U12218 (N_12218,N_11307,N_11216);
nand U12219 (N_12219,N_10041,N_11467);
and U12220 (N_12220,N_10692,N_11577);
nand U12221 (N_12221,N_10499,N_11214);
or U12222 (N_12222,N_11125,N_10371);
and U12223 (N_12223,N_11983,N_11580);
or U12224 (N_12224,N_11574,N_11616);
nor U12225 (N_12225,N_10088,N_10572);
nand U12226 (N_12226,N_10821,N_11893);
nor U12227 (N_12227,N_10031,N_11584);
xor U12228 (N_12228,N_10276,N_11755);
nand U12229 (N_12229,N_10665,N_11261);
xnor U12230 (N_12230,N_10607,N_10389);
nand U12231 (N_12231,N_10225,N_10958);
or U12232 (N_12232,N_10047,N_10742);
and U12233 (N_12233,N_11962,N_10778);
nand U12234 (N_12234,N_11390,N_10407);
xor U12235 (N_12235,N_11534,N_11256);
and U12236 (N_12236,N_11075,N_11970);
xor U12237 (N_12237,N_10044,N_11612);
nand U12238 (N_12238,N_10626,N_11487);
nor U12239 (N_12239,N_11190,N_10195);
nand U12240 (N_12240,N_10876,N_10999);
and U12241 (N_12241,N_10986,N_10497);
xnor U12242 (N_12242,N_10534,N_11775);
xnor U12243 (N_12243,N_11220,N_11280);
or U12244 (N_12244,N_11039,N_10543);
nor U12245 (N_12245,N_10904,N_11750);
nand U12246 (N_12246,N_10411,N_11648);
nand U12247 (N_12247,N_11605,N_10621);
or U12248 (N_12248,N_10256,N_11915);
xnor U12249 (N_12249,N_10916,N_10024);
xnor U12250 (N_12250,N_10341,N_11697);
nor U12251 (N_12251,N_11636,N_10347);
nor U12252 (N_12252,N_10784,N_11891);
xor U12253 (N_12253,N_11684,N_11198);
or U12254 (N_12254,N_11352,N_11798);
nor U12255 (N_12255,N_10212,N_10881);
nor U12256 (N_12256,N_10805,N_10794);
and U12257 (N_12257,N_10893,N_10432);
and U12258 (N_12258,N_10006,N_10177);
nand U12259 (N_12259,N_10731,N_10600);
nor U12260 (N_12260,N_11832,N_11508);
or U12261 (N_12261,N_10478,N_11331);
or U12262 (N_12262,N_10035,N_11005);
and U12263 (N_12263,N_11730,N_11623);
xnor U12264 (N_12264,N_10848,N_11468);
nor U12265 (N_12265,N_11441,N_10719);
or U12266 (N_12266,N_10943,N_10136);
nor U12267 (N_12267,N_11861,N_11676);
nand U12268 (N_12268,N_10598,N_10725);
and U12269 (N_12269,N_11948,N_11091);
and U12270 (N_12270,N_10123,N_11134);
and U12271 (N_12271,N_11330,N_10363);
nor U12272 (N_12272,N_10187,N_11815);
nor U12273 (N_12273,N_10685,N_10774);
nand U12274 (N_12274,N_11658,N_10511);
xnor U12275 (N_12275,N_10860,N_10545);
or U12276 (N_12276,N_10426,N_10059);
xor U12277 (N_12277,N_11530,N_11277);
or U12278 (N_12278,N_10808,N_10913);
nand U12279 (N_12279,N_10647,N_11247);
xnor U12280 (N_12280,N_10950,N_11195);
and U12281 (N_12281,N_11790,N_10099);
or U12282 (N_12282,N_11880,N_11814);
and U12283 (N_12283,N_11326,N_10892);
nand U12284 (N_12284,N_11323,N_10271);
nand U12285 (N_12285,N_11253,N_10117);
nand U12286 (N_12286,N_10966,N_10007);
xnor U12287 (N_12287,N_11858,N_10381);
and U12288 (N_12288,N_11180,N_10425);
nor U12289 (N_12289,N_10192,N_10167);
nand U12290 (N_12290,N_10924,N_10762);
nand U12291 (N_12291,N_10207,N_11391);
xor U12292 (N_12292,N_10987,N_10232);
nor U12293 (N_12293,N_11454,N_10642);
or U12294 (N_12294,N_11674,N_11800);
or U12295 (N_12295,N_11009,N_11785);
or U12296 (N_12296,N_10452,N_11728);
nor U12297 (N_12297,N_11788,N_10522);
nor U12298 (N_12298,N_11935,N_10124);
nand U12299 (N_12299,N_10610,N_10670);
xnor U12300 (N_12300,N_11076,N_11700);
xnor U12301 (N_12301,N_10306,N_11804);
xor U12302 (N_12302,N_11459,N_10272);
and U12303 (N_12303,N_10472,N_11361);
nor U12304 (N_12304,N_10161,N_10193);
or U12305 (N_12305,N_11825,N_10366);
nand U12306 (N_12306,N_10475,N_11204);
nand U12307 (N_12307,N_10064,N_11392);
xor U12308 (N_12308,N_11701,N_10144);
or U12309 (N_12309,N_10109,N_11692);
and U12310 (N_12310,N_11212,N_11952);
nor U12311 (N_12311,N_11767,N_11213);
nand U12312 (N_12312,N_10789,N_10063);
xnor U12313 (N_12313,N_11332,N_10311);
nand U12314 (N_12314,N_10011,N_10552);
nor U12315 (N_12315,N_11104,N_11938);
nand U12316 (N_12316,N_10650,N_11781);
nor U12317 (N_12317,N_10392,N_11601);
nand U12318 (N_12318,N_11475,N_11573);
or U12319 (N_12319,N_10441,N_11287);
and U12320 (N_12320,N_11747,N_11139);
or U12321 (N_12321,N_11060,N_11643);
nor U12322 (N_12322,N_11637,N_11278);
or U12323 (N_12323,N_11789,N_10528);
nor U12324 (N_12324,N_10903,N_11661);
nor U12325 (N_12325,N_10309,N_10978);
nor U12326 (N_12326,N_10151,N_11808);
xor U12327 (N_12327,N_10162,N_10901);
nand U12328 (N_12328,N_11155,N_10169);
nand U12329 (N_12329,N_10443,N_10252);
or U12330 (N_12330,N_11917,N_11327);
or U12331 (N_12331,N_11803,N_11792);
nor U12332 (N_12332,N_10673,N_10678);
nand U12333 (N_12333,N_11051,N_10457);
nor U12334 (N_12334,N_11172,N_10569);
nor U12335 (N_12335,N_11626,N_11932);
xor U12336 (N_12336,N_10948,N_10217);
nand U12337 (N_12337,N_10285,N_11557);
xor U12338 (N_12338,N_10046,N_11721);
xnor U12339 (N_12339,N_10852,N_10183);
nand U12340 (N_12340,N_11095,N_11863);
xnor U12341 (N_12341,N_11397,N_10415);
or U12342 (N_12342,N_11632,N_11768);
or U12343 (N_12343,N_10290,N_10286);
or U12344 (N_12344,N_10337,N_11849);
xnor U12345 (N_12345,N_10312,N_11279);
nor U12346 (N_12346,N_11061,N_11192);
nor U12347 (N_12347,N_11019,N_10861);
and U12348 (N_12348,N_10346,N_11654);
nor U12349 (N_12349,N_10313,N_11752);
and U12350 (N_12350,N_10640,N_11128);
nand U12351 (N_12351,N_10147,N_10139);
or U12352 (N_12352,N_10946,N_10709);
nor U12353 (N_12353,N_10612,N_11465);
and U12354 (N_12354,N_11310,N_10245);
and U12355 (N_12355,N_10605,N_10755);
and U12356 (N_12356,N_10688,N_11655);
nor U12357 (N_12357,N_10476,N_11074);
or U12358 (N_12358,N_11222,N_10775);
nor U12359 (N_12359,N_11381,N_10333);
xor U12360 (N_12360,N_10367,N_11515);
and U12361 (N_12361,N_11117,N_11933);
nor U12362 (N_12362,N_10433,N_10753);
xor U12363 (N_12363,N_10779,N_10837);
and U12364 (N_12364,N_11322,N_10853);
nand U12365 (N_12365,N_10026,N_11988);
or U12366 (N_12366,N_11946,N_10994);
or U12367 (N_12367,N_11388,N_11426);
and U12368 (N_12368,N_11365,N_10375);
nand U12369 (N_12369,N_10777,N_11089);
nor U12370 (N_12370,N_11590,N_11748);
nand U12371 (N_12371,N_11912,N_11078);
and U12372 (N_12372,N_11950,N_10745);
nor U12373 (N_12373,N_11383,N_10803);
and U12374 (N_12374,N_10530,N_10847);
nor U12375 (N_12375,N_10649,N_10298);
or U12376 (N_12376,N_11960,N_11259);
nor U12377 (N_12377,N_11065,N_11695);
or U12378 (N_12378,N_10287,N_11295);
xnor U12379 (N_12379,N_10398,N_10066);
or U12380 (N_12380,N_10076,N_10113);
or U12381 (N_12381,N_11835,N_10019);
xnor U12382 (N_12382,N_11343,N_11532);
nand U12383 (N_12383,N_10663,N_10216);
and U12384 (N_12384,N_10949,N_11671);
and U12385 (N_12385,N_11003,N_11116);
and U12386 (N_12386,N_11448,N_10625);
nand U12387 (N_12387,N_11867,N_10095);
and U12388 (N_12388,N_11667,N_11614);
or U12389 (N_12389,N_10859,N_10714);
xnor U12390 (N_12390,N_10841,N_10632);
xnor U12391 (N_12391,N_11418,N_11101);
xor U12392 (N_12392,N_10023,N_10929);
and U12393 (N_12393,N_10336,N_10661);
nor U12394 (N_12394,N_10521,N_10157);
and U12395 (N_12395,N_11283,N_11704);
or U12396 (N_12396,N_11149,N_10851);
nor U12397 (N_12397,N_11964,N_11889);
nor U12398 (N_12398,N_10672,N_11050);
and U12399 (N_12399,N_10014,N_11976);
nand U12400 (N_12400,N_10863,N_10447);
or U12401 (N_12401,N_10652,N_11201);
or U12402 (N_12402,N_10536,N_10348);
and U12403 (N_12403,N_10985,N_10444);
nor U12404 (N_12404,N_11628,N_10205);
and U12405 (N_12405,N_10083,N_11446);
nand U12406 (N_12406,N_11121,N_10369);
xnor U12407 (N_12407,N_11145,N_10251);
and U12408 (N_12408,N_10568,N_10938);
and U12409 (N_12409,N_10350,N_10428);
nor U12410 (N_12410,N_10539,N_11313);
or U12411 (N_12411,N_10733,N_11156);
and U12412 (N_12412,N_10149,N_10209);
nand U12413 (N_12413,N_10429,N_10012);
or U12414 (N_12414,N_10870,N_11576);
xnor U12415 (N_12415,N_10427,N_11469);
and U12416 (N_12416,N_11443,N_10886);
and U12417 (N_12417,N_11958,N_10760);
xor U12418 (N_12418,N_10146,N_11495);
and U12419 (N_12419,N_11743,N_11926);
or U12420 (N_12420,N_11109,N_11462);
and U12421 (N_12421,N_11120,N_11650);
nor U12422 (N_12422,N_10107,N_11558);
xnor U12423 (N_12423,N_11965,N_10206);
nand U12424 (N_12424,N_10022,N_10194);
xor U12425 (N_12425,N_11782,N_10440);
and U12426 (N_12426,N_11291,N_11439);
or U12427 (N_12427,N_10907,N_10744);
xor U12428 (N_12428,N_11396,N_11297);
and U12429 (N_12429,N_10845,N_10743);
or U12430 (N_12430,N_11890,N_11209);
and U12431 (N_12431,N_11336,N_10075);
xor U12432 (N_12432,N_11980,N_11627);
xor U12433 (N_12433,N_10111,N_10723);
and U12434 (N_12434,N_10908,N_10486);
nor U12435 (N_12435,N_10618,N_10582);
xnor U12436 (N_12436,N_10417,N_10053);
xnor U12437 (N_12437,N_10274,N_11679);
nand U12438 (N_12438,N_10166,N_11366);
nor U12439 (N_12439,N_10506,N_10514);
nand U12440 (N_12440,N_10751,N_11830);
xor U12441 (N_12441,N_11900,N_10806);
xnor U12442 (N_12442,N_11899,N_10338);
and U12443 (N_12443,N_10758,N_10378);
xor U12444 (N_12444,N_11504,N_11762);
nand U12445 (N_12445,N_11275,N_10818);
and U12446 (N_12446,N_11053,N_11127);
nand U12447 (N_12447,N_10727,N_10328);
nor U12448 (N_12448,N_10163,N_11118);
nand U12449 (N_12449,N_11466,N_10264);
nand U12450 (N_12450,N_11369,N_11028);
xnor U12451 (N_12451,N_10695,N_10683);
or U12452 (N_12452,N_11518,N_11793);
xnor U12453 (N_12453,N_10219,N_11303);
xor U12454 (N_12454,N_10937,N_11774);
xnor U12455 (N_12455,N_10073,N_10814);
or U12456 (N_12456,N_10184,N_10414);
or U12457 (N_12457,N_10874,N_11753);
nor U12458 (N_12458,N_10941,N_10523);
and U12459 (N_12459,N_10840,N_11796);
nor U12460 (N_12460,N_10302,N_10260);
nor U12461 (N_12461,N_10487,N_11449);
xnor U12462 (N_12462,N_11909,N_11132);
and U12463 (N_12463,N_11481,N_10399);
nor U12464 (N_12464,N_11707,N_10675);
nand U12465 (N_12465,N_10846,N_10448);
and U12466 (N_12466,N_11471,N_10434);
nor U12467 (N_12467,N_11739,N_10029);
nand U12468 (N_12468,N_11002,N_11666);
nor U12469 (N_12469,N_11379,N_10003);
nor U12470 (N_12470,N_10384,N_10934);
nor U12471 (N_12471,N_11778,N_11087);
xor U12472 (N_12472,N_11807,N_11990);
or U12473 (N_12473,N_11292,N_10956);
nand U12474 (N_12474,N_11077,N_11649);
or U12475 (N_12475,N_11208,N_11186);
xor U12476 (N_12476,N_11770,N_10772);
nor U12477 (N_12477,N_10490,N_10304);
xor U12478 (N_12478,N_10603,N_10288);
or U12479 (N_12479,N_10988,N_11415);
nor U12480 (N_12480,N_10679,N_10451);
nand U12481 (N_12481,N_11042,N_11203);
and U12482 (N_12482,N_11513,N_10129);
and U12483 (N_12483,N_10048,N_11073);
and U12484 (N_12484,N_11531,N_11063);
and U12485 (N_12485,N_11243,N_11772);
nand U12486 (N_12486,N_10295,N_10071);
nand U12487 (N_12487,N_11320,N_11892);
nor U12488 (N_12488,N_11680,N_11738);
xor U12489 (N_12489,N_10984,N_11547);
nor U12490 (N_12490,N_11908,N_11285);
nor U12491 (N_12491,N_11435,N_10544);
and U12492 (N_12492,N_10959,N_11827);
and U12493 (N_12493,N_11621,N_10698);
xnor U12494 (N_12494,N_11444,N_10027);
or U12495 (N_12495,N_11181,N_11507);
nor U12496 (N_12496,N_10590,N_10825);
or U12497 (N_12497,N_10517,N_10706);
xnor U12498 (N_12498,N_11232,N_10278);
xor U12499 (N_12499,N_11227,N_11148);
nor U12500 (N_12500,N_11977,N_10082);
or U12501 (N_12501,N_11898,N_11493);
xor U12502 (N_12502,N_10639,N_10492);
nor U12503 (N_12503,N_10717,N_11927);
nand U12504 (N_12504,N_11427,N_11731);
xor U12505 (N_12505,N_11540,N_11006);
and U12506 (N_12506,N_11913,N_11588);
nand U12507 (N_12507,N_10377,N_11309);
nor U12508 (N_12508,N_11773,N_10831);
or U12509 (N_12509,N_11001,N_10613);
or U12510 (N_12510,N_10121,N_10594);
nor U12511 (N_12511,N_11944,N_11812);
and U12512 (N_12512,N_11351,N_11843);
nor U12513 (N_12513,N_11822,N_10563);
or U12514 (N_12514,N_11385,N_10729);
or U12515 (N_12515,N_11918,N_11146);
nor U12516 (N_12516,N_11555,N_10382);
nor U12517 (N_12517,N_11142,N_11562);
nand U12518 (N_12518,N_10551,N_10102);
and U12519 (N_12519,N_10466,N_11606);
nand U12520 (N_12520,N_10871,N_11877);
and U12521 (N_12521,N_10180,N_10439);
xor U12522 (N_12522,N_11476,N_11267);
or U12523 (N_12523,N_10781,N_11963);
and U12524 (N_12524,N_11687,N_10479);
nand U12525 (N_12525,N_10281,N_11131);
nor U12526 (N_12526,N_10900,N_11018);
nand U12527 (N_12527,N_10021,N_10361);
nand U12528 (N_12528,N_10494,N_10965);
or U12529 (N_12529,N_10643,N_11904);
and U12530 (N_12530,N_11257,N_11568);
or U12531 (N_12531,N_10239,N_10824);
nor U12532 (N_12532,N_11344,N_11106);
nand U12533 (N_12533,N_11022,N_10883);
xnor U12534 (N_12534,N_10454,N_10100);
nor U12535 (N_12535,N_10072,N_10120);
and U12536 (N_12536,N_11410,N_10799);
nor U12537 (N_12537,N_10548,N_11265);
nand U12538 (N_12538,N_10172,N_11024);
nor U12539 (N_12539,N_11163,N_11189);
and U12540 (N_12540,N_10138,N_10084);
nor U12541 (N_12541,N_10970,N_10540);
or U12542 (N_12542,N_11372,N_11694);
or U12543 (N_12543,N_10604,N_11974);
nor U12544 (N_12544,N_10343,N_11455);
xnor U12545 (N_12545,N_11071,N_11211);
or U12546 (N_12546,N_11602,N_10259);
or U12547 (N_12547,N_11461,N_11112);
or U12548 (N_12548,N_10323,N_10508);
xor U12549 (N_12549,N_11597,N_11230);
nand U12550 (N_12550,N_10238,N_11592);
nand U12551 (N_12551,N_11742,N_10921);
or U12552 (N_12552,N_10911,N_11325);
nor U12553 (N_12553,N_11068,N_10086);
xor U12554 (N_12554,N_10445,N_11097);
xnor U12555 (N_12555,N_11609,N_10110);
and U12556 (N_12556,N_11337,N_10049);
xor U12557 (N_12557,N_11025,N_11519);
nor U12558 (N_12558,N_11378,N_10637);
nand U12559 (N_12559,N_10301,N_10009);
nand U12560 (N_12560,N_10032,N_11499);
and U12561 (N_12561,N_11920,N_11624);
or U12562 (N_12562,N_10266,N_10101);
and U12563 (N_12563,N_10738,N_10420);
or U12564 (N_12564,N_10353,N_10360);
nor U12565 (N_12565,N_11905,N_10906);
nand U12566 (N_12566,N_11248,N_10681);
and U12567 (N_12567,N_11088,N_10767);
xor U12568 (N_12568,N_10331,N_10826);
and U12569 (N_12569,N_11979,N_11064);
nand U12570 (N_12570,N_11669,N_11165);
or U12571 (N_12571,N_11517,N_11340);
nor U12572 (N_12572,N_11542,N_10442);
xnor U12573 (N_12573,N_11660,N_10495);
and U12574 (N_12574,N_10330,N_11098);
or U12575 (N_12575,N_10926,N_10535);
nor U12576 (N_12576,N_10277,N_11719);
and U12577 (N_12577,N_10577,N_10967);
nor U12578 (N_12578,N_10925,N_10030);
xor U12579 (N_12579,N_10299,N_10178);
or U12580 (N_12580,N_10237,N_10186);
xnor U12581 (N_12581,N_11154,N_10780);
or U12582 (N_12582,N_10931,N_11631);
or U12583 (N_12583,N_11021,N_11049);
or U12584 (N_12584,N_11831,N_11797);
xnor U12585 (N_12585,N_10983,N_11923);
xor U12586 (N_12586,N_11714,N_10961);
and U12587 (N_12587,N_10040,N_10092);
nand U12588 (N_12588,N_11348,N_11103);
and U12589 (N_12589,N_11834,N_11736);
nand U12590 (N_12590,N_11037,N_10408);
or U12591 (N_12591,N_11450,N_10554);
and U12592 (N_12592,N_11347,N_10746);
nor U12593 (N_12593,N_10736,N_11302);
xnor U12594 (N_12594,N_10025,N_10793);
nand U12595 (N_12595,N_11683,N_11619);
nor U12596 (N_12596,N_11706,N_10221);
nor U12597 (N_12597,N_10782,N_11015);
xnor U12598 (N_12598,N_11837,N_11272);
nor U12599 (N_12599,N_10142,N_11354);
xor U12600 (N_12600,N_11535,N_11645);
xnor U12601 (N_12601,N_10255,N_11603);
and U12602 (N_12602,N_10362,N_11846);
xor U12603 (N_12603,N_10055,N_11086);
nand U12604 (N_12604,N_10928,N_10247);
and U12605 (N_12605,N_11173,N_11196);
nand U12606 (N_12606,N_10412,N_10383);
xor U12607 (N_12607,N_11972,N_11951);
nand U12608 (N_12608,N_11973,N_11563);
nand U12609 (N_12609,N_10716,N_10595);
and U12610 (N_12610,N_11735,N_10829);
xor U12611 (N_12611,N_11445,N_11306);
xor U12612 (N_12612,N_11338,N_10635);
or U12613 (N_12613,N_10638,N_11055);
nand U12614 (N_12614,N_10198,N_11670);
and U12615 (N_12615,N_10045,N_10449);
xnor U12616 (N_12616,N_10991,N_11293);
and U12617 (N_12617,N_11566,N_11376);
nand U12618 (N_12618,N_11300,N_11610);
and U12619 (N_12619,N_11430,N_10098);
and U12620 (N_12620,N_11862,N_10899);
nor U12621 (N_12621,N_10176,N_10230);
nor U12622 (N_12622,N_10957,N_10001);
nor U12623 (N_12623,N_11185,N_10787);
nand U12624 (N_12624,N_11182,N_11763);
or U12625 (N_12625,N_10303,N_11052);
and U12626 (N_12626,N_11520,N_10693);
xor U12627 (N_12627,N_10868,N_11470);
and U12628 (N_12628,N_10502,N_11402);
xnor U12629 (N_12629,N_10843,N_11726);
nand U12630 (N_12630,N_10401,N_11818);
nor U12631 (N_12631,N_10488,N_11888);
nor U12632 (N_12632,N_11914,N_11930);
nor U12633 (N_12633,N_11969,N_10373);
and U12634 (N_12634,N_10435,N_10034);
nand U12635 (N_12635,N_11489,N_11017);
and U12636 (N_12636,N_11732,N_10537);
xnor U12637 (N_12637,N_11484,N_10220);
or U12638 (N_12638,N_10557,N_11317);
or U12639 (N_12639,N_10137,N_10982);
nand U12640 (N_12640,N_10519,N_11315);
xnor U12641 (N_12641,N_11474,N_10682);
xnor U12642 (N_12642,N_10579,N_10213);
nor U12643 (N_12643,N_11611,N_10275);
nand U12644 (N_12644,N_11883,N_11784);
xor U12645 (N_12645,N_10996,N_10261);
xnor U12646 (N_12646,N_10236,N_11368);
nor U12647 (N_12647,N_10143,N_11585);
xor U12648 (N_12648,N_10280,N_11639);
and U12649 (N_12649,N_10467,N_10325);
nor U12650 (N_12650,N_11069,N_11514);
and U12651 (N_12651,N_10935,N_11553);
nor U12652 (N_12652,N_10215,N_10253);
nand U12653 (N_12653,N_11779,N_10691);
and U12654 (N_12654,N_11399,N_10127);
nand U12655 (N_12655,N_11578,N_11225);
nand U12656 (N_12656,N_10721,N_11215);
nand U12657 (N_12657,N_11031,N_10380);
nor U12658 (N_12658,N_11852,N_10386);
nor U12659 (N_12659,N_10526,N_11894);
nand U12660 (N_12660,N_10463,N_10474);
nand U12661 (N_12661,N_10623,N_11644);
xnor U12662 (N_12662,N_11479,N_10807);
and U12663 (N_12663,N_10013,N_11512);
xnor U12664 (N_12664,N_11158,N_11638);
and U12665 (N_12665,N_11123,N_11238);
nor U12666 (N_12666,N_11539,N_10037);
nor U12667 (N_12667,N_11370,N_11183);
or U12668 (N_12668,N_10882,N_10708);
or U12669 (N_12669,N_10531,N_10866);
and U12670 (N_12670,N_10694,N_11647);
and U12671 (N_12671,N_10617,N_11129);
xnor U12672 (N_12672,N_10785,N_10969);
or U12673 (N_12673,N_11902,N_11633);
nand U12674 (N_12674,N_10856,N_11819);
and U12675 (N_12675,N_10628,N_11850);
and U12676 (N_12676,N_10170,N_11617);
xor U12677 (N_12677,N_11115,N_11771);
nor U12678 (N_12678,N_11506,N_11485);
nor U12679 (N_12679,N_10854,N_11282);
nor U12680 (N_12680,N_11703,N_10002);
nor U12681 (N_12681,N_11884,N_11685);
and U12682 (N_12682,N_10351,N_10885);
and U12683 (N_12683,N_10783,N_10397);
nor U12684 (N_12684,N_10152,N_11817);
nand U12685 (N_12685,N_11538,N_10973);
and U12686 (N_12686,N_10571,N_10791);
and U12687 (N_12687,N_10616,N_11761);
or U12688 (N_12688,N_10406,N_11067);
xor U12689 (N_12689,N_11013,N_10608);
nor U12690 (N_12690,N_11016,N_11591);
nand U12691 (N_12691,N_11829,N_10450);
or U12692 (N_12692,N_10752,N_11985);
nand U12693 (N_12693,N_11276,N_11033);
xor U12694 (N_12694,N_10822,N_11560);
and U12695 (N_12695,N_10354,N_11100);
xor U12696 (N_12696,N_11871,N_11401);
or U12697 (N_12697,N_11975,N_10079);
and U12698 (N_12698,N_10513,N_11398);
or U12699 (N_12699,N_10202,N_11873);
nor U12700 (N_12700,N_10932,N_10069);
or U12701 (N_12701,N_11490,N_10795);
nor U12702 (N_12702,N_11421,N_11311);
nand U12703 (N_12703,N_10658,N_11939);
nor U12704 (N_12704,N_10355,N_11615);
nand U12705 (N_12705,N_10696,N_11056);
nor U12706 (N_12706,N_10971,N_10017);
nand U12707 (N_12707,N_11007,N_10542);
xnor U12708 (N_12708,N_10080,N_11586);
and U12709 (N_12709,N_10686,N_10989);
nand U12710 (N_12710,N_10128,N_11550);
nor U12711 (N_12711,N_10606,N_10374);
nor U12712 (N_12712,N_10622,N_11359);
or U12713 (N_12713,N_11371,N_10116);
nor U12714 (N_12714,N_11968,N_10242);
nand U12715 (N_12715,N_11921,N_10496);
nand U12716 (N_12716,N_10561,N_11373);
or U12717 (N_12717,N_11412,N_10910);
or U12718 (N_12718,N_11855,N_10234);
or U12719 (N_12719,N_11150,N_10918);
or U12720 (N_12720,N_11864,N_10297);
xnor U12721 (N_12721,N_10684,N_10740);
nor U12722 (N_12722,N_10902,N_11733);
nand U12723 (N_12723,N_11579,N_10955);
nor U12724 (N_12724,N_11866,N_10636);
and U12725 (N_12725,N_10340,N_10244);
nor U12726 (N_12726,N_10919,N_11179);
nand U12727 (N_12727,N_10133,N_10112);
nand U12728 (N_12728,N_10173,N_10944);
nand U12729 (N_12729,N_11254,N_11982);
nand U12730 (N_12730,N_10836,N_10653);
nand U12731 (N_12731,N_10797,N_10627);
nand U12732 (N_12732,N_10891,N_11978);
xnor U12733 (N_12733,N_11160,N_10914);
nor U12734 (N_12734,N_11341,N_10587);
xnor U12735 (N_12735,N_11713,N_10315);
nand U12736 (N_12736,N_11130,N_10409);
and U12737 (N_12737,N_10997,N_10018);
and U12738 (N_12738,N_11583,N_10258);
nor U12739 (N_12739,N_11233,N_11734);
or U12740 (N_12740,N_11523,N_10096);
nand U12741 (N_12741,N_11062,N_11533);
and U12742 (N_12742,N_10196,N_10334);
xnor U12743 (N_12743,N_11618,N_11545);
nor U12744 (N_12744,N_10204,N_11879);
nand U12745 (N_12745,N_10550,N_10243);
and U12746 (N_12746,N_10458,N_10963);
xor U12747 (N_12747,N_11754,N_11874);
nor U12748 (N_12748,N_10345,N_10329);
or U12749 (N_12749,N_10179,N_10125);
nor U12750 (N_12750,N_11581,N_11054);
and U12751 (N_12751,N_11414,N_11554);
or U12752 (N_12752,N_11107,N_11460);
nand U12753 (N_12753,N_11221,N_11854);
or U12754 (N_12754,N_10455,N_10936);
nand U12755 (N_12755,N_10199,N_10051);
nand U12756 (N_12756,N_10710,N_11600);
nor U12757 (N_12757,N_10503,N_10877);
xor U12758 (N_12758,N_11147,N_11725);
xnor U12759 (N_12759,N_11301,N_10294);
and U12760 (N_12760,N_10039,N_10005);
or U12761 (N_12761,N_11229,N_11226);
xnor U12762 (N_12762,N_11389,N_11143);
or U12763 (N_12763,N_11286,N_11070);
or U12764 (N_12764,N_10827,N_11207);
xnor U12765 (N_12765,N_10815,N_11836);
and U12766 (N_12766,N_11929,N_10089);
nand U12767 (N_12767,N_10894,N_11653);
nand U12768 (N_12768,N_11500,N_11319);
and U12769 (N_12769,N_11105,N_11235);
nand U12770 (N_12770,N_11012,N_10927);
and U12771 (N_12771,N_11826,N_10228);
nor U12772 (N_12772,N_11994,N_11218);
and U12773 (N_12773,N_11672,N_10462);
or U12774 (N_12774,N_11740,N_10372);
nor U12775 (N_12775,N_10584,N_11447);
or U12776 (N_12776,N_10697,N_11681);
nand U12777 (N_12777,N_10739,N_10015);
nor U12778 (N_12778,N_10609,N_10992);
nor U12779 (N_12779,N_10830,N_11690);
nand U12780 (N_12780,N_11084,N_11166);
nor U12781 (N_12781,N_10631,N_10728);
and U12782 (N_12782,N_10889,N_10269);
or U12783 (N_12783,N_10394,N_11841);
nand U12784 (N_12784,N_11998,N_10998);
xnor U12785 (N_12785,N_11153,N_10660);
or U12786 (N_12786,N_10188,N_10344);
or U12787 (N_12787,N_11688,N_11813);
xnor U12788 (N_12788,N_11357,N_10365);
nor U12789 (N_12789,N_11795,N_10734);
and U12790 (N_12790,N_10020,N_10211);
and U12791 (N_12791,N_11034,N_11324);
or U12792 (N_12792,N_11405,N_11029);
and U12793 (N_12793,N_10993,N_10747);
nand U12794 (N_12794,N_11205,N_11250);
nor U12795 (N_12795,N_10068,N_11806);
and U12796 (N_12796,N_10480,N_11126);
or U12797 (N_12797,N_10310,N_11027);
nor U12798 (N_12798,N_10761,N_11953);
nor U12799 (N_12799,N_11544,N_11047);
nor U12800 (N_12800,N_10126,N_11543);
nor U12801 (N_12801,N_11363,N_11710);
nand U12802 (N_12802,N_10335,N_10835);
nor U12803 (N_12803,N_10776,N_11709);
nor U12804 (N_12804,N_11119,N_11408);
nor U12805 (N_12805,N_10065,N_10724);
nand U12806 (N_12806,N_10629,N_11432);
and U12807 (N_12807,N_11816,N_11708);
xor U12808 (N_12808,N_10659,N_10119);
and U12809 (N_12809,N_11757,N_10811);
or U12810 (N_12810,N_11400,N_11897);
or U12811 (N_12811,N_10469,N_10615);
nand U12812 (N_12812,N_10666,N_10181);
nand U12813 (N_12813,N_11516,N_11564);
and U12814 (N_12814,N_11811,N_11268);
nand U12815 (N_12815,N_10532,N_11613);
and U12816 (N_12816,N_11058,N_10131);
xnor U12817 (N_12817,N_10884,N_11219);
xor U12818 (N_12818,N_10766,N_10471);
or U12819 (N_12819,N_10875,N_11175);
xnor U12820 (N_12820,N_11571,N_10599);
or U12821 (N_12821,N_11057,N_10890);
xnor U12822 (N_12822,N_10873,N_11575);
nand U12823 (N_12823,N_11434,N_10284);
nand U12824 (N_12824,N_11783,N_11828);
nand U12825 (N_12825,N_11362,N_11744);
or U12826 (N_12826,N_10387,N_11595);
or U12827 (N_12827,N_11943,N_11429);
or U12828 (N_12828,N_11870,N_11966);
or U12829 (N_12829,N_11925,N_10614);
nor U12830 (N_12830,N_10390,N_10651);
nand U12831 (N_12831,N_10922,N_10671);
nor U12832 (N_12832,N_11751,N_11404);
nand U12833 (N_12833,N_11346,N_11663);
and U12834 (N_12834,N_11200,N_11240);
nand U12835 (N_12835,N_10813,N_10656);
xor U12836 (N_12836,N_10718,N_10070);
nor U12837 (N_12837,N_10754,N_10867);
xor U12838 (N_12838,N_11239,N_11038);
or U12839 (N_12839,N_11437,N_10262);
xnor U12840 (N_12840,N_10016,N_10385);
nor U12841 (N_12841,N_11594,N_11403);
xor U12842 (N_12842,N_10701,N_11171);
and U12843 (N_12843,N_11141,N_11875);
nor U12844 (N_12844,N_11174,N_10533);
or U12845 (N_12845,N_11151,N_11587);
and U12846 (N_12846,N_10689,N_10105);
nor U12847 (N_12847,N_10555,N_10043);
xor U12848 (N_12848,N_10804,N_10153);
or U12849 (N_12849,N_11787,N_10222);
nor U12850 (N_12850,N_10489,N_11842);
nor U12851 (N_12851,N_11749,N_10150);
and U12852 (N_12852,N_10620,N_10773);
or U12853 (N_12853,N_11536,N_10947);
and U12854 (N_12854,N_11741,N_10792);
nor U12855 (N_12855,N_10233,N_10832);
nand U12856 (N_12856,N_10087,N_11045);
nor U12857 (N_12857,N_10296,N_10160);
nand U12858 (N_12858,N_10185,N_11589);
nand U12859 (N_12859,N_11872,N_10737);
and U12860 (N_12860,N_10509,N_10115);
nand U12861 (N_12861,N_10000,N_10828);
nand U12862 (N_12862,N_11996,N_10008);
and U12863 (N_12863,N_11228,N_11651);
and U12864 (N_12864,N_10850,N_11177);
nand U12865 (N_12865,N_11967,N_11241);
nor U12866 (N_12866,N_10477,N_10953);
nand U12867 (N_12867,N_10707,N_10459);
and U12868 (N_12868,N_11989,N_10527);
nand U12869 (N_12869,N_11395,N_10801);
and U12870 (N_12870,N_10644,N_10470);
or U12871 (N_12871,N_11234,N_10468);
xor U12872 (N_12872,N_10456,N_11290);
xnor U12873 (N_12873,N_10191,N_10855);
and U12874 (N_12874,N_10920,N_11386);
xor U12875 (N_12875,N_10559,N_11537);
nand U12876 (N_12876,N_10541,N_10270);
or U12877 (N_12877,N_10481,N_11345);
nand U12878 (N_12878,N_10720,N_11729);
nor U12879 (N_12879,N_11678,N_11144);
nand U12880 (N_12880,N_11093,N_11756);
and U12881 (N_12881,N_11030,N_11262);
xnor U12882 (N_12882,N_10200,N_11906);
nand U12883 (N_12883,N_10878,N_10267);
xor U12884 (N_12884,N_11949,N_11111);
nor U12885 (N_12885,N_11664,N_11931);
nor U12886 (N_12886,N_11048,N_11374);
and U12887 (N_12887,N_11080,N_11483);
xor U12888 (N_12888,N_11387,N_11244);
nand U12889 (N_12889,N_11438,N_11082);
nor U12890 (N_12890,N_10122,N_11328);
xor U12891 (N_12891,N_10790,N_11745);
or U12892 (N_12892,N_10265,N_10796);
nor U12893 (N_12893,N_11202,N_10203);
xnor U12894 (N_12894,N_10424,N_11922);
nor U12895 (N_12895,N_11197,N_11524);
xor U12896 (N_12896,N_11008,N_11463);
or U12897 (N_12897,N_11957,N_10400);
xor U12898 (N_12898,N_10732,N_11046);
nor U12899 (N_12899,N_11844,N_10759);
or U12900 (N_12900,N_11284,N_10602);
nand U12901 (N_12901,N_10596,N_11656);
or U12902 (N_12902,N_11298,N_11110);
xnor U12903 (N_12903,N_11169,N_11821);
nor U12904 (N_12904,N_11847,N_11245);
nand U12905 (N_12905,N_11260,N_11251);
xor U12906 (N_12906,N_11521,N_11810);
nand U12907 (N_12907,N_10646,N_10145);
and U12908 (N_12908,N_11281,N_11599);
nor U12909 (N_12909,N_10576,N_10923);
nor U12910 (N_12910,N_11375,N_10028);
nand U12911 (N_12911,N_11596,N_10376);
or U12912 (N_12912,N_10223,N_10410);
or U12913 (N_12913,N_11838,N_10158);
or U12914 (N_12914,N_11036,N_11941);
or U12915 (N_12915,N_11456,N_10368);
nand U12916 (N_12916,N_10090,N_11270);
or U12917 (N_12917,N_10547,N_11718);
nor U12918 (N_12918,N_11407,N_10135);
and U12919 (N_12919,N_11995,N_11223);
xnor U12920 (N_12920,N_11598,N_11693);
or U12921 (N_12921,N_10314,N_11312);
and U12922 (N_12922,N_11928,N_10300);
xor U12923 (N_12923,N_10798,N_11501);
or U12924 (N_12924,N_10422,N_10437);
xor U12925 (N_12925,N_11494,N_11168);
nand U12926 (N_12926,N_11677,N_11473);
nand U12927 (N_12927,N_11522,N_10575);
or U12928 (N_12928,N_11868,N_10208);
and U12929 (N_12929,N_10104,N_10134);
xnor U12930 (N_12930,N_10976,N_10241);
nand U12931 (N_12931,N_11887,N_11486);
xnor U12932 (N_12932,N_10764,N_11711);
xnor U12933 (N_12933,N_11634,N_11801);
nand U12934 (N_12934,N_10091,N_10895);
nand U12935 (N_12935,N_11548,N_10321);
or U12936 (N_12936,N_11569,N_10108);
xor U12937 (N_12937,N_10235,N_11249);
and U12938 (N_12938,N_11296,N_11231);
xor U12939 (N_12939,N_11010,N_11604);
nand U12940 (N_12940,N_10393,N_10833);
xnor U12941 (N_12941,N_11986,N_11102);
nand U12942 (N_12942,N_11299,N_10214);
nor U12943 (N_12943,N_10730,N_10500);
or U12944 (N_12944,N_10964,N_10289);
or U12945 (N_12945,N_10842,N_11699);
xor U12946 (N_12946,N_10930,N_10396);
and U12947 (N_12947,N_10680,N_11164);
nand U12948 (N_12948,N_10227,N_11023);
nor U12949 (N_12949,N_11428,N_11956);
or U12950 (N_12950,N_10155,N_11255);
nand U12951 (N_12951,N_11765,N_10056);
xnor U12952 (N_12952,N_10954,N_11113);
xor U12953 (N_12953,N_11878,N_10085);
and U12954 (N_12954,N_11934,N_11937);
or U12955 (N_12955,N_11043,N_11094);
and U12956 (N_12956,N_10404,N_11546);
nand U12957 (N_12957,N_11099,N_10436);
xnor U12958 (N_12958,N_11853,N_11720);
xor U12959 (N_12959,N_10525,N_10349);
or U12960 (N_12960,N_11453,N_10156);
or U12961 (N_12961,N_10556,N_11440);
xnor U12962 (N_12962,N_10589,N_11712);
nand U12963 (N_12963,N_11549,N_11502);
nand U12964 (N_12964,N_11556,N_10872);
nand U12965 (N_12965,N_11237,N_10975);
or U12966 (N_12966,N_11032,N_11961);
xnor U12967 (N_12967,N_10788,N_10058);
xnor U12968 (N_12968,N_11458,N_10917);
xor U12969 (N_12969,N_10879,N_11035);
xnor U12970 (N_12970,N_11722,N_10915);
nand U12971 (N_12971,N_10418,N_11947);
and U12972 (N_12972,N_10504,N_11529);
and U12973 (N_12973,N_11417,N_10570);
nor U12974 (N_12974,N_10308,N_10898);
nand U12975 (N_12975,N_10305,N_10705);
or U12976 (N_12976,N_10268,N_11987);
nand U12977 (N_12977,N_10052,N_11274);
nor U12978 (N_12978,N_10359,N_10849);
nor U12979 (N_12979,N_10951,N_11857);
nor U12980 (N_12980,N_11138,N_10567);
and U12981 (N_12981,N_11860,N_11640);
nor U12982 (N_12982,N_11869,N_11210);
nand U12983 (N_12983,N_11083,N_10081);
nand U12984 (N_12984,N_11845,N_10741);
nand U12985 (N_12985,N_10240,N_10356);
and U12986 (N_12986,N_10857,N_10601);
nor U12987 (N_12987,N_11527,N_10722);
xnor U12988 (N_12988,N_11959,N_10942);
nor U12989 (N_12989,N_10316,N_10687);
or U12990 (N_12990,N_11377,N_11314);
nand U12991 (N_12991,N_10419,N_10461);
nor U12992 (N_12992,N_11294,N_10593);
nor U12993 (N_12993,N_11252,N_10402);
xnor U12994 (N_12994,N_11582,N_10159);
nand U12995 (N_12995,N_10464,N_11541);
nand U12996 (N_12996,N_11503,N_11264);
and U12997 (N_12997,N_10279,N_10307);
nor U12998 (N_12998,N_11096,N_10446);
or U12999 (N_12999,N_10864,N_11876);
and U13000 (N_13000,N_11816,N_11922);
xor U13001 (N_13001,N_10781,N_11483);
nand U13002 (N_13002,N_11517,N_11724);
or U13003 (N_13003,N_11678,N_11807);
or U13004 (N_13004,N_10086,N_10918);
nand U13005 (N_13005,N_10338,N_10971);
and U13006 (N_13006,N_11983,N_10970);
or U13007 (N_13007,N_10739,N_11756);
nand U13008 (N_13008,N_11608,N_10177);
nor U13009 (N_13009,N_11199,N_10799);
and U13010 (N_13010,N_10320,N_10719);
and U13011 (N_13011,N_11059,N_11603);
xnor U13012 (N_13012,N_11873,N_11844);
nor U13013 (N_13013,N_11089,N_10676);
or U13014 (N_13014,N_11196,N_10878);
and U13015 (N_13015,N_11348,N_10936);
or U13016 (N_13016,N_10341,N_10544);
nand U13017 (N_13017,N_10505,N_11278);
nor U13018 (N_13018,N_11589,N_10537);
xnor U13019 (N_13019,N_10844,N_10732);
xor U13020 (N_13020,N_11162,N_10465);
nand U13021 (N_13021,N_10056,N_11779);
xor U13022 (N_13022,N_11217,N_11608);
nor U13023 (N_13023,N_10648,N_10275);
and U13024 (N_13024,N_11532,N_10148);
and U13025 (N_13025,N_10899,N_10863);
nand U13026 (N_13026,N_11638,N_10726);
and U13027 (N_13027,N_10006,N_10346);
or U13028 (N_13028,N_11112,N_10155);
xor U13029 (N_13029,N_11665,N_10213);
and U13030 (N_13030,N_11635,N_10112);
xnor U13031 (N_13031,N_10246,N_10872);
or U13032 (N_13032,N_10346,N_11656);
and U13033 (N_13033,N_10528,N_10913);
or U13034 (N_13034,N_11936,N_10951);
or U13035 (N_13035,N_11540,N_10417);
nand U13036 (N_13036,N_11594,N_11237);
nand U13037 (N_13037,N_11240,N_10291);
and U13038 (N_13038,N_10505,N_10626);
nand U13039 (N_13039,N_11413,N_11210);
and U13040 (N_13040,N_11697,N_10025);
and U13041 (N_13041,N_10065,N_10491);
and U13042 (N_13042,N_10467,N_11890);
and U13043 (N_13043,N_10958,N_11300);
xor U13044 (N_13044,N_10915,N_10523);
nor U13045 (N_13045,N_11488,N_11138);
nor U13046 (N_13046,N_11443,N_10190);
nor U13047 (N_13047,N_10834,N_10648);
or U13048 (N_13048,N_10385,N_11066);
xnor U13049 (N_13049,N_10301,N_11474);
or U13050 (N_13050,N_11331,N_10483);
or U13051 (N_13051,N_11802,N_11028);
nor U13052 (N_13052,N_11050,N_11961);
or U13053 (N_13053,N_11725,N_10675);
nand U13054 (N_13054,N_11991,N_11932);
nor U13055 (N_13055,N_10556,N_10416);
nor U13056 (N_13056,N_11936,N_11173);
xnor U13057 (N_13057,N_11016,N_10310);
nand U13058 (N_13058,N_11504,N_11474);
xor U13059 (N_13059,N_10902,N_11268);
or U13060 (N_13060,N_11836,N_10243);
xor U13061 (N_13061,N_10369,N_11428);
nor U13062 (N_13062,N_11029,N_10953);
xor U13063 (N_13063,N_10567,N_11916);
nor U13064 (N_13064,N_10446,N_11987);
and U13065 (N_13065,N_11814,N_10563);
nand U13066 (N_13066,N_11063,N_11140);
nor U13067 (N_13067,N_10954,N_10656);
nor U13068 (N_13068,N_10453,N_11704);
xor U13069 (N_13069,N_10783,N_10560);
xor U13070 (N_13070,N_10916,N_11801);
and U13071 (N_13071,N_11988,N_10149);
and U13072 (N_13072,N_10395,N_11217);
xnor U13073 (N_13073,N_11738,N_10164);
and U13074 (N_13074,N_10730,N_11258);
nand U13075 (N_13075,N_11607,N_10676);
xnor U13076 (N_13076,N_11326,N_11013);
xnor U13077 (N_13077,N_10892,N_10574);
nand U13078 (N_13078,N_11898,N_10455);
nor U13079 (N_13079,N_11714,N_11478);
xnor U13080 (N_13080,N_10093,N_10784);
and U13081 (N_13081,N_11966,N_11278);
nor U13082 (N_13082,N_10841,N_11045);
xnor U13083 (N_13083,N_10391,N_10352);
xor U13084 (N_13084,N_10153,N_11315);
nor U13085 (N_13085,N_11184,N_10481);
nor U13086 (N_13086,N_11563,N_11136);
nor U13087 (N_13087,N_11636,N_11095);
nor U13088 (N_13088,N_11116,N_10593);
nor U13089 (N_13089,N_11541,N_10395);
xor U13090 (N_13090,N_11306,N_10407);
and U13091 (N_13091,N_11369,N_10868);
nor U13092 (N_13092,N_10052,N_11581);
xor U13093 (N_13093,N_10191,N_11463);
nor U13094 (N_13094,N_11180,N_11413);
nor U13095 (N_13095,N_10910,N_11255);
and U13096 (N_13096,N_11231,N_10073);
and U13097 (N_13097,N_11399,N_10113);
nand U13098 (N_13098,N_11358,N_11493);
or U13099 (N_13099,N_10733,N_10381);
or U13100 (N_13100,N_10773,N_10897);
xnor U13101 (N_13101,N_10564,N_11631);
and U13102 (N_13102,N_11999,N_11875);
nor U13103 (N_13103,N_11786,N_11091);
nor U13104 (N_13104,N_10315,N_10355);
nor U13105 (N_13105,N_11797,N_11689);
nand U13106 (N_13106,N_11242,N_11916);
or U13107 (N_13107,N_10739,N_11329);
xor U13108 (N_13108,N_10305,N_10460);
and U13109 (N_13109,N_11321,N_11201);
and U13110 (N_13110,N_11768,N_11117);
xnor U13111 (N_13111,N_10607,N_11312);
nor U13112 (N_13112,N_11274,N_10729);
or U13113 (N_13113,N_11839,N_10781);
nand U13114 (N_13114,N_11622,N_11011);
nor U13115 (N_13115,N_11882,N_11073);
and U13116 (N_13116,N_10978,N_10709);
nand U13117 (N_13117,N_10699,N_11715);
xnor U13118 (N_13118,N_10403,N_10948);
nor U13119 (N_13119,N_10170,N_10237);
nor U13120 (N_13120,N_11548,N_11010);
nor U13121 (N_13121,N_10595,N_11283);
nor U13122 (N_13122,N_11913,N_10820);
nor U13123 (N_13123,N_11211,N_10869);
nor U13124 (N_13124,N_10791,N_11362);
or U13125 (N_13125,N_11169,N_10827);
or U13126 (N_13126,N_11063,N_11720);
or U13127 (N_13127,N_11986,N_11838);
or U13128 (N_13128,N_10026,N_11558);
nor U13129 (N_13129,N_11310,N_11588);
xnor U13130 (N_13130,N_11061,N_10535);
xnor U13131 (N_13131,N_10380,N_11510);
or U13132 (N_13132,N_11731,N_11287);
and U13133 (N_13133,N_11265,N_10664);
nor U13134 (N_13134,N_11248,N_10241);
or U13135 (N_13135,N_10997,N_10107);
xor U13136 (N_13136,N_10075,N_11879);
xor U13137 (N_13137,N_11619,N_10062);
or U13138 (N_13138,N_11351,N_10305);
nand U13139 (N_13139,N_11959,N_11117);
nor U13140 (N_13140,N_10723,N_11399);
nand U13141 (N_13141,N_11443,N_11699);
nand U13142 (N_13142,N_11330,N_11839);
and U13143 (N_13143,N_10610,N_10823);
and U13144 (N_13144,N_11029,N_10278);
and U13145 (N_13145,N_10795,N_11919);
nor U13146 (N_13146,N_11570,N_10647);
or U13147 (N_13147,N_11985,N_10612);
xor U13148 (N_13148,N_11234,N_11877);
or U13149 (N_13149,N_10040,N_11824);
and U13150 (N_13150,N_11528,N_11120);
or U13151 (N_13151,N_11937,N_10094);
xor U13152 (N_13152,N_11420,N_11897);
or U13153 (N_13153,N_10458,N_10981);
nor U13154 (N_13154,N_10331,N_10871);
and U13155 (N_13155,N_11182,N_11798);
nor U13156 (N_13156,N_10481,N_11773);
nand U13157 (N_13157,N_10986,N_10698);
and U13158 (N_13158,N_10796,N_11130);
nand U13159 (N_13159,N_10840,N_11241);
or U13160 (N_13160,N_10213,N_10550);
nor U13161 (N_13161,N_11589,N_10942);
xnor U13162 (N_13162,N_10322,N_11668);
nand U13163 (N_13163,N_10870,N_11170);
nor U13164 (N_13164,N_11839,N_10970);
or U13165 (N_13165,N_11545,N_10161);
or U13166 (N_13166,N_11078,N_10314);
and U13167 (N_13167,N_11128,N_11335);
xor U13168 (N_13168,N_10631,N_11226);
nor U13169 (N_13169,N_10402,N_10676);
and U13170 (N_13170,N_10176,N_10864);
nand U13171 (N_13171,N_10443,N_10406);
xnor U13172 (N_13172,N_10923,N_11958);
nand U13173 (N_13173,N_10467,N_10932);
nor U13174 (N_13174,N_10536,N_10924);
nand U13175 (N_13175,N_10507,N_11482);
nor U13176 (N_13176,N_10081,N_11678);
nand U13177 (N_13177,N_11976,N_10678);
and U13178 (N_13178,N_11575,N_11977);
xnor U13179 (N_13179,N_11185,N_11141);
xnor U13180 (N_13180,N_11268,N_10199);
xnor U13181 (N_13181,N_10473,N_11236);
nor U13182 (N_13182,N_11758,N_11925);
xor U13183 (N_13183,N_11664,N_11762);
nor U13184 (N_13184,N_11831,N_11054);
and U13185 (N_13185,N_11950,N_10257);
xnor U13186 (N_13186,N_10251,N_10587);
xor U13187 (N_13187,N_10913,N_10042);
and U13188 (N_13188,N_11479,N_11441);
and U13189 (N_13189,N_11286,N_11507);
or U13190 (N_13190,N_10365,N_10370);
or U13191 (N_13191,N_11925,N_10647);
and U13192 (N_13192,N_10876,N_11088);
or U13193 (N_13193,N_11131,N_11373);
nor U13194 (N_13194,N_10225,N_11497);
or U13195 (N_13195,N_11608,N_10126);
nor U13196 (N_13196,N_11277,N_10403);
nand U13197 (N_13197,N_11388,N_11356);
nor U13198 (N_13198,N_10231,N_11392);
xor U13199 (N_13199,N_11145,N_10968);
or U13200 (N_13200,N_11899,N_10270);
nand U13201 (N_13201,N_10319,N_10110);
nand U13202 (N_13202,N_11225,N_11598);
and U13203 (N_13203,N_11421,N_10233);
nor U13204 (N_13204,N_11575,N_11524);
or U13205 (N_13205,N_11567,N_10522);
and U13206 (N_13206,N_11118,N_10498);
or U13207 (N_13207,N_10212,N_11462);
nor U13208 (N_13208,N_10981,N_11788);
xnor U13209 (N_13209,N_10373,N_11003);
nor U13210 (N_13210,N_10541,N_10104);
xnor U13211 (N_13211,N_10645,N_10488);
or U13212 (N_13212,N_10374,N_11436);
or U13213 (N_13213,N_11344,N_11997);
and U13214 (N_13214,N_11328,N_10529);
or U13215 (N_13215,N_10606,N_10448);
nand U13216 (N_13216,N_10661,N_11582);
nand U13217 (N_13217,N_11068,N_10521);
nor U13218 (N_13218,N_11296,N_11689);
or U13219 (N_13219,N_11712,N_10530);
or U13220 (N_13220,N_11577,N_10231);
and U13221 (N_13221,N_10977,N_10044);
xor U13222 (N_13222,N_10557,N_10055);
nor U13223 (N_13223,N_10249,N_10229);
and U13224 (N_13224,N_11771,N_10688);
xor U13225 (N_13225,N_11330,N_10556);
xor U13226 (N_13226,N_10779,N_11415);
or U13227 (N_13227,N_11909,N_10138);
and U13228 (N_13228,N_10965,N_10973);
or U13229 (N_13229,N_11325,N_10270);
or U13230 (N_13230,N_11463,N_10829);
or U13231 (N_13231,N_10291,N_10590);
and U13232 (N_13232,N_10767,N_11323);
xor U13233 (N_13233,N_11583,N_10620);
or U13234 (N_13234,N_11977,N_10142);
xor U13235 (N_13235,N_11978,N_11379);
and U13236 (N_13236,N_11272,N_11035);
nand U13237 (N_13237,N_10575,N_11030);
nor U13238 (N_13238,N_11395,N_10052);
nand U13239 (N_13239,N_10033,N_11246);
or U13240 (N_13240,N_11314,N_10216);
and U13241 (N_13241,N_11675,N_11790);
or U13242 (N_13242,N_11938,N_11197);
nand U13243 (N_13243,N_10070,N_10063);
nor U13244 (N_13244,N_11473,N_10045);
and U13245 (N_13245,N_10876,N_11005);
or U13246 (N_13246,N_10032,N_11363);
and U13247 (N_13247,N_11062,N_11687);
xor U13248 (N_13248,N_11011,N_11659);
nand U13249 (N_13249,N_10194,N_10500);
xor U13250 (N_13250,N_10021,N_11995);
and U13251 (N_13251,N_11445,N_11678);
nand U13252 (N_13252,N_11529,N_11691);
xor U13253 (N_13253,N_10963,N_10624);
and U13254 (N_13254,N_10492,N_10471);
and U13255 (N_13255,N_11481,N_10561);
nand U13256 (N_13256,N_11647,N_11764);
nand U13257 (N_13257,N_10521,N_10884);
nand U13258 (N_13258,N_10507,N_11604);
nor U13259 (N_13259,N_11361,N_11818);
xnor U13260 (N_13260,N_11338,N_11347);
and U13261 (N_13261,N_10633,N_11842);
xor U13262 (N_13262,N_11615,N_10448);
nor U13263 (N_13263,N_11363,N_11143);
or U13264 (N_13264,N_10919,N_11667);
nand U13265 (N_13265,N_10447,N_10064);
nor U13266 (N_13266,N_10666,N_11375);
or U13267 (N_13267,N_11925,N_11261);
nand U13268 (N_13268,N_11701,N_11829);
or U13269 (N_13269,N_10550,N_11088);
xnor U13270 (N_13270,N_10333,N_11852);
or U13271 (N_13271,N_10269,N_10206);
and U13272 (N_13272,N_11581,N_11454);
xor U13273 (N_13273,N_10008,N_11015);
or U13274 (N_13274,N_11406,N_11730);
or U13275 (N_13275,N_11421,N_11807);
or U13276 (N_13276,N_11650,N_11333);
xnor U13277 (N_13277,N_11962,N_11465);
nand U13278 (N_13278,N_11980,N_10956);
nor U13279 (N_13279,N_10625,N_11838);
nor U13280 (N_13280,N_10969,N_11101);
nor U13281 (N_13281,N_11919,N_11123);
or U13282 (N_13282,N_10595,N_11148);
xnor U13283 (N_13283,N_10189,N_10786);
nand U13284 (N_13284,N_10768,N_10994);
nor U13285 (N_13285,N_10111,N_10231);
xnor U13286 (N_13286,N_11818,N_10322);
and U13287 (N_13287,N_11988,N_10808);
nand U13288 (N_13288,N_10771,N_10179);
and U13289 (N_13289,N_11847,N_10229);
nand U13290 (N_13290,N_11593,N_10510);
or U13291 (N_13291,N_11155,N_11624);
and U13292 (N_13292,N_11041,N_10088);
xor U13293 (N_13293,N_10752,N_10716);
nand U13294 (N_13294,N_10166,N_10931);
nand U13295 (N_13295,N_10305,N_11257);
or U13296 (N_13296,N_10207,N_11256);
nand U13297 (N_13297,N_11364,N_10251);
and U13298 (N_13298,N_11827,N_11152);
nor U13299 (N_13299,N_10509,N_11122);
xnor U13300 (N_13300,N_11080,N_11558);
or U13301 (N_13301,N_10687,N_11299);
xor U13302 (N_13302,N_11018,N_11524);
xnor U13303 (N_13303,N_11571,N_11892);
nor U13304 (N_13304,N_11042,N_10207);
nand U13305 (N_13305,N_10275,N_10461);
nand U13306 (N_13306,N_11418,N_10410);
nand U13307 (N_13307,N_10305,N_11143);
xor U13308 (N_13308,N_11382,N_11000);
nand U13309 (N_13309,N_10109,N_11736);
xnor U13310 (N_13310,N_11292,N_11087);
or U13311 (N_13311,N_10951,N_10083);
or U13312 (N_13312,N_11701,N_10712);
nor U13313 (N_13313,N_10273,N_11451);
and U13314 (N_13314,N_11309,N_10693);
nand U13315 (N_13315,N_11367,N_10498);
and U13316 (N_13316,N_11874,N_11993);
xor U13317 (N_13317,N_10729,N_11445);
nor U13318 (N_13318,N_10375,N_10161);
xnor U13319 (N_13319,N_11050,N_11633);
nor U13320 (N_13320,N_10890,N_10925);
and U13321 (N_13321,N_11130,N_11942);
xnor U13322 (N_13322,N_10693,N_11697);
or U13323 (N_13323,N_11161,N_10064);
and U13324 (N_13324,N_10345,N_11010);
and U13325 (N_13325,N_11664,N_11230);
and U13326 (N_13326,N_10648,N_10539);
and U13327 (N_13327,N_11560,N_10469);
xnor U13328 (N_13328,N_10499,N_10354);
xor U13329 (N_13329,N_10823,N_11391);
or U13330 (N_13330,N_11863,N_10644);
nand U13331 (N_13331,N_10118,N_11815);
and U13332 (N_13332,N_10710,N_11555);
xor U13333 (N_13333,N_10545,N_11702);
nor U13334 (N_13334,N_11297,N_11401);
nor U13335 (N_13335,N_11771,N_10088);
nand U13336 (N_13336,N_11963,N_11032);
or U13337 (N_13337,N_10912,N_10082);
xnor U13338 (N_13338,N_10970,N_11521);
xnor U13339 (N_13339,N_11333,N_11665);
and U13340 (N_13340,N_11927,N_10808);
nand U13341 (N_13341,N_11039,N_10093);
nor U13342 (N_13342,N_11490,N_10175);
nand U13343 (N_13343,N_11883,N_10324);
or U13344 (N_13344,N_10878,N_11921);
nand U13345 (N_13345,N_11197,N_10103);
or U13346 (N_13346,N_11252,N_10479);
nor U13347 (N_13347,N_11017,N_10848);
xor U13348 (N_13348,N_11060,N_10462);
xor U13349 (N_13349,N_10018,N_10939);
nand U13350 (N_13350,N_11284,N_11098);
nand U13351 (N_13351,N_10439,N_10013);
nand U13352 (N_13352,N_10701,N_11388);
or U13353 (N_13353,N_10453,N_11723);
or U13354 (N_13354,N_11223,N_10955);
nor U13355 (N_13355,N_11058,N_10033);
nor U13356 (N_13356,N_11378,N_11465);
and U13357 (N_13357,N_11649,N_11768);
nand U13358 (N_13358,N_10292,N_10781);
and U13359 (N_13359,N_11862,N_10052);
xnor U13360 (N_13360,N_10377,N_11742);
xor U13361 (N_13361,N_10320,N_11059);
and U13362 (N_13362,N_11190,N_10484);
nor U13363 (N_13363,N_11576,N_11201);
and U13364 (N_13364,N_10900,N_11409);
nand U13365 (N_13365,N_10933,N_11346);
and U13366 (N_13366,N_11504,N_10093);
nand U13367 (N_13367,N_10288,N_11099);
xor U13368 (N_13368,N_10304,N_11669);
and U13369 (N_13369,N_10325,N_11995);
nand U13370 (N_13370,N_10700,N_10798);
or U13371 (N_13371,N_10024,N_10322);
nand U13372 (N_13372,N_11857,N_10419);
xor U13373 (N_13373,N_10554,N_11788);
xnor U13374 (N_13374,N_11806,N_11292);
nand U13375 (N_13375,N_10009,N_11866);
nand U13376 (N_13376,N_10097,N_10810);
and U13377 (N_13377,N_11108,N_10636);
nor U13378 (N_13378,N_11609,N_10930);
nand U13379 (N_13379,N_10989,N_10011);
xor U13380 (N_13380,N_10717,N_10233);
xor U13381 (N_13381,N_10426,N_11309);
xor U13382 (N_13382,N_11431,N_11067);
nor U13383 (N_13383,N_11063,N_11360);
nand U13384 (N_13384,N_10673,N_10870);
nand U13385 (N_13385,N_10755,N_11734);
nand U13386 (N_13386,N_11113,N_10866);
and U13387 (N_13387,N_11779,N_10985);
xnor U13388 (N_13388,N_10023,N_11797);
xnor U13389 (N_13389,N_10646,N_11168);
xor U13390 (N_13390,N_10416,N_11222);
and U13391 (N_13391,N_11200,N_11237);
or U13392 (N_13392,N_10202,N_11332);
xor U13393 (N_13393,N_10895,N_10388);
nor U13394 (N_13394,N_10161,N_10248);
nand U13395 (N_13395,N_11040,N_10179);
or U13396 (N_13396,N_10092,N_10259);
nor U13397 (N_13397,N_11609,N_11950);
or U13398 (N_13398,N_10427,N_10520);
or U13399 (N_13399,N_11918,N_11175);
or U13400 (N_13400,N_10426,N_11575);
xnor U13401 (N_13401,N_10433,N_11944);
or U13402 (N_13402,N_11281,N_10077);
or U13403 (N_13403,N_11852,N_10416);
xor U13404 (N_13404,N_10874,N_10272);
nor U13405 (N_13405,N_10472,N_11766);
and U13406 (N_13406,N_11158,N_11194);
nand U13407 (N_13407,N_11994,N_11965);
or U13408 (N_13408,N_10005,N_11728);
xor U13409 (N_13409,N_10115,N_10935);
and U13410 (N_13410,N_10299,N_11359);
and U13411 (N_13411,N_11204,N_11107);
and U13412 (N_13412,N_10656,N_11750);
nor U13413 (N_13413,N_10287,N_11858);
nand U13414 (N_13414,N_11363,N_11497);
xor U13415 (N_13415,N_11231,N_11089);
or U13416 (N_13416,N_11887,N_10228);
or U13417 (N_13417,N_11371,N_10074);
or U13418 (N_13418,N_10552,N_11421);
nor U13419 (N_13419,N_11732,N_10787);
and U13420 (N_13420,N_11634,N_11794);
xor U13421 (N_13421,N_10968,N_10883);
and U13422 (N_13422,N_11360,N_11652);
nand U13423 (N_13423,N_10184,N_10362);
xor U13424 (N_13424,N_10264,N_10554);
xnor U13425 (N_13425,N_10725,N_11270);
nor U13426 (N_13426,N_10937,N_10702);
nor U13427 (N_13427,N_10221,N_10137);
nand U13428 (N_13428,N_11879,N_10913);
and U13429 (N_13429,N_11787,N_11124);
and U13430 (N_13430,N_10573,N_11409);
nand U13431 (N_13431,N_11716,N_10053);
nand U13432 (N_13432,N_11390,N_11078);
nor U13433 (N_13433,N_10796,N_10313);
or U13434 (N_13434,N_11247,N_11428);
and U13435 (N_13435,N_10689,N_10092);
nor U13436 (N_13436,N_10785,N_10354);
nand U13437 (N_13437,N_11526,N_11402);
and U13438 (N_13438,N_10501,N_10053);
nand U13439 (N_13439,N_10055,N_10355);
nor U13440 (N_13440,N_10172,N_10203);
nor U13441 (N_13441,N_10357,N_11791);
nor U13442 (N_13442,N_11777,N_10639);
nand U13443 (N_13443,N_10720,N_10377);
nor U13444 (N_13444,N_10837,N_10836);
xnor U13445 (N_13445,N_11304,N_10549);
nand U13446 (N_13446,N_10477,N_11825);
nor U13447 (N_13447,N_10853,N_10799);
nand U13448 (N_13448,N_11308,N_10621);
nand U13449 (N_13449,N_11065,N_11214);
xnor U13450 (N_13450,N_11852,N_11302);
or U13451 (N_13451,N_10655,N_11066);
or U13452 (N_13452,N_11421,N_11935);
and U13453 (N_13453,N_10201,N_11258);
and U13454 (N_13454,N_10413,N_10211);
or U13455 (N_13455,N_10773,N_11778);
xnor U13456 (N_13456,N_10920,N_11404);
xor U13457 (N_13457,N_11811,N_11353);
nor U13458 (N_13458,N_11991,N_10999);
and U13459 (N_13459,N_11851,N_10963);
and U13460 (N_13460,N_10783,N_11145);
and U13461 (N_13461,N_11692,N_11679);
nor U13462 (N_13462,N_10895,N_10962);
nand U13463 (N_13463,N_10166,N_11053);
or U13464 (N_13464,N_11409,N_11024);
nor U13465 (N_13465,N_10269,N_10166);
xor U13466 (N_13466,N_11788,N_10261);
nor U13467 (N_13467,N_11619,N_11558);
and U13468 (N_13468,N_11320,N_11645);
or U13469 (N_13469,N_10870,N_10232);
xnor U13470 (N_13470,N_11728,N_10811);
nand U13471 (N_13471,N_11922,N_10838);
nor U13472 (N_13472,N_11774,N_11869);
xnor U13473 (N_13473,N_11110,N_10919);
nor U13474 (N_13474,N_10196,N_10855);
nor U13475 (N_13475,N_10876,N_11670);
nand U13476 (N_13476,N_10499,N_11829);
nor U13477 (N_13477,N_11623,N_11904);
or U13478 (N_13478,N_11774,N_10435);
nand U13479 (N_13479,N_11066,N_11819);
nor U13480 (N_13480,N_10953,N_10608);
or U13481 (N_13481,N_10089,N_11736);
or U13482 (N_13482,N_10831,N_10126);
and U13483 (N_13483,N_11024,N_10794);
or U13484 (N_13484,N_10093,N_11082);
nor U13485 (N_13485,N_11984,N_10520);
nand U13486 (N_13486,N_11848,N_10638);
or U13487 (N_13487,N_11591,N_10158);
or U13488 (N_13488,N_10339,N_10855);
nand U13489 (N_13489,N_11945,N_10663);
nor U13490 (N_13490,N_11256,N_10310);
xnor U13491 (N_13491,N_10526,N_10034);
nor U13492 (N_13492,N_11234,N_11102);
xnor U13493 (N_13493,N_10369,N_11211);
nand U13494 (N_13494,N_11392,N_10934);
nand U13495 (N_13495,N_10221,N_10533);
xnor U13496 (N_13496,N_10216,N_11123);
nor U13497 (N_13497,N_10921,N_11021);
or U13498 (N_13498,N_11952,N_11946);
xor U13499 (N_13499,N_10058,N_11632);
nor U13500 (N_13500,N_10778,N_11520);
xor U13501 (N_13501,N_10928,N_11293);
nor U13502 (N_13502,N_11304,N_11311);
nand U13503 (N_13503,N_11766,N_10190);
nor U13504 (N_13504,N_10579,N_11744);
and U13505 (N_13505,N_10340,N_10032);
nand U13506 (N_13506,N_11468,N_11346);
nand U13507 (N_13507,N_10833,N_11807);
nand U13508 (N_13508,N_10397,N_11536);
and U13509 (N_13509,N_11728,N_11021);
nand U13510 (N_13510,N_11088,N_11733);
and U13511 (N_13511,N_10920,N_11713);
or U13512 (N_13512,N_10421,N_11078);
and U13513 (N_13513,N_10128,N_10104);
xnor U13514 (N_13514,N_11350,N_10476);
or U13515 (N_13515,N_10600,N_11738);
nor U13516 (N_13516,N_10728,N_10347);
nand U13517 (N_13517,N_11479,N_11207);
xnor U13518 (N_13518,N_11513,N_11582);
nand U13519 (N_13519,N_10805,N_11158);
nor U13520 (N_13520,N_11993,N_10157);
and U13521 (N_13521,N_10984,N_10968);
xnor U13522 (N_13522,N_10403,N_11454);
nor U13523 (N_13523,N_11602,N_11564);
nor U13524 (N_13524,N_11121,N_11821);
and U13525 (N_13525,N_11347,N_10439);
nand U13526 (N_13526,N_10372,N_11011);
and U13527 (N_13527,N_10065,N_11877);
nand U13528 (N_13528,N_11224,N_11686);
or U13529 (N_13529,N_10211,N_11862);
nand U13530 (N_13530,N_11600,N_11780);
or U13531 (N_13531,N_10483,N_10771);
xnor U13532 (N_13532,N_10194,N_11192);
xor U13533 (N_13533,N_10199,N_10725);
nor U13534 (N_13534,N_11626,N_11020);
and U13535 (N_13535,N_10819,N_10479);
and U13536 (N_13536,N_10740,N_11854);
xor U13537 (N_13537,N_10491,N_10487);
and U13538 (N_13538,N_10003,N_11435);
nand U13539 (N_13539,N_11674,N_10823);
nor U13540 (N_13540,N_11542,N_10960);
or U13541 (N_13541,N_10743,N_10926);
and U13542 (N_13542,N_11394,N_10410);
nor U13543 (N_13543,N_11567,N_11351);
nor U13544 (N_13544,N_10459,N_10590);
nand U13545 (N_13545,N_10252,N_11608);
nor U13546 (N_13546,N_10028,N_11899);
and U13547 (N_13547,N_10950,N_11324);
or U13548 (N_13548,N_11611,N_10263);
and U13549 (N_13549,N_11116,N_11566);
nor U13550 (N_13550,N_11903,N_10089);
nor U13551 (N_13551,N_11297,N_11826);
and U13552 (N_13552,N_11776,N_11247);
nor U13553 (N_13553,N_11817,N_11765);
xnor U13554 (N_13554,N_10002,N_10495);
xor U13555 (N_13555,N_11524,N_11393);
nor U13556 (N_13556,N_10620,N_11902);
or U13557 (N_13557,N_10076,N_11225);
nor U13558 (N_13558,N_11318,N_11455);
and U13559 (N_13559,N_11196,N_11686);
nor U13560 (N_13560,N_10979,N_11784);
nand U13561 (N_13561,N_10507,N_10234);
or U13562 (N_13562,N_10981,N_11226);
nand U13563 (N_13563,N_11860,N_10238);
or U13564 (N_13564,N_10488,N_11502);
xor U13565 (N_13565,N_11692,N_10693);
nand U13566 (N_13566,N_10135,N_11578);
nand U13567 (N_13567,N_10079,N_10797);
nand U13568 (N_13568,N_11463,N_11771);
xor U13569 (N_13569,N_11489,N_10501);
nor U13570 (N_13570,N_10654,N_10483);
xnor U13571 (N_13571,N_11494,N_11964);
or U13572 (N_13572,N_11045,N_11047);
nor U13573 (N_13573,N_10963,N_10693);
nand U13574 (N_13574,N_11312,N_10656);
nor U13575 (N_13575,N_11095,N_11865);
nand U13576 (N_13576,N_11366,N_10375);
and U13577 (N_13577,N_11310,N_11199);
xor U13578 (N_13578,N_10068,N_11060);
nand U13579 (N_13579,N_11554,N_10176);
nor U13580 (N_13580,N_11948,N_10036);
nor U13581 (N_13581,N_11921,N_11901);
or U13582 (N_13582,N_11404,N_11622);
nand U13583 (N_13583,N_11293,N_10624);
nand U13584 (N_13584,N_10452,N_11965);
nand U13585 (N_13585,N_10986,N_10808);
or U13586 (N_13586,N_10747,N_11009);
xnor U13587 (N_13587,N_10119,N_11488);
nand U13588 (N_13588,N_10244,N_11858);
xor U13589 (N_13589,N_10064,N_11205);
xor U13590 (N_13590,N_10046,N_10337);
nor U13591 (N_13591,N_10645,N_10822);
xnor U13592 (N_13592,N_10842,N_11570);
nand U13593 (N_13593,N_10317,N_11801);
or U13594 (N_13594,N_10375,N_11181);
and U13595 (N_13595,N_10357,N_10407);
xor U13596 (N_13596,N_10365,N_10442);
and U13597 (N_13597,N_11305,N_10912);
xnor U13598 (N_13598,N_11048,N_10547);
and U13599 (N_13599,N_10085,N_11147);
or U13600 (N_13600,N_10138,N_10181);
nand U13601 (N_13601,N_11442,N_11617);
or U13602 (N_13602,N_11560,N_10222);
and U13603 (N_13603,N_11424,N_10344);
or U13604 (N_13604,N_11881,N_10862);
or U13605 (N_13605,N_11786,N_11051);
nand U13606 (N_13606,N_10898,N_10566);
xor U13607 (N_13607,N_11562,N_10151);
and U13608 (N_13608,N_10242,N_10813);
nand U13609 (N_13609,N_10274,N_10743);
nor U13610 (N_13610,N_11240,N_11503);
nand U13611 (N_13611,N_10630,N_11955);
and U13612 (N_13612,N_10239,N_11375);
xor U13613 (N_13613,N_11035,N_11843);
and U13614 (N_13614,N_10228,N_11073);
nor U13615 (N_13615,N_11571,N_10574);
nand U13616 (N_13616,N_11940,N_10261);
nor U13617 (N_13617,N_11607,N_10334);
xor U13618 (N_13618,N_11125,N_10173);
nor U13619 (N_13619,N_10278,N_10904);
nor U13620 (N_13620,N_11659,N_10417);
xor U13621 (N_13621,N_10599,N_11110);
and U13622 (N_13622,N_11020,N_10109);
and U13623 (N_13623,N_10871,N_11286);
or U13624 (N_13624,N_10824,N_10028);
or U13625 (N_13625,N_10597,N_10660);
xnor U13626 (N_13626,N_10196,N_11048);
nand U13627 (N_13627,N_10111,N_10423);
nor U13628 (N_13628,N_10551,N_11052);
nor U13629 (N_13629,N_10423,N_11378);
nand U13630 (N_13630,N_10247,N_11365);
or U13631 (N_13631,N_11279,N_11101);
nand U13632 (N_13632,N_11275,N_10349);
nand U13633 (N_13633,N_11021,N_11762);
xnor U13634 (N_13634,N_10004,N_10440);
and U13635 (N_13635,N_11924,N_10164);
xnor U13636 (N_13636,N_11670,N_11578);
or U13637 (N_13637,N_11002,N_10819);
or U13638 (N_13638,N_11964,N_10920);
xor U13639 (N_13639,N_11741,N_11833);
or U13640 (N_13640,N_11840,N_11335);
nand U13641 (N_13641,N_10749,N_10384);
nand U13642 (N_13642,N_11965,N_10555);
xnor U13643 (N_13643,N_11338,N_11320);
and U13644 (N_13644,N_11780,N_11888);
nor U13645 (N_13645,N_11752,N_11795);
xnor U13646 (N_13646,N_10167,N_10883);
xnor U13647 (N_13647,N_11936,N_10830);
xnor U13648 (N_13648,N_11301,N_10104);
nor U13649 (N_13649,N_11660,N_11772);
and U13650 (N_13650,N_10588,N_10145);
nand U13651 (N_13651,N_11639,N_10602);
or U13652 (N_13652,N_10271,N_11236);
or U13653 (N_13653,N_10735,N_10497);
and U13654 (N_13654,N_11188,N_10192);
nand U13655 (N_13655,N_11316,N_11200);
nor U13656 (N_13656,N_10755,N_11284);
nand U13657 (N_13657,N_10772,N_10954);
nor U13658 (N_13658,N_11205,N_10290);
and U13659 (N_13659,N_10330,N_11367);
xor U13660 (N_13660,N_10154,N_11985);
or U13661 (N_13661,N_11157,N_10801);
or U13662 (N_13662,N_10974,N_11362);
xor U13663 (N_13663,N_11538,N_10265);
or U13664 (N_13664,N_10085,N_11899);
nand U13665 (N_13665,N_10496,N_11804);
and U13666 (N_13666,N_11359,N_11008);
or U13667 (N_13667,N_11510,N_11562);
nand U13668 (N_13668,N_10724,N_11428);
or U13669 (N_13669,N_11806,N_10964);
and U13670 (N_13670,N_11882,N_10927);
or U13671 (N_13671,N_11216,N_10317);
nor U13672 (N_13672,N_10110,N_10381);
nor U13673 (N_13673,N_11816,N_10683);
nand U13674 (N_13674,N_10296,N_11684);
nand U13675 (N_13675,N_11744,N_11681);
xor U13676 (N_13676,N_10327,N_11746);
nand U13677 (N_13677,N_10061,N_11208);
or U13678 (N_13678,N_11679,N_11642);
xor U13679 (N_13679,N_11417,N_10140);
nor U13680 (N_13680,N_10327,N_11756);
xnor U13681 (N_13681,N_11512,N_10705);
nor U13682 (N_13682,N_11846,N_11774);
or U13683 (N_13683,N_11824,N_10779);
or U13684 (N_13684,N_10581,N_10966);
nor U13685 (N_13685,N_11370,N_10553);
xor U13686 (N_13686,N_10088,N_10483);
nor U13687 (N_13687,N_10997,N_10702);
or U13688 (N_13688,N_11272,N_11481);
xnor U13689 (N_13689,N_11644,N_11692);
nor U13690 (N_13690,N_11993,N_11177);
nand U13691 (N_13691,N_11270,N_11128);
and U13692 (N_13692,N_10852,N_11889);
or U13693 (N_13693,N_10059,N_10217);
or U13694 (N_13694,N_10615,N_11468);
and U13695 (N_13695,N_10625,N_10197);
nor U13696 (N_13696,N_11087,N_11131);
xor U13697 (N_13697,N_10169,N_10348);
xor U13698 (N_13698,N_10097,N_11193);
xnor U13699 (N_13699,N_10815,N_11276);
or U13700 (N_13700,N_10203,N_10374);
or U13701 (N_13701,N_11308,N_10015);
or U13702 (N_13702,N_10663,N_11952);
or U13703 (N_13703,N_10807,N_10988);
or U13704 (N_13704,N_10516,N_11107);
xnor U13705 (N_13705,N_10406,N_10881);
xnor U13706 (N_13706,N_11843,N_11648);
and U13707 (N_13707,N_10288,N_11974);
and U13708 (N_13708,N_11163,N_11049);
xnor U13709 (N_13709,N_11084,N_10548);
and U13710 (N_13710,N_11699,N_10501);
xnor U13711 (N_13711,N_10907,N_10215);
nor U13712 (N_13712,N_11768,N_11867);
xor U13713 (N_13713,N_10895,N_10084);
or U13714 (N_13714,N_11005,N_11398);
nand U13715 (N_13715,N_11271,N_11444);
nor U13716 (N_13716,N_10864,N_10628);
nor U13717 (N_13717,N_10715,N_11792);
or U13718 (N_13718,N_11914,N_10434);
nand U13719 (N_13719,N_11120,N_10864);
and U13720 (N_13720,N_11712,N_10861);
nand U13721 (N_13721,N_10504,N_11938);
nand U13722 (N_13722,N_10538,N_11699);
nor U13723 (N_13723,N_10916,N_11816);
and U13724 (N_13724,N_11357,N_10599);
nor U13725 (N_13725,N_11141,N_10665);
or U13726 (N_13726,N_11142,N_10502);
nand U13727 (N_13727,N_11204,N_11962);
and U13728 (N_13728,N_10343,N_11132);
nor U13729 (N_13729,N_11992,N_11970);
or U13730 (N_13730,N_10699,N_11686);
and U13731 (N_13731,N_11611,N_11982);
or U13732 (N_13732,N_10986,N_11548);
nand U13733 (N_13733,N_10350,N_10928);
nand U13734 (N_13734,N_10980,N_11634);
nand U13735 (N_13735,N_10219,N_11474);
nand U13736 (N_13736,N_10868,N_10377);
or U13737 (N_13737,N_11333,N_10359);
and U13738 (N_13738,N_10130,N_11514);
or U13739 (N_13739,N_11584,N_11168);
nand U13740 (N_13740,N_11138,N_10372);
nor U13741 (N_13741,N_11432,N_11163);
and U13742 (N_13742,N_10740,N_10519);
xnor U13743 (N_13743,N_10064,N_10748);
xnor U13744 (N_13744,N_11951,N_11606);
nor U13745 (N_13745,N_11985,N_11446);
xor U13746 (N_13746,N_10741,N_10203);
or U13747 (N_13747,N_10365,N_10696);
nand U13748 (N_13748,N_10681,N_11719);
and U13749 (N_13749,N_10429,N_11732);
nand U13750 (N_13750,N_11867,N_11656);
or U13751 (N_13751,N_10206,N_10180);
nand U13752 (N_13752,N_11848,N_11126);
and U13753 (N_13753,N_10448,N_10178);
or U13754 (N_13754,N_11658,N_10002);
nor U13755 (N_13755,N_10393,N_11498);
or U13756 (N_13756,N_10514,N_10143);
or U13757 (N_13757,N_11972,N_11909);
or U13758 (N_13758,N_11129,N_11176);
and U13759 (N_13759,N_11188,N_10457);
nor U13760 (N_13760,N_11992,N_10332);
and U13761 (N_13761,N_10593,N_11468);
nor U13762 (N_13762,N_11012,N_11746);
and U13763 (N_13763,N_10417,N_10685);
xnor U13764 (N_13764,N_11888,N_10054);
nor U13765 (N_13765,N_11899,N_11307);
nor U13766 (N_13766,N_10181,N_11952);
nor U13767 (N_13767,N_10848,N_11645);
and U13768 (N_13768,N_10341,N_11271);
or U13769 (N_13769,N_10892,N_11271);
nor U13770 (N_13770,N_11637,N_11749);
nand U13771 (N_13771,N_11665,N_10901);
xor U13772 (N_13772,N_10727,N_10584);
nand U13773 (N_13773,N_11303,N_11935);
and U13774 (N_13774,N_10238,N_10740);
nand U13775 (N_13775,N_10692,N_10153);
xnor U13776 (N_13776,N_10195,N_10677);
xnor U13777 (N_13777,N_11708,N_10979);
xor U13778 (N_13778,N_10001,N_10886);
or U13779 (N_13779,N_10916,N_11564);
nand U13780 (N_13780,N_11584,N_10207);
nor U13781 (N_13781,N_11883,N_11301);
xnor U13782 (N_13782,N_10109,N_11700);
or U13783 (N_13783,N_10336,N_11904);
nand U13784 (N_13784,N_10059,N_10671);
nor U13785 (N_13785,N_10702,N_11846);
or U13786 (N_13786,N_11353,N_11973);
nor U13787 (N_13787,N_10922,N_10492);
nand U13788 (N_13788,N_11072,N_10799);
or U13789 (N_13789,N_11657,N_11409);
or U13790 (N_13790,N_11823,N_10877);
or U13791 (N_13791,N_11879,N_11841);
nand U13792 (N_13792,N_11829,N_10687);
nand U13793 (N_13793,N_11211,N_10888);
nand U13794 (N_13794,N_10709,N_11653);
and U13795 (N_13795,N_10245,N_11532);
nand U13796 (N_13796,N_11646,N_10024);
or U13797 (N_13797,N_11843,N_10740);
or U13798 (N_13798,N_11661,N_10838);
nand U13799 (N_13799,N_10952,N_11719);
xor U13800 (N_13800,N_10172,N_10562);
xor U13801 (N_13801,N_10601,N_11640);
nor U13802 (N_13802,N_11513,N_10062);
and U13803 (N_13803,N_11602,N_10897);
or U13804 (N_13804,N_10258,N_11252);
nor U13805 (N_13805,N_11011,N_10972);
nor U13806 (N_13806,N_10671,N_11354);
and U13807 (N_13807,N_11171,N_10082);
or U13808 (N_13808,N_11513,N_10326);
or U13809 (N_13809,N_10624,N_10841);
nor U13810 (N_13810,N_10949,N_10111);
nor U13811 (N_13811,N_11305,N_11432);
xor U13812 (N_13812,N_11756,N_10798);
xnor U13813 (N_13813,N_10252,N_11623);
and U13814 (N_13814,N_10977,N_11902);
and U13815 (N_13815,N_10794,N_11070);
xor U13816 (N_13816,N_11158,N_11866);
or U13817 (N_13817,N_10071,N_10932);
and U13818 (N_13818,N_11489,N_11087);
nand U13819 (N_13819,N_11199,N_11392);
nor U13820 (N_13820,N_11642,N_11097);
nor U13821 (N_13821,N_11496,N_10846);
and U13822 (N_13822,N_10969,N_11617);
and U13823 (N_13823,N_10349,N_11655);
nand U13824 (N_13824,N_11717,N_11961);
and U13825 (N_13825,N_10435,N_10294);
nor U13826 (N_13826,N_10649,N_10619);
nor U13827 (N_13827,N_11906,N_10765);
or U13828 (N_13828,N_10874,N_10744);
and U13829 (N_13829,N_11130,N_11987);
or U13830 (N_13830,N_11500,N_10152);
and U13831 (N_13831,N_11069,N_11818);
nor U13832 (N_13832,N_10173,N_11192);
xor U13833 (N_13833,N_11226,N_10033);
and U13834 (N_13834,N_11815,N_11835);
nor U13835 (N_13835,N_10950,N_11311);
xnor U13836 (N_13836,N_10444,N_10994);
or U13837 (N_13837,N_10001,N_10504);
and U13838 (N_13838,N_11393,N_10847);
or U13839 (N_13839,N_10832,N_11139);
nor U13840 (N_13840,N_10140,N_11618);
xor U13841 (N_13841,N_10867,N_11898);
nand U13842 (N_13842,N_10180,N_11711);
or U13843 (N_13843,N_11464,N_10881);
and U13844 (N_13844,N_10522,N_10706);
and U13845 (N_13845,N_11127,N_11756);
nand U13846 (N_13846,N_11710,N_10309);
nand U13847 (N_13847,N_10886,N_11753);
or U13848 (N_13848,N_11386,N_11687);
nand U13849 (N_13849,N_11468,N_11811);
nand U13850 (N_13850,N_10268,N_11320);
or U13851 (N_13851,N_10877,N_10904);
or U13852 (N_13852,N_10101,N_11635);
xor U13853 (N_13853,N_11654,N_11709);
xnor U13854 (N_13854,N_10440,N_11401);
and U13855 (N_13855,N_11076,N_10520);
nand U13856 (N_13856,N_10969,N_11416);
xor U13857 (N_13857,N_11715,N_10036);
nor U13858 (N_13858,N_11567,N_10856);
nand U13859 (N_13859,N_11824,N_11684);
nand U13860 (N_13860,N_10404,N_11044);
xnor U13861 (N_13861,N_11305,N_10019);
or U13862 (N_13862,N_10972,N_10683);
nor U13863 (N_13863,N_10010,N_10466);
nand U13864 (N_13864,N_10662,N_11601);
nand U13865 (N_13865,N_11321,N_10469);
xnor U13866 (N_13866,N_11347,N_10893);
nand U13867 (N_13867,N_11645,N_10069);
nand U13868 (N_13868,N_10382,N_10423);
or U13869 (N_13869,N_10221,N_11501);
and U13870 (N_13870,N_10104,N_11392);
xor U13871 (N_13871,N_11272,N_10436);
or U13872 (N_13872,N_11877,N_11210);
xnor U13873 (N_13873,N_11113,N_10998);
nor U13874 (N_13874,N_10575,N_11603);
nor U13875 (N_13875,N_11881,N_10008);
nor U13876 (N_13876,N_11024,N_10656);
nor U13877 (N_13877,N_10636,N_11767);
and U13878 (N_13878,N_10042,N_10488);
and U13879 (N_13879,N_10336,N_11879);
nand U13880 (N_13880,N_10208,N_11715);
or U13881 (N_13881,N_10210,N_11988);
and U13882 (N_13882,N_11948,N_11837);
or U13883 (N_13883,N_11373,N_10702);
nor U13884 (N_13884,N_11759,N_10299);
and U13885 (N_13885,N_11619,N_11940);
nand U13886 (N_13886,N_11893,N_10901);
and U13887 (N_13887,N_10929,N_11673);
or U13888 (N_13888,N_11997,N_11133);
nor U13889 (N_13889,N_11649,N_10638);
or U13890 (N_13890,N_11920,N_10221);
and U13891 (N_13891,N_11333,N_11661);
or U13892 (N_13892,N_10735,N_10464);
nand U13893 (N_13893,N_10510,N_10322);
and U13894 (N_13894,N_10182,N_11701);
nand U13895 (N_13895,N_11154,N_10814);
xnor U13896 (N_13896,N_10573,N_10947);
and U13897 (N_13897,N_10662,N_10188);
or U13898 (N_13898,N_10393,N_11074);
nor U13899 (N_13899,N_11719,N_10137);
or U13900 (N_13900,N_11231,N_11887);
xnor U13901 (N_13901,N_10237,N_10872);
xnor U13902 (N_13902,N_11288,N_11149);
xnor U13903 (N_13903,N_11865,N_11743);
nor U13904 (N_13904,N_10346,N_10975);
and U13905 (N_13905,N_11891,N_11537);
and U13906 (N_13906,N_11224,N_11296);
nand U13907 (N_13907,N_10588,N_10976);
or U13908 (N_13908,N_10214,N_11899);
or U13909 (N_13909,N_10402,N_11775);
and U13910 (N_13910,N_10890,N_10633);
or U13911 (N_13911,N_10289,N_10458);
or U13912 (N_13912,N_10437,N_11707);
nand U13913 (N_13913,N_10273,N_11116);
nor U13914 (N_13914,N_11965,N_11052);
or U13915 (N_13915,N_10257,N_11995);
nor U13916 (N_13916,N_11661,N_10322);
xor U13917 (N_13917,N_10000,N_11034);
nand U13918 (N_13918,N_11330,N_11950);
xnor U13919 (N_13919,N_11575,N_11158);
or U13920 (N_13920,N_10470,N_10271);
and U13921 (N_13921,N_11736,N_10723);
nand U13922 (N_13922,N_11150,N_11739);
and U13923 (N_13923,N_10536,N_11271);
xnor U13924 (N_13924,N_11247,N_10427);
or U13925 (N_13925,N_10548,N_10077);
or U13926 (N_13926,N_11626,N_11393);
xnor U13927 (N_13927,N_10749,N_11866);
xor U13928 (N_13928,N_10570,N_10266);
or U13929 (N_13929,N_11016,N_11283);
and U13930 (N_13930,N_11385,N_11019);
and U13931 (N_13931,N_10567,N_10896);
xnor U13932 (N_13932,N_10349,N_11916);
and U13933 (N_13933,N_10481,N_10021);
nor U13934 (N_13934,N_11494,N_11882);
nor U13935 (N_13935,N_10481,N_10823);
nand U13936 (N_13936,N_10166,N_11308);
xor U13937 (N_13937,N_11196,N_10838);
xor U13938 (N_13938,N_10592,N_11417);
nor U13939 (N_13939,N_11430,N_11154);
or U13940 (N_13940,N_11085,N_10686);
nand U13941 (N_13941,N_11446,N_11079);
nand U13942 (N_13942,N_11267,N_10144);
or U13943 (N_13943,N_11160,N_10811);
or U13944 (N_13944,N_10188,N_11557);
nor U13945 (N_13945,N_11756,N_11371);
and U13946 (N_13946,N_10426,N_11047);
nand U13947 (N_13947,N_11260,N_10444);
nor U13948 (N_13948,N_10703,N_10072);
nor U13949 (N_13949,N_10988,N_11421);
nor U13950 (N_13950,N_10358,N_11596);
nand U13951 (N_13951,N_10796,N_10575);
or U13952 (N_13952,N_11041,N_11023);
and U13953 (N_13953,N_10746,N_11666);
nor U13954 (N_13954,N_11082,N_10879);
nor U13955 (N_13955,N_10205,N_10086);
nor U13956 (N_13956,N_11202,N_10234);
and U13957 (N_13957,N_10548,N_10326);
or U13958 (N_13958,N_10158,N_10950);
nand U13959 (N_13959,N_10616,N_10119);
or U13960 (N_13960,N_11131,N_10302);
nor U13961 (N_13961,N_11391,N_11401);
xor U13962 (N_13962,N_10473,N_11705);
nand U13963 (N_13963,N_11124,N_10396);
or U13964 (N_13964,N_11973,N_11214);
nand U13965 (N_13965,N_10766,N_10452);
xor U13966 (N_13966,N_10464,N_10064);
or U13967 (N_13967,N_10785,N_11075);
and U13968 (N_13968,N_11740,N_11042);
and U13969 (N_13969,N_10641,N_11005);
or U13970 (N_13970,N_10276,N_11767);
nand U13971 (N_13971,N_11522,N_10715);
and U13972 (N_13972,N_11643,N_10381);
nor U13973 (N_13973,N_11533,N_10078);
and U13974 (N_13974,N_10143,N_11234);
xor U13975 (N_13975,N_11288,N_10950);
and U13976 (N_13976,N_11386,N_10004);
and U13977 (N_13977,N_10151,N_10261);
nand U13978 (N_13978,N_11654,N_11129);
xor U13979 (N_13979,N_11505,N_10307);
nand U13980 (N_13980,N_11020,N_10942);
or U13981 (N_13981,N_11377,N_11326);
nand U13982 (N_13982,N_11764,N_11903);
or U13983 (N_13983,N_10007,N_11079);
xnor U13984 (N_13984,N_10315,N_11938);
nor U13985 (N_13985,N_10093,N_10440);
and U13986 (N_13986,N_10485,N_11852);
and U13987 (N_13987,N_11202,N_11847);
or U13988 (N_13988,N_11624,N_10132);
nand U13989 (N_13989,N_10796,N_10211);
nand U13990 (N_13990,N_11925,N_10931);
and U13991 (N_13991,N_11854,N_10515);
or U13992 (N_13992,N_10994,N_11072);
xor U13993 (N_13993,N_11610,N_10138);
and U13994 (N_13994,N_11641,N_10024);
nor U13995 (N_13995,N_11205,N_11925);
nor U13996 (N_13996,N_11517,N_11037);
and U13997 (N_13997,N_11371,N_11613);
xor U13998 (N_13998,N_11245,N_10905);
or U13999 (N_13999,N_11655,N_10678);
xor U14000 (N_14000,N_12343,N_12227);
or U14001 (N_14001,N_12741,N_13288);
nor U14002 (N_14002,N_12915,N_12099);
nor U14003 (N_14003,N_12554,N_13159);
xnor U14004 (N_14004,N_13353,N_12053);
nand U14005 (N_14005,N_13139,N_12941);
nor U14006 (N_14006,N_12972,N_13201);
and U14007 (N_14007,N_13213,N_12035);
nor U14008 (N_14008,N_12073,N_13348);
nand U14009 (N_14009,N_13758,N_12120);
nand U14010 (N_14010,N_13927,N_12057);
xor U14011 (N_14011,N_12874,N_12883);
and U14012 (N_14012,N_12397,N_12748);
and U14013 (N_14013,N_12720,N_13311);
and U14014 (N_14014,N_12802,N_12846);
and U14015 (N_14015,N_12785,N_13218);
nand U14016 (N_14016,N_13732,N_13893);
and U14017 (N_14017,N_12418,N_12641);
nand U14018 (N_14018,N_12970,N_13250);
nand U14019 (N_14019,N_13793,N_12012);
nand U14020 (N_14020,N_12228,N_13798);
nor U14021 (N_14021,N_13546,N_13053);
or U14022 (N_14022,N_12632,N_12516);
xor U14023 (N_14023,N_13601,N_13235);
xnor U14024 (N_14024,N_12047,N_13572);
nand U14025 (N_14025,N_12617,N_13292);
nand U14026 (N_14026,N_12364,N_12833);
nor U14027 (N_14027,N_13778,N_13521);
nor U14028 (N_14028,N_13960,N_12649);
nand U14029 (N_14029,N_12929,N_12960);
xor U14030 (N_14030,N_12985,N_13228);
xnor U14031 (N_14031,N_12181,N_12147);
or U14032 (N_14032,N_12605,N_12962);
nor U14033 (N_14033,N_13285,N_13144);
and U14034 (N_14034,N_12310,N_12019);
nor U14035 (N_14035,N_12030,N_13796);
nor U14036 (N_14036,N_13323,N_12913);
and U14037 (N_14037,N_12443,N_13882);
nand U14038 (N_14038,N_13909,N_12995);
and U14039 (N_14039,N_12560,N_12008);
nand U14040 (N_14040,N_12010,N_12188);
nand U14041 (N_14041,N_13907,N_12623);
or U14042 (N_14042,N_12897,N_13189);
and U14043 (N_14043,N_12451,N_12644);
and U14044 (N_14044,N_12286,N_13522);
xnor U14045 (N_14045,N_13097,N_13983);
xnor U14046 (N_14046,N_13341,N_12569);
nand U14047 (N_14047,N_12432,N_12570);
and U14048 (N_14048,N_12378,N_12412);
or U14049 (N_14049,N_12584,N_12021);
or U14050 (N_14050,N_13004,N_13608);
and U14051 (N_14051,N_12187,N_13272);
xnor U14052 (N_14052,N_12629,N_13221);
and U14053 (N_14053,N_12555,N_12730);
xnor U14054 (N_14054,N_12202,N_12052);
and U14055 (N_14055,N_13722,N_13185);
or U14056 (N_14056,N_12164,N_12182);
nand U14057 (N_14057,N_13008,N_13889);
nor U14058 (N_14058,N_13901,N_13950);
nand U14059 (N_14059,N_13503,N_12337);
nor U14060 (N_14060,N_13112,N_13611);
nand U14061 (N_14061,N_13880,N_13985);
or U14062 (N_14062,N_13484,N_12018);
nor U14063 (N_14063,N_12464,N_13707);
nor U14064 (N_14064,N_12705,N_12184);
xnor U14065 (N_14065,N_12390,N_13931);
nor U14066 (N_14066,N_13766,N_13324);
xnor U14067 (N_14067,N_13036,N_13895);
nand U14068 (N_14068,N_12075,N_12868);
nand U14069 (N_14069,N_12621,N_13647);
and U14070 (N_14070,N_13455,N_12814);
nor U14071 (N_14071,N_13307,N_13493);
xor U14072 (N_14072,N_12321,N_12471);
xor U14073 (N_14073,N_12449,N_13232);
nor U14074 (N_14074,N_13795,N_13850);
xor U14075 (N_14075,N_13849,N_13634);
and U14076 (N_14076,N_13073,N_12331);
nand U14077 (N_14077,N_13343,N_13171);
nand U14078 (N_14078,N_13859,N_12093);
and U14079 (N_14079,N_13309,N_12658);
and U14080 (N_14080,N_13587,N_12266);
or U14081 (N_14081,N_12582,N_13439);
and U14082 (N_14082,N_12664,N_12747);
and U14083 (N_14083,N_13891,N_13765);
nor U14084 (N_14084,N_12681,N_12152);
nand U14085 (N_14085,N_13266,N_12521);
nand U14086 (N_14086,N_13822,N_12971);
xnor U14087 (N_14087,N_12279,N_12540);
or U14088 (N_14088,N_12460,N_13061);
and U14089 (N_14089,N_13701,N_12701);
nor U14090 (N_14090,N_12514,N_12739);
nand U14091 (N_14091,N_12771,N_13888);
and U14092 (N_14092,N_13590,N_12637);
xor U14093 (N_14093,N_12952,N_13517);
nand U14094 (N_14094,N_12190,N_13468);
or U14095 (N_14095,N_12282,N_13957);
nor U14096 (N_14096,N_13267,N_13500);
or U14097 (N_14097,N_13453,N_12657);
nand U14098 (N_14098,N_13858,N_13204);
nor U14099 (N_14099,N_13083,N_13033);
nor U14100 (N_14100,N_12209,N_13496);
and U14101 (N_14101,N_13440,N_13801);
xor U14102 (N_14102,N_13562,N_12502);
and U14103 (N_14103,N_13072,N_13642);
or U14104 (N_14104,N_12326,N_13052);
and U14105 (N_14105,N_12945,N_13188);
xor U14106 (N_14106,N_12625,N_12411);
nor U14107 (N_14107,N_13238,N_12236);
xnor U14108 (N_14108,N_12065,N_12595);
or U14109 (N_14109,N_12261,N_13620);
xor U14110 (N_14110,N_12684,N_13833);
nor U14111 (N_14111,N_13239,N_12303);
or U14112 (N_14112,N_13205,N_12238);
nand U14113 (N_14113,N_13812,N_13320);
nor U14114 (N_14114,N_13436,N_13691);
nor U14115 (N_14115,N_12288,N_12284);
or U14116 (N_14116,N_13283,N_13720);
xor U14117 (N_14117,N_12043,N_13193);
nand U14118 (N_14118,N_12153,N_13945);
nand U14119 (N_14119,N_12338,N_13943);
xor U14120 (N_14120,N_13593,N_12342);
nor U14121 (N_14121,N_12636,N_12148);
nor U14122 (N_14122,N_12702,N_13099);
nand U14123 (N_14123,N_12054,N_13698);
or U14124 (N_14124,N_13750,N_12685);
and U14125 (N_14125,N_13915,N_12185);
and U14126 (N_14126,N_12507,N_12653);
and U14127 (N_14127,N_13686,N_13489);
xor U14128 (N_14128,N_13437,N_13016);
xnor U14129 (N_14129,N_13695,N_13531);
and U14130 (N_14130,N_13013,N_13081);
nand U14131 (N_14131,N_13740,N_13080);
nor U14132 (N_14132,N_13044,N_13234);
nand U14133 (N_14133,N_13923,N_13295);
or U14134 (N_14134,N_12927,N_13119);
or U14135 (N_14135,N_13474,N_12103);
or U14136 (N_14136,N_12956,N_12999);
nand U14137 (N_14137,N_13363,N_12839);
xnor U14138 (N_14138,N_12254,N_13598);
and U14139 (N_14139,N_12575,N_12643);
or U14140 (N_14140,N_13856,N_13871);
or U14141 (N_14141,N_12132,N_13490);
xor U14142 (N_14142,N_13303,N_13336);
xor U14143 (N_14143,N_13526,N_13946);
or U14144 (N_14144,N_12170,N_13739);
or U14145 (N_14145,N_12580,N_13212);
nand U14146 (N_14146,N_12843,N_13567);
nor U14147 (N_14147,N_12368,N_13196);
nand U14148 (N_14148,N_12611,N_12167);
xnor U14149 (N_14149,N_12224,N_13499);
or U14150 (N_14150,N_12698,N_12647);
and U14151 (N_14151,N_13675,N_13625);
xnor U14152 (N_14152,N_13141,N_13865);
nand U14153 (N_14153,N_12352,N_13709);
or U14154 (N_14154,N_13971,N_12886);
and U14155 (N_14155,N_13254,N_13300);
or U14156 (N_14156,N_13605,N_13580);
or U14157 (N_14157,N_13784,N_13289);
nand U14158 (N_14158,N_12026,N_12417);
or U14159 (N_14159,N_12781,N_12078);
xnor U14160 (N_14160,N_13592,N_13211);
and U14161 (N_14161,N_12854,N_13098);
nand U14162 (N_14162,N_13414,N_13892);
nor U14163 (N_14163,N_12646,N_12004);
nor U14164 (N_14164,N_12572,N_13617);
or U14165 (N_14165,N_13225,N_12955);
and U14166 (N_14166,N_13970,N_12539);
and U14167 (N_14167,N_12299,N_13138);
or U14168 (N_14168,N_12574,N_13821);
nor U14169 (N_14169,N_12718,N_13578);
nor U14170 (N_14170,N_12434,N_12322);
nor U14171 (N_14171,N_12003,N_12244);
and U14172 (N_14172,N_12064,N_12353);
and U14173 (N_14173,N_13006,N_13077);
nand U14174 (N_14174,N_13207,N_13905);
and U14175 (N_14175,N_13543,N_13071);
and U14176 (N_14176,N_12461,N_12892);
and U14177 (N_14177,N_13120,N_13480);
or U14178 (N_14178,N_13021,N_13153);
nand U14179 (N_14179,N_12553,N_13354);
nor U14180 (N_14180,N_13248,N_13019);
xor U14181 (N_14181,N_12424,N_12069);
nor U14182 (N_14182,N_12376,N_12504);
xor U14183 (N_14183,N_12174,N_13506);
nor U14184 (N_14184,N_12896,N_12682);
nand U14185 (N_14185,N_13262,N_13017);
xnor U14186 (N_14186,N_13824,N_12964);
and U14187 (N_14187,N_12158,N_12013);
nor U14188 (N_14188,N_12585,N_13461);
nor U14189 (N_14189,N_13242,N_12109);
xor U14190 (N_14190,N_12752,N_12440);
or U14191 (N_14191,N_13552,N_13948);
or U14192 (N_14192,N_13007,N_13651);
nor U14193 (N_14193,N_13803,N_13229);
nor U14194 (N_14194,N_12976,N_13210);
xor U14195 (N_14195,N_12577,N_12719);
and U14196 (N_14196,N_12478,N_12648);
and U14197 (N_14197,N_12058,N_12690);
nor U14198 (N_14198,N_12932,N_13975);
or U14199 (N_14199,N_12051,N_13917);
xor U14200 (N_14200,N_13419,N_12459);
or U14201 (N_14201,N_12361,N_12815);
and U14202 (N_14202,N_12216,N_12499);
nor U14203 (N_14203,N_13163,N_13752);
nand U14204 (N_14204,N_13676,N_13402);
xor U14205 (N_14205,N_13743,N_13847);
nor U14206 (N_14206,N_12757,N_12373);
or U14207 (N_14207,N_12393,N_12127);
nand U14208 (N_14208,N_13902,N_13060);
nor U14209 (N_14209,N_13733,N_12317);
xor U14210 (N_14210,N_13403,N_13757);
and U14211 (N_14211,N_13249,N_12490);
and U14212 (N_14212,N_12769,N_13866);
and U14213 (N_14213,N_13360,N_13559);
nand U14214 (N_14214,N_13337,N_12339);
nand U14215 (N_14215,N_13881,N_13938);
and U14216 (N_14216,N_13906,N_12211);
and U14217 (N_14217,N_13922,N_12340);
nor U14218 (N_14218,N_13633,N_13184);
and U14219 (N_14219,N_12234,N_13529);
xnor U14220 (N_14220,N_12509,N_12172);
and U14221 (N_14221,N_12660,N_12257);
xor U14222 (N_14222,N_13683,N_13125);
nor U14223 (N_14223,N_12674,N_13084);
nand U14224 (N_14224,N_12845,N_12294);
or U14225 (N_14225,N_13934,N_12639);
nor U14226 (N_14226,N_13181,N_13152);
or U14227 (N_14227,N_12655,N_12865);
xor U14228 (N_14228,N_12931,N_13622);
nor U14229 (N_14229,N_13199,N_12667);
xor U14230 (N_14230,N_13227,N_12409);
nand U14231 (N_14231,N_13776,N_12037);
or U14232 (N_14232,N_12709,N_12670);
nor U14233 (N_14233,N_12413,N_12953);
and U14234 (N_14234,N_13400,N_12711);
nand U14235 (N_14235,N_13838,N_13668);
nand U14236 (N_14236,N_12259,N_13510);
xnor U14237 (N_14237,N_13714,N_13308);
nor U14238 (N_14238,N_13845,N_12716);
xnor U14239 (N_14239,N_12028,N_13420);
or U14240 (N_14240,N_13550,N_13515);
nand U14241 (N_14241,N_12818,N_13771);
xor U14242 (N_14242,N_12036,N_12903);
xnor U14243 (N_14243,N_12697,N_12095);
xor U14244 (N_14244,N_12797,N_12163);
nand U14245 (N_14245,N_13870,N_12768);
nand U14246 (N_14246,N_13460,N_12899);
nor U14247 (N_14247,N_13672,N_13756);
nor U14248 (N_14248,N_13466,N_12488);
nand U14249 (N_14249,N_12689,N_12056);
or U14250 (N_14250,N_13217,N_12094);
and U14251 (N_14251,N_13802,N_12810);
nand U14252 (N_14252,N_13101,N_13685);
nand U14253 (N_14253,N_12816,N_12363);
and U14254 (N_14254,N_12830,N_12793);
and U14255 (N_14255,N_12477,N_13327);
or U14256 (N_14256,N_13987,N_12300);
xnor U14257 (N_14257,N_12407,N_12497);
and U14258 (N_14258,N_13694,N_12602);
xnor U14259 (N_14259,N_12842,N_13155);
nor U14260 (N_14260,N_12848,N_13147);
xnor U14261 (N_14261,N_13222,N_13753);
xor U14262 (N_14262,N_12077,N_13240);
and U14263 (N_14263,N_13724,N_12622);
nor U14264 (N_14264,N_12751,N_13376);
or U14265 (N_14265,N_12517,N_13407);
nor U14266 (N_14266,N_12450,N_13245);
nor U14267 (N_14267,N_12136,N_13048);
nor U14268 (N_14268,N_12744,N_13602);
and U14269 (N_14269,N_12811,N_12391);
and U14270 (N_14270,N_13162,N_12954);
or U14271 (N_14271,N_12694,N_13998);
xnor U14272 (N_14272,N_12448,N_12386);
nor U14273 (N_14273,N_13322,N_12676);
or U14274 (N_14274,N_12776,N_13842);
xor U14275 (N_14275,N_13145,N_12360);
or U14276 (N_14276,N_13257,N_12023);
xnor U14277 (N_14277,N_13825,N_13887);
nor U14278 (N_14278,N_12834,N_13105);
or U14279 (N_14279,N_13610,N_12594);
or U14280 (N_14280,N_13716,N_12963);
xnor U14281 (N_14281,N_13638,N_13131);
nand U14282 (N_14282,N_12290,N_12958);
nand U14283 (N_14283,N_13172,N_13467);
nand U14284 (N_14284,N_13456,N_12472);
nand U14285 (N_14285,N_12015,N_13367);
xor U14286 (N_14286,N_13346,N_13606);
or U14287 (N_14287,N_12453,N_13596);
xnor U14288 (N_14288,N_13462,N_13342);
xor U14289 (N_14289,N_13860,N_12197);
nor U14290 (N_14290,N_13956,N_13664);
and U14291 (N_14291,N_12923,N_12989);
xnor U14292 (N_14292,N_13852,N_12792);
xnor U14293 (N_14293,N_13565,N_12910);
xor U14294 (N_14294,N_13713,N_13165);
nor U14295 (N_14295,N_12729,N_13657);
or U14296 (N_14296,N_13444,N_12157);
nor U14297 (N_14297,N_12520,N_13412);
nor U14298 (N_14298,N_13113,N_12559);
and U14299 (N_14299,N_13696,N_13644);
xnor U14300 (N_14300,N_13382,N_13140);
or U14301 (N_14301,N_12366,N_13059);
and U14302 (N_14302,N_12947,N_12587);
nand U14303 (N_14303,N_13573,N_13555);
xor U14304 (N_14304,N_12176,N_13667);
and U14305 (N_14305,N_12548,N_12505);
nand U14306 (N_14306,N_12777,N_12341);
and U14307 (N_14307,N_13237,N_13769);
or U14308 (N_14308,N_12873,N_13886);
nand U14309 (N_14309,N_13800,N_12154);
or U14310 (N_14310,N_12269,N_13949);
or U14311 (N_14311,N_12600,N_13779);
or U14312 (N_14312,N_13645,N_12467);
or U14313 (N_14313,N_12351,N_12966);
or U14314 (N_14314,N_12610,N_12083);
nand U14315 (N_14315,N_13215,N_13107);
or U14316 (N_14316,N_13994,N_13198);
nand U14317 (N_14317,N_12260,N_13340);
and U14318 (N_14318,N_13111,N_12313);
and U14319 (N_14319,N_12809,N_13941);
nand U14320 (N_14320,N_12765,N_12276);
nand U14321 (N_14321,N_13754,N_13973);
nor U14322 (N_14322,N_12060,N_12822);
or U14323 (N_14323,N_13995,N_12404);
xnor U14324 (N_14324,N_12885,N_12597);
nor U14325 (N_14325,N_13326,N_12606);
nand U14326 (N_14326,N_12129,N_13532);
or U14327 (N_14327,N_12346,N_13330);
or U14328 (N_14328,N_13169,N_13999);
and U14329 (N_14329,N_13160,N_12663);
xor U14330 (N_14330,N_12289,N_13093);
or U14331 (N_14331,N_13557,N_12905);
or U14332 (N_14332,N_13604,N_13851);
nand U14333 (N_14333,N_13966,N_13132);
nand U14334 (N_14334,N_12370,N_13434);
nand U14335 (N_14335,N_13361,N_13536);
and U14336 (N_14336,N_13737,N_13030);
xnor U14337 (N_14337,N_13810,N_12344);
xor U14338 (N_14338,N_13066,N_12151);
nor U14339 (N_14339,N_13435,N_12389);
xor U14340 (N_14340,N_13829,N_12220);
nand U14341 (N_14341,N_12588,N_12609);
nand U14342 (N_14342,N_12925,N_13524);
xnor U14343 (N_14343,N_13780,N_13942);
nor U14344 (N_14344,N_12237,N_13314);
xor U14345 (N_14345,N_13380,N_13054);
xnor U14346 (N_14346,N_13231,N_13561);
nand U14347 (N_14347,N_12975,N_13261);
xnor U14348 (N_14348,N_12480,N_12482);
or U14349 (N_14349,N_13002,N_13725);
nor U14350 (N_14350,N_12889,N_12466);
and U14351 (N_14351,N_13287,N_12433);
nand U14352 (N_14352,N_13398,N_13772);
nor U14353 (N_14353,N_13449,N_13318);
nand U14354 (N_14354,N_13424,N_12495);
and U14355 (N_14355,N_13377,N_13595);
and U14356 (N_14356,N_13986,N_12543);
nand U14357 (N_14357,N_12055,N_12025);
and U14358 (N_14358,N_13589,N_13355);
and U14359 (N_14359,N_13932,N_12193);
xnor U14360 (N_14360,N_12435,N_13495);
nand U14361 (N_14361,N_13386,N_12596);
and U14362 (N_14362,N_12076,N_13432);
nand U14363 (N_14363,N_12252,N_12746);
nand U14364 (N_14364,N_12071,N_13661);
or U14365 (N_14365,N_12579,N_12961);
and U14366 (N_14366,N_13274,N_13627);
and U14367 (N_14367,N_13178,N_13834);
and U14368 (N_14368,N_13264,N_12959);
or U14369 (N_14369,N_12473,N_12369);
nand U14370 (N_14370,N_13777,N_13259);
nand U14371 (N_14371,N_12142,N_13936);
or U14372 (N_14372,N_12319,N_13418);
nand U14373 (N_14373,N_12911,N_13206);
or U14374 (N_14374,N_13290,N_13840);
nand U14375 (N_14375,N_12463,N_12535);
or U14376 (N_14376,N_12624,N_12108);
xnor U14377 (N_14377,N_12562,N_12233);
xnor U14378 (N_14378,N_12264,N_13678);
xor U14379 (N_14379,N_12908,N_13304);
xnor U14380 (N_14380,N_12307,N_13136);
xor U14381 (N_14381,N_12620,N_12855);
nor U14382 (N_14382,N_12715,N_12862);
nor U14383 (N_14383,N_12997,N_12662);
nor U14384 (N_14384,N_13397,N_13142);
nor U14385 (N_14385,N_12032,N_12919);
nand U14386 (N_14386,N_13547,N_13747);
nand U14387 (N_14387,N_12223,N_13183);
nand U14388 (N_14388,N_13626,N_12526);
nor U14389 (N_14389,N_12029,N_12101);
xnor U14390 (N_14390,N_12468,N_13738);
and U14391 (N_14391,N_12280,N_13646);
xor U14392 (N_14392,N_13051,N_13884);
or U14393 (N_14393,N_12766,N_13862);
and U14394 (N_14394,N_12978,N_12949);
or U14395 (N_14395,N_13214,N_12330);
nand U14396 (N_14396,N_12248,N_13997);
or U14397 (N_14397,N_13269,N_13003);
nor U14398 (N_14398,N_12189,N_13996);
nor U14399 (N_14399,N_12727,N_13293);
and U14400 (N_14400,N_13670,N_13122);
nand U14401 (N_14401,N_13538,N_13182);
nor U14402 (N_14402,N_12375,N_13746);
or U14403 (N_14403,N_12844,N_12401);
or U14404 (N_14404,N_13279,N_13579);
nor U14405 (N_14405,N_13074,N_13175);
or U14406 (N_14406,N_13442,N_13086);
nand U14407 (N_14407,N_12686,N_12563);
and U14408 (N_14408,N_13711,N_13425);
nor U14409 (N_14409,N_13421,N_12105);
nand U14410 (N_14410,N_12381,N_12489);
or U14411 (N_14411,N_13513,N_12011);
and U14412 (N_14412,N_12519,N_13878);
nand U14413 (N_14413,N_13063,N_12324);
xor U14414 (N_14414,N_13256,N_12091);
nor U14415 (N_14415,N_12270,N_12256);
and U14416 (N_14416,N_13154,N_13090);
nor U14417 (N_14417,N_13548,N_12239);
nand U14418 (N_14418,N_12576,N_12828);
xnor U14419 (N_14419,N_13628,N_13268);
or U14420 (N_14420,N_13118,N_13270);
nor U14421 (N_14421,N_13416,N_12683);
nand U14422 (N_14422,N_13704,N_13486);
or U14423 (N_14423,N_12027,N_12942);
and U14424 (N_14424,N_12863,N_13116);
nor U14425 (N_14425,N_12869,N_12982);
xnor U14426 (N_14426,N_12112,N_13788);
nand U14427 (N_14427,N_13088,N_13273);
nor U14428 (N_14428,N_13177,N_12302);
nand U14429 (N_14429,N_12017,N_12618);
or U14430 (N_14430,N_12628,N_12529);
xor U14431 (N_14431,N_12309,N_13639);
nor U14432 (N_14432,N_12819,N_12426);
xor U14433 (N_14433,N_13673,N_12118);
nand U14434 (N_14434,N_13399,N_13869);
and U14435 (N_14435,N_12673,N_13069);
nor U14436 (N_14436,N_12329,N_13528);
and U14437 (N_14437,N_12125,N_12175);
or U14438 (N_14438,N_13102,N_13762);
xnor U14439 (N_14439,N_13702,N_12183);
nand U14440 (N_14440,N_12084,N_13523);
xnor U14441 (N_14441,N_13364,N_13065);
xnor U14442 (N_14442,N_12327,N_12422);
xor U14443 (N_14443,N_13167,N_13982);
nor U14444 (N_14444,N_13001,N_12967);
nand U14445 (N_14445,N_13961,N_13959);
and U14446 (N_14446,N_12804,N_12528);
or U14447 (N_14447,N_12651,N_13876);
and U14448 (N_14448,N_13582,N_12573);
and U14449 (N_14449,N_13904,N_12046);
xor U14450 (N_14450,N_13542,N_13451);
or U14451 (N_14451,N_13700,N_13504);
nand U14452 (N_14452,N_12511,N_13569);
or U14453 (N_14453,N_12799,N_13134);
xor U14454 (N_14454,N_12496,N_12492);
xor U14455 (N_14455,N_12130,N_13368);
or U14456 (N_14456,N_13393,N_12801);
xor U14457 (N_14457,N_12392,N_13475);
xnor U14458 (N_14458,N_13710,N_12441);
and U14459 (N_14459,N_12838,N_12522);
nor U14460 (N_14460,N_13058,N_12455);
and U14461 (N_14461,N_12824,N_13637);
nand U14462 (N_14462,N_13839,N_12537);
xnor U14463 (N_14463,N_12042,N_12458);
nor U14464 (N_14464,N_12107,N_13962);
or U14465 (N_14465,N_12387,N_13457);
nand U14466 (N_14466,N_12494,N_13085);
and U14467 (N_14467,N_13223,N_13362);
and U14468 (N_14468,N_13166,N_12123);
nand U14469 (N_14469,N_13458,N_12832);
nor U14470 (N_14470,N_13665,N_13417);
nor U14471 (N_14471,N_13133,N_13446);
nand U14472 (N_14472,N_13817,N_12110);
nand U14473 (N_14473,N_13813,N_12456);
nor U14474 (N_14474,N_13284,N_13908);
nand U14475 (N_14475,N_12857,N_13345);
and U14476 (N_14476,N_13321,N_13681);
nor U14477 (N_14477,N_13023,N_12837);
nand U14478 (N_14478,N_12699,N_13662);
or U14479 (N_14479,N_13600,N_12968);
nor U14480 (N_14480,N_13978,N_12275);
nand U14481 (N_14481,N_13649,N_13791);
nand U14482 (N_14482,N_12550,N_12476);
nor U14483 (N_14483,N_13459,N_12831);
or U14484 (N_14484,N_13050,N_12423);
and U14485 (N_14485,N_12858,N_12583);
nand U14486 (N_14486,N_13990,N_13352);
xor U14487 (N_14487,N_12631,N_12040);
xor U14488 (N_14488,N_12734,N_13616);
and U14489 (N_14489,N_13040,N_12079);
nor U14490 (N_14490,N_13751,N_12316);
or U14491 (N_14491,N_12613,N_13447);
or U14492 (N_14492,N_12470,N_12592);
or U14493 (N_14493,N_12336,N_13310);
nor U14494 (N_14494,N_13034,N_12936);
or U14495 (N_14495,N_12780,N_13247);
or U14496 (N_14496,N_12388,N_13615);
nor U14497 (N_14497,N_13674,N_13693);
or U14498 (N_14498,N_12820,N_13599);
or U14499 (N_14499,N_13263,N_13096);
and U14500 (N_14500,N_13518,N_12988);
nor U14501 (N_14501,N_12934,N_13554);
and U14502 (N_14502,N_13507,N_12180);
nand U14503 (N_14503,N_13854,N_12738);
and U14504 (N_14504,N_12098,N_13075);
xnor U14505 (N_14505,N_12138,N_13656);
or U14506 (N_14506,N_13325,N_13551);
and U14507 (N_14507,N_12090,N_13390);
nor U14508 (N_14508,N_13282,N_13233);
xor U14509 (N_14509,N_13150,N_13375);
and U14510 (N_14510,N_12914,N_13603);
xnor U14511 (N_14511,N_12285,N_13984);
nor U14512 (N_14512,N_13339,N_12263);
nor U14513 (N_14513,N_12800,N_12474);
or U14514 (N_14514,N_13022,N_13764);
nand U14515 (N_14515,N_12222,N_12208);
or U14516 (N_14516,N_12436,N_13335);
xor U14517 (N_14517,N_12700,N_12928);
and U14518 (N_14518,N_13875,N_13655);
xnor U14519 (N_14519,N_12249,N_12638);
and U14520 (N_14520,N_12372,N_12578);
or U14521 (N_14521,N_12566,N_12045);
nor U14522 (N_14522,N_12939,N_12612);
or U14523 (N_14523,N_12437,N_13597);
xnor U14524 (N_14524,N_12117,N_13815);
nor U14525 (N_14525,N_13928,N_13613);
nor U14526 (N_14526,N_13168,N_13715);
nand U14527 (N_14527,N_13512,N_13879);
or U14528 (N_14528,N_13498,N_12139);
nor U14529 (N_14529,N_12323,N_13514);
nor U14530 (N_14530,N_12195,N_13089);
xor U14531 (N_14531,N_13607,N_12778);
nor U14532 (N_14532,N_12201,N_12994);
or U14533 (N_14533,N_12813,N_13843);
or U14534 (N_14534,N_12640,N_13527);
or U14535 (N_14535,N_12671,N_13736);
xor U14536 (N_14536,N_13497,N_13180);
nand U14537 (N_14537,N_12419,N_13035);
xnor U14538 (N_14538,N_13079,N_12798);
and U14539 (N_14539,N_13430,N_13391);
or U14540 (N_14540,N_13024,N_12710);
nand U14541 (N_14541,N_13848,N_13690);
nand U14542 (N_14542,N_12096,N_13963);
or U14543 (N_14543,N_12794,N_13900);
or U14544 (N_14544,N_13808,N_12367);
nand U14545 (N_14545,N_12005,N_13621);
and U14546 (N_14546,N_12213,N_13916);
nor U14547 (N_14547,N_12416,N_12050);
nand U14548 (N_14548,N_13319,N_13785);
or U14549 (N_14549,N_12704,N_13979);
nor U14550 (N_14550,N_13703,N_13291);
or U14551 (N_14551,N_13076,N_12541);
and U14552 (N_14552,N_13988,N_13164);
nand U14553 (N_14553,N_12827,N_13545);
or U14554 (N_14554,N_13799,N_13563);
and U14555 (N_14555,N_13768,N_12775);
xnor U14556 (N_14556,N_12615,N_12733);
nor U14557 (N_14557,N_13826,N_12067);
and U14558 (N_14558,N_13899,N_12898);
nand U14559 (N_14559,N_12991,N_12246);
xnor U14560 (N_14560,N_12135,N_12242);
xnor U14561 (N_14561,N_13438,N_13200);
xor U14562 (N_14562,N_12374,N_13143);
or U14563 (N_14563,N_12770,N_13408);
or U14564 (N_14564,N_12735,N_12758);
or U14565 (N_14565,N_12803,N_12930);
or U14566 (N_14566,N_12714,N_12616);
nor U14567 (N_14567,N_13806,N_13539);
nand U14568 (N_14568,N_12909,N_12552);
or U14569 (N_14569,N_13315,N_12214);
and U14570 (N_14570,N_12755,N_12283);
nand U14571 (N_14571,N_13684,N_12483);
xnor U14572 (N_14572,N_12666,N_12203);
nand U14573 (N_14573,N_13958,N_13057);
and U14574 (N_14574,N_13811,N_13091);
or U14575 (N_14575,N_13574,N_12022);
and U14576 (N_14576,N_13903,N_13654);
and U14577 (N_14577,N_12603,N_12133);
or U14578 (N_14578,N_13260,N_13508);
or U14579 (N_14579,N_13464,N_13078);
nor U14580 (N_14580,N_12221,N_13465);
xnor U14581 (N_14581,N_12841,N_13049);
and U14582 (N_14582,N_13005,N_12268);
nand U14583 (N_14583,N_12406,N_13014);
xnor U14584 (N_14584,N_13357,N_13919);
nor U14585 (N_14585,N_13056,N_13535);
and U14586 (N_14586,N_13594,N_13426);
nor U14587 (N_14587,N_13742,N_13191);
nand U14588 (N_14588,N_13404,N_12565);
xor U14589 (N_14589,N_13470,N_13192);
or U14590 (N_14590,N_13026,N_12836);
or U14591 (N_14591,N_12503,N_12431);
nand U14592 (N_14592,N_12493,N_12038);
nand U14593 (N_14593,N_13735,N_13045);
nor U14594 (N_14594,N_12088,N_12062);
and U14595 (N_14595,N_13965,N_12124);
or U14596 (N_14596,N_12900,N_13383);
or U14597 (N_14597,N_12253,N_12979);
nand U14598 (N_14598,N_13993,N_13429);
xnor U14599 (N_14599,N_12024,N_13659);
nand U14600 (N_14600,N_12335,N_12295);
nand U14601 (N_14601,N_12267,N_13038);
nor U14602 (N_14602,N_12557,N_13632);
and U14603 (N_14603,N_12205,N_13989);
nand U14604 (N_14604,N_12675,N_12287);
xnor U14605 (N_14605,N_12879,N_12262);
nor U14606 (N_14606,N_12542,N_13197);
nor U14607 (N_14607,N_13925,N_12764);
nand U14608 (N_14608,N_12512,N_13835);
nand U14609 (N_14609,N_13276,N_12231);
or U14610 (N_14610,N_12115,N_13062);
nor U14611 (N_14611,N_13415,N_12498);
and U14612 (N_14612,N_12332,N_13441);
and U14613 (N_14613,N_12782,N_12888);
or U14614 (N_14614,N_13469,N_13012);
nor U14615 (N_14615,N_12325,N_12767);
or U14616 (N_14616,N_12131,N_13146);
or U14617 (N_14617,N_12547,N_13964);
nor U14618 (N_14618,N_13820,N_12111);
xor U14619 (N_14619,N_12365,N_12410);
or U14620 (N_14620,N_12281,N_13623);
nand U14621 (N_14621,N_13501,N_12977);
or U14622 (N_14622,N_12935,N_13669);
or U14623 (N_14623,N_13396,N_12912);
and U14624 (N_14624,N_12679,N_12795);
or U14625 (N_14625,N_13280,N_13770);
or U14626 (N_14626,N_12867,N_12875);
or U14627 (N_14627,N_12271,N_12049);
or U14628 (N_14628,N_13478,N_13570);
nor U14629 (N_14629,N_12922,N_13618);
xor U14630 (N_14630,N_12159,N_12604);
xor U14631 (N_14631,N_12880,N_12992);
nor U14632 (N_14632,N_13443,N_12402);
and U14633 (N_14633,N_13334,N_12128);
xnor U14634 (N_14634,N_12784,N_13298);
nand U14635 (N_14635,N_13203,N_13874);
and U14636 (N_14636,N_13405,N_13070);
and U14637 (N_14637,N_12166,N_13190);
xor U14638 (N_14638,N_12400,N_12591);
xor U14639 (N_14639,N_12523,N_13109);
nand U14640 (N_14640,N_12835,N_12696);
nand U14641 (N_14641,N_13636,N_13135);
or U14642 (N_14642,N_12173,N_12354);
and U14643 (N_14643,N_12786,N_13186);
and U14644 (N_14644,N_13873,N_13481);
xor U14645 (N_14645,N_13389,N_13741);
nand U14646 (N_14646,N_12851,N_12318);
or U14647 (N_14647,N_13373,N_12590);
xnor U14648 (N_14648,N_12487,N_13299);
or U14649 (N_14649,N_12371,N_12619);
and U14650 (N_14650,N_13855,N_13688);
nor U14651 (N_14651,N_12186,N_12864);
xnor U14652 (N_14652,N_12298,N_13540);
nor U14653 (N_14653,N_13028,N_13156);
nor U14654 (N_14654,N_13055,N_13920);
or U14655 (N_14655,N_12439,N_12462);
or U14656 (N_14656,N_13585,N_12427);
xor U14657 (N_14657,N_13387,N_13179);
and U14658 (N_14658,N_12215,N_12444);
nor U14659 (N_14659,N_13525,N_12177);
and U14660 (N_14660,N_13365,N_13652);
and U14661 (N_14661,N_12066,N_12893);
xnor U14662 (N_14662,N_12693,N_13374);
nor U14663 (N_14663,N_13823,N_12745);
xnor U14664 (N_14664,N_13553,N_12041);
nor U14665 (N_14665,N_12904,N_13872);
and U14666 (N_14666,N_13129,N_12395);
or U14667 (N_14667,N_12532,N_12856);
nand U14668 (N_14668,N_13100,N_13609);
or U14669 (N_14669,N_12974,N_12876);
and U14670 (N_14670,N_13413,N_12944);
nand U14671 (N_14671,N_13104,N_12847);
nand U14672 (N_14672,N_13473,N_13729);
nand U14673 (N_14673,N_12633,N_13641);
or U14674 (N_14674,N_13488,N_12382);
xnor U14675 (N_14675,N_12454,N_12506);
xor U14676 (N_14676,N_13680,N_13723);
nor U14677 (N_14677,N_12415,N_12383);
nand U14678 (N_14678,N_12272,N_12551);
and U14679 (N_14679,N_13763,N_12940);
xor U14680 (N_14680,N_13744,N_13816);
xor U14681 (N_14681,N_12447,N_12920);
or U14682 (N_14682,N_13974,N_13043);
or U14683 (N_14683,N_12304,N_13082);
xnor U14684 (N_14684,N_13819,N_12122);
nor U14685 (N_14685,N_12359,N_12082);
nand U14686 (N_14686,N_12345,N_12853);
nor U14687 (N_14687,N_12510,N_13479);
nor U14688 (N_14688,N_13094,N_12840);
or U14689 (N_14689,N_13560,N_12891);
nand U14690 (N_14690,N_12726,N_12951);
or U14691 (N_14691,N_12396,N_12308);
xor U14692 (N_14692,N_13846,N_12219);
xor U14693 (N_14693,N_12750,N_12980);
nand U14694 (N_14694,N_13805,N_13472);
xor U14695 (N_14695,N_12821,N_12772);
xnor U14696 (N_14696,N_13313,N_12059);
and U14697 (N_14697,N_12538,N_12773);
nand U14698 (N_14698,N_12198,N_13395);
xnor U14699 (N_14699,N_12116,N_13195);
nor U14700 (N_14700,N_13556,N_12162);
nor U14701 (N_14701,N_13381,N_12212);
nor U14702 (N_14702,N_13316,N_13252);
xnor U14703 (N_14703,N_13760,N_13505);
xor U14704 (N_14704,N_13614,N_13794);
or U14705 (N_14705,N_13924,N_12278);
and U14706 (N_14706,N_13452,N_12950);
nand U14707 (N_14707,N_13857,N_12002);
xnor U14708 (N_14708,N_13127,N_13828);
nand U14709 (N_14709,N_12790,N_12328);
or U14710 (N_14710,N_12206,N_12677);
nor U14711 (N_14711,N_13110,N_13581);
nand U14712 (N_14712,N_12140,N_12420);
or U14713 (N_14713,N_13544,N_13761);
nand U14714 (N_14714,N_13445,N_12469);
nand U14715 (N_14715,N_12501,N_12034);
nand U14716 (N_14716,N_13448,N_12063);
nand U14717 (N_14717,N_12627,N_13114);
nand U14718 (N_14718,N_12742,N_13861);
nand U14719 (N_14719,N_13658,N_12812);
or U14720 (N_14720,N_13450,N_12760);
nand U14721 (N_14721,N_12906,N_13000);
and U14722 (N_14722,N_13329,N_13302);
and U14723 (N_14723,N_12121,N_13566);
xnor U14724 (N_14724,N_12204,N_13896);
nor U14725 (N_14725,N_13378,N_13951);
nor U14726 (N_14726,N_12001,N_12146);
and U14727 (N_14727,N_12688,N_13992);
and U14728 (N_14728,N_13115,N_12783);
or U14729 (N_14729,N_13394,N_12986);
nor U14730 (N_14730,N_12762,N_13286);
xnor U14731 (N_14731,N_13630,N_13161);
xor U14732 (N_14732,N_12334,N_12866);
and U14733 (N_14733,N_12513,N_13726);
xor U14734 (N_14734,N_12006,N_13583);
or U14735 (N_14735,N_12475,N_13106);
nor U14736 (N_14736,N_13124,N_13047);
and U14737 (N_14737,N_12225,N_12104);
nor U14738 (N_14738,N_13277,N_12301);
xor U14739 (N_14739,N_13251,N_13660);
or U14740 (N_14740,N_13575,N_13671);
nand U14741 (N_14741,N_12134,N_12086);
nor U14742 (N_14742,N_12881,N_12884);
nand U14743 (N_14743,N_13792,N_13520);
and U14744 (N_14744,N_13864,N_12984);
or U14745 (N_14745,N_13831,N_13305);
and U14746 (N_14746,N_12531,N_13379);
nand U14747 (N_14747,N_13037,N_12442);
xor U14748 (N_14748,N_13366,N_13980);
xor U14749 (N_14749,N_13258,N_12007);
nand U14750 (N_14750,N_12870,N_13369);
nor U14751 (N_14751,N_12527,N_13372);
or U14752 (N_14752,N_12740,N_13954);
nand U14753 (N_14753,N_13631,N_13392);
nand U14754 (N_14754,N_13410,N_12403);
xor U14755 (N_14755,N_12882,N_12349);
xor U14756 (N_14756,N_12946,N_12787);
and U14757 (N_14757,N_13549,N_12564);
and U14758 (N_14758,N_12545,N_12530);
nand U14759 (N_14759,N_12274,N_13677);
nand U14760 (N_14760,N_12515,N_12161);
and U14761 (N_14761,N_12965,N_13911);
xnor U14762 (N_14762,N_12273,N_13748);
or U14763 (N_14763,N_13431,N_12571);
nor U14764 (N_14764,N_13868,N_13216);
and U14765 (N_14765,N_12917,N_12706);
and U14766 (N_14766,N_12508,N_13883);
and U14767 (N_14767,N_12825,N_12191);
xnor U14768 (N_14768,N_13041,N_13929);
xor U14769 (N_14769,N_12428,N_13087);
xnor U14770 (N_14770,N_13509,N_12763);
nand U14771 (N_14771,N_12394,N_12072);
or U14772 (N_14772,N_12241,N_12430);
nor U14773 (N_14773,N_12355,N_13491);
nand U14774 (N_14774,N_13624,N_12296);
nand U14775 (N_14775,N_13428,N_12305);
and U14776 (N_14776,N_12518,N_13371);
nor U14777 (N_14777,N_13485,N_13255);
and U14778 (N_14778,N_12721,N_12168);
and U14779 (N_14779,N_12779,N_12315);
nand U14780 (N_14780,N_13433,N_12996);
nor U14781 (N_14781,N_12070,N_13253);
nor U14782 (N_14782,N_13663,N_13734);
or U14783 (N_14783,N_12149,N_13344);
or U14784 (N_14784,N_13697,N_12544);
nor U14785 (N_14785,N_13981,N_12081);
nor U14786 (N_14786,N_12258,N_13349);
nand U14787 (N_14787,N_13347,N_13356);
xnor U14788 (N_14788,N_12533,N_12421);
nor U14789 (N_14789,N_13867,N_12672);
xnor U14790 (N_14790,N_13219,N_13727);
nand U14791 (N_14791,N_12556,N_13243);
and U14792 (N_14792,N_13830,N_13220);
xor U14793 (N_14793,N_12907,N_13281);
or U14794 (N_14794,N_13804,N_13388);
nand U14795 (N_14795,N_12218,N_13328);
nand U14796 (N_14796,N_12306,N_13786);
nand U14797 (N_14797,N_13730,N_13967);
xor U14798 (N_14798,N_13914,N_13351);
nor U14799 (N_14799,N_13137,N_12333);
nor U14800 (N_14800,N_12000,N_12080);
and U14801 (N_14801,N_13121,N_12044);
or U14802 (N_14802,N_12826,N_12399);
nor U14803 (N_14803,N_12805,N_12481);
or U14804 (N_14804,N_13708,N_13149);
or U14805 (N_14805,N_13679,N_12860);
xor U14806 (N_14806,N_13358,N_13797);
or U14807 (N_14807,N_12379,N_12635);
nor U14808 (N_14808,N_12969,N_12806);
nand U14809 (N_14809,N_13385,N_12348);
xor U14810 (N_14810,N_12500,N_13534);
xnor U14811 (N_14811,N_13406,N_12320);
nor U14812 (N_14812,N_13236,N_12250);
nor U14813 (N_14813,N_12534,N_12479);
nor U14814 (N_14814,N_12634,N_12723);
and U14815 (N_14815,N_12484,N_13775);
nor U14816 (N_14816,N_13643,N_13926);
nand U14817 (N_14817,N_12717,N_12169);
and U14818 (N_14818,N_13687,N_13719);
xnor U14819 (N_14819,N_13230,N_12119);
and U14820 (N_14820,N_13728,N_12092);
or U14821 (N_14821,N_13092,N_12926);
and U14822 (N_14822,N_13209,N_12895);
and U14823 (N_14823,N_13296,N_12918);
nand U14824 (N_14824,N_13818,N_13333);
xor U14825 (N_14825,N_12156,N_12761);
and U14826 (N_14826,N_12987,N_12887);
xor U14827 (N_14827,N_13068,N_13126);
or U14828 (N_14828,N_12446,N_12247);
or U14829 (N_14829,N_13477,N_12292);
nor U14830 (N_14830,N_12277,N_12014);
xnor U14831 (N_14831,N_13718,N_13294);
or U14832 (N_14832,N_13568,N_12438);
xor U14833 (N_14833,N_12039,N_12668);
nor U14834 (N_14834,N_13411,N_12141);
xor U14835 (N_14835,N_13947,N_13749);
nand U14836 (N_14836,N_12567,N_12645);
xnor U14837 (N_14837,N_12665,N_13844);
nor U14838 (N_14838,N_12691,N_12728);
and U14839 (N_14839,N_12990,N_13029);
or U14840 (N_14840,N_12106,N_12491);
xor U14841 (N_14841,N_12485,N_12921);
nand U14842 (N_14842,N_13009,N_12314);
nor U14843 (N_14843,N_12957,N_12085);
and U14844 (N_14844,N_13564,N_12877);
or U14845 (N_14845,N_13454,N_12265);
and U14846 (N_14846,N_12722,N_12255);
or U14847 (N_14847,N_13912,N_13095);
and U14848 (N_14848,N_12425,N_13666);
or U14849 (N_14849,N_12650,N_12524);
nor U14850 (N_14850,N_12377,N_13721);
and U14851 (N_14851,N_12938,N_13067);
nor U14852 (N_14852,N_12724,N_12350);
nand U14853 (N_14853,N_12210,N_13913);
nand U14854 (N_14854,N_12031,N_13194);
nor U14855 (N_14855,N_13894,N_12731);
nand U14856 (N_14856,N_13619,N_13588);
nand U14857 (N_14857,N_12823,N_13699);
xnor U14858 (N_14858,N_13148,N_12708);
nand U14859 (N_14859,N_12293,N_13241);
xor U14860 (N_14860,N_13492,N_12235);
nor U14861 (N_14861,N_12196,N_12598);
xnor U14862 (N_14862,N_13511,N_13032);
and U14863 (N_14863,N_12126,N_13031);
xnor U14864 (N_14864,N_12901,N_12145);
or U14865 (N_14865,N_13301,N_12737);
nor U14866 (N_14866,N_12357,N_12245);
nand U14867 (N_14867,N_13576,N_13046);
and U14868 (N_14868,N_12150,N_12144);
and U14869 (N_14869,N_13955,N_13359);
xor U14870 (N_14870,N_12902,N_13706);
xnor U14871 (N_14871,N_13275,N_12097);
nand U14872 (N_14872,N_12347,N_12754);
nand U14873 (N_14873,N_12561,N_12192);
nor U14874 (N_14874,N_12380,N_13841);
nand U14875 (N_14875,N_13494,N_12998);
or U14876 (N_14876,N_13306,N_13692);
or U14877 (N_14877,N_13331,N_13640);
and U14878 (N_14878,N_12626,N_13897);
xnor U14879 (N_14879,N_12749,N_12654);
and U14880 (N_14880,N_12016,N_13271);
xor U14881 (N_14881,N_13837,N_12849);
nor U14882 (N_14882,N_12973,N_13937);
xnor U14883 (N_14883,N_13558,N_12788);
xnor U14884 (N_14884,N_13863,N_12852);
xnor U14885 (N_14885,N_13409,N_13427);
nand U14886 (N_14886,N_12102,N_13853);
or U14887 (N_14887,N_13025,N_12549);
nor U14888 (N_14888,N_12362,N_12948);
nand U14889 (N_14889,N_13635,N_12074);
xor U14890 (N_14890,N_13571,N_12593);
nor U14891 (N_14891,N_12894,N_13944);
xnor U14892 (N_14892,N_13705,N_12695);
xnor U14893 (N_14893,N_12405,N_12703);
or U14894 (N_14894,N_13530,N_13972);
nor U14895 (N_14895,N_12179,N_12385);
and U14896 (N_14896,N_13332,N_12398);
nor U14897 (N_14897,N_12546,N_13463);
and U14898 (N_14898,N_12155,N_12871);
nand U14899 (N_14899,N_13117,N_12652);
or U14900 (N_14900,N_13629,N_13278);
nand U14901 (N_14901,N_12568,N_13773);
nor U14902 (N_14902,N_12068,N_12680);
and U14903 (N_14903,N_12607,N_13755);
or U14904 (N_14904,N_13782,N_12217);
nor U14905 (N_14905,N_12113,N_12890);
nand U14906 (N_14906,N_13158,N_12356);
xor U14907 (N_14907,N_12291,N_12981);
nand U14908 (N_14908,N_13653,N_12009);
xnor U14909 (N_14909,N_12358,N_13930);
and U14910 (N_14910,N_12789,N_13952);
nand U14911 (N_14911,N_12589,N_12207);
and U14912 (N_14912,N_12736,N_12659);
nand U14913 (N_14913,N_13586,N_12687);
nor U14914 (N_14914,N_12586,N_12137);
nand U14915 (N_14915,N_12486,N_13370);
and U14916 (N_14916,N_12933,N_13176);
or U14917 (N_14917,N_12712,N_13890);
or U14918 (N_14918,N_13537,N_13921);
and U14919 (N_14919,N_12656,N_12143);
and U14920 (N_14920,N_12756,N_13064);
nand U14921 (N_14921,N_13297,N_13682);
nand U14922 (N_14922,N_12408,N_13898);
nand U14923 (N_14923,N_13712,N_13173);
nand U14924 (N_14924,N_12114,N_13244);
and U14925 (N_14925,N_13533,N_13591);
xor U14926 (N_14926,N_12924,N_12807);
or U14927 (N_14927,N_13745,N_12829);
and U14928 (N_14928,N_12457,N_13789);
nand U14929 (N_14929,N_13039,N_12601);
xor U14930 (N_14930,N_13027,N_13783);
nand U14931 (N_14931,N_12311,N_12859);
and U14932 (N_14932,N_13933,N_13108);
nor U14933 (N_14933,N_12414,N_12817);
nand U14934 (N_14934,N_12725,N_13877);
nand U14935 (N_14935,N_12916,N_13717);
or U14936 (N_14936,N_13018,N_12943);
nand U14937 (N_14937,N_13969,N_13010);
and U14938 (N_14938,N_13471,N_12240);
or U14939 (N_14939,N_13423,N_13885);
or U14940 (N_14940,N_13103,N_12536);
nand U14941 (N_14941,N_13759,N_12100);
or U14942 (N_14942,N_13968,N_12743);
or U14943 (N_14943,N_12608,N_12230);
or U14944 (N_14944,N_12226,N_13809);
xor U14945 (N_14945,N_12243,N_12312);
or U14946 (N_14946,N_13918,N_13689);
xor U14947 (N_14947,N_13787,N_12200);
or U14948 (N_14948,N_13584,N_13128);
or U14949 (N_14949,N_13541,N_12774);
nand U14950 (N_14950,N_13187,N_13731);
nor U14951 (N_14951,N_13224,N_12692);
and U14952 (N_14952,N_12048,N_12229);
or U14953 (N_14953,N_13910,N_12872);
and U14954 (N_14954,N_13774,N_12661);
and U14955 (N_14955,N_13042,N_12993);
nand U14956 (N_14956,N_12707,N_13130);
nor U14957 (N_14957,N_13781,N_12642);
and U14958 (N_14958,N_12808,N_12165);
or U14959 (N_14959,N_12581,N_13935);
or U14960 (N_14960,N_13350,N_12791);
or U14961 (N_14961,N_13174,N_13650);
nand U14962 (N_14962,N_12232,N_12251);
xnor U14963 (N_14963,N_13502,N_13648);
xnor U14964 (N_14964,N_13516,N_12061);
or U14965 (N_14965,N_13939,N_12850);
nor U14966 (N_14966,N_12878,N_13170);
xnor U14967 (N_14967,N_13836,N_13157);
xnor U14968 (N_14968,N_13977,N_12171);
nand U14969 (N_14969,N_13953,N_12525);
and U14970 (N_14970,N_12713,N_12465);
nor U14971 (N_14971,N_12558,N_12983);
and U14972 (N_14972,N_13577,N_13483);
nand U14973 (N_14973,N_13384,N_13827);
nand U14974 (N_14974,N_12937,N_13246);
nand U14975 (N_14975,N_13487,N_12199);
and U14976 (N_14976,N_12297,N_12445);
nand U14977 (N_14977,N_13476,N_13976);
nor U14978 (N_14978,N_12759,N_13151);
or U14979 (N_14979,N_13612,N_13422);
and U14980 (N_14980,N_12087,N_13123);
xor U14981 (N_14981,N_12020,N_12160);
or U14982 (N_14982,N_13020,N_13011);
nand U14983 (N_14983,N_13519,N_13312);
or U14984 (N_14984,N_13226,N_13940);
xnor U14985 (N_14985,N_12599,N_12384);
and U14986 (N_14986,N_13208,N_12669);
nand U14987 (N_14987,N_12630,N_13482);
nand U14988 (N_14988,N_12614,N_12732);
or U14989 (N_14989,N_13832,N_13202);
nor U14990 (N_14990,N_13265,N_12033);
nor U14991 (N_14991,N_13338,N_13814);
xor U14992 (N_14992,N_12861,N_12178);
nor U14993 (N_14993,N_13767,N_13317);
nor U14994 (N_14994,N_13991,N_12678);
nand U14995 (N_14995,N_13401,N_13790);
nand U14996 (N_14996,N_12194,N_12753);
nor U14997 (N_14997,N_12796,N_13015);
nand U14998 (N_14998,N_12429,N_12452);
or U14999 (N_14999,N_13807,N_12089);
xor U15000 (N_15000,N_13061,N_12546);
and U15001 (N_15001,N_13135,N_12097);
nand U15002 (N_15002,N_12824,N_12626);
and U15003 (N_15003,N_13771,N_12372);
and U15004 (N_15004,N_13126,N_12769);
xor U15005 (N_15005,N_12919,N_12134);
xor U15006 (N_15006,N_12060,N_13346);
nor U15007 (N_15007,N_12132,N_12185);
nand U15008 (N_15008,N_12328,N_13361);
and U15009 (N_15009,N_12283,N_12077);
or U15010 (N_15010,N_13966,N_12477);
nand U15011 (N_15011,N_12866,N_13696);
nand U15012 (N_15012,N_12519,N_12241);
nor U15013 (N_15013,N_13076,N_13541);
nand U15014 (N_15014,N_13973,N_12589);
and U15015 (N_15015,N_13708,N_13648);
nor U15016 (N_15016,N_13292,N_12911);
and U15017 (N_15017,N_13027,N_13601);
or U15018 (N_15018,N_13431,N_13288);
or U15019 (N_15019,N_12869,N_12304);
xnor U15020 (N_15020,N_12808,N_12895);
xnor U15021 (N_15021,N_12608,N_12059);
nor U15022 (N_15022,N_12550,N_12719);
and U15023 (N_15023,N_13839,N_13505);
nand U15024 (N_15024,N_12628,N_13209);
or U15025 (N_15025,N_12322,N_13768);
or U15026 (N_15026,N_12722,N_12937);
or U15027 (N_15027,N_12092,N_12765);
nand U15028 (N_15028,N_12568,N_13091);
nor U15029 (N_15029,N_12157,N_12105);
and U15030 (N_15030,N_13861,N_12297);
and U15031 (N_15031,N_12314,N_12500);
xor U15032 (N_15032,N_12550,N_13052);
nor U15033 (N_15033,N_12171,N_13311);
or U15034 (N_15034,N_13217,N_13703);
or U15035 (N_15035,N_12463,N_12874);
and U15036 (N_15036,N_12757,N_13358);
nand U15037 (N_15037,N_12334,N_12602);
and U15038 (N_15038,N_13890,N_13539);
xnor U15039 (N_15039,N_12401,N_12909);
xor U15040 (N_15040,N_12644,N_13741);
and U15041 (N_15041,N_12525,N_12043);
nand U15042 (N_15042,N_12438,N_13684);
nand U15043 (N_15043,N_13988,N_12047);
nand U15044 (N_15044,N_13015,N_12419);
nor U15045 (N_15045,N_12927,N_12071);
nand U15046 (N_15046,N_13513,N_13946);
and U15047 (N_15047,N_13148,N_13717);
nor U15048 (N_15048,N_13306,N_12711);
xnor U15049 (N_15049,N_12453,N_13495);
or U15050 (N_15050,N_12298,N_12434);
nand U15051 (N_15051,N_12838,N_12040);
or U15052 (N_15052,N_12931,N_12769);
and U15053 (N_15053,N_13974,N_12592);
xor U15054 (N_15054,N_13430,N_13572);
nand U15055 (N_15055,N_12129,N_13486);
and U15056 (N_15056,N_12358,N_13888);
and U15057 (N_15057,N_12696,N_12041);
or U15058 (N_15058,N_13413,N_13903);
nand U15059 (N_15059,N_12312,N_12860);
or U15060 (N_15060,N_12656,N_12982);
nand U15061 (N_15061,N_13299,N_12810);
nand U15062 (N_15062,N_13087,N_13444);
nor U15063 (N_15063,N_12239,N_12105);
and U15064 (N_15064,N_12783,N_12553);
and U15065 (N_15065,N_12836,N_12960);
or U15066 (N_15066,N_12326,N_12460);
and U15067 (N_15067,N_13455,N_13597);
nor U15068 (N_15068,N_13801,N_12342);
nor U15069 (N_15069,N_13564,N_13421);
nor U15070 (N_15070,N_13172,N_13632);
or U15071 (N_15071,N_13481,N_13494);
nor U15072 (N_15072,N_12820,N_12951);
xnor U15073 (N_15073,N_13580,N_12374);
nor U15074 (N_15074,N_12268,N_12271);
xnor U15075 (N_15075,N_12334,N_12590);
nor U15076 (N_15076,N_12430,N_12072);
or U15077 (N_15077,N_12691,N_12426);
or U15078 (N_15078,N_13301,N_12064);
or U15079 (N_15079,N_12185,N_13899);
nand U15080 (N_15080,N_13736,N_12495);
and U15081 (N_15081,N_13686,N_13139);
and U15082 (N_15082,N_12269,N_12087);
or U15083 (N_15083,N_13713,N_12299);
nor U15084 (N_15084,N_12359,N_12762);
or U15085 (N_15085,N_12699,N_13601);
or U15086 (N_15086,N_12313,N_13775);
and U15087 (N_15087,N_12892,N_12691);
nand U15088 (N_15088,N_12464,N_13351);
and U15089 (N_15089,N_12355,N_12926);
nand U15090 (N_15090,N_12844,N_12437);
xor U15091 (N_15091,N_13273,N_13575);
or U15092 (N_15092,N_12054,N_12053);
and U15093 (N_15093,N_13460,N_12704);
or U15094 (N_15094,N_13243,N_12464);
and U15095 (N_15095,N_12874,N_13587);
nand U15096 (N_15096,N_13621,N_12152);
or U15097 (N_15097,N_13739,N_12082);
or U15098 (N_15098,N_12449,N_12822);
nor U15099 (N_15099,N_12391,N_13536);
xor U15100 (N_15100,N_13087,N_12516);
nand U15101 (N_15101,N_13293,N_13230);
xnor U15102 (N_15102,N_12684,N_12242);
or U15103 (N_15103,N_12816,N_12191);
nor U15104 (N_15104,N_12462,N_12980);
or U15105 (N_15105,N_13015,N_12739);
or U15106 (N_15106,N_13075,N_12259);
nor U15107 (N_15107,N_12232,N_12373);
or U15108 (N_15108,N_13316,N_13699);
xnor U15109 (N_15109,N_12153,N_13324);
nand U15110 (N_15110,N_12351,N_13747);
and U15111 (N_15111,N_12670,N_12525);
nor U15112 (N_15112,N_12345,N_13613);
nand U15113 (N_15113,N_13239,N_12697);
xnor U15114 (N_15114,N_13918,N_13283);
nand U15115 (N_15115,N_13161,N_13486);
and U15116 (N_15116,N_12678,N_12039);
nand U15117 (N_15117,N_12664,N_13879);
and U15118 (N_15118,N_13833,N_12143);
nand U15119 (N_15119,N_13704,N_13727);
and U15120 (N_15120,N_13785,N_13900);
xor U15121 (N_15121,N_12118,N_13608);
nand U15122 (N_15122,N_12746,N_13415);
or U15123 (N_15123,N_13080,N_13044);
nand U15124 (N_15124,N_12288,N_13132);
nor U15125 (N_15125,N_12491,N_12323);
nor U15126 (N_15126,N_13803,N_12334);
nand U15127 (N_15127,N_13798,N_13396);
xnor U15128 (N_15128,N_12295,N_13739);
nor U15129 (N_15129,N_13052,N_12542);
nor U15130 (N_15130,N_12311,N_13166);
nor U15131 (N_15131,N_13855,N_13279);
or U15132 (N_15132,N_13949,N_13421);
and U15133 (N_15133,N_13919,N_13321);
or U15134 (N_15134,N_13275,N_12869);
xnor U15135 (N_15135,N_13181,N_13372);
nand U15136 (N_15136,N_13709,N_12219);
xor U15137 (N_15137,N_12853,N_12679);
or U15138 (N_15138,N_13450,N_12731);
or U15139 (N_15139,N_13101,N_13476);
nand U15140 (N_15140,N_13695,N_12349);
nor U15141 (N_15141,N_13342,N_13310);
or U15142 (N_15142,N_13323,N_12379);
or U15143 (N_15143,N_13540,N_12323);
xnor U15144 (N_15144,N_13881,N_13105);
xnor U15145 (N_15145,N_13822,N_13151);
nand U15146 (N_15146,N_13163,N_12743);
or U15147 (N_15147,N_12861,N_12256);
and U15148 (N_15148,N_12005,N_13385);
and U15149 (N_15149,N_12216,N_13391);
xnor U15150 (N_15150,N_13625,N_13665);
xnor U15151 (N_15151,N_12053,N_13522);
nand U15152 (N_15152,N_12790,N_12714);
nor U15153 (N_15153,N_12160,N_13185);
or U15154 (N_15154,N_12263,N_13053);
nand U15155 (N_15155,N_12102,N_12746);
and U15156 (N_15156,N_12545,N_12122);
nand U15157 (N_15157,N_12650,N_12221);
and U15158 (N_15158,N_12357,N_12940);
and U15159 (N_15159,N_12867,N_13166);
or U15160 (N_15160,N_12104,N_13028);
or U15161 (N_15161,N_13479,N_12905);
nor U15162 (N_15162,N_12983,N_12706);
and U15163 (N_15163,N_12167,N_13577);
xnor U15164 (N_15164,N_12127,N_12397);
or U15165 (N_15165,N_12833,N_13443);
and U15166 (N_15166,N_12821,N_12287);
xor U15167 (N_15167,N_12242,N_12454);
and U15168 (N_15168,N_12943,N_12413);
xnor U15169 (N_15169,N_12634,N_12384);
and U15170 (N_15170,N_12638,N_12215);
nand U15171 (N_15171,N_12682,N_12375);
nor U15172 (N_15172,N_13421,N_12613);
nand U15173 (N_15173,N_13798,N_13962);
nand U15174 (N_15174,N_13382,N_12645);
xnor U15175 (N_15175,N_13839,N_12941);
and U15176 (N_15176,N_12137,N_13650);
xor U15177 (N_15177,N_13107,N_12488);
xor U15178 (N_15178,N_13797,N_13240);
or U15179 (N_15179,N_13234,N_13577);
xor U15180 (N_15180,N_13520,N_12485);
nor U15181 (N_15181,N_13492,N_13207);
and U15182 (N_15182,N_13940,N_13259);
xor U15183 (N_15183,N_12633,N_13999);
xnor U15184 (N_15184,N_13920,N_12279);
nor U15185 (N_15185,N_13266,N_12682);
nand U15186 (N_15186,N_13768,N_13929);
and U15187 (N_15187,N_12031,N_12442);
or U15188 (N_15188,N_12222,N_12618);
and U15189 (N_15189,N_12261,N_12143);
and U15190 (N_15190,N_13368,N_12725);
or U15191 (N_15191,N_12974,N_12406);
nor U15192 (N_15192,N_12630,N_12543);
xor U15193 (N_15193,N_13372,N_13420);
or U15194 (N_15194,N_13866,N_12837);
and U15195 (N_15195,N_13045,N_13027);
nor U15196 (N_15196,N_13276,N_13677);
nand U15197 (N_15197,N_13824,N_13248);
xor U15198 (N_15198,N_12116,N_12856);
nand U15199 (N_15199,N_12013,N_12313);
nand U15200 (N_15200,N_13666,N_12472);
or U15201 (N_15201,N_13335,N_13158);
nor U15202 (N_15202,N_12908,N_12261);
xnor U15203 (N_15203,N_12257,N_13275);
nand U15204 (N_15204,N_12137,N_13299);
xnor U15205 (N_15205,N_13959,N_13821);
nand U15206 (N_15206,N_13013,N_13182);
and U15207 (N_15207,N_13216,N_13902);
and U15208 (N_15208,N_12211,N_12476);
nor U15209 (N_15209,N_12332,N_12138);
and U15210 (N_15210,N_12646,N_13517);
nand U15211 (N_15211,N_13135,N_12377);
nand U15212 (N_15212,N_12565,N_12079);
nor U15213 (N_15213,N_13601,N_13494);
xnor U15214 (N_15214,N_12984,N_13403);
or U15215 (N_15215,N_12711,N_12141);
nand U15216 (N_15216,N_13145,N_13202);
xnor U15217 (N_15217,N_13864,N_13705);
nor U15218 (N_15218,N_13307,N_13871);
nor U15219 (N_15219,N_13699,N_13805);
xnor U15220 (N_15220,N_13754,N_12336);
or U15221 (N_15221,N_12890,N_12169);
nand U15222 (N_15222,N_13022,N_12252);
nand U15223 (N_15223,N_13261,N_12647);
nand U15224 (N_15224,N_12726,N_12844);
nor U15225 (N_15225,N_13409,N_13689);
or U15226 (N_15226,N_13117,N_13058);
nand U15227 (N_15227,N_13073,N_13216);
nand U15228 (N_15228,N_12658,N_13545);
nor U15229 (N_15229,N_12245,N_13397);
xnor U15230 (N_15230,N_12348,N_12577);
and U15231 (N_15231,N_13794,N_12765);
xor U15232 (N_15232,N_12759,N_12684);
and U15233 (N_15233,N_13465,N_12173);
nand U15234 (N_15234,N_13857,N_13743);
or U15235 (N_15235,N_13582,N_12319);
or U15236 (N_15236,N_12984,N_12691);
xnor U15237 (N_15237,N_12307,N_13509);
and U15238 (N_15238,N_12093,N_12150);
nor U15239 (N_15239,N_13968,N_13001);
or U15240 (N_15240,N_12336,N_12398);
nor U15241 (N_15241,N_12740,N_12516);
nand U15242 (N_15242,N_13580,N_12270);
xor U15243 (N_15243,N_13177,N_12303);
nor U15244 (N_15244,N_12468,N_12016);
xnor U15245 (N_15245,N_13274,N_12037);
nor U15246 (N_15246,N_13843,N_12211);
and U15247 (N_15247,N_13877,N_12300);
nand U15248 (N_15248,N_12711,N_12994);
xor U15249 (N_15249,N_13596,N_13500);
nand U15250 (N_15250,N_13680,N_12594);
xor U15251 (N_15251,N_13908,N_13899);
xnor U15252 (N_15252,N_12083,N_12005);
and U15253 (N_15253,N_12247,N_13859);
xnor U15254 (N_15254,N_13874,N_13862);
nand U15255 (N_15255,N_12323,N_13303);
nor U15256 (N_15256,N_12387,N_13319);
xor U15257 (N_15257,N_12682,N_12086);
or U15258 (N_15258,N_12640,N_12987);
or U15259 (N_15259,N_12255,N_13752);
xor U15260 (N_15260,N_13392,N_13147);
or U15261 (N_15261,N_12703,N_13709);
and U15262 (N_15262,N_13564,N_13978);
nand U15263 (N_15263,N_12500,N_13707);
xor U15264 (N_15264,N_13544,N_13978);
nand U15265 (N_15265,N_13827,N_12235);
and U15266 (N_15266,N_13635,N_12935);
or U15267 (N_15267,N_12377,N_13593);
xnor U15268 (N_15268,N_12229,N_12991);
and U15269 (N_15269,N_12901,N_12879);
and U15270 (N_15270,N_12223,N_13533);
xor U15271 (N_15271,N_13841,N_13576);
or U15272 (N_15272,N_12458,N_12700);
or U15273 (N_15273,N_12948,N_12776);
xor U15274 (N_15274,N_12628,N_13836);
or U15275 (N_15275,N_13446,N_12347);
nor U15276 (N_15276,N_13531,N_13082);
and U15277 (N_15277,N_12721,N_12845);
and U15278 (N_15278,N_12219,N_13909);
xnor U15279 (N_15279,N_13162,N_12701);
and U15280 (N_15280,N_12179,N_12730);
and U15281 (N_15281,N_12485,N_12351);
and U15282 (N_15282,N_13969,N_12144);
and U15283 (N_15283,N_13450,N_12548);
or U15284 (N_15284,N_12854,N_12443);
and U15285 (N_15285,N_13361,N_12784);
nor U15286 (N_15286,N_12987,N_12709);
or U15287 (N_15287,N_12230,N_13936);
or U15288 (N_15288,N_13722,N_13956);
nand U15289 (N_15289,N_12218,N_12242);
and U15290 (N_15290,N_13265,N_13766);
xor U15291 (N_15291,N_12493,N_13268);
nor U15292 (N_15292,N_13151,N_12400);
nand U15293 (N_15293,N_13552,N_13664);
xnor U15294 (N_15294,N_12269,N_13094);
nor U15295 (N_15295,N_13326,N_13126);
and U15296 (N_15296,N_13649,N_12032);
and U15297 (N_15297,N_12489,N_13365);
or U15298 (N_15298,N_12813,N_12540);
and U15299 (N_15299,N_13836,N_12584);
nand U15300 (N_15300,N_13282,N_13332);
and U15301 (N_15301,N_13758,N_13412);
nor U15302 (N_15302,N_12100,N_12312);
xor U15303 (N_15303,N_13290,N_12128);
and U15304 (N_15304,N_13995,N_13996);
xnor U15305 (N_15305,N_12184,N_13259);
xnor U15306 (N_15306,N_13057,N_12408);
or U15307 (N_15307,N_13693,N_12822);
nor U15308 (N_15308,N_13669,N_13004);
and U15309 (N_15309,N_12898,N_12285);
nand U15310 (N_15310,N_13111,N_13789);
xnor U15311 (N_15311,N_13623,N_12259);
nor U15312 (N_15312,N_12904,N_13014);
and U15313 (N_15313,N_12157,N_12209);
and U15314 (N_15314,N_13275,N_13038);
or U15315 (N_15315,N_12393,N_12903);
or U15316 (N_15316,N_12601,N_12732);
and U15317 (N_15317,N_12224,N_13529);
nor U15318 (N_15318,N_12225,N_12277);
nand U15319 (N_15319,N_12838,N_12561);
nor U15320 (N_15320,N_13237,N_12723);
and U15321 (N_15321,N_13510,N_13586);
nand U15322 (N_15322,N_13156,N_13200);
or U15323 (N_15323,N_12538,N_12895);
nand U15324 (N_15324,N_13064,N_12250);
nand U15325 (N_15325,N_12154,N_13617);
and U15326 (N_15326,N_13893,N_13236);
and U15327 (N_15327,N_12169,N_13713);
nor U15328 (N_15328,N_13041,N_13786);
nor U15329 (N_15329,N_13327,N_13865);
or U15330 (N_15330,N_12198,N_13389);
nor U15331 (N_15331,N_13940,N_12054);
and U15332 (N_15332,N_13360,N_13068);
and U15333 (N_15333,N_13283,N_12608);
or U15334 (N_15334,N_13682,N_12256);
xor U15335 (N_15335,N_13403,N_13194);
nand U15336 (N_15336,N_13270,N_13887);
xor U15337 (N_15337,N_12419,N_12402);
or U15338 (N_15338,N_12853,N_12340);
nor U15339 (N_15339,N_13840,N_13287);
or U15340 (N_15340,N_12703,N_12376);
and U15341 (N_15341,N_12091,N_13177);
nor U15342 (N_15342,N_12769,N_13646);
nor U15343 (N_15343,N_12852,N_12915);
and U15344 (N_15344,N_13449,N_12627);
and U15345 (N_15345,N_13727,N_12871);
nor U15346 (N_15346,N_13041,N_13457);
or U15347 (N_15347,N_13563,N_13074);
and U15348 (N_15348,N_13041,N_12832);
or U15349 (N_15349,N_13875,N_13135);
nor U15350 (N_15350,N_12381,N_13326);
nand U15351 (N_15351,N_13590,N_13466);
and U15352 (N_15352,N_12351,N_12659);
or U15353 (N_15353,N_13184,N_13914);
nor U15354 (N_15354,N_13675,N_12780);
and U15355 (N_15355,N_13279,N_13287);
xnor U15356 (N_15356,N_12740,N_13249);
and U15357 (N_15357,N_13899,N_13952);
xnor U15358 (N_15358,N_12819,N_12565);
or U15359 (N_15359,N_12109,N_13582);
nor U15360 (N_15360,N_13108,N_12755);
nand U15361 (N_15361,N_12408,N_13037);
or U15362 (N_15362,N_13179,N_13272);
and U15363 (N_15363,N_12623,N_13120);
nand U15364 (N_15364,N_12694,N_12565);
nand U15365 (N_15365,N_12803,N_13957);
nor U15366 (N_15366,N_13326,N_13856);
or U15367 (N_15367,N_12330,N_13301);
nor U15368 (N_15368,N_12865,N_13731);
nand U15369 (N_15369,N_12771,N_13723);
nor U15370 (N_15370,N_13832,N_12867);
nand U15371 (N_15371,N_13788,N_12707);
nand U15372 (N_15372,N_12707,N_13600);
and U15373 (N_15373,N_13315,N_12997);
xor U15374 (N_15374,N_13089,N_12170);
xor U15375 (N_15375,N_12610,N_13798);
and U15376 (N_15376,N_12281,N_12951);
nand U15377 (N_15377,N_13610,N_12778);
and U15378 (N_15378,N_13946,N_13830);
or U15379 (N_15379,N_13970,N_13549);
nand U15380 (N_15380,N_12938,N_13167);
or U15381 (N_15381,N_12580,N_12422);
nor U15382 (N_15382,N_13130,N_13026);
or U15383 (N_15383,N_12993,N_13872);
or U15384 (N_15384,N_12623,N_12862);
nor U15385 (N_15385,N_12174,N_12980);
nand U15386 (N_15386,N_13063,N_13916);
and U15387 (N_15387,N_13533,N_13687);
and U15388 (N_15388,N_13521,N_13592);
nand U15389 (N_15389,N_12843,N_12848);
nor U15390 (N_15390,N_13384,N_13687);
and U15391 (N_15391,N_13630,N_13418);
or U15392 (N_15392,N_12841,N_13122);
or U15393 (N_15393,N_13664,N_12237);
or U15394 (N_15394,N_13150,N_12173);
xor U15395 (N_15395,N_13928,N_13996);
xnor U15396 (N_15396,N_13987,N_13423);
nor U15397 (N_15397,N_13654,N_12535);
nand U15398 (N_15398,N_12046,N_12695);
nand U15399 (N_15399,N_13363,N_13961);
or U15400 (N_15400,N_12541,N_12559);
nand U15401 (N_15401,N_12975,N_12876);
or U15402 (N_15402,N_12343,N_13451);
and U15403 (N_15403,N_12703,N_13665);
nor U15404 (N_15404,N_13674,N_13444);
or U15405 (N_15405,N_12432,N_12198);
nor U15406 (N_15406,N_12516,N_12142);
nor U15407 (N_15407,N_13330,N_13859);
or U15408 (N_15408,N_13387,N_13270);
nand U15409 (N_15409,N_13187,N_12251);
and U15410 (N_15410,N_12102,N_13930);
or U15411 (N_15411,N_12029,N_12116);
xnor U15412 (N_15412,N_13385,N_12658);
and U15413 (N_15413,N_13228,N_12641);
or U15414 (N_15414,N_12100,N_12738);
nand U15415 (N_15415,N_12183,N_12120);
nor U15416 (N_15416,N_12456,N_12117);
nor U15417 (N_15417,N_13510,N_13089);
or U15418 (N_15418,N_13448,N_13658);
or U15419 (N_15419,N_13251,N_12223);
and U15420 (N_15420,N_13567,N_13893);
nand U15421 (N_15421,N_12203,N_12893);
and U15422 (N_15422,N_12870,N_13921);
xnor U15423 (N_15423,N_13010,N_13824);
or U15424 (N_15424,N_12051,N_12939);
or U15425 (N_15425,N_13834,N_12921);
xnor U15426 (N_15426,N_13017,N_12582);
and U15427 (N_15427,N_13272,N_12996);
nor U15428 (N_15428,N_12766,N_12333);
or U15429 (N_15429,N_13597,N_12758);
nor U15430 (N_15430,N_12376,N_12941);
xor U15431 (N_15431,N_12107,N_13328);
nor U15432 (N_15432,N_13464,N_13874);
nor U15433 (N_15433,N_13253,N_12038);
or U15434 (N_15434,N_13200,N_13868);
or U15435 (N_15435,N_13912,N_13213);
nor U15436 (N_15436,N_13977,N_13884);
nand U15437 (N_15437,N_12408,N_13952);
nor U15438 (N_15438,N_13489,N_12258);
or U15439 (N_15439,N_13589,N_13648);
and U15440 (N_15440,N_12299,N_12480);
or U15441 (N_15441,N_13256,N_12197);
xor U15442 (N_15442,N_12126,N_12950);
xnor U15443 (N_15443,N_13864,N_12374);
or U15444 (N_15444,N_12935,N_13419);
nor U15445 (N_15445,N_13119,N_13783);
or U15446 (N_15446,N_13366,N_12996);
and U15447 (N_15447,N_12370,N_13827);
nand U15448 (N_15448,N_13611,N_12422);
xor U15449 (N_15449,N_12870,N_12755);
xor U15450 (N_15450,N_12657,N_13112);
xor U15451 (N_15451,N_13631,N_12370);
xnor U15452 (N_15452,N_12020,N_13314);
nor U15453 (N_15453,N_12923,N_13845);
nor U15454 (N_15454,N_13875,N_13826);
and U15455 (N_15455,N_12815,N_12056);
and U15456 (N_15456,N_13972,N_12210);
nor U15457 (N_15457,N_12459,N_12811);
nand U15458 (N_15458,N_12313,N_13759);
and U15459 (N_15459,N_12011,N_13297);
xnor U15460 (N_15460,N_12649,N_12060);
xor U15461 (N_15461,N_13185,N_13059);
or U15462 (N_15462,N_12325,N_13394);
nand U15463 (N_15463,N_12497,N_13395);
or U15464 (N_15464,N_12239,N_13038);
nor U15465 (N_15465,N_12341,N_13536);
and U15466 (N_15466,N_12022,N_13700);
nor U15467 (N_15467,N_12866,N_13913);
and U15468 (N_15468,N_13055,N_12874);
xor U15469 (N_15469,N_12118,N_12508);
xor U15470 (N_15470,N_12186,N_13672);
nor U15471 (N_15471,N_12224,N_12622);
and U15472 (N_15472,N_12447,N_13751);
nand U15473 (N_15473,N_12735,N_13723);
or U15474 (N_15474,N_12098,N_13480);
or U15475 (N_15475,N_12124,N_13665);
or U15476 (N_15476,N_13239,N_12785);
nand U15477 (N_15477,N_12343,N_12618);
nor U15478 (N_15478,N_13566,N_12161);
and U15479 (N_15479,N_13889,N_13386);
nor U15480 (N_15480,N_13990,N_12071);
and U15481 (N_15481,N_13185,N_12791);
xnor U15482 (N_15482,N_12676,N_13745);
xor U15483 (N_15483,N_13638,N_13158);
nor U15484 (N_15484,N_12338,N_12155);
or U15485 (N_15485,N_12429,N_13488);
or U15486 (N_15486,N_12643,N_13238);
and U15487 (N_15487,N_13631,N_13624);
and U15488 (N_15488,N_12738,N_13137);
nand U15489 (N_15489,N_13930,N_13518);
nand U15490 (N_15490,N_12008,N_12038);
xnor U15491 (N_15491,N_12425,N_12750);
xor U15492 (N_15492,N_13690,N_13416);
or U15493 (N_15493,N_12920,N_13161);
or U15494 (N_15494,N_12992,N_13757);
nor U15495 (N_15495,N_12811,N_12595);
nand U15496 (N_15496,N_13541,N_12836);
or U15497 (N_15497,N_13829,N_12813);
or U15498 (N_15498,N_13598,N_12299);
xor U15499 (N_15499,N_13261,N_13651);
nor U15500 (N_15500,N_13031,N_12728);
xnor U15501 (N_15501,N_12671,N_12801);
and U15502 (N_15502,N_13167,N_13270);
and U15503 (N_15503,N_12603,N_12467);
or U15504 (N_15504,N_12855,N_12460);
and U15505 (N_15505,N_13856,N_13963);
or U15506 (N_15506,N_13864,N_12086);
nand U15507 (N_15507,N_13505,N_12810);
and U15508 (N_15508,N_13829,N_13804);
nor U15509 (N_15509,N_13368,N_13297);
nand U15510 (N_15510,N_12305,N_12841);
and U15511 (N_15511,N_13309,N_12913);
nor U15512 (N_15512,N_12608,N_13407);
nand U15513 (N_15513,N_12464,N_13793);
xnor U15514 (N_15514,N_13550,N_13714);
nor U15515 (N_15515,N_12566,N_13075);
nor U15516 (N_15516,N_12217,N_12469);
and U15517 (N_15517,N_12044,N_13166);
xor U15518 (N_15518,N_13018,N_13869);
nor U15519 (N_15519,N_13236,N_13378);
nand U15520 (N_15520,N_12717,N_13306);
nand U15521 (N_15521,N_13175,N_13922);
and U15522 (N_15522,N_13776,N_12157);
and U15523 (N_15523,N_12144,N_12323);
xor U15524 (N_15524,N_12969,N_12856);
and U15525 (N_15525,N_13698,N_13161);
or U15526 (N_15526,N_12642,N_12984);
nor U15527 (N_15527,N_12455,N_13814);
nor U15528 (N_15528,N_13260,N_13180);
or U15529 (N_15529,N_12350,N_13995);
nand U15530 (N_15530,N_12107,N_12512);
xor U15531 (N_15531,N_13721,N_13339);
nor U15532 (N_15532,N_13551,N_12313);
or U15533 (N_15533,N_12186,N_12996);
or U15534 (N_15534,N_13608,N_13698);
or U15535 (N_15535,N_12347,N_12403);
nand U15536 (N_15536,N_12886,N_12868);
nor U15537 (N_15537,N_12104,N_13768);
nor U15538 (N_15538,N_12407,N_13057);
or U15539 (N_15539,N_12012,N_13146);
nand U15540 (N_15540,N_12432,N_12828);
or U15541 (N_15541,N_12067,N_13467);
and U15542 (N_15542,N_12426,N_12353);
nand U15543 (N_15543,N_13602,N_13898);
and U15544 (N_15544,N_13039,N_12329);
and U15545 (N_15545,N_13400,N_12104);
nor U15546 (N_15546,N_12833,N_13302);
and U15547 (N_15547,N_12794,N_12089);
nand U15548 (N_15548,N_12881,N_13559);
nand U15549 (N_15549,N_13701,N_12071);
and U15550 (N_15550,N_13198,N_13322);
or U15551 (N_15551,N_13106,N_13196);
xor U15552 (N_15552,N_12091,N_12172);
or U15553 (N_15553,N_12639,N_12940);
nand U15554 (N_15554,N_12633,N_13794);
nor U15555 (N_15555,N_13834,N_12159);
xnor U15556 (N_15556,N_12415,N_12341);
nor U15557 (N_15557,N_13017,N_13255);
or U15558 (N_15558,N_13563,N_12883);
nand U15559 (N_15559,N_12026,N_13897);
or U15560 (N_15560,N_13298,N_12172);
and U15561 (N_15561,N_12794,N_12966);
xnor U15562 (N_15562,N_13951,N_13475);
and U15563 (N_15563,N_12885,N_12246);
or U15564 (N_15564,N_13171,N_13450);
and U15565 (N_15565,N_12312,N_13754);
or U15566 (N_15566,N_12427,N_12356);
nand U15567 (N_15567,N_12866,N_12475);
or U15568 (N_15568,N_13638,N_13834);
and U15569 (N_15569,N_12117,N_13040);
and U15570 (N_15570,N_12889,N_13129);
nor U15571 (N_15571,N_12354,N_13249);
or U15572 (N_15572,N_12652,N_12764);
or U15573 (N_15573,N_12882,N_13315);
xor U15574 (N_15574,N_12891,N_12170);
and U15575 (N_15575,N_13085,N_12682);
nor U15576 (N_15576,N_12542,N_13037);
xnor U15577 (N_15577,N_13649,N_13724);
nand U15578 (N_15578,N_13326,N_12412);
nor U15579 (N_15579,N_12972,N_13575);
xnor U15580 (N_15580,N_13010,N_12560);
nor U15581 (N_15581,N_13469,N_13452);
xnor U15582 (N_15582,N_13579,N_13771);
xor U15583 (N_15583,N_12877,N_13412);
or U15584 (N_15584,N_13777,N_13203);
nand U15585 (N_15585,N_12425,N_13314);
nand U15586 (N_15586,N_13243,N_13612);
and U15587 (N_15587,N_12849,N_12679);
and U15588 (N_15588,N_12644,N_13161);
or U15589 (N_15589,N_12204,N_12698);
nor U15590 (N_15590,N_12445,N_12449);
nor U15591 (N_15591,N_13103,N_13058);
xnor U15592 (N_15592,N_12785,N_12183);
nand U15593 (N_15593,N_13052,N_12351);
or U15594 (N_15594,N_13546,N_13624);
nor U15595 (N_15595,N_13736,N_13441);
nor U15596 (N_15596,N_12981,N_13589);
xnor U15597 (N_15597,N_12718,N_13339);
nand U15598 (N_15598,N_12091,N_12823);
or U15599 (N_15599,N_13474,N_13182);
and U15600 (N_15600,N_13234,N_13384);
nand U15601 (N_15601,N_13767,N_13279);
or U15602 (N_15602,N_12140,N_13031);
xor U15603 (N_15603,N_13673,N_12430);
nand U15604 (N_15604,N_12207,N_13094);
nor U15605 (N_15605,N_12753,N_13434);
nand U15606 (N_15606,N_12271,N_13671);
nand U15607 (N_15607,N_13994,N_12212);
nand U15608 (N_15608,N_13961,N_12170);
nor U15609 (N_15609,N_13918,N_13267);
xnor U15610 (N_15610,N_13499,N_12722);
nand U15611 (N_15611,N_12738,N_12930);
xnor U15612 (N_15612,N_12450,N_12647);
and U15613 (N_15613,N_13294,N_12297);
xnor U15614 (N_15614,N_12465,N_12605);
nand U15615 (N_15615,N_13322,N_13496);
xnor U15616 (N_15616,N_13528,N_12908);
and U15617 (N_15617,N_13111,N_13604);
nor U15618 (N_15618,N_13821,N_12292);
xnor U15619 (N_15619,N_13066,N_13334);
or U15620 (N_15620,N_12373,N_12854);
and U15621 (N_15621,N_12213,N_12768);
and U15622 (N_15622,N_13090,N_12894);
nor U15623 (N_15623,N_12468,N_13083);
xnor U15624 (N_15624,N_13069,N_12044);
xnor U15625 (N_15625,N_13844,N_13100);
and U15626 (N_15626,N_13440,N_13713);
xor U15627 (N_15627,N_13176,N_12167);
nand U15628 (N_15628,N_12768,N_12338);
and U15629 (N_15629,N_12313,N_13455);
xor U15630 (N_15630,N_12673,N_12345);
nor U15631 (N_15631,N_12198,N_13551);
or U15632 (N_15632,N_13245,N_13211);
nand U15633 (N_15633,N_12214,N_12023);
or U15634 (N_15634,N_13066,N_13979);
and U15635 (N_15635,N_13217,N_13687);
and U15636 (N_15636,N_12637,N_12429);
or U15637 (N_15637,N_12723,N_12037);
xor U15638 (N_15638,N_12147,N_13211);
and U15639 (N_15639,N_13349,N_13684);
and U15640 (N_15640,N_13484,N_13102);
nand U15641 (N_15641,N_13538,N_13949);
xor U15642 (N_15642,N_13206,N_12421);
nor U15643 (N_15643,N_12282,N_12523);
nor U15644 (N_15644,N_13617,N_12511);
or U15645 (N_15645,N_13087,N_13780);
nand U15646 (N_15646,N_13707,N_13317);
nor U15647 (N_15647,N_12784,N_13612);
xnor U15648 (N_15648,N_13494,N_12563);
and U15649 (N_15649,N_13804,N_12158);
nor U15650 (N_15650,N_12157,N_13117);
nor U15651 (N_15651,N_13804,N_13338);
nor U15652 (N_15652,N_13650,N_12727);
nor U15653 (N_15653,N_13334,N_12821);
or U15654 (N_15654,N_13186,N_13362);
and U15655 (N_15655,N_13129,N_12905);
and U15656 (N_15656,N_12890,N_13122);
or U15657 (N_15657,N_13260,N_12788);
xor U15658 (N_15658,N_12045,N_13564);
nand U15659 (N_15659,N_12186,N_12580);
nor U15660 (N_15660,N_12971,N_12241);
and U15661 (N_15661,N_13138,N_13605);
and U15662 (N_15662,N_13477,N_13873);
xor U15663 (N_15663,N_12338,N_13187);
and U15664 (N_15664,N_13869,N_12388);
or U15665 (N_15665,N_12152,N_13200);
and U15666 (N_15666,N_13546,N_13523);
nor U15667 (N_15667,N_13723,N_12307);
nor U15668 (N_15668,N_13883,N_13285);
and U15669 (N_15669,N_12604,N_12667);
nand U15670 (N_15670,N_12405,N_13877);
and U15671 (N_15671,N_12890,N_13205);
nand U15672 (N_15672,N_13225,N_12221);
xor U15673 (N_15673,N_12059,N_13464);
xor U15674 (N_15674,N_12818,N_12728);
xnor U15675 (N_15675,N_12456,N_12179);
or U15676 (N_15676,N_12990,N_13501);
or U15677 (N_15677,N_12669,N_12577);
and U15678 (N_15678,N_12628,N_13615);
xor U15679 (N_15679,N_12207,N_13977);
nor U15680 (N_15680,N_12292,N_12537);
nor U15681 (N_15681,N_13625,N_12936);
and U15682 (N_15682,N_12034,N_13322);
nor U15683 (N_15683,N_12559,N_12569);
xnor U15684 (N_15684,N_13113,N_13409);
or U15685 (N_15685,N_12310,N_12046);
xor U15686 (N_15686,N_13802,N_13466);
or U15687 (N_15687,N_13735,N_13381);
xnor U15688 (N_15688,N_12336,N_12813);
and U15689 (N_15689,N_13011,N_13136);
xnor U15690 (N_15690,N_12549,N_12961);
nand U15691 (N_15691,N_12084,N_12711);
and U15692 (N_15692,N_13151,N_13601);
and U15693 (N_15693,N_12115,N_13993);
nand U15694 (N_15694,N_13672,N_12178);
nand U15695 (N_15695,N_13545,N_13862);
or U15696 (N_15696,N_12390,N_13816);
nand U15697 (N_15697,N_13744,N_12176);
nor U15698 (N_15698,N_12497,N_12526);
nor U15699 (N_15699,N_12211,N_13152);
or U15700 (N_15700,N_12191,N_12201);
nand U15701 (N_15701,N_13583,N_13288);
and U15702 (N_15702,N_13627,N_13898);
xor U15703 (N_15703,N_12971,N_13831);
or U15704 (N_15704,N_13039,N_13387);
nand U15705 (N_15705,N_13535,N_12011);
and U15706 (N_15706,N_13314,N_12785);
xor U15707 (N_15707,N_13442,N_13167);
xnor U15708 (N_15708,N_13052,N_13681);
and U15709 (N_15709,N_12217,N_13507);
nor U15710 (N_15710,N_13389,N_12781);
and U15711 (N_15711,N_12719,N_12381);
and U15712 (N_15712,N_13496,N_12003);
and U15713 (N_15713,N_13352,N_12617);
or U15714 (N_15714,N_13241,N_13724);
and U15715 (N_15715,N_12036,N_12775);
or U15716 (N_15716,N_13075,N_13715);
or U15717 (N_15717,N_12469,N_13142);
or U15718 (N_15718,N_13290,N_12956);
and U15719 (N_15719,N_12969,N_13145);
nand U15720 (N_15720,N_12793,N_12729);
or U15721 (N_15721,N_13621,N_13944);
or U15722 (N_15722,N_12918,N_12192);
and U15723 (N_15723,N_12633,N_13516);
nand U15724 (N_15724,N_12715,N_12516);
and U15725 (N_15725,N_12877,N_13616);
xor U15726 (N_15726,N_13874,N_12575);
nand U15727 (N_15727,N_13907,N_12255);
xor U15728 (N_15728,N_12369,N_13095);
nand U15729 (N_15729,N_13170,N_13163);
nand U15730 (N_15730,N_13487,N_12423);
nor U15731 (N_15731,N_12155,N_13055);
nor U15732 (N_15732,N_13172,N_13001);
nand U15733 (N_15733,N_12116,N_12177);
xor U15734 (N_15734,N_13294,N_13048);
nor U15735 (N_15735,N_12406,N_13695);
xnor U15736 (N_15736,N_12253,N_13880);
nand U15737 (N_15737,N_12927,N_13843);
xnor U15738 (N_15738,N_12089,N_13089);
and U15739 (N_15739,N_13434,N_12589);
or U15740 (N_15740,N_13241,N_13807);
or U15741 (N_15741,N_13147,N_12347);
and U15742 (N_15742,N_13418,N_13542);
xor U15743 (N_15743,N_13992,N_13076);
nand U15744 (N_15744,N_12300,N_13703);
nand U15745 (N_15745,N_12244,N_12975);
and U15746 (N_15746,N_13346,N_13134);
or U15747 (N_15747,N_13414,N_13856);
xor U15748 (N_15748,N_13112,N_12648);
or U15749 (N_15749,N_13850,N_13359);
nand U15750 (N_15750,N_13113,N_13243);
and U15751 (N_15751,N_13877,N_13852);
or U15752 (N_15752,N_12623,N_13923);
nand U15753 (N_15753,N_12530,N_13618);
nor U15754 (N_15754,N_12713,N_12546);
xnor U15755 (N_15755,N_12460,N_13657);
nor U15756 (N_15756,N_13509,N_12051);
xor U15757 (N_15757,N_13307,N_13593);
or U15758 (N_15758,N_13101,N_12903);
and U15759 (N_15759,N_13945,N_13448);
nand U15760 (N_15760,N_13121,N_13769);
or U15761 (N_15761,N_13422,N_12548);
or U15762 (N_15762,N_13457,N_12567);
or U15763 (N_15763,N_13608,N_12567);
and U15764 (N_15764,N_13298,N_13497);
or U15765 (N_15765,N_13354,N_13585);
or U15766 (N_15766,N_13939,N_12985);
and U15767 (N_15767,N_13432,N_13840);
xnor U15768 (N_15768,N_12837,N_13099);
nor U15769 (N_15769,N_12216,N_12093);
or U15770 (N_15770,N_13960,N_13592);
nor U15771 (N_15771,N_12687,N_13447);
nand U15772 (N_15772,N_13736,N_12140);
nor U15773 (N_15773,N_12201,N_13994);
or U15774 (N_15774,N_13029,N_13837);
and U15775 (N_15775,N_13021,N_12361);
nand U15776 (N_15776,N_12059,N_13358);
nor U15777 (N_15777,N_13746,N_13335);
nor U15778 (N_15778,N_13285,N_13809);
and U15779 (N_15779,N_13076,N_13392);
nand U15780 (N_15780,N_13842,N_12783);
xor U15781 (N_15781,N_13398,N_13776);
xnor U15782 (N_15782,N_13841,N_12563);
nand U15783 (N_15783,N_13726,N_12253);
xor U15784 (N_15784,N_13189,N_12187);
xor U15785 (N_15785,N_13387,N_12272);
xor U15786 (N_15786,N_12240,N_12596);
nand U15787 (N_15787,N_13562,N_13308);
nand U15788 (N_15788,N_12508,N_12364);
xor U15789 (N_15789,N_12708,N_13013);
and U15790 (N_15790,N_12848,N_13204);
and U15791 (N_15791,N_13799,N_12417);
xor U15792 (N_15792,N_12090,N_12928);
xnor U15793 (N_15793,N_12620,N_12130);
xor U15794 (N_15794,N_12701,N_12035);
xor U15795 (N_15795,N_12271,N_12242);
nor U15796 (N_15796,N_12987,N_13962);
nor U15797 (N_15797,N_12820,N_13573);
or U15798 (N_15798,N_12044,N_13714);
xnor U15799 (N_15799,N_12004,N_12275);
nand U15800 (N_15800,N_12764,N_13370);
nor U15801 (N_15801,N_12379,N_13336);
nand U15802 (N_15802,N_13375,N_13516);
and U15803 (N_15803,N_12496,N_12353);
and U15804 (N_15804,N_12907,N_13591);
nand U15805 (N_15805,N_13076,N_13802);
xnor U15806 (N_15806,N_13621,N_13172);
xnor U15807 (N_15807,N_12943,N_13914);
xor U15808 (N_15808,N_13794,N_12651);
nand U15809 (N_15809,N_13686,N_13400);
and U15810 (N_15810,N_12855,N_13540);
or U15811 (N_15811,N_13068,N_13270);
nand U15812 (N_15812,N_12147,N_12581);
and U15813 (N_15813,N_13257,N_12498);
xor U15814 (N_15814,N_13388,N_13154);
and U15815 (N_15815,N_12992,N_12994);
or U15816 (N_15816,N_13364,N_13932);
or U15817 (N_15817,N_13286,N_12361);
nand U15818 (N_15818,N_13960,N_13393);
nor U15819 (N_15819,N_13482,N_12221);
and U15820 (N_15820,N_13675,N_12202);
nand U15821 (N_15821,N_12960,N_13319);
nand U15822 (N_15822,N_12280,N_13127);
and U15823 (N_15823,N_13701,N_12000);
and U15824 (N_15824,N_12097,N_13270);
nor U15825 (N_15825,N_12923,N_12394);
nor U15826 (N_15826,N_12287,N_13558);
nand U15827 (N_15827,N_13167,N_13295);
xnor U15828 (N_15828,N_12834,N_13902);
nand U15829 (N_15829,N_13868,N_13847);
and U15830 (N_15830,N_13625,N_12609);
or U15831 (N_15831,N_13164,N_12264);
nor U15832 (N_15832,N_13870,N_12993);
or U15833 (N_15833,N_12564,N_12591);
and U15834 (N_15834,N_12169,N_12136);
or U15835 (N_15835,N_13291,N_13966);
nand U15836 (N_15836,N_13701,N_12024);
or U15837 (N_15837,N_13934,N_12530);
and U15838 (N_15838,N_13633,N_12139);
or U15839 (N_15839,N_12624,N_12760);
or U15840 (N_15840,N_12988,N_12511);
and U15841 (N_15841,N_12400,N_12551);
nor U15842 (N_15842,N_12467,N_13498);
nand U15843 (N_15843,N_13074,N_12816);
nand U15844 (N_15844,N_13517,N_12612);
nor U15845 (N_15845,N_12973,N_12355);
or U15846 (N_15846,N_13134,N_13030);
or U15847 (N_15847,N_12638,N_13327);
nand U15848 (N_15848,N_13574,N_12626);
or U15849 (N_15849,N_13071,N_12138);
or U15850 (N_15850,N_12189,N_13546);
xor U15851 (N_15851,N_13762,N_12524);
and U15852 (N_15852,N_12680,N_12868);
xnor U15853 (N_15853,N_12955,N_12561);
nor U15854 (N_15854,N_13816,N_13654);
and U15855 (N_15855,N_12302,N_13886);
nor U15856 (N_15856,N_13399,N_13004);
and U15857 (N_15857,N_13904,N_12653);
or U15858 (N_15858,N_13493,N_13078);
or U15859 (N_15859,N_12544,N_12976);
xor U15860 (N_15860,N_13621,N_13014);
xnor U15861 (N_15861,N_13773,N_13559);
nand U15862 (N_15862,N_13603,N_12706);
xor U15863 (N_15863,N_12565,N_12850);
or U15864 (N_15864,N_12704,N_13282);
nor U15865 (N_15865,N_12568,N_13207);
xnor U15866 (N_15866,N_12855,N_13155);
xnor U15867 (N_15867,N_13301,N_12480);
xor U15868 (N_15868,N_13412,N_13349);
nand U15869 (N_15869,N_13089,N_13188);
xnor U15870 (N_15870,N_13581,N_13983);
nand U15871 (N_15871,N_12034,N_13117);
nor U15872 (N_15872,N_13602,N_13062);
nor U15873 (N_15873,N_12679,N_13761);
xnor U15874 (N_15874,N_13486,N_12549);
nand U15875 (N_15875,N_13733,N_13593);
or U15876 (N_15876,N_13119,N_13361);
or U15877 (N_15877,N_13205,N_13515);
and U15878 (N_15878,N_12804,N_12930);
and U15879 (N_15879,N_12793,N_12600);
xnor U15880 (N_15880,N_12792,N_13126);
nand U15881 (N_15881,N_13371,N_12260);
or U15882 (N_15882,N_13346,N_12471);
nand U15883 (N_15883,N_12897,N_12584);
and U15884 (N_15884,N_13368,N_13416);
nor U15885 (N_15885,N_12445,N_12524);
and U15886 (N_15886,N_12465,N_12175);
xnor U15887 (N_15887,N_13030,N_13753);
xnor U15888 (N_15888,N_12454,N_12177);
or U15889 (N_15889,N_12841,N_13512);
nand U15890 (N_15890,N_12520,N_13598);
xnor U15891 (N_15891,N_12043,N_13911);
and U15892 (N_15892,N_13452,N_13985);
and U15893 (N_15893,N_12133,N_12963);
nor U15894 (N_15894,N_13151,N_13204);
or U15895 (N_15895,N_12535,N_12114);
or U15896 (N_15896,N_12923,N_12859);
nand U15897 (N_15897,N_13980,N_12052);
xnor U15898 (N_15898,N_12606,N_12823);
nor U15899 (N_15899,N_12154,N_13275);
nor U15900 (N_15900,N_13848,N_12289);
nand U15901 (N_15901,N_13770,N_13109);
and U15902 (N_15902,N_12744,N_13954);
xor U15903 (N_15903,N_12355,N_12196);
or U15904 (N_15904,N_13491,N_13169);
nand U15905 (N_15905,N_13497,N_13990);
xor U15906 (N_15906,N_13122,N_13809);
nand U15907 (N_15907,N_13237,N_13137);
or U15908 (N_15908,N_12153,N_12720);
nand U15909 (N_15909,N_13555,N_13178);
or U15910 (N_15910,N_13013,N_13576);
xor U15911 (N_15911,N_12070,N_12336);
or U15912 (N_15912,N_12633,N_13627);
nor U15913 (N_15913,N_12576,N_12649);
or U15914 (N_15914,N_13661,N_12603);
nor U15915 (N_15915,N_12870,N_13936);
nor U15916 (N_15916,N_12887,N_12472);
or U15917 (N_15917,N_12278,N_12419);
and U15918 (N_15918,N_12325,N_12040);
xnor U15919 (N_15919,N_12229,N_13384);
or U15920 (N_15920,N_12846,N_13302);
xor U15921 (N_15921,N_12906,N_12184);
or U15922 (N_15922,N_13520,N_13702);
xor U15923 (N_15923,N_12282,N_13485);
xnor U15924 (N_15924,N_13386,N_13012);
nand U15925 (N_15925,N_13643,N_13160);
and U15926 (N_15926,N_12033,N_13740);
xor U15927 (N_15927,N_13325,N_12909);
or U15928 (N_15928,N_12554,N_12388);
xnor U15929 (N_15929,N_12634,N_12264);
nor U15930 (N_15930,N_12337,N_12611);
xor U15931 (N_15931,N_12841,N_13846);
xor U15932 (N_15932,N_12940,N_12433);
xnor U15933 (N_15933,N_12555,N_12557);
nor U15934 (N_15934,N_12619,N_12991);
and U15935 (N_15935,N_12895,N_13014);
nor U15936 (N_15936,N_12407,N_12188);
xnor U15937 (N_15937,N_13387,N_12755);
and U15938 (N_15938,N_13401,N_13479);
nand U15939 (N_15939,N_12279,N_13230);
and U15940 (N_15940,N_12506,N_12390);
and U15941 (N_15941,N_13458,N_13104);
xnor U15942 (N_15942,N_12463,N_12926);
xnor U15943 (N_15943,N_12188,N_12893);
nand U15944 (N_15944,N_12612,N_12619);
nand U15945 (N_15945,N_12078,N_12836);
and U15946 (N_15946,N_12032,N_13328);
xnor U15947 (N_15947,N_13340,N_12723);
nand U15948 (N_15948,N_12770,N_13606);
and U15949 (N_15949,N_13655,N_12767);
xor U15950 (N_15950,N_12923,N_12678);
xnor U15951 (N_15951,N_12106,N_13440);
xor U15952 (N_15952,N_13653,N_12060);
and U15953 (N_15953,N_13823,N_13068);
or U15954 (N_15954,N_12223,N_13489);
nand U15955 (N_15955,N_13484,N_13167);
and U15956 (N_15956,N_12909,N_13746);
and U15957 (N_15957,N_12099,N_12575);
xor U15958 (N_15958,N_12241,N_13677);
nor U15959 (N_15959,N_12439,N_13618);
nand U15960 (N_15960,N_13451,N_13030);
nand U15961 (N_15961,N_12933,N_12989);
and U15962 (N_15962,N_12877,N_12405);
nor U15963 (N_15963,N_12679,N_13739);
and U15964 (N_15964,N_13991,N_13635);
or U15965 (N_15965,N_13960,N_13346);
nand U15966 (N_15966,N_12494,N_12590);
or U15967 (N_15967,N_13023,N_12900);
and U15968 (N_15968,N_12153,N_13225);
nand U15969 (N_15969,N_13197,N_13951);
nand U15970 (N_15970,N_13369,N_12066);
xor U15971 (N_15971,N_13609,N_12661);
and U15972 (N_15972,N_13199,N_13228);
nor U15973 (N_15973,N_12695,N_12521);
or U15974 (N_15974,N_13985,N_12224);
nor U15975 (N_15975,N_13232,N_13654);
xor U15976 (N_15976,N_13605,N_12788);
or U15977 (N_15977,N_12783,N_12117);
or U15978 (N_15978,N_13176,N_12659);
and U15979 (N_15979,N_13898,N_13949);
and U15980 (N_15980,N_13226,N_12632);
nor U15981 (N_15981,N_12818,N_13108);
xnor U15982 (N_15982,N_12104,N_12907);
or U15983 (N_15983,N_13381,N_12818);
or U15984 (N_15984,N_13539,N_12165);
nand U15985 (N_15985,N_12461,N_12228);
nor U15986 (N_15986,N_13654,N_13046);
or U15987 (N_15987,N_12121,N_12103);
or U15988 (N_15988,N_12010,N_13742);
xor U15989 (N_15989,N_12062,N_13525);
or U15990 (N_15990,N_12853,N_12747);
or U15991 (N_15991,N_12293,N_13302);
nor U15992 (N_15992,N_12826,N_13773);
and U15993 (N_15993,N_13171,N_13036);
xor U15994 (N_15994,N_12182,N_12687);
nand U15995 (N_15995,N_13461,N_13967);
xor U15996 (N_15996,N_13573,N_13645);
nand U15997 (N_15997,N_12056,N_12036);
xor U15998 (N_15998,N_13565,N_13686);
nand U15999 (N_15999,N_12741,N_13139);
and U16000 (N_16000,N_15356,N_15308);
or U16001 (N_16001,N_14887,N_14404);
and U16002 (N_16002,N_14791,N_15320);
and U16003 (N_16003,N_15892,N_14129);
nand U16004 (N_16004,N_14581,N_14606);
or U16005 (N_16005,N_14039,N_14910);
xnor U16006 (N_16006,N_15298,N_14725);
xnor U16007 (N_16007,N_14455,N_14999);
nand U16008 (N_16008,N_14665,N_14403);
nor U16009 (N_16009,N_14584,N_15691);
and U16010 (N_16010,N_14079,N_14456);
and U16011 (N_16011,N_14257,N_14513);
nor U16012 (N_16012,N_14767,N_15056);
or U16013 (N_16013,N_15515,N_14476);
nor U16014 (N_16014,N_14831,N_15381);
and U16015 (N_16015,N_14097,N_15879);
or U16016 (N_16016,N_14934,N_15862);
and U16017 (N_16017,N_14422,N_15583);
nand U16018 (N_16018,N_15251,N_14912);
or U16019 (N_16019,N_14120,N_14130);
nand U16020 (N_16020,N_15528,N_14571);
xor U16021 (N_16021,N_14537,N_14304);
nand U16022 (N_16022,N_15058,N_15881);
and U16023 (N_16023,N_15970,N_14516);
and U16024 (N_16024,N_14994,N_14902);
xnor U16025 (N_16025,N_15947,N_14405);
nor U16026 (N_16026,N_15034,N_15632);
nor U16027 (N_16027,N_14534,N_14815);
xnor U16028 (N_16028,N_15804,N_14260);
or U16029 (N_16029,N_14917,N_14427);
and U16030 (N_16030,N_15309,N_14923);
or U16031 (N_16031,N_14166,N_15290);
and U16032 (N_16032,N_15452,N_15702);
nor U16033 (N_16033,N_14546,N_14685);
xnor U16034 (N_16034,N_15374,N_15730);
xor U16035 (N_16035,N_14470,N_15326);
xnor U16036 (N_16036,N_15018,N_14245);
nor U16037 (N_16037,N_15624,N_14701);
and U16038 (N_16038,N_15194,N_15030);
nor U16039 (N_16039,N_14749,N_14351);
nand U16040 (N_16040,N_15671,N_15407);
xor U16041 (N_16041,N_15650,N_15176);
nand U16042 (N_16042,N_15763,N_15753);
nor U16043 (N_16043,N_15435,N_15080);
nand U16044 (N_16044,N_14515,N_15684);
xor U16045 (N_16045,N_14191,N_15395);
or U16046 (N_16046,N_15443,N_15111);
nand U16047 (N_16047,N_14609,N_14564);
and U16048 (N_16048,N_14909,N_15346);
xor U16049 (N_16049,N_14291,N_15166);
and U16050 (N_16050,N_15835,N_15504);
nand U16051 (N_16051,N_15561,N_14213);
xor U16052 (N_16052,N_15483,N_15345);
nor U16053 (N_16053,N_15061,N_14635);
nor U16054 (N_16054,N_15682,N_15066);
and U16055 (N_16055,N_15226,N_15805);
nor U16056 (N_16056,N_15826,N_14139);
or U16057 (N_16057,N_14598,N_14179);
and U16058 (N_16058,N_15410,N_14349);
and U16059 (N_16059,N_15943,N_14672);
or U16060 (N_16060,N_14886,N_15453);
nor U16061 (N_16061,N_14919,N_15052);
xor U16062 (N_16062,N_14868,N_14880);
or U16063 (N_16063,N_14094,N_14849);
and U16064 (N_16064,N_14223,N_14485);
xor U16065 (N_16065,N_14569,N_14484);
or U16066 (N_16066,N_15225,N_15797);
xnor U16067 (N_16067,N_14420,N_14595);
and U16068 (N_16068,N_14864,N_15032);
xor U16069 (N_16069,N_15602,N_15460);
and U16070 (N_16070,N_14350,N_15084);
nor U16071 (N_16071,N_14675,N_15690);
or U16072 (N_16072,N_15623,N_14463);
xnor U16073 (N_16073,N_15422,N_15743);
xnor U16074 (N_16074,N_15161,N_15289);
xnor U16075 (N_16075,N_15609,N_14652);
xnor U16076 (N_16076,N_15698,N_15924);
nand U16077 (N_16077,N_14861,N_14242);
or U16078 (N_16078,N_14222,N_15649);
and U16079 (N_16079,N_14268,N_14826);
and U16080 (N_16080,N_15051,N_14360);
and U16081 (N_16081,N_15180,N_14765);
nand U16082 (N_16082,N_14869,N_15020);
or U16083 (N_16083,N_14807,N_14804);
nor U16084 (N_16084,N_14353,N_15488);
nor U16085 (N_16085,N_14649,N_15704);
xnor U16086 (N_16086,N_15847,N_14981);
and U16087 (N_16087,N_15096,N_14611);
or U16088 (N_16088,N_15431,N_15342);
nor U16089 (N_16089,N_15614,N_15127);
or U16090 (N_16090,N_14036,N_14789);
nand U16091 (N_16091,N_14633,N_15503);
nand U16092 (N_16092,N_15575,N_14644);
nand U16093 (N_16093,N_14095,N_14107);
xor U16094 (N_16094,N_14338,N_15105);
or U16095 (N_16095,N_15274,N_14785);
nor U16096 (N_16096,N_15249,N_15604);
and U16097 (N_16097,N_15037,N_14555);
nor U16098 (N_16098,N_14916,N_14385);
and U16099 (N_16099,N_15258,N_15792);
and U16100 (N_16100,N_14946,N_15386);
xor U16101 (N_16101,N_14751,N_14339);
or U16102 (N_16102,N_14656,N_15198);
xnor U16103 (N_16103,N_15236,N_14173);
xor U16104 (N_16104,N_15578,N_15424);
or U16105 (N_16105,N_15736,N_15855);
xnor U16106 (N_16106,N_14823,N_15116);
and U16107 (N_16107,N_15134,N_15783);
and U16108 (N_16108,N_15364,N_14926);
or U16109 (N_16109,N_14828,N_14706);
or U16110 (N_16110,N_14538,N_14871);
nand U16111 (N_16111,N_15551,N_15284);
nand U16112 (N_16112,N_14400,N_14276);
nand U16113 (N_16113,N_15762,N_14745);
or U16114 (N_16114,N_15789,N_15667);
nor U16115 (N_16115,N_15296,N_15715);
nor U16116 (N_16116,N_15574,N_14145);
nand U16117 (N_16117,N_15206,N_15347);
and U16118 (N_16118,N_14763,N_15843);
nand U16119 (N_16119,N_14087,N_14881);
nor U16120 (N_16120,N_14956,N_15660);
or U16121 (N_16121,N_14592,N_15800);
nand U16122 (N_16122,N_14048,N_14387);
xnor U16123 (N_16123,N_15746,N_14374);
and U16124 (N_16124,N_15509,N_15669);
nor U16125 (N_16125,N_14324,N_15335);
or U16126 (N_16126,N_14272,N_14773);
or U16127 (N_16127,N_15268,N_14188);
nand U16128 (N_16128,N_14195,N_14068);
and U16129 (N_16129,N_14168,N_14215);
nand U16130 (N_16130,N_14895,N_14972);
nor U16131 (N_16131,N_14281,N_15190);
or U16132 (N_16132,N_14838,N_14174);
and U16133 (N_16133,N_15982,N_14586);
nor U16134 (N_16134,N_14110,N_15189);
xnor U16135 (N_16135,N_14551,N_14529);
nand U16136 (N_16136,N_15334,N_15617);
xor U16137 (N_16137,N_14875,N_15586);
and U16138 (N_16138,N_15240,N_14704);
nor U16139 (N_16139,N_15067,N_15007);
nand U16140 (N_16140,N_14983,N_15998);
xnor U16141 (N_16141,N_14031,N_15780);
nand U16142 (N_16142,N_14090,N_14713);
nand U16143 (N_16143,N_15670,N_14348);
and U16144 (N_16144,N_15512,N_14066);
nand U16145 (N_16145,N_15192,N_15566);
nand U16146 (N_16146,N_14140,N_14892);
nand U16147 (N_16147,N_14311,N_14296);
nor U16148 (N_16148,N_14793,N_14820);
or U16149 (N_16149,N_15465,N_14734);
and U16150 (N_16150,N_14308,N_15295);
xor U16151 (N_16151,N_14002,N_14993);
or U16152 (N_16152,N_15112,N_15680);
nand U16153 (N_16153,N_14459,N_15491);
nor U16154 (N_16154,N_14824,N_14677);
nand U16155 (N_16155,N_14716,N_15960);
xnor U16156 (N_16156,N_15215,N_14949);
and U16157 (N_16157,N_15315,N_15338);
nor U16158 (N_16158,N_15014,N_15807);
nor U16159 (N_16159,N_14426,N_15956);
nor U16160 (N_16160,N_15462,N_15911);
nand U16161 (N_16161,N_15310,N_15322);
nor U16162 (N_16162,N_15776,N_15884);
nor U16163 (N_16163,N_15729,N_14358);
and U16164 (N_16164,N_15177,N_15380);
or U16165 (N_16165,N_15661,N_14444);
xor U16166 (N_16166,N_15477,N_14844);
and U16167 (N_16167,N_15203,N_15328);
nand U16168 (N_16168,N_14112,N_15231);
or U16169 (N_16169,N_14812,N_15044);
xnor U16170 (N_16170,N_14720,N_15209);
and U16171 (N_16171,N_15664,N_15471);
nand U16172 (N_16172,N_14769,N_14989);
nand U16173 (N_16173,N_15159,N_14991);
xnor U16174 (N_16174,N_15849,N_14375);
xnor U16175 (N_16175,N_15731,N_14380);
nand U16176 (N_16176,N_15695,N_15842);
xor U16177 (N_16177,N_15354,N_14181);
or U16178 (N_16178,N_14498,N_14445);
and U16179 (N_16179,N_14448,N_14264);
xor U16180 (N_16180,N_15820,N_15863);
nand U16181 (N_16181,N_15097,N_14719);
xnor U16182 (N_16182,N_15217,N_14128);
or U16183 (N_16183,N_14968,N_15565);
nand U16184 (N_16184,N_15658,N_14214);
xnor U16185 (N_16185,N_14980,N_15406);
xnor U16186 (N_16186,N_15631,N_15875);
or U16187 (N_16187,N_15841,N_14646);
nand U16188 (N_16188,N_15358,N_15360);
nand U16189 (N_16189,N_14654,N_14152);
or U16190 (N_16190,N_15557,N_14561);
nand U16191 (N_16191,N_15644,N_15076);
and U16192 (N_16192,N_14176,N_14735);
and U16193 (N_16193,N_15511,N_14616);
xor U16194 (N_16194,N_15155,N_14398);
or U16195 (N_16195,N_15492,N_14787);
and U16196 (N_16196,N_15179,N_15742);
and U16197 (N_16197,N_14056,N_15539);
nand U16198 (N_16198,N_14285,N_15031);
nor U16199 (N_16199,N_14494,N_15321);
and U16200 (N_16200,N_14325,N_15140);
nor U16201 (N_16201,N_14340,N_15141);
nand U16202 (N_16202,N_15094,N_15750);
xor U16203 (N_16203,N_15461,N_14370);
nand U16204 (N_16204,N_14939,N_15784);
xor U16205 (N_16205,N_14841,N_15005);
and U16206 (N_16206,N_14805,N_14146);
xnor U16207 (N_16207,N_15950,N_14940);
nand U16208 (N_16208,N_14199,N_14477);
and U16209 (N_16209,N_14987,N_15778);
nor U16210 (N_16210,N_15832,N_14573);
nor U16211 (N_16211,N_14707,N_15377);
or U16212 (N_16212,N_14373,N_15425);
and U16213 (N_16213,N_14723,N_15603);
nand U16214 (N_16214,N_14362,N_15764);
nor U16215 (N_16215,N_14776,N_15917);
and U16216 (N_16216,N_14618,N_14167);
and U16217 (N_16217,N_14539,N_15683);
nand U16218 (N_16218,N_14071,N_14729);
xnor U16219 (N_16219,N_14627,N_14419);
and U16220 (N_16220,N_14591,N_15754);
or U16221 (N_16221,N_15716,N_15556);
nor U16222 (N_16222,N_14950,N_14920);
and U16223 (N_16223,N_14877,N_15560);
nor U16224 (N_16224,N_14552,N_14064);
nand U16225 (N_16225,N_15919,N_14377);
nor U16226 (N_16226,N_14599,N_14842);
xor U16227 (N_16227,N_15212,N_14741);
xor U16228 (N_16228,N_14479,N_15009);
nor U16229 (N_16229,N_14102,N_14737);
or U16230 (N_16230,N_15874,N_14417);
xnor U16231 (N_16231,N_15933,N_14990);
xor U16232 (N_16232,N_15057,N_15876);
nand U16233 (N_16233,N_14367,N_14261);
or U16234 (N_16234,N_15630,N_14022);
and U16235 (N_16235,N_14286,N_15339);
xnor U16236 (N_16236,N_15314,N_14298);
nor U16237 (N_16237,N_14423,N_14683);
xor U16238 (N_16238,N_14021,N_14921);
and U16239 (N_16239,N_15330,N_14744);
or U16240 (N_16240,N_15077,N_14495);
nor U16241 (N_16241,N_15999,N_14857);
nor U16242 (N_16242,N_15908,N_14535);
xor U16243 (N_16243,N_15962,N_15043);
and U16244 (N_16244,N_14297,N_15813);
or U16245 (N_16245,N_14088,N_15629);
nand U16246 (N_16246,N_14288,N_14446);
nand U16247 (N_16247,N_14813,N_14858);
xor U16248 (N_16248,N_14834,N_15829);
xnor U16249 (N_16249,N_14634,N_14307);
or U16250 (N_16250,N_15101,N_15655);
or U16251 (N_16251,N_15168,N_15756);
nand U16252 (N_16252,N_15571,N_14526);
xor U16253 (N_16253,N_14392,N_15517);
and U16254 (N_16254,N_14708,N_15376);
or U16255 (N_16255,N_14044,N_14696);
nand U16256 (N_16256,N_15902,N_15865);
and U16257 (N_16257,N_14415,N_14251);
or U16258 (N_16258,N_15098,N_14846);
nor U16259 (N_16259,N_15459,N_14918);
nor U16260 (N_16260,N_15259,N_14180);
xor U16261 (N_16261,N_14436,N_14275);
nor U16262 (N_16262,N_14086,N_15899);
xnor U16263 (N_16263,N_15191,N_14657);
and U16264 (N_16264,N_15622,N_14396);
nor U16265 (N_16265,N_14142,N_15955);
nand U16266 (N_16266,N_15234,N_14442);
xor U16267 (N_16267,N_14234,N_15648);
and U16268 (N_16268,N_14575,N_15078);
nand U16269 (N_16269,N_14277,N_14560);
and U16270 (N_16270,N_15872,N_14397);
or U16271 (N_16271,N_14010,N_14366);
xor U16272 (N_16272,N_14029,N_14045);
and U16273 (N_16273,N_14664,N_14619);
nand U16274 (N_16274,N_15208,N_14289);
nand U16275 (N_16275,N_14421,N_14012);
xnor U16276 (N_16276,N_14760,N_14579);
xnor U16277 (N_16277,N_15589,N_14492);
and U16278 (N_16278,N_14658,N_14621);
nand U16279 (N_16279,N_15861,N_15516);
or U16280 (N_16280,N_14384,N_15361);
or U16281 (N_16281,N_15352,N_14714);
xnor U16282 (N_16282,N_15547,N_15705);
xor U16283 (N_16283,N_15499,N_15988);
xor U16284 (N_16284,N_15696,N_14305);
xnor U16285 (N_16285,N_14015,N_14628);
and U16286 (N_16286,N_14578,N_15653);
nand U16287 (N_16287,N_15106,N_15312);
nand U16288 (N_16288,N_14401,N_14080);
nand U16289 (N_16289,N_15454,N_15264);
or U16290 (N_16290,N_14389,N_15935);
or U16291 (N_16291,N_15638,N_14085);
nand U16292 (N_16292,N_15184,N_14493);
nand U16293 (N_16293,N_14184,N_14355);
or U16294 (N_16294,N_15286,N_14393);
nand U16295 (N_16295,N_15430,N_14705);
or U16296 (N_16296,N_15333,N_14489);
xor U16297 (N_16297,N_14574,N_15230);
xnor U16298 (N_16298,N_14078,N_14301);
nand U16299 (N_16299,N_14057,N_15439);
nand U16300 (N_16300,N_14237,N_15302);
nand U16301 (N_16301,N_14155,N_15319);
nand U16302 (N_16302,N_14660,N_15441);
nor U16303 (N_16303,N_15666,N_14866);
and U16304 (N_16304,N_15091,N_15866);
xnor U16305 (N_16305,N_15541,N_15652);
nor U16306 (N_16306,N_15010,N_14164);
nand U16307 (N_16307,N_14638,N_15344);
or U16308 (N_16308,N_14931,N_14810);
and U16309 (N_16309,N_15596,N_15785);
and U16310 (N_16310,N_14679,N_14718);
and U16311 (N_16311,N_15062,N_14648);
nor U16312 (N_16312,N_15971,N_14160);
and U16313 (N_16313,N_14863,N_14511);
and U16314 (N_16314,N_14783,N_15553);
or U16315 (N_16315,N_15129,N_15378);
or U16316 (N_16316,N_14799,N_15484);
or U16317 (N_16317,N_14369,N_14502);
nor U16318 (N_16318,N_14792,N_14957);
and U16319 (N_16319,N_14964,N_14522);
nor U16320 (N_16320,N_15979,N_14282);
nand U16321 (N_16321,N_15697,N_14548);
xor U16322 (N_16322,N_15688,N_14279);
nand U16323 (N_16323,N_14471,N_14811);
xor U16324 (N_16324,N_15469,N_14684);
and U16325 (N_16325,N_14196,N_15054);
or U16326 (N_16326,N_14778,N_14017);
and U16327 (N_16327,N_15564,N_14009);
or U16328 (N_16328,N_15858,N_15996);
nand U16329 (N_16329,N_14608,N_14466);
or U16330 (N_16330,N_14676,N_14135);
xor U16331 (N_16331,N_15535,N_15385);
xnor U16332 (N_16332,N_14441,N_14273);
or U16333 (N_16333,N_14819,N_14204);
or U16334 (N_16334,N_15167,N_14333);
or U16335 (N_16335,N_15411,N_15994);
nand U16336 (N_16336,N_14035,N_14536);
or U16337 (N_16337,N_15513,N_14236);
nor U16338 (N_16338,N_14216,N_15252);
nor U16339 (N_16339,N_15288,N_15827);
and U16340 (N_16340,N_15867,N_15109);
xnor U16341 (N_16341,N_14814,N_14637);
nand U16342 (N_16342,N_15022,N_14689);
and U16343 (N_16343,N_14092,N_14406);
nand U16344 (N_16344,N_15771,N_15337);
or U16345 (N_16345,N_14726,N_15397);
and U16346 (N_16346,N_14583,N_15145);
xnor U16347 (N_16347,N_14318,N_15903);
nand U16348 (N_16348,N_14118,N_14890);
or U16349 (N_16349,N_15393,N_14106);
nor U16350 (N_16350,N_14727,N_14030);
xor U16351 (N_16351,N_14801,N_14506);
nor U16352 (N_16352,N_14817,N_15654);
nor U16353 (N_16353,N_14472,N_14996);
nor U16354 (N_16354,N_14944,N_15375);
and U16355 (N_16355,N_15498,N_14596);
nor U16356 (N_16356,N_14651,N_15779);
and U16357 (N_16357,N_15362,N_14224);
or U16358 (N_16358,N_14465,N_14076);
nand U16359 (N_16359,N_14985,N_15836);
nor U16360 (N_16360,N_15703,N_14321);
xor U16361 (N_16361,N_14225,N_14556);
xnor U16362 (N_16362,N_15174,N_15087);
xor U16363 (N_16363,N_14518,N_14133);
nand U16364 (N_16364,N_14109,N_15297);
xor U16365 (N_16365,N_15404,N_14661);
nand U16366 (N_16366,N_14319,N_14019);
xnor U16367 (N_16367,N_15173,N_14461);
xor U16368 (N_16368,N_15772,N_14037);
and U16369 (N_16369,N_15635,N_15977);
xnor U16370 (N_16370,N_15668,N_14692);
and U16371 (N_16371,N_14310,N_15687);
nor U16372 (N_16372,N_14103,N_14900);
nand U16373 (N_16373,N_14433,N_15823);
xnor U16374 (N_16374,N_14945,N_15235);
nor U16375 (N_16375,N_14149,N_14460);
or U16376 (N_16376,N_15068,N_14005);
nand U16377 (N_16377,N_15972,N_14452);
and U16378 (N_16378,N_15110,N_14893);
and U16379 (N_16379,N_15341,N_14653);
xnor U16380 (N_16380,N_15608,N_14150);
nand U16381 (N_16381,N_15382,N_14532);
nand U16382 (N_16382,N_15317,N_14270);
or U16383 (N_16383,N_15373,N_15572);
and U16384 (N_16384,N_14328,N_15525);
nand U16385 (N_16385,N_14054,N_15142);
xor U16386 (N_16386,N_15612,N_14632);
nand U16387 (N_16387,N_14577,N_14700);
or U16388 (N_16388,N_14941,N_15391);
nor U16389 (N_16389,N_14848,N_15081);
or U16390 (N_16390,N_15915,N_14986);
or U16391 (N_16391,N_15082,N_15355);
nand U16392 (N_16392,N_15639,N_15976);
nor U16393 (N_16393,N_14185,N_15214);
nand U16394 (N_16394,N_15103,N_15003);
xor U16395 (N_16395,N_15895,N_15398);
xnor U16396 (N_16396,N_15348,N_14607);
nor U16397 (N_16397,N_15967,N_14739);
nand U16398 (N_16398,N_15961,N_15121);
nor U16399 (N_16399,N_14306,N_15790);
and U16400 (N_16400,N_15228,N_14201);
nor U16401 (N_16401,N_14528,N_14356);
nor U16402 (N_16402,N_15047,N_14903);
or U16403 (N_16403,N_14901,N_14709);
or U16404 (N_16404,N_14229,N_14963);
nor U16405 (N_16405,N_15301,N_14099);
or U16406 (N_16406,N_14250,N_14984);
xnor U16407 (N_16407,N_15197,N_15239);
and U16408 (N_16408,N_15942,N_15673);
xor U16409 (N_16409,N_15611,N_14069);
xor U16410 (N_16410,N_15545,N_14721);
nor U16411 (N_16411,N_14100,N_14138);
or U16412 (N_16412,N_15267,N_14780);
and U16413 (N_16413,N_15216,N_15283);
nor U16414 (N_16414,N_15048,N_14323);
or U16415 (N_16415,N_15672,N_14077);
nor U16416 (N_16416,N_15389,N_14190);
nor U16417 (N_16417,N_14854,N_14835);
nand U16418 (N_16418,N_15907,N_15852);
xor U16419 (N_16419,N_14205,N_15130);
and U16420 (N_16420,N_14797,N_14898);
nand U16421 (N_16421,N_15542,N_14915);
or U16422 (N_16422,N_14309,N_15923);
nor U16423 (N_16423,N_14695,N_14239);
xor U16424 (N_16424,N_15456,N_15429);
nor U16425 (N_16425,N_14170,N_14211);
xor U16426 (N_16426,N_14932,N_15299);
nand U16427 (N_16427,N_14694,N_15250);
or U16428 (N_16428,N_15038,N_14897);
or U16429 (N_16429,N_15263,N_14425);
nand U16430 (N_16430,N_15475,N_15725);
nand U16431 (N_16431,N_15412,N_15464);
xnor U16432 (N_16432,N_15615,N_14557);
nand U16433 (N_16433,N_14975,N_15605);
xor U16434 (N_16434,N_15944,N_15567);
or U16435 (N_16435,N_14065,N_15722);
nor U16436 (N_16436,N_14175,N_14473);
and U16437 (N_16437,N_14733,N_15679);
nor U16438 (N_16438,N_14759,N_14962);
xor U16439 (N_16439,N_15147,N_15436);
xor U16440 (N_16440,N_14105,N_14488);
and U16441 (N_16441,N_14979,N_15597);
xor U16442 (N_16442,N_14645,N_14060);
xnor U16443 (N_16443,N_14860,N_14597);
nand U16444 (N_16444,N_15914,N_14717);
nand U16445 (N_16445,N_15645,N_15266);
and U16446 (N_16446,N_14025,N_14883);
or U16447 (N_16447,N_14171,N_14050);
or U16448 (N_16448,N_15675,N_15659);
xor U16449 (N_16449,N_15403,N_14402);
or U16450 (N_16450,N_14073,N_14383);
and U16451 (N_16451,N_14391,N_15647);
nand U16452 (N_16452,N_15808,N_15773);
and U16453 (N_16453,N_14702,N_15898);
nor U16454 (N_16454,N_15628,N_14197);
nor U16455 (N_16455,N_15201,N_14259);
xor U16456 (N_16456,N_14263,N_15793);
nand U16457 (N_16457,N_14547,N_15794);
and U16458 (N_16458,N_14331,N_14499);
or U16459 (N_16459,N_15276,N_15621);
nor U16460 (N_16460,N_15025,N_15195);
nor U16461 (N_16461,N_14958,N_14008);
nand U16462 (N_16462,N_15026,N_15363);
xor U16463 (N_16463,N_15522,N_15428);
nand U16464 (N_16464,N_15749,N_14988);
nor U16465 (N_16465,N_14662,N_14302);
and U16466 (N_16466,N_14469,N_15969);
nor U16467 (N_16467,N_14666,N_15012);
or U16468 (N_16468,N_15995,N_14514);
xor U16469 (N_16469,N_14407,N_15965);
and U16470 (N_16470,N_15726,N_15712);
nor U16471 (N_16471,N_14040,N_15782);
xnor U16472 (N_16472,N_14951,N_15856);
and U16473 (N_16473,N_14137,N_14033);
xnor U16474 (N_16474,N_15952,N_15633);
nand U16475 (N_16475,N_15706,N_15934);
xnor U16476 (N_16476,N_15951,N_14746);
nor U16477 (N_16477,N_15592,N_14788);
xnor U16478 (N_16478,N_15757,N_15246);
and U16479 (N_16479,N_15088,N_14750);
xor U16480 (N_16480,N_15126,N_14559);
nor U16481 (N_16481,N_14589,N_15293);
and U16482 (N_16482,N_14284,N_15839);
or U16483 (N_16483,N_15627,N_14856);
nor U16484 (N_16484,N_15538,N_14954);
nand U16485 (N_16485,N_15885,N_14061);
nor U16486 (N_16486,N_15304,N_15311);
nor U16487 (N_16487,N_14935,N_15905);
nor U16488 (N_16488,N_14313,N_14889);
and U16489 (N_16489,N_14192,N_14254);
nor U16490 (N_16490,N_14113,N_15708);
or U16491 (N_16491,N_14620,N_14122);
nand U16492 (N_16492,N_15767,N_15759);
and U16493 (N_16493,N_14642,N_15143);
nand U16494 (N_16494,N_15562,N_14710);
nor U16495 (N_16495,N_15984,N_14067);
nor U16496 (N_16496,N_15906,N_15457);
nand U16497 (N_16497,N_15591,N_15946);
or U16498 (N_16498,N_14491,N_14582);
nand U16499 (N_16499,N_15626,N_15990);
and U16500 (N_16500,N_14378,N_15711);
nor U16501 (N_16501,N_14347,N_14879);
xnor U16502 (N_16502,N_15149,N_14059);
nor U16503 (N_16503,N_15928,N_15519);
nor U16504 (N_16504,N_15744,N_14255);
xor U16505 (N_16505,N_15501,N_15848);
nor U16506 (N_16506,N_14292,N_15818);
nor U16507 (N_16507,N_14359,N_15401);
xnor U16508 (N_16508,N_14154,N_14217);
and U16509 (N_16509,N_14243,N_15663);
nand U16510 (N_16510,N_15985,N_15340);
nor U16511 (N_16511,N_15482,N_14630);
nor U16512 (N_16512,N_15882,N_14959);
xnor U16513 (N_16513,N_14198,N_15493);
and U16514 (N_16514,N_15193,N_15300);
nand U16515 (N_16515,N_15183,N_14640);
nand U16516 (N_16516,N_14394,N_15940);
and U16517 (N_16517,N_15154,N_15616);
xnor U16518 (N_16518,N_15458,N_15497);
and U16519 (N_16519,N_14024,N_14833);
or U16520 (N_16520,N_14438,N_15728);
nor U16521 (N_16521,N_14558,N_14411);
or U16522 (N_16522,N_14669,N_14527);
nand U16523 (N_16523,N_15791,N_15527);
xnor U16524 (N_16524,N_14468,N_15641);
xor U16525 (N_16525,N_14743,N_15368);
nand U16526 (N_16526,N_15383,N_15825);
or U16527 (N_16527,N_15799,N_15978);
xor U16528 (N_16528,N_14249,N_15137);
xnor U16529 (N_16529,N_15074,N_14907);
nor U16530 (N_16530,N_15280,N_15864);
nand U16531 (N_16531,N_14790,N_15421);
or U16532 (N_16532,N_14742,N_15816);
xnor U16533 (N_16533,N_15163,N_15886);
nand U16534 (N_16534,N_15774,N_14416);
or U16535 (N_16535,N_14376,N_14796);
or U16536 (N_16536,N_14567,N_15507);
xnor U16537 (N_16537,N_14462,N_14730);
nor U16538 (N_16538,N_14451,N_15253);
nor U16539 (N_16539,N_14995,N_14906);
xor U16540 (N_16540,N_14523,N_14722);
nor U16541 (N_16541,N_15303,N_15029);
nor U16542 (N_16542,N_15532,N_14207);
nand U16543 (N_16543,N_14091,N_14872);
nand U16544 (N_16544,N_14014,N_15255);
xnor U16545 (N_16545,N_15563,N_14905);
and U16546 (N_16546,N_15218,N_15438);
or U16547 (N_16547,N_15086,N_14613);
nor U16548 (N_16548,N_15957,N_15247);
xnor U16549 (N_16549,N_15981,N_15170);
nor U16550 (N_16550,N_15305,N_15099);
xor U16551 (N_16551,N_15686,N_15442);
xnor U16552 (N_16552,N_14101,N_15598);
nand U16553 (N_16553,N_15090,N_14178);
nor U16554 (N_16554,N_15256,N_15758);
nor U16555 (N_16555,N_14531,N_14287);
and U16556 (N_16556,N_15402,N_14413);
nand U16557 (N_16557,N_15104,N_15795);
nand U16558 (N_16558,N_14299,N_14280);
nor U16559 (N_16559,N_15041,N_15569);
xor U16560 (N_16560,N_14314,N_15162);
and U16561 (N_16561,N_15755,N_15287);
or U16562 (N_16562,N_14117,N_14052);
xor U16563 (N_16563,N_14303,N_14157);
or U16564 (N_16564,N_14342,N_14784);
nand U16565 (N_16565,N_15426,N_15927);
xor U16566 (N_16566,N_15815,N_15113);
or U16567 (N_16567,N_15446,N_14757);
nor U16568 (N_16568,N_14221,N_14697);
nor U16569 (N_16569,N_14617,N_15871);
or U16570 (N_16570,N_15693,N_15814);
and U16571 (N_16571,N_15964,N_14603);
and U16572 (N_16572,N_15107,N_14588);
nand U16573 (N_16573,N_15419,N_14554);
and U16574 (N_16574,N_14690,N_15001);
nand U16575 (N_16575,N_15577,N_14625);
and U16576 (N_16576,N_15570,N_14346);
or U16577 (N_16577,N_14978,N_15432);
xnor U16578 (N_16578,N_14326,N_15900);
nor U16579 (N_16579,N_15336,N_14165);
nand U16580 (N_16580,N_14293,N_15024);
nand U16581 (N_16581,N_14159,N_15987);
and U16582 (N_16582,N_15479,N_14731);
or U16583 (N_16583,N_15039,N_15042);
nand U16584 (N_16584,N_14832,N_15467);
and U16585 (N_16585,N_15323,N_14115);
or U16586 (N_16586,N_15543,N_15781);
xnor U16587 (N_16587,N_14952,N_15242);
xor U16588 (N_16588,N_14141,N_15139);
nor U16589 (N_16589,N_15991,N_15656);
nor U16590 (N_16590,N_15824,N_15440);
nor U16591 (N_16591,N_14212,N_15445);
nor U16592 (N_16592,N_14521,N_14930);
nor U16593 (N_16593,N_14712,N_14836);
xnor U16594 (N_16594,N_15701,N_15500);
nor U16595 (N_16595,N_15548,N_14758);
or U16596 (N_16596,N_14691,N_14437);
nor U16597 (N_16597,N_15860,N_15496);
or U16598 (N_16598,N_15822,N_14233);
nor U16599 (N_16599,N_15600,N_14023);
and U16600 (N_16600,N_15692,N_15365);
xor U16601 (N_16601,N_15260,N_14885);
and U16602 (N_16602,N_14363,N_15877);
nand U16603 (N_16603,N_14051,N_15444);
xnor U16604 (N_16604,N_14294,N_15285);
or U16605 (N_16605,N_15601,N_14253);
nor U16606 (N_16606,N_14779,N_15476);
and U16607 (N_16607,N_14075,N_15963);
nand U16608 (N_16608,N_15085,N_14982);
xnor U16609 (N_16609,N_14258,N_15409);
xnor U16610 (N_16610,N_14206,N_14246);
nor U16611 (N_16611,N_15221,N_15396);
or U16612 (N_16612,N_15138,N_14381);
nor U16613 (N_16613,N_15169,N_14770);
xor U16614 (N_16614,N_14283,N_15366);
or U16615 (N_16615,N_15806,N_14929);
nor U16616 (N_16616,N_14967,N_14566);
and U16617 (N_16617,N_15219,N_14317);
or U16618 (N_16618,N_15490,N_15853);
or U16619 (N_16619,N_14247,N_15451);
nand U16620 (N_16620,N_14533,N_14668);
and U16621 (N_16621,N_14084,N_14803);
xnor U16622 (N_16622,N_14777,N_14732);
nand U16623 (N_16623,N_15017,N_15745);
xor U16624 (N_16624,N_15405,N_15040);
nand U16625 (N_16625,N_15738,N_14687);
nand U16626 (N_16626,N_15844,N_15894);
nand U16627 (N_16627,N_15033,N_15222);
xnor U16628 (N_16628,N_14818,N_14063);
xnor U16629 (N_16629,N_14177,N_15677);
or U16630 (N_16630,N_14808,N_15721);
nand U16631 (N_16631,N_15837,N_15470);
nor U16632 (N_16632,N_15920,N_15117);
nor U16633 (N_16633,N_14386,N_15092);
xnor U16634 (N_16634,N_15854,N_15157);
nor U16635 (N_16635,N_14379,N_14925);
xor U16636 (N_16636,N_14601,N_15619);
nor U16637 (N_16637,N_14938,N_15651);
or U16638 (N_16638,N_14703,N_15939);
and U16639 (N_16639,N_15699,N_14781);
nor U16640 (N_16640,N_14344,N_14865);
xor U16641 (N_16641,N_15119,N_15261);
or U16642 (N_16642,N_15420,N_14997);
and U16643 (N_16643,N_14368,N_14123);
nor U16644 (N_16644,N_14332,N_15188);
and U16645 (N_16645,N_15646,N_14114);
nand U16646 (N_16646,N_15148,N_15733);
or U16647 (N_16647,N_14336,N_15741);
nand U16648 (N_16648,N_14134,N_15248);
xnor U16649 (N_16649,N_15727,N_15118);
nand U16650 (N_16650,N_15153,N_15271);
and U16651 (N_16651,N_14335,N_14354);
nor U16652 (N_16652,N_15384,N_15909);
nand U16653 (N_16653,N_14412,N_14775);
and U16654 (N_16654,N_15593,N_15739);
and U16655 (N_16655,N_15945,N_15948);
or U16656 (N_16656,N_14698,N_15700);
xor U16657 (N_16657,N_14663,N_14768);
nand U16658 (N_16658,N_15819,N_14312);
and U16659 (N_16659,N_14867,N_14434);
and U16660 (N_16660,N_15887,N_14161);
nand U16661 (N_16661,N_14058,N_15747);
xnor U16662 (N_16662,N_14248,N_15584);
and U16663 (N_16663,N_14372,N_14568);
and U16664 (N_16664,N_15307,N_15114);
and U16665 (N_16665,N_14007,N_14062);
nor U16666 (N_16666,N_14458,N_14673);
nand U16667 (N_16667,N_14474,N_14837);
or U16668 (N_16668,N_15502,N_14827);
nand U16669 (N_16669,N_15473,N_14517);
nor U16670 (N_16670,N_14267,N_15463);
or U16671 (N_16671,N_14125,N_14976);
xnor U16672 (N_16672,N_14512,N_14816);
xor U16673 (N_16673,N_15595,N_14821);
nor U16674 (N_16674,N_14795,N_14410);
xor U16675 (N_16675,N_15369,N_14852);
and U16676 (N_16676,N_15046,N_14576);
or U16677 (N_16677,N_15599,N_14647);
xor U16678 (N_16678,N_15851,N_15124);
and U16679 (N_16679,N_14913,N_15555);
nand U16680 (N_16680,N_14316,N_14878);
nor U16681 (N_16681,N_14262,N_14859);
nor U16682 (N_16682,N_15833,N_15158);
nor U16683 (N_16683,N_14933,N_14525);
or U16684 (N_16684,N_15417,N_14928);
nand U16685 (N_16685,N_14728,N_15359);
nand U16686 (N_16686,N_15685,N_14553);
xnor U16687 (N_16687,N_15850,N_14936);
nor U16688 (N_16688,N_15845,N_14449);
and U16689 (N_16689,N_14266,N_15912);
xnor U16690 (N_16690,N_15164,N_14418);
xor U16691 (N_16691,N_15857,N_14042);
and U16692 (N_16692,N_14208,N_14830);
xnor U16693 (N_16693,N_15922,N_15171);
xor U16694 (N_16694,N_14424,N_14432);
nand U16695 (N_16695,N_15270,N_15021);
nor U16696 (N_16696,N_15986,N_15787);
or U16697 (N_16697,N_15580,N_14011);
and U16698 (N_16698,N_15802,N_15229);
nand U16699 (N_16699,N_15766,N_15279);
and U16700 (N_16700,N_15678,N_15576);
nand U16701 (N_16701,N_14622,N_15643);
or U16702 (N_16702,N_14428,N_14688);
nand U16703 (N_16703,N_14341,N_15869);
nand U16704 (N_16704,N_15714,N_14970);
and U16705 (N_16705,N_14960,N_14414);
and U16706 (N_16706,N_15798,N_15053);
nor U16707 (N_16707,N_15520,N_14467);
nor U16708 (N_16708,N_14156,N_14670);
nand U16709 (N_16709,N_15204,N_14047);
nand U16710 (N_16710,N_14043,N_14829);
xnor U16711 (N_16711,N_14218,N_14131);
and U16712 (N_16712,N_14390,N_14256);
and U16713 (N_16713,N_15408,N_14240);
nor U16714 (N_16714,N_15072,N_15132);
or U16715 (N_16715,N_15834,N_15954);
xnor U16716 (N_16716,N_15752,N_14070);
xor U16717 (N_16717,N_15510,N_15810);
and U16718 (N_16718,N_14501,N_14230);
nor U16719 (N_16719,N_15400,N_14503);
nand U16720 (N_16720,N_15064,N_14235);
nor U16721 (N_16721,N_14565,N_15594);
or U16722 (N_16722,N_15093,N_15275);
nor U16723 (N_16723,N_14636,N_15257);
xor U16724 (N_16724,N_15524,N_14334);
xnor U16725 (N_16725,N_15466,N_15870);
or U16726 (N_16726,N_15050,N_15587);
and U16727 (N_16727,N_15075,N_14330);
xor U16728 (N_16728,N_14200,N_14158);
and U16729 (N_16729,N_15172,N_15156);
nor U16730 (N_16730,N_15796,N_15182);
and U16731 (N_16731,N_14371,N_14111);
or U16732 (N_16732,N_15045,N_14602);
or U16733 (N_16733,N_14026,N_14626);
and U16734 (N_16734,N_14116,N_14911);
nand U16735 (N_16735,N_15573,N_14032);
or U16736 (N_16736,N_14480,N_14443);
or U16737 (N_16737,N_14269,N_14943);
nor U16738 (N_16738,N_15175,N_14643);
nor U16739 (N_16739,N_14600,N_15243);
or U16740 (N_16740,N_15232,N_15019);
nor U16741 (N_16741,N_14352,N_15449);
nand U16742 (N_16742,N_15331,N_15786);
or U16743 (N_16743,N_15989,N_15568);
and U16744 (N_16744,N_15828,N_15925);
nor U16745 (N_16745,N_14193,N_15069);
nand U16746 (N_16746,N_14226,N_15505);
or U16747 (N_16747,N_15122,N_15968);
xor U16748 (N_16748,N_14151,N_14231);
nand U16749 (N_16749,N_15238,N_14210);
nand U16750 (N_16750,N_14509,N_15450);
or U16751 (N_16751,N_14585,N_15100);
nor U16752 (N_16752,N_15327,N_15478);
xnor U16753 (N_16753,N_15588,N_15060);
nor U16754 (N_16754,N_14096,N_14182);
xnor U16755 (N_16755,N_14082,N_15868);
xor U16756 (N_16756,N_14153,N_15748);
or U16757 (N_16757,N_14771,N_15717);
nor U16758 (N_16758,N_15735,N_14464);
xor U16759 (N_16759,N_14650,N_15151);
and U16760 (N_16760,N_15723,N_15846);
or U16761 (N_16761,N_15891,N_15681);
nor U16762 (N_16762,N_14974,N_14755);
xnor U16763 (N_16763,N_14274,N_14049);
xor U16764 (N_16764,N_15079,N_14322);
and U16765 (N_16765,N_15620,N_14530);
nor U16766 (N_16766,N_15893,N_15637);
and U16767 (N_16767,N_15199,N_14873);
and U16768 (N_16768,N_15272,N_15073);
and U16769 (N_16769,N_14922,N_14550);
and U16770 (N_16770,N_15625,N_14753);
or U16771 (N_16771,N_14290,N_15332);
nand U16772 (N_16772,N_15761,N_14388);
nor U16773 (N_16773,N_15202,N_15719);
xor U16774 (N_16774,N_15415,N_15812);
or U16775 (N_16775,N_14870,N_15936);
nand U16776 (N_16776,N_15904,N_15371);
and U16777 (N_16777,N_15133,N_14549);
nand U16778 (N_16778,N_15838,N_14300);
nor U16779 (N_16779,N_15262,N_15146);
nor U16780 (N_16780,N_14053,N_15889);
and U16781 (N_16781,N_15494,N_14454);
xnor U16782 (N_16782,N_15485,N_14641);
and U16783 (N_16783,N_14631,N_14680);
or U16784 (N_16784,N_15351,N_15992);
nor U16785 (N_16785,N_15136,N_14612);
nor U16786 (N_16786,N_14343,N_15737);
or U16787 (N_16787,N_15241,N_14853);
nor U16788 (N_16788,N_15049,N_14271);
xor U16789 (N_16789,N_14614,N_14678);
nor U16790 (N_16790,N_15953,N_15379);
nor U16791 (N_16791,N_15526,N_15486);
and U16792 (N_16792,N_15634,N_15277);
nor U16793 (N_16793,N_14924,N_14855);
xor U16794 (N_16794,N_14754,N_14093);
and U16795 (N_16795,N_15770,N_15803);
or U16796 (N_16796,N_15809,N_15120);
or U16797 (N_16797,N_14659,N_14481);
and U16798 (N_16798,N_15938,N_14439);
or U16799 (N_16799,N_15233,N_14430);
xnor U16800 (N_16800,N_14738,N_15941);
and U16801 (N_16801,N_14232,N_15546);
xnor U16802 (N_16802,N_15811,N_15394);
nand U16803 (N_16803,N_15227,N_14562);
nor U16804 (N_16804,N_14891,N_14147);
and U16805 (N_16805,N_15533,N_15581);
nand U16806 (N_16806,N_15294,N_15196);
and U16807 (N_16807,N_15537,N_14519);
xor U16808 (N_16808,N_14020,N_15890);
nand U16809 (N_16809,N_15178,N_15552);
and U16810 (N_16810,N_14524,N_15185);
nand U16811 (N_16811,N_14961,N_14003);
nor U16812 (N_16812,N_14089,N_15329);
nand U16813 (N_16813,N_14038,N_15518);
xor U16814 (N_16814,N_15775,N_15931);
or U16815 (N_16815,N_14590,N_15662);
and U16816 (N_16816,N_14041,N_15896);
or U16817 (N_16817,N_15063,N_15102);
nand U16818 (N_16818,N_15387,N_14593);
nand U16819 (N_16819,N_15220,N_14948);
nand U16820 (N_16820,N_14006,N_14508);
nand U16821 (N_16821,N_15059,N_15544);
nand U16822 (N_16822,N_15281,N_15455);
xnor U16823 (N_16823,N_14840,N_15926);
xor U16824 (N_16824,N_14357,N_15718);
nor U16825 (N_16825,N_15244,N_14850);
or U16826 (N_16826,N_15531,N_15187);
xor U16827 (N_16827,N_15474,N_14126);
nand U16828 (N_16828,N_15674,N_14971);
nor U16829 (N_16829,N_14711,N_14018);
and U16830 (N_16830,N_14748,N_15413);
nand U16831 (N_16831,N_14629,N_14822);
nor U16832 (N_16832,N_14252,N_14800);
or U16833 (N_16833,N_15388,N_15540);
or U16834 (N_16834,N_14942,N_14899);
nand U16835 (N_16835,N_14000,N_14163);
xnor U16836 (N_16836,N_15447,N_14543);
nand U16837 (N_16837,N_15558,N_14605);
or U16838 (N_16838,N_14496,N_15740);
nor U16839 (N_16839,N_14655,N_14762);
nor U16840 (N_16840,N_15610,N_14594);
nand U16841 (N_16841,N_14973,N_15713);
xnor U16842 (N_16842,N_14570,N_14202);
xnor U16843 (N_16843,N_15036,N_14752);
and U16844 (N_16844,N_15636,N_14786);
xor U16845 (N_16845,N_15210,N_15313);
nand U16846 (N_16846,N_14927,N_14013);
and U16847 (N_16847,N_15414,N_14862);
nand U16848 (N_16848,N_15318,N_14327);
nor U16849 (N_16849,N_15974,N_14992);
and U16850 (N_16850,N_14794,N_14074);
nand U16851 (N_16851,N_15237,N_15028);
nor U16852 (N_16852,N_15487,N_15004);
and U16853 (N_16853,N_14409,N_15160);
xor U16854 (N_16854,N_14265,N_14241);
or U16855 (N_16855,N_15165,N_15980);
nor U16856 (N_16856,N_14072,N_14295);
xor U16857 (N_16857,N_15910,N_14806);
xor U16858 (N_16858,N_14483,N_15152);
xnor U16859 (N_16859,N_14674,N_14623);
nor U16860 (N_16860,N_14510,N_15427);
xnor U16861 (N_16861,N_15665,N_15929);
xor U16862 (N_16862,N_15211,N_14144);
nand U16863 (N_16863,N_14203,N_15769);
xor U16864 (N_16864,N_14027,N_15390);
nor U16865 (N_16865,N_15095,N_15123);
and U16866 (N_16866,N_14847,N_15523);
nand U16867 (N_16867,N_15357,N_15489);
or U16868 (N_16868,N_15416,N_14486);
or U16869 (N_16869,N_14046,N_15224);
and U16870 (N_16870,N_14337,N_15181);
and U16871 (N_16871,N_14440,N_14540);
nor U16872 (N_16872,N_14487,N_15657);
or U16873 (N_16873,N_15873,N_14894);
nor U16874 (N_16874,N_14004,N_14186);
nor U16875 (N_16875,N_15125,N_14450);
xor U16876 (N_16876,N_15554,N_14747);
and U16877 (N_16877,N_14604,N_14364);
and U16878 (N_16878,N_14194,N_15959);
or U16879 (N_16879,N_15035,N_15128);
or U16880 (N_16880,N_14132,N_15997);
nand U16881 (N_16881,N_14953,N_14772);
nand U16882 (N_16882,N_15521,N_15324);
xor U16883 (N_16883,N_14715,N_15027);
or U16884 (N_16884,N_14851,N_15720);
nand U16885 (N_16885,N_15343,N_14908);
and U16886 (N_16886,N_14693,N_14162);
or U16887 (N_16887,N_15751,N_14977);
xor U16888 (N_16888,N_15901,N_15734);
or U16889 (N_16889,N_15536,N_14034);
or U16890 (N_16890,N_15506,N_14520);
xor U16891 (N_16891,N_15011,N_14969);
and U16892 (N_16892,N_15200,N_15878);
xnor U16893 (N_16893,N_14724,N_15777);
and U16894 (N_16894,N_15707,N_15694);
nor U16895 (N_16895,N_14435,N_15590);
nor U16896 (N_16896,N_15724,N_14966);
nand U16897 (N_16897,N_14624,N_15370);
nor U16898 (N_16898,N_14055,N_15131);
or U16899 (N_16899,N_14104,N_14782);
or U16900 (N_16900,N_15821,N_14169);
nand U16901 (N_16901,N_15089,N_14172);
nor U16902 (N_16902,N_14809,N_14083);
or U16903 (N_16903,N_14127,N_15399);
nand U16904 (N_16904,N_14955,N_14802);
or U16905 (N_16905,N_15930,N_15083);
nor U16906 (N_16906,N_14447,N_15514);
and U16907 (N_16907,N_14843,N_15002);
nand U16908 (N_16908,N_15481,N_15423);
and U16909 (N_16909,N_14615,N_15367);
xor U16910 (N_16910,N_14587,N_15640);
nand U16911 (N_16911,N_15186,N_15015);
nor U16912 (N_16912,N_15448,N_14839);
nand U16913 (N_16913,N_15205,N_15830);
nand U16914 (N_16914,N_15306,N_14542);
nand U16915 (N_16915,N_14497,N_15291);
nor U16916 (N_16916,N_15316,N_14361);
and U16917 (N_16917,N_15559,N_14189);
nor U16918 (N_16918,N_15606,N_14028);
or U16919 (N_16919,N_14227,N_15788);
xor U16920 (N_16920,N_14736,N_14507);
or U16921 (N_16921,N_14682,N_14845);
nor U16922 (N_16922,N_14315,N_14937);
or U16923 (N_16923,N_14884,N_14278);
and U16924 (N_16924,N_14882,N_15245);
and U16925 (N_16925,N_15966,N_15065);
and U16926 (N_16926,N_14228,N_14238);
xnor U16927 (N_16927,N_14431,N_15000);
xor U16928 (N_16928,N_15055,N_14429);
and U16929 (N_16929,N_15150,N_15618);
nor U16930 (N_16930,N_14671,N_15392);
xnor U16931 (N_16931,N_15254,N_15709);
nor U16932 (N_16932,N_15353,N_15549);
xnor U16933 (N_16933,N_15883,N_15434);
and U16934 (N_16934,N_15472,N_14219);
nand U16935 (N_16935,N_15958,N_15418);
nor U16936 (N_16936,N_14563,N_15676);
or U16937 (N_16937,N_15710,N_15765);
nor U16938 (N_16938,N_14998,N_15585);
or U16939 (N_16939,N_15372,N_15983);
nor U16940 (N_16940,N_14667,N_15768);
xor U16941 (N_16941,N_15530,N_15880);
nor U16942 (N_16942,N_15859,N_14639);
nand U16943 (N_16943,N_14888,N_15529);
or U16944 (N_16944,N_14124,N_15433);
xor U16945 (N_16945,N_15071,N_14965);
nor U16946 (N_16946,N_14016,N_15115);
nand U16947 (N_16947,N_14774,N_15207);
nor U16948 (N_16948,N_14408,N_14382);
nand U16949 (N_16949,N_15937,N_14320);
and U16950 (N_16950,N_14395,N_15817);
and U16951 (N_16951,N_15265,N_14098);
xor U16952 (N_16952,N_15325,N_14761);
xnor U16953 (N_16953,N_14081,N_15993);
xor U16954 (N_16954,N_15292,N_14482);
or U16955 (N_16955,N_15918,N_14183);
xnor U16956 (N_16956,N_14545,N_14686);
and U16957 (N_16957,N_15732,N_14244);
nand U16958 (N_16958,N_15223,N_14544);
and U16959 (N_16959,N_15508,N_14500);
nand U16960 (N_16960,N_15760,N_14108);
or U16961 (N_16961,N_15349,N_15213);
and U16962 (N_16962,N_15840,N_14825);
nor U16963 (N_16963,N_14504,N_15269);
nand U16964 (N_16964,N_15534,N_15932);
and U16965 (N_16965,N_15495,N_14399);
nand U16966 (N_16966,N_15108,N_14580);
or U16967 (N_16967,N_15278,N_14610);
xor U16968 (N_16968,N_14136,N_15468);
xor U16969 (N_16969,N_15613,N_15023);
and U16970 (N_16970,N_15921,N_15135);
xnor U16971 (N_16971,N_14329,N_15144);
or U16972 (N_16972,N_14874,N_14209);
nand U16973 (N_16973,N_14478,N_14766);
or U16974 (N_16974,N_14505,N_14475);
nor U16975 (N_16975,N_14365,N_14904);
nor U16976 (N_16976,N_15013,N_15016);
nor U16977 (N_16977,N_15008,N_15913);
or U16978 (N_16978,N_15897,N_14681);
nor U16979 (N_16979,N_14699,N_15480);
xor U16980 (N_16980,N_15006,N_15582);
nand U16981 (N_16981,N_14220,N_15579);
nor U16982 (N_16982,N_14764,N_15689);
nor U16983 (N_16983,N_15550,N_14490);
nor U16984 (N_16984,N_15437,N_15916);
xor U16985 (N_16985,N_15070,N_14148);
and U16986 (N_16986,N_15273,N_14453);
nor U16987 (N_16987,N_14457,N_14798);
and U16988 (N_16988,N_14143,N_14187);
or U16989 (N_16989,N_15801,N_15350);
nand U16990 (N_16990,N_15888,N_15642);
nand U16991 (N_16991,N_14896,N_15975);
or U16992 (N_16992,N_15282,N_14121);
nand U16993 (N_16993,N_15831,N_15949);
nand U16994 (N_16994,N_15973,N_14541);
and U16995 (N_16995,N_14876,N_14756);
or U16996 (N_16996,N_14914,N_14740);
nand U16997 (N_16997,N_14119,N_14572);
nand U16998 (N_16998,N_15607,N_14001);
xor U16999 (N_16999,N_14947,N_14345);
nand U17000 (N_17000,N_14117,N_15538);
nor U17001 (N_17001,N_15503,N_14962);
and U17002 (N_17002,N_14329,N_14050);
or U17003 (N_17003,N_15019,N_15192);
and U17004 (N_17004,N_15276,N_15720);
xnor U17005 (N_17005,N_14227,N_14179);
or U17006 (N_17006,N_15650,N_15729);
xnor U17007 (N_17007,N_15388,N_15916);
or U17008 (N_17008,N_14194,N_14031);
xnor U17009 (N_17009,N_15358,N_14223);
nor U17010 (N_17010,N_15837,N_15651);
or U17011 (N_17011,N_14680,N_14049);
nand U17012 (N_17012,N_14203,N_15092);
and U17013 (N_17013,N_15575,N_14744);
nand U17014 (N_17014,N_14117,N_15783);
nor U17015 (N_17015,N_15249,N_14886);
xor U17016 (N_17016,N_15310,N_15806);
nand U17017 (N_17017,N_14729,N_15949);
nor U17018 (N_17018,N_15430,N_15598);
or U17019 (N_17019,N_15094,N_15226);
nor U17020 (N_17020,N_15782,N_14709);
and U17021 (N_17021,N_15878,N_14327);
nor U17022 (N_17022,N_15230,N_15565);
nand U17023 (N_17023,N_14399,N_14760);
nand U17024 (N_17024,N_14270,N_15552);
nand U17025 (N_17025,N_14019,N_15687);
or U17026 (N_17026,N_14322,N_15024);
nor U17027 (N_17027,N_15956,N_15155);
and U17028 (N_17028,N_14942,N_15061);
or U17029 (N_17029,N_15736,N_15648);
and U17030 (N_17030,N_14997,N_14320);
nor U17031 (N_17031,N_14966,N_15043);
nand U17032 (N_17032,N_14708,N_14393);
nor U17033 (N_17033,N_15583,N_15787);
and U17034 (N_17034,N_15577,N_15221);
xor U17035 (N_17035,N_15729,N_15468);
xnor U17036 (N_17036,N_14463,N_14540);
and U17037 (N_17037,N_15307,N_15287);
and U17038 (N_17038,N_15416,N_14140);
xnor U17039 (N_17039,N_14046,N_14549);
or U17040 (N_17040,N_15131,N_15435);
or U17041 (N_17041,N_14526,N_14021);
nand U17042 (N_17042,N_14860,N_14286);
nand U17043 (N_17043,N_15056,N_14484);
xnor U17044 (N_17044,N_15475,N_15287);
nand U17045 (N_17045,N_15047,N_14831);
or U17046 (N_17046,N_15289,N_15518);
or U17047 (N_17047,N_15369,N_15187);
nand U17048 (N_17048,N_15405,N_15714);
xor U17049 (N_17049,N_14168,N_15885);
xnor U17050 (N_17050,N_15363,N_14623);
or U17051 (N_17051,N_14924,N_15560);
or U17052 (N_17052,N_15992,N_14172);
or U17053 (N_17053,N_15643,N_15347);
or U17054 (N_17054,N_15539,N_14427);
nor U17055 (N_17055,N_15689,N_15867);
nor U17056 (N_17056,N_15529,N_15686);
nor U17057 (N_17057,N_15371,N_15437);
xor U17058 (N_17058,N_14219,N_14975);
xnor U17059 (N_17059,N_14634,N_15535);
xnor U17060 (N_17060,N_15341,N_15161);
xor U17061 (N_17061,N_15196,N_15987);
nor U17062 (N_17062,N_15543,N_15998);
nand U17063 (N_17063,N_15584,N_14626);
nand U17064 (N_17064,N_14960,N_15477);
nor U17065 (N_17065,N_14780,N_14834);
nand U17066 (N_17066,N_14023,N_15976);
xor U17067 (N_17067,N_15372,N_14032);
xnor U17068 (N_17068,N_15128,N_14460);
and U17069 (N_17069,N_15509,N_14957);
and U17070 (N_17070,N_15475,N_14293);
or U17071 (N_17071,N_15868,N_15811);
nor U17072 (N_17072,N_15189,N_14578);
or U17073 (N_17073,N_14793,N_14418);
nand U17074 (N_17074,N_14610,N_14266);
nor U17075 (N_17075,N_15757,N_14264);
nand U17076 (N_17076,N_14435,N_15221);
nand U17077 (N_17077,N_15637,N_15397);
and U17078 (N_17078,N_15553,N_14217);
nand U17079 (N_17079,N_14163,N_15313);
xor U17080 (N_17080,N_15311,N_15454);
nand U17081 (N_17081,N_14463,N_14522);
and U17082 (N_17082,N_14439,N_15028);
or U17083 (N_17083,N_15094,N_14078);
xor U17084 (N_17084,N_15439,N_15455);
and U17085 (N_17085,N_15557,N_15453);
nor U17086 (N_17086,N_14528,N_14415);
or U17087 (N_17087,N_14414,N_14364);
and U17088 (N_17088,N_14516,N_14979);
nor U17089 (N_17089,N_14082,N_14416);
or U17090 (N_17090,N_14410,N_14177);
or U17091 (N_17091,N_14052,N_15982);
nor U17092 (N_17092,N_15050,N_14441);
or U17093 (N_17093,N_15658,N_14338);
or U17094 (N_17094,N_15003,N_14625);
xnor U17095 (N_17095,N_14349,N_14762);
and U17096 (N_17096,N_14668,N_14035);
or U17097 (N_17097,N_15262,N_15903);
and U17098 (N_17098,N_15035,N_15662);
nor U17099 (N_17099,N_14296,N_15958);
nand U17100 (N_17100,N_15254,N_14154);
and U17101 (N_17101,N_14297,N_15891);
or U17102 (N_17102,N_15801,N_14044);
xnor U17103 (N_17103,N_15085,N_14515);
nand U17104 (N_17104,N_15525,N_15654);
xnor U17105 (N_17105,N_14741,N_15376);
nor U17106 (N_17106,N_15461,N_14317);
nor U17107 (N_17107,N_15099,N_14854);
nor U17108 (N_17108,N_14023,N_15342);
xnor U17109 (N_17109,N_15704,N_14285);
or U17110 (N_17110,N_15913,N_14515);
nor U17111 (N_17111,N_15243,N_15907);
or U17112 (N_17112,N_14307,N_15603);
nor U17113 (N_17113,N_14092,N_14935);
xor U17114 (N_17114,N_15856,N_15025);
xnor U17115 (N_17115,N_15369,N_14715);
and U17116 (N_17116,N_14597,N_14341);
nor U17117 (N_17117,N_15221,N_14219);
and U17118 (N_17118,N_15584,N_15643);
and U17119 (N_17119,N_15556,N_14017);
nor U17120 (N_17120,N_14587,N_15697);
and U17121 (N_17121,N_15115,N_14143);
and U17122 (N_17122,N_15884,N_14557);
nand U17123 (N_17123,N_14705,N_14440);
or U17124 (N_17124,N_15457,N_15709);
and U17125 (N_17125,N_15351,N_14384);
or U17126 (N_17126,N_15717,N_15416);
or U17127 (N_17127,N_14762,N_15884);
xnor U17128 (N_17128,N_14940,N_15597);
or U17129 (N_17129,N_15001,N_14874);
xor U17130 (N_17130,N_15037,N_15744);
xor U17131 (N_17131,N_14351,N_14597);
or U17132 (N_17132,N_15330,N_14310);
and U17133 (N_17133,N_15779,N_14521);
xor U17134 (N_17134,N_14084,N_14071);
xnor U17135 (N_17135,N_15709,N_15729);
or U17136 (N_17136,N_14563,N_14984);
nand U17137 (N_17137,N_14597,N_15256);
and U17138 (N_17138,N_14711,N_15432);
nand U17139 (N_17139,N_14872,N_14699);
or U17140 (N_17140,N_14252,N_14335);
xor U17141 (N_17141,N_14138,N_15160);
nand U17142 (N_17142,N_14464,N_15675);
nor U17143 (N_17143,N_15780,N_14013);
nand U17144 (N_17144,N_14663,N_15959);
or U17145 (N_17145,N_15720,N_14594);
or U17146 (N_17146,N_15246,N_15324);
and U17147 (N_17147,N_14986,N_15021);
nand U17148 (N_17148,N_15356,N_14122);
or U17149 (N_17149,N_14428,N_15211);
or U17150 (N_17150,N_15962,N_14874);
nor U17151 (N_17151,N_15932,N_15637);
nor U17152 (N_17152,N_14011,N_14541);
nand U17153 (N_17153,N_14119,N_15838);
nor U17154 (N_17154,N_15139,N_14301);
xor U17155 (N_17155,N_15110,N_14091);
or U17156 (N_17156,N_14570,N_15644);
xnor U17157 (N_17157,N_14450,N_15996);
and U17158 (N_17158,N_14409,N_15919);
nor U17159 (N_17159,N_14427,N_15488);
nor U17160 (N_17160,N_14438,N_14497);
and U17161 (N_17161,N_15328,N_14315);
nor U17162 (N_17162,N_14070,N_14362);
nand U17163 (N_17163,N_15706,N_15922);
and U17164 (N_17164,N_15454,N_15385);
nor U17165 (N_17165,N_15073,N_15432);
xnor U17166 (N_17166,N_14012,N_14841);
and U17167 (N_17167,N_14553,N_14882);
or U17168 (N_17168,N_14923,N_15798);
nand U17169 (N_17169,N_15209,N_15435);
and U17170 (N_17170,N_15842,N_15097);
or U17171 (N_17171,N_15484,N_15349);
or U17172 (N_17172,N_15492,N_15051);
or U17173 (N_17173,N_15111,N_14978);
nand U17174 (N_17174,N_15864,N_15255);
nand U17175 (N_17175,N_14691,N_14589);
xnor U17176 (N_17176,N_15381,N_15063);
nor U17177 (N_17177,N_15281,N_15567);
xnor U17178 (N_17178,N_14462,N_14863);
xnor U17179 (N_17179,N_15049,N_14428);
nand U17180 (N_17180,N_15534,N_15454);
nor U17181 (N_17181,N_15688,N_15807);
xor U17182 (N_17182,N_15749,N_15485);
or U17183 (N_17183,N_14916,N_15925);
xor U17184 (N_17184,N_14572,N_14557);
and U17185 (N_17185,N_14139,N_14970);
nand U17186 (N_17186,N_15679,N_14737);
xnor U17187 (N_17187,N_14251,N_15890);
xor U17188 (N_17188,N_14158,N_14323);
or U17189 (N_17189,N_14509,N_15347);
nand U17190 (N_17190,N_14903,N_14841);
and U17191 (N_17191,N_15851,N_14185);
nor U17192 (N_17192,N_14921,N_14438);
nor U17193 (N_17193,N_14159,N_15681);
or U17194 (N_17194,N_14657,N_15012);
nor U17195 (N_17195,N_14727,N_15678);
xor U17196 (N_17196,N_15598,N_15471);
nand U17197 (N_17197,N_15724,N_15188);
or U17198 (N_17198,N_15693,N_14660);
xor U17199 (N_17199,N_15836,N_14923);
nand U17200 (N_17200,N_14090,N_15070);
xnor U17201 (N_17201,N_15367,N_14844);
or U17202 (N_17202,N_15290,N_15565);
nor U17203 (N_17203,N_15317,N_14912);
and U17204 (N_17204,N_15482,N_14102);
nand U17205 (N_17205,N_15659,N_14658);
xor U17206 (N_17206,N_15688,N_15433);
or U17207 (N_17207,N_15782,N_14292);
nand U17208 (N_17208,N_14694,N_15018);
xor U17209 (N_17209,N_15689,N_15365);
xor U17210 (N_17210,N_14069,N_14678);
xor U17211 (N_17211,N_15305,N_15384);
or U17212 (N_17212,N_14155,N_14335);
and U17213 (N_17213,N_15724,N_15603);
and U17214 (N_17214,N_14633,N_14486);
and U17215 (N_17215,N_14470,N_14317);
nand U17216 (N_17216,N_14158,N_14623);
xor U17217 (N_17217,N_15016,N_14050);
and U17218 (N_17218,N_14492,N_14083);
xor U17219 (N_17219,N_15721,N_15941);
nand U17220 (N_17220,N_15206,N_14336);
nand U17221 (N_17221,N_15297,N_14410);
and U17222 (N_17222,N_15130,N_15383);
or U17223 (N_17223,N_14435,N_14793);
or U17224 (N_17224,N_14785,N_14834);
or U17225 (N_17225,N_14928,N_15816);
nand U17226 (N_17226,N_14954,N_14664);
xnor U17227 (N_17227,N_14518,N_15167);
or U17228 (N_17228,N_14648,N_15426);
and U17229 (N_17229,N_14821,N_14627);
and U17230 (N_17230,N_15461,N_14099);
and U17231 (N_17231,N_15254,N_14119);
or U17232 (N_17232,N_15344,N_15796);
or U17233 (N_17233,N_15575,N_15111);
nor U17234 (N_17234,N_15099,N_14714);
and U17235 (N_17235,N_14792,N_15150);
or U17236 (N_17236,N_14800,N_14209);
nand U17237 (N_17237,N_15037,N_14021);
or U17238 (N_17238,N_14393,N_14772);
nand U17239 (N_17239,N_14232,N_14503);
xor U17240 (N_17240,N_15234,N_14734);
nor U17241 (N_17241,N_15095,N_15192);
and U17242 (N_17242,N_14177,N_15726);
nand U17243 (N_17243,N_14834,N_14207);
nand U17244 (N_17244,N_14663,N_14923);
xor U17245 (N_17245,N_14015,N_15526);
nand U17246 (N_17246,N_15947,N_14559);
xor U17247 (N_17247,N_14604,N_14991);
nor U17248 (N_17248,N_15388,N_15231);
nor U17249 (N_17249,N_14475,N_14130);
and U17250 (N_17250,N_15955,N_15211);
nand U17251 (N_17251,N_15565,N_14166);
nor U17252 (N_17252,N_14546,N_14033);
xor U17253 (N_17253,N_15352,N_14874);
xnor U17254 (N_17254,N_15580,N_14086);
and U17255 (N_17255,N_14577,N_15103);
xor U17256 (N_17256,N_14884,N_15820);
nor U17257 (N_17257,N_15447,N_15661);
nand U17258 (N_17258,N_14389,N_15530);
nand U17259 (N_17259,N_14935,N_14666);
nor U17260 (N_17260,N_15842,N_15870);
xor U17261 (N_17261,N_15065,N_14354);
nand U17262 (N_17262,N_14520,N_15923);
and U17263 (N_17263,N_14455,N_15904);
xnor U17264 (N_17264,N_15035,N_14964);
nand U17265 (N_17265,N_15106,N_15630);
nor U17266 (N_17266,N_15169,N_14097);
and U17267 (N_17267,N_14149,N_15815);
and U17268 (N_17268,N_15080,N_15040);
nor U17269 (N_17269,N_15916,N_14894);
and U17270 (N_17270,N_15780,N_14650);
or U17271 (N_17271,N_14598,N_15049);
or U17272 (N_17272,N_14547,N_15125);
nand U17273 (N_17273,N_15718,N_15562);
nor U17274 (N_17274,N_14354,N_15485);
nor U17275 (N_17275,N_14043,N_14835);
and U17276 (N_17276,N_15512,N_14986);
xnor U17277 (N_17277,N_15119,N_15761);
nor U17278 (N_17278,N_15167,N_15212);
and U17279 (N_17279,N_14117,N_15585);
nand U17280 (N_17280,N_15401,N_14722);
nor U17281 (N_17281,N_14983,N_15648);
nand U17282 (N_17282,N_15517,N_14522);
and U17283 (N_17283,N_15484,N_15544);
xnor U17284 (N_17284,N_15638,N_15312);
nor U17285 (N_17285,N_15149,N_15726);
xnor U17286 (N_17286,N_14042,N_15128);
or U17287 (N_17287,N_14764,N_14485);
xor U17288 (N_17288,N_15720,N_14494);
nor U17289 (N_17289,N_15102,N_14147);
or U17290 (N_17290,N_14689,N_15337);
and U17291 (N_17291,N_14320,N_15748);
or U17292 (N_17292,N_15296,N_14785);
nand U17293 (N_17293,N_14507,N_14383);
or U17294 (N_17294,N_14841,N_15415);
nand U17295 (N_17295,N_15410,N_15878);
nor U17296 (N_17296,N_14114,N_14851);
and U17297 (N_17297,N_14045,N_15884);
xor U17298 (N_17298,N_14580,N_15506);
and U17299 (N_17299,N_15572,N_15216);
or U17300 (N_17300,N_15266,N_14101);
xor U17301 (N_17301,N_15410,N_15117);
nand U17302 (N_17302,N_15927,N_15111);
xnor U17303 (N_17303,N_15599,N_14673);
nand U17304 (N_17304,N_15212,N_15670);
and U17305 (N_17305,N_14172,N_14328);
nor U17306 (N_17306,N_14263,N_15050);
and U17307 (N_17307,N_15680,N_15579);
and U17308 (N_17308,N_14381,N_15494);
nand U17309 (N_17309,N_15064,N_14430);
or U17310 (N_17310,N_15556,N_15788);
and U17311 (N_17311,N_14153,N_15037);
nor U17312 (N_17312,N_15340,N_14193);
and U17313 (N_17313,N_14054,N_15777);
nand U17314 (N_17314,N_15135,N_14170);
or U17315 (N_17315,N_15038,N_15498);
nor U17316 (N_17316,N_14292,N_15584);
and U17317 (N_17317,N_14707,N_15919);
nor U17318 (N_17318,N_15418,N_15755);
nor U17319 (N_17319,N_14067,N_14838);
or U17320 (N_17320,N_14684,N_14329);
nand U17321 (N_17321,N_14854,N_14659);
xor U17322 (N_17322,N_14610,N_15805);
or U17323 (N_17323,N_14634,N_14179);
or U17324 (N_17324,N_15050,N_14363);
xnor U17325 (N_17325,N_14297,N_15433);
xor U17326 (N_17326,N_14351,N_15455);
xor U17327 (N_17327,N_15672,N_14226);
and U17328 (N_17328,N_15206,N_15730);
nand U17329 (N_17329,N_14620,N_14561);
nor U17330 (N_17330,N_15484,N_14238);
nand U17331 (N_17331,N_14264,N_14977);
and U17332 (N_17332,N_14132,N_14621);
and U17333 (N_17333,N_15050,N_14850);
and U17334 (N_17334,N_15364,N_14188);
or U17335 (N_17335,N_15813,N_15543);
nor U17336 (N_17336,N_15594,N_14359);
nand U17337 (N_17337,N_15588,N_14485);
and U17338 (N_17338,N_15117,N_15445);
nor U17339 (N_17339,N_14727,N_15133);
nor U17340 (N_17340,N_14526,N_14961);
or U17341 (N_17341,N_15334,N_15045);
nand U17342 (N_17342,N_14764,N_15407);
nand U17343 (N_17343,N_15889,N_15243);
nor U17344 (N_17344,N_15780,N_15590);
nand U17345 (N_17345,N_14056,N_14672);
nand U17346 (N_17346,N_15721,N_14940);
nor U17347 (N_17347,N_14526,N_14423);
nor U17348 (N_17348,N_14297,N_15387);
nor U17349 (N_17349,N_14367,N_15459);
or U17350 (N_17350,N_15811,N_15517);
nor U17351 (N_17351,N_15901,N_14328);
nor U17352 (N_17352,N_14769,N_15576);
nor U17353 (N_17353,N_14529,N_14955);
and U17354 (N_17354,N_15917,N_15857);
and U17355 (N_17355,N_15978,N_14932);
or U17356 (N_17356,N_14465,N_15196);
nor U17357 (N_17357,N_14020,N_15686);
nor U17358 (N_17358,N_14465,N_15555);
xor U17359 (N_17359,N_14297,N_14062);
nor U17360 (N_17360,N_15330,N_14894);
nor U17361 (N_17361,N_15533,N_15622);
nor U17362 (N_17362,N_14637,N_15018);
or U17363 (N_17363,N_15182,N_14089);
or U17364 (N_17364,N_15104,N_14528);
nand U17365 (N_17365,N_14578,N_15203);
or U17366 (N_17366,N_15223,N_15129);
nand U17367 (N_17367,N_15030,N_15531);
nand U17368 (N_17368,N_14404,N_15655);
and U17369 (N_17369,N_14717,N_14644);
xnor U17370 (N_17370,N_14139,N_15152);
xnor U17371 (N_17371,N_15665,N_15304);
nand U17372 (N_17372,N_14159,N_15081);
or U17373 (N_17373,N_14417,N_15062);
nand U17374 (N_17374,N_14189,N_14008);
and U17375 (N_17375,N_15975,N_15512);
xor U17376 (N_17376,N_14677,N_14590);
and U17377 (N_17377,N_14719,N_15765);
and U17378 (N_17378,N_15430,N_15075);
nor U17379 (N_17379,N_14214,N_15297);
nor U17380 (N_17380,N_15999,N_14606);
nand U17381 (N_17381,N_14838,N_14307);
and U17382 (N_17382,N_14192,N_14154);
xor U17383 (N_17383,N_14935,N_15553);
nor U17384 (N_17384,N_15416,N_14703);
and U17385 (N_17385,N_14214,N_15630);
nor U17386 (N_17386,N_14620,N_14129);
xnor U17387 (N_17387,N_14599,N_14003);
nand U17388 (N_17388,N_15643,N_15878);
nand U17389 (N_17389,N_15305,N_14278);
and U17390 (N_17390,N_15803,N_14440);
nor U17391 (N_17391,N_14049,N_15267);
nor U17392 (N_17392,N_14821,N_15452);
and U17393 (N_17393,N_15577,N_14372);
and U17394 (N_17394,N_15562,N_15432);
nor U17395 (N_17395,N_15508,N_14830);
or U17396 (N_17396,N_14646,N_15761);
nand U17397 (N_17397,N_14875,N_14841);
and U17398 (N_17398,N_15921,N_15865);
nand U17399 (N_17399,N_15885,N_15981);
or U17400 (N_17400,N_15335,N_15783);
or U17401 (N_17401,N_14797,N_15460);
nand U17402 (N_17402,N_15458,N_15704);
xnor U17403 (N_17403,N_15187,N_14123);
or U17404 (N_17404,N_14712,N_15571);
nor U17405 (N_17405,N_15904,N_14480);
nor U17406 (N_17406,N_15167,N_14167);
nor U17407 (N_17407,N_14471,N_14039);
or U17408 (N_17408,N_14187,N_14272);
nand U17409 (N_17409,N_15471,N_14638);
xnor U17410 (N_17410,N_15348,N_14816);
nor U17411 (N_17411,N_15671,N_15563);
and U17412 (N_17412,N_14386,N_14582);
xor U17413 (N_17413,N_15919,N_15530);
nor U17414 (N_17414,N_15372,N_15943);
xor U17415 (N_17415,N_15738,N_15108);
and U17416 (N_17416,N_15611,N_14706);
nand U17417 (N_17417,N_14502,N_14317);
or U17418 (N_17418,N_15068,N_14982);
nor U17419 (N_17419,N_14739,N_14354);
and U17420 (N_17420,N_14677,N_15905);
nor U17421 (N_17421,N_15033,N_15528);
nor U17422 (N_17422,N_14215,N_15775);
nor U17423 (N_17423,N_14318,N_15201);
nor U17424 (N_17424,N_15395,N_15913);
or U17425 (N_17425,N_14098,N_14813);
nand U17426 (N_17426,N_15131,N_14515);
nor U17427 (N_17427,N_15348,N_15697);
and U17428 (N_17428,N_15798,N_15107);
or U17429 (N_17429,N_15282,N_14179);
nor U17430 (N_17430,N_14911,N_15691);
and U17431 (N_17431,N_15480,N_15792);
xnor U17432 (N_17432,N_15719,N_14287);
nand U17433 (N_17433,N_15273,N_14212);
xnor U17434 (N_17434,N_14871,N_14881);
and U17435 (N_17435,N_14118,N_14597);
nand U17436 (N_17436,N_15580,N_14360);
nor U17437 (N_17437,N_15923,N_14892);
and U17438 (N_17438,N_15969,N_15307);
and U17439 (N_17439,N_15021,N_14883);
xnor U17440 (N_17440,N_14655,N_14241);
and U17441 (N_17441,N_14169,N_15074);
and U17442 (N_17442,N_15945,N_14975);
xor U17443 (N_17443,N_14575,N_15812);
xnor U17444 (N_17444,N_14163,N_15993);
nand U17445 (N_17445,N_14086,N_15204);
xnor U17446 (N_17446,N_14189,N_14561);
and U17447 (N_17447,N_14475,N_15500);
xnor U17448 (N_17448,N_14272,N_14718);
xor U17449 (N_17449,N_14861,N_14989);
nand U17450 (N_17450,N_15967,N_15915);
nand U17451 (N_17451,N_14617,N_15142);
and U17452 (N_17452,N_14469,N_14924);
and U17453 (N_17453,N_14010,N_14570);
nand U17454 (N_17454,N_15351,N_15458);
and U17455 (N_17455,N_15707,N_15658);
nor U17456 (N_17456,N_15416,N_14158);
or U17457 (N_17457,N_15053,N_15095);
and U17458 (N_17458,N_14399,N_14679);
nand U17459 (N_17459,N_15676,N_15210);
or U17460 (N_17460,N_15337,N_14591);
or U17461 (N_17461,N_15911,N_15578);
nand U17462 (N_17462,N_15842,N_15768);
nor U17463 (N_17463,N_14266,N_15026);
or U17464 (N_17464,N_15292,N_14450);
and U17465 (N_17465,N_14062,N_14998);
and U17466 (N_17466,N_14934,N_15198);
and U17467 (N_17467,N_14423,N_14442);
and U17468 (N_17468,N_15391,N_15289);
xnor U17469 (N_17469,N_14427,N_14125);
nand U17470 (N_17470,N_14994,N_15215);
xnor U17471 (N_17471,N_14469,N_14519);
nand U17472 (N_17472,N_14478,N_15833);
and U17473 (N_17473,N_15317,N_14987);
nor U17474 (N_17474,N_15512,N_14078);
nor U17475 (N_17475,N_14054,N_15059);
xnor U17476 (N_17476,N_14081,N_14696);
nor U17477 (N_17477,N_15570,N_14159);
and U17478 (N_17478,N_15230,N_14309);
nand U17479 (N_17479,N_15739,N_15738);
and U17480 (N_17480,N_14383,N_15661);
xnor U17481 (N_17481,N_14256,N_15866);
and U17482 (N_17482,N_15703,N_15624);
nand U17483 (N_17483,N_15053,N_14258);
nand U17484 (N_17484,N_15036,N_14370);
or U17485 (N_17485,N_14943,N_14027);
nor U17486 (N_17486,N_15419,N_14145);
and U17487 (N_17487,N_15429,N_15984);
nand U17488 (N_17488,N_14527,N_15219);
and U17489 (N_17489,N_15721,N_15718);
or U17490 (N_17490,N_14357,N_15124);
nor U17491 (N_17491,N_14286,N_14464);
and U17492 (N_17492,N_14730,N_14486);
or U17493 (N_17493,N_15846,N_14604);
nor U17494 (N_17494,N_14098,N_14368);
nor U17495 (N_17495,N_15968,N_14910);
and U17496 (N_17496,N_14790,N_15047);
or U17497 (N_17497,N_15375,N_14420);
xnor U17498 (N_17498,N_14048,N_15396);
xor U17499 (N_17499,N_14170,N_15464);
nor U17500 (N_17500,N_14711,N_14851);
nor U17501 (N_17501,N_15623,N_14845);
nand U17502 (N_17502,N_14858,N_15244);
nand U17503 (N_17503,N_15945,N_14814);
or U17504 (N_17504,N_14174,N_14305);
nor U17505 (N_17505,N_15648,N_15749);
nor U17506 (N_17506,N_15815,N_14832);
or U17507 (N_17507,N_14838,N_14619);
or U17508 (N_17508,N_15093,N_14706);
nor U17509 (N_17509,N_15184,N_14098);
and U17510 (N_17510,N_15846,N_15699);
nand U17511 (N_17511,N_14633,N_15699);
xor U17512 (N_17512,N_15906,N_14177);
and U17513 (N_17513,N_15455,N_15071);
xor U17514 (N_17514,N_14955,N_14244);
xnor U17515 (N_17515,N_15427,N_15371);
nor U17516 (N_17516,N_15376,N_14339);
nor U17517 (N_17517,N_14806,N_15199);
nor U17518 (N_17518,N_15108,N_15439);
nor U17519 (N_17519,N_14166,N_14470);
nor U17520 (N_17520,N_15787,N_14632);
or U17521 (N_17521,N_14544,N_15554);
nand U17522 (N_17522,N_15872,N_14553);
or U17523 (N_17523,N_15846,N_15147);
xnor U17524 (N_17524,N_15932,N_15907);
xnor U17525 (N_17525,N_14334,N_14589);
nand U17526 (N_17526,N_14755,N_15365);
nand U17527 (N_17527,N_15205,N_14577);
nor U17528 (N_17528,N_14361,N_15275);
nor U17529 (N_17529,N_15679,N_15377);
nor U17530 (N_17530,N_15842,N_15828);
xor U17531 (N_17531,N_14148,N_14061);
xnor U17532 (N_17532,N_15803,N_14263);
nand U17533 (N_17533,N_15535,N_14034);
nor U17534 (N_17534,N_15408,N_15276);
nor U17535 (N_17535,N_14100,N_15450);
xor U17536 (N_17536,N_14017,N_14244);
nand U17537 (N_17537,N_14980,N_15913);
nor U17538 (N_17538,N_15642,N_14716);
nand U17539 (N_17539,N_14083,N_15840);
nor U17540 (N_17540,N_14880,N_15012);
nor U17541 (N_17541,N_14672,N_14750);
and U17542 (N_17542,N_14016,N_15935);
xnor U17543 (N_17543,N_14417,N_15427);
and U17544 (N_17544,N_15017,N_15715);
xor U17545 (N_17545,N_14990,N_14926);
nand U17546 (N_17546,N_15641,N_14737);
or U17547 (N_17547,N_15653,N_14142);
or U17548 (N_17548,N_14567,N_14277);
and U17549 (N_17549,N_14117,N_15780);
nand U17550 (N_17550,N_14536,N_14480);
or U17551 (N_17551,N_15206,N_15772);
xnor U17552 (N_17552,N_15066,N_15881);
nand U17553 (N_17553,N_14845,N_15599);
or U17554 (N_17554,N_14740,N_14579);
nand U17555 (N_17555,N_15325,N_15428);
xnor U17556 (N_17556,N_15399,N_14287);
nand U17557 (N_17557,N_15311,N_14235);
nand U17558 (N_17558,N_15138,N_15061);
xor U17559 (N_17559,N_15074,N_15755);
and U17560 (N_17560,N_15543,N_14972);
nand U17561 (N_17561,N_15859,N_14797);
nand U17562 (N_17562,N_14119,N_14619);
and U17563 (N_17563,N_14551,N_15105);
xnor U17564 (N_17564,N_15129,N_15183);
and U17565 (N_17565,N_15975,N_14913);
or U17566 (N_17566,N_14183,N_15719);
nor U17567 (N_17567,N_15558,N_15872);
nor U17568 (N_17568,N_14192,N_14330);
nand U17569 (N_17569,N_15795,N_15233);
nor U17570 (N_17570,N_15972,N_14047);
or U17571 (N_17571,N_14694,N_15488);
xnor U17572 (N_17572,N_15245,N_15667);
xor U17573 (N_17573,N_14866,N_14071);
nand U17574 (N_17574,N_14349,N_15801);
xor U17575 (N_17575,N_15223,N_15847);
nand U17576 (N_17576,N_15806,N_14253);
and U17577 (N_17577,N_14510,N_15344);
and U17578 (N_17578,N_14126,N_15482);
or U17579 (N_17579,N_14998,N_15519);
or U17580 (N_17580,N_14648,N_14907);
and U17581 (N_17581,N_14894,N_14194);
xor U17582 (N_17582,N_14753,N_15530);
and U17583 (N_17583,N_15215,N_14073);
xnor U17584 (N_17584,N_14316,N_14346);
or U17585 (N_17585,N_14694,N_14060);
xor U17586 (N_17586,N_14661,N_14374);
xnor U17587 (N_17587,N_15447,N_14035);
nand U17588 (N_17588,N_14419,N_15493);
or U17589 (N_17589,N_15367,N_14422);
xnor U17590 (N_17590,N_14943,N_15822);
nand U17591 (N_17591,N_14915,N_14289);
nor U17592 (N_17592,N_15620,N_14593);
or U17593 (N_17593,N_15686,N_15239);
xnor U17594 (N_17594,N_15259,N_15326);
nand U17595 (N_17595,N_14151,N_14230);
nand U17596 (N_17596,N_14163,N_14344);
nor U17597 (N_17597,N_15644,N_15352);
xor U17598 (N_17598,N_14430,N_15155);
xor U17599 (N_17599,N_15723,N_15803);
nor U17600 (N_17600,N_15423,N_14971);
and U17601 (N_17601,N_14973,N_15692);
or U17602 (N_17602,N_14215,N_15143);
or U17603 (N_17603,N_15807,N_14235);
nor U17604 (N_17604,N_14540,N_14258);
xor U17605 (N_17605,N_14315,N_15545);
nor U17606 (N_17606,N_15889,N_14325);
nor U17607 (N_17607,N_14934,N_15733);
xnor U17608 (N_17608,N_14769,N_15792);
nand U17609 (N_17609,N_15385,N_15400);
or U17610 (N_17610,N_14655,N_14228);
and U17611 (N_17611,N_15285,N_14640);
xor U17612 (N_17612,N_15180,N_15653);
and U17613 (N_17613,N_14865,N_15071);
and U17614 (N_17614,N_14703,N_15859);
nor U17615 (N_17615,N_14840,N_15587);
nand U17616 (N_17616,N_14103,N_15028);
nand U17617 (N_17617,N_14796,N_14413);
nand U17618 (N_17618,N_14069,N_15417);
xnor U17619 (N_17619,N_15882,N_15649);
or U17620 (N_17620,N_15619,N_15811);
nor U17621 (N_17621,N_15545,N_14688);
xor U17622 (N_17622,N_14560,N_14147);
and U17623 (N_17623,N_14621,N_15938);
nor U17624 (N_17624,N_15815,N_15792);
xnor U17625 (N_17625,N_14705,N_14985);
nor U17626 (N_17626,N_15208,N_14526);
nand U17627 (N_17627,N_14125,N_15537);
nor U17628 (N_17628,N_15795,N_14522);
or U17629 (N_17629,N_14388,N_14845);
xor U17630 (N_17630,N_14103,N_15193);
or U17631 (N_17631,N_14393,N_14811);
and U17632 (N_17632,N_14191,N_14651);
nor U17633 (N_17633,N_15382,N_15591);
xnor U17634 (N_17634,N_15299,N_14256);
and U17635 (N_17635,N_14839,N_15755);
nor U17636 (N_17636,N_14613,N_15539);
and U17637 (N_17637,N_15001,N_14713);
nand U17638 (N_17638,N_15510,N_14634);
nor U17639 (N_17639,N_14867,N_15436);
and U17640 (N_17640,N_14318,N_14999);
and U17641 (N_17641,N_14126,N_14646);
xor U17642 (N_17642,N_15443,N_15416);
nor U17643 (N_17643,N_15307,N_15526);
or U17644 (N_17644,N_15589,N_15971);
or U17645 (N_17645,N_15484,N_15457);
xnor U17646 (N_17646,N_14841,N_15124);
nand U17647 (N_17647,N_14058,N_14475);
xnor U17648 (N_17648,N_15006,N_14938);
xnor U17649 (N_17649,N_14156,N_15089);
nor U17650 (N_17650,N_14481,N_15916);
and U17651 (N_17651,N_15892,N_14646);
or U17652 (N_17652,N_15816,N_14456);
or U17653 (N_17653,N_15928,N_14040);
nor U17654 (N_17654,N_14497,N_15113);
nand U17655 (N_17655,N_14030,N_14271);
and U17656 (N_17656,N_14948,N_15258);
xnor U17657 (N_17657,N_14352,N_15516);
xor U17658 (N_17658,N_14590,N_14826);
and U17659 (N_17659,N_14421,N_15470);
nand U17660 (N_17660,N_14053,N_14364);
and U17661 (N_17661,N_15493,N_15298);
nand U17662 (N_17662,N_14844,N_15050);
nand U17663 (N_17663,N_14538,N_15921);
or U17664 (N_17664,N_15713,N_14155);
xor U17665 (N_17665,N_15135,N_14589);
xor U17666 (N_17666,N_15450,N_15890);
xnor U17667 (N_17667,N_15060,N_14089);
nand U17668 (N_17668,N_15222,N_15507);
xor U17669 (N_17669,N_15561,N_15569);
and U17670 (N_17670,N_15277,N_14776);
nand U17671 (N_17671,N_15986,N_15665);
and U17672 (N_17672,N_14100,N_15907);
xor U17673 (N_17673,N_14388,N_15693);
or U17674 (N_17674,N_15957,N_15802);
nor U17675 (N_17675,N_14523,N_15490);
nor U17676 (N_17676,N_15393,N_14644);
nand U17677 (N_17677,N_15754,N_14889);
nand U17678 (N_17678,N_14010,N_15296);
and U17679 (N_17679,N_14944,N_14420);
or U17680 (N_17680,N_14889,N_14127);
xor U17681 (N_17681,N_14208,N_14801);
nor U17682 (N_17682,N_14177,N_14830);
xor U17683 (N_17683,N_15507,N_14855);
nor U17684 (N_17684,N_15225,N_14604);
xor U17685 (N_17685,N_15845,N_14635);
or U17686 (N_17686,N_15682,N_15608);
nor U17687 (N_17687,N_14117,N_15088);
xor U17688 (N_17688,N_14036,N_14678);
xor U17689 (N_17689,N_15285,N_15027);
nor U17690 (N_17690,N_15201,N_15074);
nand U17691 (N_17691,N_14520,N_14477);
xor U17692 (N_17692,N_15043,N_14525);
nand U17693 (N_17693,N_14114,N_14207);
and U17694 (N_17694,N_15332,N_15385);
nor U17695 (N_17695,N_14296,N_14114);
xnor U17696 (N_17696,N_14127,N_14108);
nor U17697 (N_17697,N_15777,N_14058);
or U17698 (N_17698,N_14441,N_14323);
and U17699 (N_17699,N_14146,N_14852);
xnor U17700 (N_17700,N_15236,N_15971);
nor U17701 (N_17701,N_15539,N_15404);
and U17702 (N_17702,N_14287,N_14181);
xnor U17703 (N_17703,N_15410,N_14123);
nand U17704 (N_17704,N_15037,N_14884);
or U17705 (N_17705,N_14259,N_15963);
or U17706 (N_17706,N_14255,N_14958);
and U17707 (N_17707,N_15837,N_15801);
xor U17708 (N_17708,N_14076,N_14010);
and U17709 (N_17709,N_14380,N_15873);
and U17710 (N_17710,N_14741,N_15941);
xnor U17711 (N_17711,N_15502,N_14123);
nand U17712 (N_17712,N_14262,N_14535);
and U17713 (N_17713,N_14948,N_14382);
nor U17714 (N_17714,N_15904,N_15554);
nor U17715 (N_17715,N_15159,N_14374);
and U17716 (N_17716,N_14737,N_14736);
or U17717 (N_17717,N_15541,N_14162);
or U17718 (N_17718,N_14581,N_15669);
nand U17719 (N_17719,N_15683,N_14886);
xor U17720 (N_17720,N_15619,N_14274);
nand U17721 (N_17721,N_14775,N_15883);
xor U17722 (N_17722,N_15590,N_15671);
and U17723 (N_17723,N_15140,N_15375);
xor U17724 (N_17724,N_15360,N_15415);
nand U17725 (N_17725,N_14152,N_14151);
or U17726 (N_17726,N_15003,N_14835);
and U17727 (N_17727,N_14127,N_14167);
or U17728 (N_17728,N_14633,N_14662);
nor U17729 (N_17729,N_15665,N_14476);
nor U17730 (N_17730,N_15633,N_14733);
and U17731 (N_17731,N_14364,N_15730);
or U17732 (N_17732,N_14833,N_15183);
and U17733 (N_17733,N_14317,N_14276);
xor U17734 (N_17734,N_14840,N_15215);
xnor U17735 (N_17735,N_15259,N_14711);
and U17736 (N_17736,N_15074,N_14380);
xnor U17737 (N_17737,N_15995,N_15182);
xor U17738 (N_17738,N_14406,N_14389);
xor U17739 (N_17739,N_14868,N_14265);
nor U17740 (N_17740,N_14820,N_14353);
xor U17741 (N_17741,N_14667,N_15454);
xnor U17742 (N_17742,N_14709,N_14750);
and U17743 (N_17743,N_14316,N_15055);
nor U17744 (N_17744,N_15336,N_15875);
xor U17745 (N_17745,N_14190,N_15750);
xnor U17746 (N_17746,N_15755,N_14276);
and U17747 (N_17747,N_14483,N_14373);
xor U17748 (N_17748,N_15465,N_14957);
nor U17749 (N_17749,N_14651,N_15866);
xor U17750 (N_17750,N_15392,N_15478);
nor U17751 (N_17751,N_14811,N_14676);
xor U17752 (N_17752,N_15026,N_15683);
and U17753 (N_17753,N_14860,N_15444);
nor U17754 (N_17754,N_14354,N_14119);
nor U17755 (N_17755,N_14194,N_14217);
and U17756 (N_17756,N_15225,N_15270);
or U17757 (N_17757,N_14444,N_15172);
and U17758 (N_17758,N_15872,N_14568);
nor U17759 (N_17759,N_14660,N_14385);
xor U17760 (N_17760,N_15127,N_14509);
xnor U17761 (N_17761,N_15206,N_14459);
nand U17762 (N_17762,N_15198,N_14263);
xor U17763 (N_17763,N_15196,N_14498);
and U17764 (N_17764,N_14621,N_15792);
xnor U17765 (N_17765,N_15659,N_14179);
xnor U17766 (N_17766,N_14722,N_15573);
and U17767 (N_17767,N_14249,N_15545);
nand U17768 (N_17768,N_15674,N_14111);
nand U17769 (N_17769,N_14820,N_15290);
and U17770 (N_17770,N_15040,N_15222);
xor U17771 (N_17771,N_15626,N_14557);
nor U17772 (N_17772,N_14748,N_14092);
and U17773 (N_17773,N_15697,N_15565);
xor U17774 (N_17774,N_15941,N_14632);
nand U17775 (N_17775,N_14954,N_15078);
or U17776 (N_17776,N_15485,N_15676);
nor U17777 (N_17777,N_14719,N_14907);
or U17778 (N_17778,N_15959,N_14286);
nor U17779 (N_17779,N_15907,N_14791);
xor U17780 (N_17780,N_15567,N_15950);
xor U17781 (N_17781,N_14464,N_15214);
and U17782 (N_17782,N_15790,N_14403);
nand U17783 (N_17783,N_15868,N_15619);
or U17784 (N_17784,N_14956,N_14498);
nor U17785 (N_17785,N_15227,N_15952);
or U17786 (N_17786,N_14684,N_15851);
xor U17787 (N_17787,N_15897,N_14701);
or U17788 (N_17788,N_14212,N_15018);
xor U17789 (N_17789,N_14476,N_15675);
and U17790 (N_17790,N_14563,N_14370);
or U17791 (N_17791,N_15141,N_14732);
nor U17792 (N_17792,N_14322,N_14905);
nor U17793 (N_17793,N_15647,N_15194);
nor U17794 (N_17794,N_14814,N_15136);
or U17795 (N_17795,N_14621,N_14989);
nand U17796 (N_17796,N_14598,N_14348);
xor U17797 (N_17797,N_15173,N_14765);
or U17798 (N_17798,N_14283,N_14277);
xor U17799 (N_17799,N_14878,N_14495);
nor U17800 (N_17800,N_15308,N_14964);
nor U17801 (N_17801,N_15047,N_15906);
and U17802 (N_17802,N_15449,N_15971);
nand U17803 (N_17803,N_14899,N_14177);
nor U17804 (N_17804,N_14946,N_15252);
or U17805 (N_17805,N_15712,N_14600);
nand U17806 (N_17806,N_15376,N_15689);
nor U17807 (N_17807,N_14539,N_15859);
or U17808 (N_17808,N_14714,N_15195);
or U17809 (N_17809,N_14925,N_14868);
nand U17810 (N_17810,N_14963,N_14824);
and U17811 (N_17811,N_14930,N_14085);
nand U17812 (N_17812,N_14501,N_14161);
nand U17813 (N_17813,N_15336,N_14506);
nand U17814 (N_17814,N_14908,N_14477);
xnor U17815 (N_17815,N_15938,N_14124);
xnor U17816 (N_17816,N_14643,N_14305);
xnor U17817 (N_17817,N_15248,N_15118);
nand U17818 (N_17818,N_15297,N_15555);
and U17819 (N_17819,N_15356,N_14153);
and U17820 (N_17820,N_15491,N_14833);
or U17821 (N_17821,N_14146,N_15727);
or U17822 (N_17822,N_15455,N_15468);
xor U17823 (N_17823,N_15399,N_14996);
nand U17824 (N_17824,N_14930,N_14166);
and U17825 (N_17825,N_14664,N_15530);
and U17826 (N_17826,N_15625,N_14360);
nand U17827 (N_17827,N_14544,N_14270);
or U17828 (N_17828,N_15866,N_14889);
xnor U17829 (N_17829,N_14845,N_15743);
or U17830 (N_17830,N_15098,N_14023);
nand U17831 (N_17831,N_14736,N_15417);
nor U17832 (N_17832,N_15751,N_15604);
nand U17833 (N_17833,N_14631,N_15762);
and U17834 (N_17834,N_15908,N_15321);
nand U17835 (N_17835,N_14508,N_15086);
nand U17836 (N_17836,N_15147,N_15967);
and U17837 (N_17837,N_14728,N_14156);
nor U17838 (N_17838,N_14772,N_15542);
xnor U17839 (N_17839,N_14506,N_14414);
and U17840 (N_17840,N_14573,N_14079);
nor U17841 (N_17841,N_14985,N_14232);
nand U17842 (N_17842,N_15125,N_14923);
nor U17843 (N_17843,N_15977,N_14328);
xor U17844 (N_17844,N_14798,N_15569);
xor U17845 (N_17845,N_15396,N_15327);
nor U17846 (N_17846,N_14821,N_15689);
or U17847 (N_17847,N_14005,N_14064);
nor U17848 (N_17848,N_14454,N_14803);
and U17849 (N_17849,N_15180,N_14842);
xor U17850 (N_17850,N_15901,N_15132);
xor U17851 (N_17851,N_14244,N_15693);
and U17852 (N_17852,N_15772,N_15021);
xnor U17853 (N_17853,N_15618,N_15909);
nor U17854 (N_17854,N_14068,N_15463);
and U17855 (N_17855,N_15633,N_15732);
or U17856 (N_17856,N_14373,N_15292);
or U17857 (N_17857,N_15268,N_14653);
or U17858 (N_17858,N_14098,N_14217);
and U17859 (N_17859,N_15810,N_14144);
nor U17860 (N_17860,N_14319,N_14130);
or U17861 (N_17861,N_15434,N_15737);
nor U17862 (N_17862,N_14299,N_14122);
nand U17863 (N_17863,N_15949,N_14740);
nor U17864 (N_17864,N_15476,N_15173);
nand U17865 (N_17865,N_15382,N_14551);
xnor U17866 (N_17866,N_14976,N_14704);
or U17867 (N_17867,N_15226,N_14631);
or U17868 (N_17868,N_15076,N_14413);
or U17869 (N_17869,N_15288,N_14287);
xnor U17870 (N_17870,N_14891,N_14057);
xnor U17871 (N_17871,N_14010,N_14100);
nand U17872 (N_17872,N_15298,N_15213);
nand U17873 (N_17873,N_15148,N_14315);
xor U17874 (N_17874,N_15287,N_14653);
and U17875 (N_17875,N_14460,N_15160);
xor U17876 (N_17876,N_14072,N_14200);
nor U17877 (N_17877,N_15514,N_15102);
or U17878 (N_17878,N_14841,N_14307);
nor U17879 (N_17879,N_15149,N_15336);
and U17880 (N_17880,N_14407,N_15613);
and U17881 (N_17881,N_14543,N_14046);
xor U17882 (N_17882,N_15716,N_14961);
or U17883 (N_17883,N_15993,N_15752);
nor U17884 (N_17884,N_14830,N_14734);
xnor U17885 (N_17885,N_14860,N_14560);
nand U17886 (N_17886,N_15543,N_15104);
or U17887 (N_17887,N_14889,N_15801);
nor U17888 (N_17888,N_15196,N_14826);
nor U17889 (N_17889,N_14195,N_14520);
or U17890 (N_17890,N_15690,N_15320);
and U17891 (N_17891,N_14010,N_15194);
xor U17892 (N_17892,N_14227,N_15323);
nand U17893 (N_17893,N_15517,N_14677);
and U17894 (N_17894,N_14594,N_15022);
xor U17895 (N_17895,N_14894,N_14313);
xnor U17896 (N_17896,N_14541,N_14871);
nand U17897 (N_17897,N_14863,N_14473);
nor U17898 (N_17898,N_14860,N_14319);
nand U17899 (N_17899,N_15171,N_15970);
nor U17900 (N_17900,N_14119,N_14847);
or U17901 (N_17901,N_15610,N_14356);
nor U17902 (N_17902,N_15390,N_15585);
nor U17903 (N_17903,N_14434,N_15709);
and U17904 (N_17904,N_15338,N_14924);
and U17905 (N_17905,N_14530,N_15175);
nand U17906 (N_17906,N_15684,N_15166);
and U17907 (N_17907,N_15071,N_15694);
nand U17908 (N_17908,N_15236,N_15130);
xnor U17909 (N_17909,N_14016,N_14923);
and U17910 (N_17910,N_14794,N_14325);
nand U17911 (N_17911,N_14773,N_15042);
xor U17912 (N_17912,N_15186,N_14423);
or U17913 (N_17913,N_15645,N_14840);
nor U17914 (N_17914,N_15319,N_15281);
and U17915 (N_17915,N_14245,N_15660);
nor U17916 (N_17916,N_15024,N_14792);
or U17917 (N_17917,N_15298,N_15441);
nor U17918 (N_17918,N_14871,N_14936);
xnor U17919 (N_17919,N_14125,N_14610);
xnor U17920 (N_17920,N_14213,N_14147);
or U17921 (N_17921,N_15737,N_14665);
or U17922 (N_17922,N_14786,N_15641);
or U17923 (N_17923,N_15272,N_15739);
nand U17924 (N_17924,N_15616,N_15209);
nor U17925 (N_17925,N_14693,N_15981);
xor U17926 (N_17926,N_15668,N_15703);
nand U17927 (N_17927,N_15590,N_15379);
xnor U17928 (N_17928,N_15513,N_14109);
and U17929 (N_17929,N_15342,N_14359);
xnor U17930 (N_17930,N_15294,N_14759);
or U17931 (N_17931,N_15781,N_15325);
xnor U17932 (N_17932,N_14018,N_15125);
nand U17933 (N_17933,N_15275,N_15165);
and U17934 (N_17934,N_14533,N_14429);
nor U17935 (N_17935,N_14122,N_14647);
or U17936 (N_17936,N_15507,N_14710);
xnor U17937 (N_17937,N_15108,N_15380);
or U17938 (N_17938,N_15958,N_15066);
xor U17939 (N_17939,N_15821,N_15455);
nor U17940 (N_17940,N_15819,N_14261);
and U17941 (N_17941,N_14712,N_14134);
nand U17942 (N_17942,N_15353,N_14664);
nand U17943 (N_17943,N_14849,N_15747);
xor U17944 (N_17944,N_14373,N_15075);
nor U17945 (N_17945,N_14975,N_15301);
and U17946 (N_17946,N_14758,N_15728);
nand U17947 (N_17947,N_14915,N_15790);
nand U17948 (N_17948,N_14899,N_15474);
xor U17949 (N_17949,N_15427,N_15912);
xnor U17950 (N_17950,N_14602,N_14790);
and U17951 (N_17951,N_15273,N_15024);
xnor U17952 (N_17952,N_14455,N_15064);
and U17953 (N_17953,N_15836,N_14640);
or U17954 (N_17954,N_15955,N_14354);
nor U17955 (N_17955,N_14147,N_14608);
nor U17956 (N_17956,N_15138,N_15706);
nor U17957 (N_17957,N_15743,N_15267);
xnor U17958 (N_17958,N_14399,N_14070);
nand U17959 (N_17959,N_14380,N_14038);
nand U17960 (N_17960,N_14927,N_14472);
or U17961 (N_17961,N_15164,N_14527);
or U17962 (N_17962,N_14534,N_15792);
or U17963 (N_17963,N_14640,N_14289);
xor U17964 (N_17964,N_15958,N_15013);
nand U17965 (N_17965,N_15253,N_15101);
or U17966 (N_17966,N_14909,N_14249);
or U17967 (N_17967,N_14518,N_14872);
xnor U17968 (N_17968,N_15131,N_14418);
nand U17969 (N_17969,N_15633,N_15783);
or U17970 (N_17970,N_14427,N_15808);
xnor U17971 (N_17971,N_15748,N_15939);
or U17972 (N_17972,N_15831,N_14901);
nand U17973 (N_17973,N_15847,N_14188);
xnor U17974 (N_17974,N_15932,N_14014);
or U17975 (N_17975,N_15973,N_14058);
and U17976 (N_17976,N_15224,N_15768);
or U17977 (N_17977,N_15168,N_15147);
nor U17978 (N_17978,N_15240,N_15653);
nor U17979 (N_17979,N_15222,N_14638);
and U17980 (N_17980,N_14454,N_14152);
and U17981 (N_17981,N_14609,N_15844);
and U17982 (N_17982,N_15833,N_14835);
xnor U17983 (N_17983,N_15567,N_14376);
xor U17984 (N_17984,N_15699,N_15616);
nand U17985 (N_17985,N_14085,N_14670);
nor U17986 (N_17986,N_15623,N_15999);
nand U17987 (N_17987,N_15990,N_14989);
xnor U17988 (N_17988,N_15378,N_15136);
or U17989 (N_17989,N_14572,N_15127);
nand U17990 (N_17990,N_14190,N_14336);
nand U17991 (N_17991,N_15497,N_15726);
and U17992 (N_17992,N_15989,N_14175);
and U17993 (N_17993,N_15201,N_15006);
xnor U17994 (N_17994,N_15855,N_15575);
xnor U17995 (N_17995,N_15963,N_14844);
or U17996 (N_17996,N_15729,N_15574);
xnor U17997 (N_17997,N_14620,N_15408);
xor U17998 (N_17998,N_14376,N_14171);
nand U17999 (N_17999,N_15558,N_15113);
or U18000 (N_18000,N_16065,N_16559);
xnor U18001 (N_18001,N_17473,N_17756);
or U18002 (N_18002,N_17511,N_16438);
and U18003 (N_18003,N_16641,N_16134);
nand U18004 (N_18004,N_17692,N_16150);
xnor U18005 (N_18005,N_16864,N_17388);
or U18006 (N_18006,N_17361,N_17804);
nor U18007 (N_18007,N_17063,N_17409);
nor U18008 (N_18008,N_16849,N_16482);
and U18009 (N_18009,N_16330,N_16887);
nand U18010 (N_18010,N_16106,N_17151);
and U18011 (N_18011,N_17449,N_17205);
and U18012 (N_18012,N_16934,N_16143);
and U18013 (N_18013,N_16568,N_16374);
nor U18014 (N_18014,N_16349,N_16229);
nand U18015 (N_18015,N_16920,N_16021);
or U18016 (N_18016,N_16178,N_17288);
nand U18017 (N_18017,N_17874,N_17013);
nor U18018 (N_18018,N_16933,N_17610);
nor U18019 (N_18019,N_16790,N_16671);
nor U18020 (N_18020,N_16263,N_17172);
nor U18021 (N_18021,N_17836,N_16453);
or U18022 (N_18022,N_17625,N_16596);
nor U18023 (N_18023,N_17468,N_17408);
nand U18024 (N_18024,N_16385,N_16504);
and U18025 (N_18025,N_17180,N_16310);
or U18026 (N_18026,N_16648,N_17275);
or U18027 (N_18027,N_16771,N_16042);
nor U18028 (N_18028,N_16830,N_17111);
or U18029 (N_18029,N_17157,N_16114);
and U18030 (N_18030,N_16531,N_16617);
xor U18031 (N_18031,N_16649,N_16287);
and U18032 (N_18032,N_16160,N_17305);
nor U18033 (N_18033,N_16490,N_17261);
nand U18034 (N_18034,N_17947,N_16600);
nand U18035 (N_18035,N_16081,N_16045);
or U18036 (N_18036,N_16866,N_16799);
or U18037 (N_18037,N_17389,N_16534);
nor U18038 (N_18038,N_17097,N_16540);
nand U18039 (N_18039,N_16867,N_17679);
or U18040 (N_18040,N_17726,N_16392);
or U18041 (N_18041,N_16204,N_16828);
nand U18042 (N_18042,N_17778,N_17474);
or U18043 (N_18043,N_16888,N_16476);
nand U18044 (N_18044,N_17050,N_16917);
nor U18045 (N_18045,N_17149,N_16121);
nand U18046 (N_18046,N_17764,N_16004);
or U18047 (N_18047,N_16789,N_16355);
or U18048 (N_18048,N_17426,N_16581);
nand U18049 (N_18049,N_16039,N_17696);
and U18050 (N_18050,N_17020,N_17958);
nand U18051 (N_18051,N_17249,N_16657);
nand U18052 (N_18052,N_17035,N_17752);
and U18053 (N_18053,N_16492,N_17347);
nand U18054 (N_18054,N_16725,N_16926);
or U18055 (N_18055,N_17533,N_16272);
nor U18056 (N_18056,N_17278,N_17216);
nor U18057 (N_18057,N_17255,N_17646);
nand U18058 (N_18058,N_17030,N_16523);
or U18059 (N_18059,N_16532,N_17173);
nor U18060 (N_18060,N_17319,N_17066);
and U18061 (N_18061,N_16970,N_17462);
xnor U18062 (N_18062,N_17669,N_16773);
or U18063 (N_18063,N_16136,N_17870);
or U18064 (N_18064,N_17745,N_17315);
and U18065 (N_18065,N_17605,N_17008);
xnor U18066 (N_18066,N_16881,N_17177);
or U18067 (N_18067,N_17144,N_16792);
nor U18068 (N_18068,N_16661,N_17419);
or U18069 (N_18069,N_17276,N_16459);
and U18070 (N_18070,N_17776,N_16687);
nand U18071 (N_18071,N_17964,N_16951);
and U18072 (N_18072,N_17711,N_17952);
or U18073 (N_18073,N_17951,N_17314);
nor U18074 (N_18074,N_17795,N_17913);
or U18075 (N_18075,N_17195,N_16109);
or U18076 (N_18076,N_17139,N_16537);
and U18077 (N_18077,N_16986,N_17940);
xnor U18078 (N_18078,N_16710,N_16588);
or U18079 (N_18079,N_17155,N_16611);
or U18080 (N_18080,N_17143,N_17790);
and U18081 (N_18081,N_17211,N_16550);
nand U18082 (N_18082,N_16275,N_16288);
xnor U18083 (N_18083,N_17571,N_17576);
nor U18084 (N_18084,N_17110,N_16095);
nand U18085 (N_18085,N_16479,N_17203);
or U18086 (N_18086,N_17443,N_17192);
nand U18087 (N_18087,N_17678,N_17023);
and U18088 (N_18088,N_16604,N_16696);
nand U18089 (N_18089,N_16026,N_16918);
nor U18090 (N_18090,N_16111,N_17971);
or U18091 (N_18091,N_17350,N_16505);
and U18092 (N_18092,N_17966,N_17675);
xor U18093 (N_18093,N_16660,N_17585);
and U18094 (N_18094,N_16521,N_17835);
or U18095 (N_18095,N_17648,N_16359);
nor U18096 (N_18096,N_16775,N_17842);
and U18097 (N_18097,N_17187,N_17374);
xor U18098 (N_18098,N_16304,N_16798);
nor U18099 (N_18099,N_16651,N_16421);
nand U18100 (N_18100,N_16590,N_16025);
nand U18101 (N_18101,N_16712,N_16836);
nor U18102 (N_18102,N_17580,N_16627);
nand U18103 (N_18103,N_17793,N_17346);
nand U18104 (N_18104,N_16736,N_16414);
nand U18105 (N_18105,N_16578,N_17717);
xor U18106 (N_18106,N_17472,N_16670);
nand U18107 (N_18107,N_17456,N_16742);
nor U18108 (N_18108,N_17856,N_17233);
nor U18109 (N_18109,N_16399,N_17201);
nor U18110 (N_18110,N_16658,N_17165);
xor U18111 (N_18111,N_17397,N_17674);
or U18112 (N_18112,N_17269,N_16442);
xnor U18113 (N_18113,N_16960,N_17744);
or U18114 (N_18114,N_16612,N_16377);
or U18115 (N_18115,N_17619,N_17991);
nand U18116 (N_18116,N_17093,N_16739);
xnor U18117 (N_18117,N_16577,N_17170);
nor U18118 (N_18118,N_17036,N_16211);
or U18119 (N_18119,N_16829,N_16549);
and U18120 (N_18120,N_16086,N_16890);
or U18121 (N_18121,N_16464,N_17943);
nand U18122 (N_18122,N_17916,N_16806);
and U18123 (N_18123,N_16312,N_17718);
xnor U18124 (N_18124,N_17125,N_17312);
xnor U18125 (N_18125,N_17156,N_16583);
xor U18126 (N_18126,N_16693,N_17387);
nand U18127 (N_18127,N_16551,N_16205);
and U18128 (N_18128,N_16754,N_17891);
or U18129 (N_18129,N_17207,N_16036);
and U18130 (N_18130,N_17961,N_17041);
nor U18131 (N_18131,N_17003,N_16848);
nor U18132 (N_18132,N_16198,N_16099);
or U18133 (N_18133,N_16524,N_17309);
and U18134 (N_18134,N_16619,N_16939);
nor U18135 (N_18135,N_16393,N_16560);
xnor U18136 (N_18136,N_17663,N_16317);
and U18137 (N_18137,N_16076,N_16984);
xnor U18138 (N_18138,N_16498,N_16292);
xor U18139 (N_18139,N_17955,N_17534);
xor U18140 (N_18140,N_17837,N_16652);
nand U18141 (N_18141,N_17875,N_17546);
or U18142 (N_18142,N_16512,N_16668);
nor U18143 (N_18143,N_16838,N_17911);
and U18144 (N_18144,N_17182,N_17828);
and U18145 (N_18145,N_16883,N_17059);
nand U18146 (N_18146,N_17259,N_16885);
nor U18147 (N_18147,N_16757,N_16700);
and U18148 (N_18148,N_16435,N_17236);
nor U18149 (N_18149,N_17591,N_17983);
xor U18150 (N_18150,N_17781,N_17672);
nand U18151 (N_18151,N_16235,N_16237);
nor U18152 (N_18152,N_16935,N_17789);
nor U18153 (N_18153,N_16842,N_17119);
xor U18154 (N_18154,N_16519,N_17649);
nor U18155 (N_18155,N_16470,N_17981);
nor U18156 (N_18156,N_16232,N_16103);
or U18157 (N_18157,N_17996,N_16751);
or U18158 (N_18158,N_17896,N_17611);
xnor U18159 (N_18159,N_16472,N_16118);
xnor U18160 (N_18160,N_17498,N_17355);
or U18161 (N_18161,N_17827,N_16953);
xor U18162 (N_18162,N_16930,N_16437);
and U18163 (N_18163,N_16663,N_17299);
nand U18164 (N_18164,N_17291,N_16522);
nand U18165 (N_18165,N_16796,N_17416);
and U18166 (N_18166,N_16625,N_17061);
nand U18167 (N_18167,N_16357,N_16572);
nand U18168 (N_18168,N_17710,N_17751);
nor U18169 (N_18169,N_16667,N_17936);
and U18170 (N_18170,N_17308,N_17514);
nor U18171 (N_18171,N_17923,N_17774);
nor U18172 (N_18172,N_17713,N_17666);
xor U18173 (N_18173,N_16616,N_16916);
or U18174 (N_18174,N_16394,N_16202);
nor U18175 (N_18175,N_17818,N_17258);
nand U18176 (N_18176,N_17920,N_17682);
xnor U18177 (N_18177,N_16869,N_17453);
nor U18178 (N_18178,N_17786,N_16213);
nand U18179 (N_18179,N_17163,N_17731);
and U18180 (N_18180,N_17454,N_16878);
and U18181 (N_18181,N_16297,N_17739);
xor U18182 (N_18182,N_16206,N_17803);
and U18183 (N_18183,N_16269,N_16159);
nand U18184 (N_18184,N_16173,N_16501);
nor U18185 (N_18185,N_16231,N_16078);
nor U18186 (N_18186,N_17242,N_16116);
xnor U18187 (N_18187,N_17171,N_16456);
nor U18188 (N_18188,N_17325,N_16928);
or U18189 (N_18189,N_16436,N_17014);
and U18190 (N_18190,N_16841,N_16937);
nand U18191 (N_18191,N_16580,N_17054);
xnor U18192 (N_18192,N_17104,N_17767);
or U18193 (N_18193,N_17274,N_16943);
and U18194 (N_18194,N_16419,N_16546);
nand U18195 (N_18195,N_16779,N_16098);
nand U18196 (N_18196,N_17244,N_16638);
nor U18197 (N_18197,N_17011,N_17915);
nor U18198 (N_18198,N_16452,N_16242);
nor U18199 (N_18199,N_16956,N_17892);
nand U18200 (N_18200,N_16728,N_16650);
xnor U18201 (N_18201,N_16972,N_16424);
nor U18202 (N_18202,N_17181,N_16791);
nor U18203 (N_18203,N_17503,N_16262);
or U18204 (N_18204,N_16711,N_17825);
xor U18205 (N_18205,N_16644,N_17372);
xnor U18206 (N_18206,N_17190,N_17526);
and U18207 (N_18207,N_16046,N_17425);
nand U18208 (N_18208,N_16748,N_17967);
or U18209 (N_18209,N_16276,N_16784);
nor U18210 (N_18210,N_16607,N_16759);
or U18211 (N_18211,N_17026,N_17217);
nand U18212 (N_18212,N_17561,N_16676);
nor U18213 (N_18213,N_16397,N_16915);
or U18214 (N_18214,N_17256,N_16138);
and U18215 (N_18215,N_17247,N_16019);
xor U18216 (N_18216,N_16450,N_17004);
and U18217 (N_18217,N_16162,N_16966);
nand U18218 (N_18218,N_17748,N_17266);
xor U18219 (N_18219,N_16383,N_16024);
and U18220 (N_18220,N_17525,N_16955);
xnor U18221 (N_18221,N_16015,N_16183);
xnor U18222 (N_18222,N_17229,N_16724);
nor U18223 (N_18223,N_16469,N_16620);
xor U18224 (N_18224,N_16738,N_17114);
nor U18225 (N_18225,N_16815,N_17701);
and U18226 (N_18226,N_16055,N_17475);
or U18227 (N_18227,N_16695,N_17343);
and U18228 (N_18228,N_17427,N_17019);
nand U18229 (N_18229,N_17279,N_16203);
xor U18230 (N_18230,N_17366,N_16694);
nor U18231 (N_18231,N_17001,N_16454);
xnor U18232 (N_18232,N_17594,N_16012);
nor U18233 (N_18233,N_17984,N_16431);
nor U18234 (N_18234,N_16023,N_16803);
nor U18235 (N_18235,N_17327,N_17841);
nor U18236 (N_18236,N_16264,N_16072);
nand U18237 (N_18237,N_17687,N_16413);
and U18238 (N_18238,N_17185,N_16073);
nor U18239 (N_18239,N_17307,N_16463);
xor U18240 (N_18240,N_16952,N_16518);
nand U18241 (N_18241,N_16043,N_17224);
or U18242 (N_18242,N_17417,N_17615);
nand U18243 (N_18243,N_16063,N_16749);
xnor U18244 (N_18244,N_17959,N_16455);
xor U18245 (N_18245,N_17942,N_17765);
and U18246 (N_18246,N_16767,N_16718);
xor U18247 (N_18247,N_17740,N_17862);
or U18248 (N_18248,N_16513,N_17385);
nor U18249 (N_18249,N_16682,N_16250);
xor U18250 (N_18250,N_16101,N_16837);
xnor U18251 (N_18251,N_16558,N_17147);
xnor U18252 (N_18252,N_16233,N_17694);
xnor U18253 (N_18253,N_16475,N_17797);
or U18254 (N_18254,N_17868,N_17444);
nand U18255 (N_18255,N_16684,N_17887);
xnor U18256 (N_18256,N_16416,N_17547);
xor U18257 (N_18257,N_17762,N_16007);
nor U18258 (N_18258,N_16904,N_17792);
xor U18259 (N_18259,N_16761,N_17895);
nor U18260 (N_18260,N_16851,N_16222);
and U18261 (N_18261,N_16329,N_16388);
xor U18262 (N_18262,N_16555,N_17714);
nor U18263 (N_18263,N_16339,N_16247);
nand U18264 (N_18264,N_16158,N_16514);
or U18265 (N_18265,N_17115,N_16702);
or U18266 (N_18266,N_16129,N_17685);
nand U18267 (N_18267,N_17016,N_17623);
nand U18268 (N_18268,N_16940,N_17654);
and U18269 (N_18269,N_17045,N_16253);
nor U18270 (N_18270,N_17065,N_17336);
or U18271 (N_18271,N_16566,N_16369);
or U18272 (N_18272,N_16654,N_17091);
nand U18273 (N_18273,N_17763,N_16239);
or U18274 (N_18274,N_16192,N_16786);
xor U18275 (N_18275,N_16194,N_16674);
or U18276 (N_18276,N_16112,N_17956);
nor U18277 (N_18277,N_16591,N_16238);
nor U18278 (N_18278,N_16876,N_16283);
nand U18279 (N_18279,N_17141,N_17396);
xor U18280 (N_18280,N_17878,N_17548);
nor U18281 (N_18281,N_16685,N_17301);
xnor U18282 (N_18282,N_16130,N_16857);
xnor U18283 (N_18283,N_16985,N_17791);
xnor U18284 (N_18284,N_17550,N_17889);
xor U18285 (N_18285,N_17829,N_16922);
xor U18286 (N_18286,N_16686,N_16659);
nor U18287 (N_18287,N_16066,N_17415);
or U18288 (N_18288,N_16995,N_16057);
xnor U18289 (N_18289,N_17912,N_17863);
nand U18290 (N_18290,N_16062,N_16166);
xnor U18291 (N_18291,N_17902,N_16161);
nor U18292 (N_18292,N_17502,N_16488);
and U18293 (N_18293,N_17549,N_16900);
and U18294 (N_18294,N_17824,N_16240);
and U18295 (N_18295,N_17189,N_16860);
nor U18296 (N_18296,N_16894,N_17957);
nor U18297 (N_18297,N_16809,N_17584);
and U18298 (N_18298,N_17176,N_16449);
nand U18299 (N_18299,N_17142,N_16755);
nor U18300 (N_18300,N_16919,N_16107);
and U18301 (N_18301,N_16533,N_17438);
nand U18302 (N_18302,N_16557,N_17819);
nand U18303 (N_18303,N_17706,N_17062);
and U18304 (N_18304,N_16389,N_17465);
or U18305 (N_18305,N_16426,N_16760);
nor U18306 (N_18306,N_17292,N_17908);
and U18307 (N_18307,N_17130,N_16365);
xor U18308 (N_18308,N_16884,N_16974);
and U18309 (N_18309,N_16647,N_17394);
nor U18310 (N_18310,N_16331,N_17976);
nand U18311 (N_18311,N_16945,N_17658);
nor U18312 (N_18312,N_17689,N_16681);
nand U18313 (N_18313,N_16520,N_16010);
or U18314 (N_18314,N_17127,N_16305);
or U18315 (N_18315,N_17496,N_16642);
nand U18316 (N_18316,N_16586,N_16959);
and U18317 (N_18317,N_16294,N_17643);
or U18318 (N_18318,N_17467,N_17169);
nor U18319 (N_18319,N_16669,N_17568);
or U18320 (N_18320,N_16003,N_17742);
and U18321 (N_18321,N_17563,N_17064);
nand U18322 (N_18322,N_17469,N_16993);
nor U18323 (N_18323,N_16144,N_17126);
nor U18324 (N_18324,N_16268,N_16741);
or U18325 (N_18325,N_16853,N_16373);
or U18326 (N_18326,N_17872,N_16541);
xor U18327 (N_18327,N_17633,N_17564);
nor U18328 (N_18328,N_17933,N_16207);
xnor U18329 (N_18329,N_16224,N_16196);
or U18330 (N_18330,N_16858,N_17452);
and U18331 (N_18331,N_17459,N_17608);
nor U18332 (N_18332,N_16195,N_16376);
nor U18333 (N_18333,N_16875,N_16177);
nand U18334 (N_18334,N_17284,N_17531);
xnor U18335 (N_18335,N_16054,N_17403);
xor U18336 (N_18336,N_16309,N_16047);
nor U18337 (N_18337,N_17593,N_16124);
nand U18338 (N_18338,N_16298,N_17962);
and U18339 (N_18339,N_16096,N_16163);
nand U18340 (N_18340,N_17510,N_17321);
or U18341 (N_18341,N_17414,N_16530);
nor U18342 (N_18342,N_16108,N_17929);
or U18343 (N_18343,N_17652,N_17138);
or U18344 (N_18344,N_16913,N_16731);
nand U18345 (N_18345,N_16418,N_17709);
xor U18346 (N_18346,N_17477,N_16484);
and U18347 (N_18347,N_17491,N_16936);
xor U18348 (N_18348,N_17822,N_16636);
nand U18349 (N_18349,N_17077,N_17831);
nand U18350 (N_18350,N_17551,N_17458);
nor U18351 (N_18351,N_17049,N_17555);
or U18352 (N_18352,N_16574,N_17304);
nand U18353 (N_18353,N_16990,N_17302);
or U18354 (N_18354,N_16303,N_16545);
or U18355 (N_18355,N_16104,N_16209);
and U18356 (N_18356,N_17941,N_16016);
xor U18357 (N_18357,N_17112,N_17069);
nand U18358 (N_18358,N_17690,N_16286);
nand U18359 (N_18359,N_16139,N_17293);
and U18360 (N_18360,N_16634,N_16631);
or U18361 (N_18361,N_16221,N_16698);
and U18362 (N_18362,N_16968,N_16274);
nor U18363 (N_18363,N_17864,N_16353);
or U18364 (N_18364,N_17349,N_16733);
or U18365 (N_18365,N_17683,N_16148);
nand U18366 (N_18366,N_16125,N_17365);
or U18367 (N_18367,N_17681,N_17528);
nand U18368 (N_18368,N_16181,N_17047);
or U18369 (N_18369,N_16461,N_17447);
or U18370 (N_18370,N_16400,N_17174);
and U18371 (N_18371,N_16527,N_17807);
or U18372 (N_18372,N_17716,N_16844);
nor U18373 (N_18373,N_16034,N_16987);
xnor U18374 (N_18374,N_17746,N_16780);
and U18375 (N_18375,N_16074,N_17727);
and U18376 (N_18376,N_17486,N_16637);
or U18377 (N_18377,N_16325,N_16079);
nor U18378 (N_18378,N_17676,N_16903);
nor U18379 (N_18379,N_16914,N_16979);
xnor U18380 (N_18380,N_17046,N_16680);
and U18381 (N_18381,N_16190,N_16525);
xor U18382 (N_18382,N_17344,N_17303);
nor U18383 (N_18383,N_17659,N_17434);
nand U18384 (N_18384,N_17768,N_16156);
or U18385 (N_18385,N_17404,N_17544);
or U18386 (N_18386,N_17741,N_17154);
xor U18387 (N_18387,N_17965,N_17210);
nor U18388 (N_18388,N_17482,N_17973);
xor U18389 (N_18389,N_16535,N_17858);
or U18390 (N_18390,N_17759,N_16147);
nand U18391 (N_18391,N_17116,N_17038);
xor U18392 (N_18392,N_16092,N_17530);
or U18393 (N_18393,N_17131,N_16234);
nand U18394 (N_18394,N_17113,N_17720);
nand U18395 (N_18395,N_17437,N_16941);
and U18396 (N_18396,N_16982,N_16061);
xor U18397 (N_18397,N_17384,N_16592);
nand U18398 (N_18398,N_17993,N_17616);
and U18399 (N_18399,N_17053,N_17285);
nand U18400 (N_18400,N_17442,N_17529);
nor U18401 (N_18401,N_16152,N_16191);
xnor U18402 (N_18402,N_17721,N_16998);
xor U18403 (N_18403,N_16944,N_17243);
nor U18404 (N_18404,N_16091,N_16422);
nand U18405 (N_18405,N_16093,N_17847);
and U18406 (N_18406,N_17796,N_17369);
and U18407 (N_18407,N_17802,N_16656);
nand U18408 (N_18408,N_17260,N_16494);
nor U18409 (N_18409,N_16745,N_17934);
and U18410 (N_18410,N_17843,N_16486);
or U18411 (N_18411,N_17927,N_16967);
or U18412 (N_18412,N_16141,N_16323);
xor U18413 (N_18413,N_17101,N_16510);
nand U18414 (N_18414,N_16688,N_16151);
or U18415 (N_18415,N_17150,N_16322);
and U18416 (N_18416,N_16599,N_16316);
xnor U18417 (N_18417,N_16006,N_16333);
nand U18418 (N_18418,N_16335,N_17281);
nand U18419 (N_18419,N_17160,N_16013);
and U18420 (N_18420,N_16897,N_16145);
xor U18421 (N_18421,N_17630,N_16149);
xnor U18422 (N_18422,N_17939,N_16477);
nand U18423 (N_18423,N_17579,N_16737);
and U18424 (N_18424,N_17245,N_16140);
nor U18425 (N_18425,N_16816,N_16610);
or U18426 (N_18426,N_16613,N_17928);
xor U18427 (N_18427,N_16794,N_17488);
and U18428 (N_18428,N_16905,N_17618);
nor U18429 (N_18429,N_16705,N_16585);
nand U18430 (N_18430,N_17029,N_17431);
or U18431 (N_18431,N_16179,N_17411);
or U18432 (N_18432,N_17950,N_16722);
xor U18433 (N_18433,N_17317,N_17846);
xor U18434 (N_18434,N_17167,N_17805);
and U18435 (N_18435,N_17515,N_17298);
nor U18436 (N_18436,N_17821,N_16495);
nand U18437 (N_18437,N_17267,N_17645);
xnor U18438 (N_18438,N_16182,N_16348);
or U18439 (N_18439,N_16785,N_16906);
xnor U18440 (N_18440,N_16689,N_17784);
nand U18441 (N_18441,N_17820,N_17446);
xor U18442 (N_18442,N_17607,N_16840);
nor U18443 (N_18443,N_16401,N_16227);
nand U18444 (N_18444,N_17271,N_17405);
or U18445 (N_18445,N_16030,N_17379);
and U18446 (N_18446,N_17068,N_17206);
xor U18447 (N_18447,N_16843,N_17704);
nand U18448 (N_18448,N_16931,N_16100);
or U18449 (N_18449,N_17575,N_16764);
nor U18450 (N_18450,N_17082,N_16817);
nand U18451 (N_18451,N_16254,N_16542);
nand U18452 (N_18452,N_17345,N_17117);
nand U18453 (N_18453,N_16340,N_16259);
and U18454 (N_18454,N_17280,N_16087);
nand U18455 (N_18455,N_17183,N_16506);
and U18456 (N_18456,N_16278,N_17883);
and U18457 (N_18457,N_17680,N_16833);
xnor U18458 (N_18458,N_16969,N_17376);
xor U18459 (N_18459,N_16902,N_17322);
and U18460 (N_18460,N_17103,N_17225);
or U18461 (N_18461,N_17371,N_17910);
nor U18462 (N_18462,N_16266,N_16180);
or U18463 (N_18463,N_16726,N_16037);
and U18464 (N_18464,N_16528,N_16723);
nand U18465 (N_18465,N_16466,N_17034);
and U18466 (N_18466,N_16556,N_17277);
nand U18467 (N_18467,N_16306,N_17987);
and U18468 (N_18468,N_17476,N_17351);
nor U18469 (N_18469,N_16293,N_17702);
or U18470 (N_18470,N_16430,N_17614);
xor U18471 (N_18471,N_17677,N_17234);
and U18472 (N_18472,N_16014,N_17478);
xnor U18473 (N_18473,N_17257,N_17455);
nor U18474 (N_18474,N_17471,N_16199);
and U18475 (N_18475,N_17199,N_17581);
and U18476 (N_18476,N_17262,N_17900);
nor U18477 (N_18477,N_17090,N_17760);
or U18478 (N_18478,N_16153,N_17754);
nand U18479 (N_18479,N_17650,N_17209);
or U18480 (N_18480,N_17081,N_16420);
nor U18481 (N_18481,N_17200,N_17306);
nor U18482 (N_18482,N_16075,N_16407);
and U18483 (N_18483,N_16801,N_16802);
nand U18484 (N_18484,N_17644,N_17897);
nand U18485 (N_18485,N_17620,N_17129);
or U18486 (N_18486,N_17202,N_16788);
nor U18487 (N_18487,N_17159,N_17342);
xor U18488 (N_18488,N_16334,N_17226);
or U18489 (N_18489,N_16009,N_17048);
nor U18490 (N_18490,N_17118,N_17461);
nand U18491 (N_18491,N_17076,N_17894);
or U18492 (N_18492,N_16097,N_17250);
xor U18493 (N_18493,N_16408,N_17052);
and U18494 (N_18494,N_16579,N_17595);
nor U18495 (N_18495,N_17901,N_16635);
and U18496 (N_18496,N_16172,N_16753);
or U18497 (N_18497,N_16500,N_16999);
nor U18498 (N_18498,N_17918,N_17823);
and U18499 (N_18499,N_16811,N_17073);
and U18500 (N_18500,N_16508,N_16908);
or U18501 (N_18501,N_17757,N_17494);
and U18502 (N_18502,N_16548,N_17589);
xor U18503 (N_18503,N_17215,N_17990);
nor U18504 (N_18504,N_17241,N_17191);
xor U18505 (N_18505,N_16871,N_16370);
nand U18506 (N_18506,N_16352,N_16314);
and U18507 (N_18507,N_16621,N_17148);
and U18508 (N_18508,N_16793,N_17535);
nand U18509 (N_18509,N_17158,N_17231);
and U18510 (N_18510,N_16228,N_16384);
and U18511 (N_18511,N_17641,N_17134);
or U18512 (N_18512,N_17930,N_17882);
or U18513 (N_18513,N_17656,N_17286);
xor U18514 (N_18514,N_16119,N_16497);
xnor U18515 (N_18515,N_16398,N_16448);
nand U18516 (N_18516,N_17088,N_16996);
and U18517 (N_18517,N_16976,N_17135);
nor U18518 (N_18518,N_17833,N_16822);
and U18519 (N_18519,N_16200,N_17783);
nand U18520 (N_18520,N_17310,N_17647);
xnor U18521 (N_18521,N_16746,N_16861);
or U18522 (N_18522,N_17755,N_16703);
nand U18523 (N_18523,N_17060,N_16664);
and U18524 (N_18524,N_17031,N_17507);
nor U18525 (N_18525,N_16102,N_16992);
xnor U18526 (N_18526,N_17377,N_16038);
nor U18527 (N_18527,N_16699,N_16845);
xnor U18528 (N_18528,N_16117,N_17339);
and U18529 (N_18529,N_17697,N_16445);
nand U18530 (N_18530,N_16640,N_17320);
nor U18531 (N_18531,N_17490,N_16701);
and U18532 (N_18532,N_17992,N_16320);
or U18533 (N_18533,N_17265,N_16502);
xnor U18534 (N_18534,N_17985,N_17809);
and U18535 (N_18535,N_16423,N_16257);
and U18536 (N_18536,N_16245,N_16769);
or U18537 (N_18537,N_17075,N_16110);
and U18538 (N_18538,N_16938,N_17164);
xor U18539 (N_18539,N_17588,N_16538);
nor U18540 (N_18540,N_17067,N_17880);
or U18541 (N_18541,N_17410,N_17089);
or U18542 (N_18542,N_16243,N_17705);
and U18543 (N_18543,N_16319,N_17290);
or U18544 (N_18544,N_17179,N_16364);
nor U18545 (N_18545,N_16387,N_17532);
or U18546 (N_18546,N_16573,N_17998);
xor U18547 (N_18547,N_16882,N_16781);
nor U18548 (N_18548,N_17812,N_16481);
xor U18549 (N_18549,N_17855,N_17204);
or U18550 (N_18550,N_16290,N_16336);
or U18551 (N_18551,N_17566,N_16032);
or U18552 (N_18552,N_17657,N_17660);
or U18553 (N_18553,N_16035,N_16929);
or U18554 (N_18554,N_17899,N_16561);
nand U18555 (N_18555,N_16899,N_16517);
nand U18556 (N_18556,N_17033,N_16361);
xor U18557 (N_18557,N_16175,N_17738);
or U18558 (N_18558,N_16017,N_17300);
nand U18559 (N_18559,N_17363,N_16212);
and U18560 (N_18560,N_17634,N_17295);
or U18561 (N_18561,N_16261,N_17428);
and U18562 (N_18562,N_17196,N_16311);
and U18563 (N_18563,N_16872,N_16544);
xor U18564 (N_18564,N_17642,N_16427);
and U18565 (N_18565,N_17775,N_16576);
xnor U18566 (N_18566,N_17166,N_17251);
xnor U18567 (N_18567,N_17334,N_16618);
and U18568 (N_18568,N_16975,N_17673);
and U18569 (N_18569,N_17771,N_16084);
nor U18570 (N_18570,N_16965,N_16346);
or U18571 (N_18571,N_17095,N_17924);
and U18572 (N_18572,N_17968,N_17516);
nor U18573 (N_18573,N_16351,N_17273);
xnor U18574 (N_18574,N_16868,N_17423);
and U18575 (N_18575,N_16244,N_16391);
nor U18576 (N_18576,N_16282,N_17736);
xnor U18577 (N_18577,N_17145,N_16342);
and U18578 (N_18578,N_17235,N_17734);
and U18579 (N_18579,N_17794,N_17570);
nor U18580 (N_18580,N_17380,N_16825);
nand U18581 (N_18581,N_16923,N_17867);
or U18582 (N_18582,N_17331,N_17671);
nand U18583 (N_18583,N_17422,N_16302);
nor U18584 (N_18584,N_16344,N_16814);
or U18585 (N_18585,N_16059,N_17944);
nand U18586 (N_18586,N_16473,N_16020);
or U18587 (N_18587,N_17629,N_17626);
and U18588 (N_18588,N_17395,N_17813);
xor U18589 (N_18589,N_16214,N_16605);
or U18590 (N_18590,N_17071,N_17606);
xor U18591 (N_18591,N_17636,N_17092);
or U18592 (N_18592,N_16327,N_16947);
or U18593 (N_18593,N_16717,N_16819);
or U18594 (N_18594,N_16249,N_17335);
xnor U18595 (N_18595,N_17028,N_17826);
or U18596 (N_18596,N_16308,N_17518);
nand U18597 (N_18597,N_16337,N_17337);
or U18598 (N_18598,N_16950,N_17982);
nor U18599 (N_18599,N_16375,N_17960);
and U18600 (N_18600,N_17137,N_16405);
nor U18601 (N_18601,N_16614,N_16273);
or U18602 (N_18602,N_16324,N_17613);
xnor U18603 (N_18603,N_16571,N_16584);
xnor U18604 (N_18604,N_17859,N_17798);
and U18605 (N_18605,N_17246,N_16491);
or U18606 (N_18606,N_17024,N_16973);
or U18607 (N_18607,N_17451,N_17107);
nand U18608 (N_18608,N_16690,N_17378);
nand U18609 (N_18609,N_17788,N_17429);
nor U18610 (N_18610,N_17501,N_17087);
xnor U18611 (N_18611,N_17832,N_17583);
or U18612 (N_18612,N_17040,N_16877);
nor U18613 (N_18613,N_17815,N_17773);
and U18614 (N_18614,N_16123,N_17945);
nor U18615 (N_18615,N_16406,N_16256);
xnor U18616 (N_18616,N_16127,N_16957);
or U18617 (N_18617,N_17356,N_17055);
nand U18618 (N_18618,N_17333,N_17070);
nand U18619 (N_18619,N_17599,N_16083);
nand U18620 (N_18620,N_16763,N_17208);
or U18621 (N_18621,N_16208,N_17979);
nor U18622 (N_18622,N_16778,N_17421);
or U18623 (N_18623,N_17230,N_17313);
or U18624 (N_18624,N_17402,N_17420);
nand U18625 (N_18625,N_16608,N_17512);
xor U18626 (N_18626,N_17707,N_17106);
nand U18627 (N_18627,N_16632,N_17995);
nand U18628 (N_18628,N_16168,N_16265);
and U18629 (N_18629,N_17464,N_17905);
nand U18630 (N_18630,N_16425,N_16457);
and U18631 (N_18631,N_17027,N_16187);
or U18632 (N_18632,N_17785,N_16409);
xnor U18633 (N_18633,N_16859,N_17359);
nand U18634 (N_18634,N_16909,N_17133);
nor U18635 (N_18635,N_16289,N_16332);
or U18636 (N_18636,N_16411,N_16105);
xnor U18637 (N_18637,N_17537,N_17670);
or U18638 (N_18638,N_17348,N_17484);
and U18639 (N_18639,N_17032,N_16810);
or U18640 (N_18640,N_16465,N_17949);
xnor U18641 (N_18641,N_16033,N_16721);
nand U18642 (N_18642,N_17724,N_16041);
nand U18643 (N_18643,N_17043,N_17198);
nand U18644 (N_18644,N_17424,N_17919);
and U18645 (N_18645,N_16665,N_17590);
and U18646 (N_18646,N_16709,N_17853);
and U18647 (N_18647,N_17640,N_16891);
nand U18648 (N_18648,N_17552,N_16028);
or U18649 (N_18649,N_16994,N_17220);
or U18650 (N_18650,N_16932,N_16715);
or U18651 (N_18651,N_17485,N_17539);
nor U18652 (N_18652,N_17597,N_16164);
xnor U18653 (N_18653,N_16053,N_17044);
xnor U18654 (N_18654,N_17770,N_17617);
nand U18655 (N_18655,N_16051,N_17898);
nand U18656 (N_18656,N_17074,N_17098);
and U18657 (N_18657,N_16443,N_17362);
nand U18658 (N_18658,N_17997,N_16615);
or U18659 (N_18659,N_16485,N_17686);
nor U18660 (N_18660,N_16729,N_16886);
xnor U18661 (N_18661,N_17638,N_17750);
or U18662 (N_18662,N_17691,N_17289);
or U18663 (N_18663,N_16318,N_16085);
nand U18664 (N_18664,N_16270,N_16018);
or U18665 (N_18665,N_17850,N_17457);
or U18666 (N_18666,N_17886,N_17609);
nor U18667 (N_18667,N_16328,N_17407);
nand U18668 (N_18668,N_16458,N_17536);
or U18669 (N_18669,N_16673,N_16772);
nand U18670 (N_18670,N_17972,N_16730);
nand U18671 (N_18671,N_16402,N_16743);
or U18672 (N_18672,N_16515,N_17401);
or U18673 (N_18673,N_16971,N_17466);
or U18674 (N_18674,N_17221,N_16839);
and U18675 (N_18675,N_16706,N_16593);
nor U18676 (N_18676,N_16727,N_17161);
or U18677 (N_18677,N_17651,N_17695);
nor U18678 (N_18678,N_16201,N_16587);
and U18679 (N_18679,N_17329,N_16386);
nor U18680 (N_18680,N_17057,N_16852);
or U18681 (N_18681,N_16804,N_17099);
or U18682 (N_18682,N_16291,N_17747);
nor U18683 (N_18683,N_16474,N_17481);
xor U18684 (N_18684,N_17730,N_16241);
nor U18685 (N_18685,N_17931,N_16027);
or U18686 (N_18686,N_17914,N_16582);
nand U18687 (N_18687,N_16856,N_17974);
xor U18688 (N_18688,N_16029,N_16142);
and U18689 (N_18689,N_16553,N_16662);
xor U18690 (N_18690,N_16218,N_16855);
and U18691 (N_18691,N_16089,N_17123);
nand U18692 (N_18692,N_17932,N_17096);
nand U18693 (N_18693,N_17392,N_17338);
or U18694 (N_18694,N_16624,N_17136);
xor U18695 (N_18695,N_17296,N_16367);
nand U18696 (N_18696,N_17777,N_16874);
xor U18697 (N_18697,N_16893,N_17375);
nand U18698 (N_18698,N_16354,N_16835);
or U18699 (N_18699,N_17574,N_16850);
or U18700 (N_18700,N_17884,N_16050);
nor U18701 (N_18701,N_17018,N_16372);
nand U18702 (N_18702,N_17569,N_17592);
and U18703 (N_18703,N_17294,N_17497);
nand U18704 (N_18704,N_16734,N_16444);
nand U18705 (N_18705,N_16429,N_16981);
nor U18706 (N_18706,N_17653,N_16441);
nand U18707 (N_18707,N_17523,N_17400);
nor U18708 (N_18708,N_16820,N_17688);
xnor U18709 (N_18709,N_17753,N_16338);
and U18710 (N_18710,N_17435,N_17876);
and U18711 (N_18711,N_16921,N_16925);
nand U18712 (N_18712,N_17860,N_16363);
and U18713 (N_18713,N_16765,N_17439);
and U18714 (N_18714,N_17852,N_17857);
nand U18715 (N_18715,N_17237,N_17975);
nand U18716 (N_18716,N_17223,N_16251);
nor U18717 (N_18717,N_16776,N_17100);
xnor U18718 (N_18718,N_17080,N_16978);
xnor U18719 (N_18719,N_17184,N_17360);
nand U18720 (N_18720,N_16708,N_17668);
and U18721 (N_18721,N_16911,N_16447);
and U18722 (N_18722,N_17287,N_17328);
or U18723 (N_18723,N_16417,N_17854);
and U18724 (N_18724,N_17661,N_17513);
and U18725 (N_18725,N_16653,N_17504);
and U18726 (N_18726,N_17330,N_16948);
xnor U18727 (N_18727,N_17479,N_16060);
and U18728 (N_18728,N_17922,N_16747);
nand U18729 (N_18729,N_17463,N_16539);
xnor U18730 (N_18730,N_17086,N_17567);
or U18731 (N_18731,N_16783,N_17282);
xnor U18732 (N_18732,N_16345,N_16439);
xor U18733 (N_18733,N_17072,N_16193);
or U18734 (N_18734,N_17554,N_17540);
xor U18735 (N_18735,N_17627,N_17977);
and U18736 (N_18736,N_17937,N_17586);
or U18737 (N_18737,N_17413,N_17037);
nor U18738 (N_18738,N_17885,N_17212);
or U18739 (N_18739,N_16296,N_16863);
nand U18740 (N_18740,N_16483,N_16122);
xor U18741 (N_18741,N_17398,N_16752);
xor U18742 (N_18742,N_16895,N_17861);
xor U18743 (N_18743,N_16350,N_17505);
nand U18744 (N_18744,N_16719,N_17005);
or U18745 (N_18745,N_16892,N_17712);
xor U18746 (N_18746,N_17527,N_16901);
xnor U18747 (N_18747,N_17194,N_16639);
and U18748 (N_18748,N_17079,N_17025);
and U18749 (N_18749,N_17839,N_17412);
nor U18750 (N_18750,N_17357,N_16570);
and U18751 (N_18751,N_16720,N_17723);
and U18752 (N_18752,N_17628,N_16924);
nand U18753 (N_18753,N_17140,N_17522);
nor U18754 (N_18754,N_16044,N_16646);
or U18755 (N_18755,N_16285,N_17782);
or U18756 (N_18756,N_16382,N_17228);
nor U18757 (N_18757,N_17178,N_16766);
or U18758 (N_18758,N_17509,N_17602);
and U18759 (N_18759,N_17830,N_17051);
nor U18760 (N_18760,N_17382,N_17297);
and U18761 (N_18761,N_16225,N_17543);
and U18762 (N_18762,N_17572,N_16380);
and U18763 (N_18763,N_17058,N_17881);
nor U18764 (N_18764,N_17909,N_16167);
xor U18765 (N_18765,N_17197,N_17268);
nor U18766 (N_18766,N_17703,N_16489);
and U18767 (N_18767,N_16602,N_16378);
nand U18768 (N_18768,N_17520,N_16679);
or U18769 (N_18769,N_17399,N_17903);
nand U18770 (N_18770,N_17352,N_16758);
nand U18771 (N_18771,N_17598,N_16001);
nor U18772 (N_18772,N_16565,N_17441);
nand U18773 (N_18773,N_17728,N_16997);
xor U18774 (N_18774,N_17175,N_17541);
and U18775 (N_18775,N_17370,N_16008);
nand U18776 (N_18776,N_16462,N_17917);
nor U18777 (N_18777,N_17573,N_16567);
and U18778 (N_18778,N_16597,N_17326);
nor U18779 (N_18779,N_17925,N_16655);
nor U18780 (N_18780,N_17948,N_16821);
nor U18781 (N_18781,N_16390,N_16300);
xor U18782 (N_18782,N_16326,N_16188);
nand U18783 (N_18783,N_17582,N_16064);
and U18784 (N_18784,N_16433,N_16547);
nor U18785 (N_18785,N_16942,N_17105);
or U18786 (N_18786,N_17729,N_17816);
or U18787 (N_18787,N_17907,N_16280);
and U18788 (N_18788,N_16299,N_17779);
xor U18789 (N_18789,N_16499,N_17042);
nand U18790 (N_18790,N_17538,N_16236);
and U18791 (N_18791,N_16000,N_17733);
nand U18792 (N_18792,N_17921,N_16011);
nand U18793 (N_18793,N_16487,N_17364);
or U18794 (N_18794,N_17935,N_17631);
nand U18795 (N_18795,N_17562,N_16467);
nor U18796 (N_18796,N_16807,N_17844);
nand U18797 (N_18797,N_17213,N_17808);
xnor U18798 (N_18798,N_16626,N_16230);
and U18799 (N_18799,N_17272,N_16220);
xor U18800 (N_18800,N_16603,N_16165);
and U18801 (N_18801,N_17508,N_16137);
and U18802 (N_18802,N_17698,N_17009);
xnor U18803 (N_18803,N_16898,N_16410);
xnor U18804 (N_18804,N_17871,N_16113);
and U18805 (N_18805,N_17980,N_16770);
and U18806 (N_18806,N_16434,N_16315);
nand U18807 (N_18807,N_16049,N_16284);
or U18808 (N_18808,N_16048,N_17799);
or U18809 (N_18809,N_16912,N_16403);
nand U18810 (N_18810,N_16077,N_17153);
xor U18811 (N_18811,N_16562,N_17084);
xor U18812 (N_18812,N_16983,N_16865);
and U18813 (N_18813,N_17848,N_16279);
or U18814 (N_18814,N_16080,N_17021);
and U18815 (N_18815,N_16927,N_16088);
nor U18816 (N_18816,N_17010,N_16307);
and U18817 (N_18817,N_16347,N_16831);
xnor U18818 (N_18818,N_16554,N_16126);
nand U18819 (N_18819,N_17239,N_16823);
nand U18820 (N_18820,N_17056,N_17367);
nand U18821 (N_18821,N_16509,N_16002);
nand U18822 (N_18822,N_16255,N_17227);
or U18823 (N_18823,N_16478,N_16451);
or U18824 (N_18824,N_17719,N_16946);
xor U18825 (N_18825,N_16988,N_16609);
or U18826 (N_18826,N_16082,N_17083);
nor U18827 (N_18827,N_16963,N_17323);
or U18828 (N_18828,N_16832,N_17146);
nor U18829 (N_18829,N_16468,N_16341);
nand U18830 (N_18830,N_16252,N_17109);
or U18831 (N_18831,N_17078,N_17761);
nand U18832 (N_18832,N_17332,N_17904);
xnor U18833 (N_18833,N_16511,N_17122);
nand U18834 (N_18834,N_16896,N_17865);
and U18835 (N_18835,N_17906,N_16873);
nor U18836 (N_18836,N_16379,N_17749);
nor U18837 (N_18837,N_16713,N_17604);
or U18838 (N_18838,N_17708,N_16630);
and U18839 (N_18839,N_17232,N_17926);
nor U18840 (N_18840,N_16827,N_16977);
and U18841 (N_18841,N_17684,N_17811);
nand U18842 (N_18842,N_16677,N_16750);
or U18843 (N_18843,N_17186,N_17787);
xnor U18844 (N_18844,N_16589,N_17430);
and U18845 (N_18845,N_16575,N_17386);
nand U18846 (N_18846,N_17565,N_17621);
nand U18847 (N_18847,N_17094,N_17810);
and U18848 (N_18848,N_17664,N_16381);
nor U18849 (N_18849,N_17869,N_17715);
xnor U18850 (N_18850,N_17596,N_17521);
xor U18851 (N_18851,N_16128,N_16629);
nor U18852 (N_18852,N_17358,N_17600);
and U18853 (N_18853,N_16716,N_16735);
nor U18854 (N_18854,N_16362,N_17637);
xor U18855 (N_18855,N_17834,N_16756);
or U18856 (N_18856,N_17017,N_16185);
nand U18857 (N_18857,N_17460,N_17743);
nor U18858 (N_18858,N_17890,N_16846);
nand U18859 (N_18859,N_17487,N_16170);
nand U18860 (N_18860,N_16090,N_16503);
or U18861 (N_18861,N_16601,N_17986);
or U18862 (N_18862,N_17102,N_16672);
or U18863 (N_18863,N_16782,N_17383);
xor U18864 (N_18864,N_17353,N_17524);
nand U18865 (N_18865,N_17601,N_16697);
xnor U18866 (N_18866,N_17492,N_17969);
and U18867 (N_18867,N_17493,N_17851);
and U18868 (N_18868,N_17354,N_16186);
or U18869 (N_18869,N_17222,N_17622);
nor U18870 (N_18870,N_16847,N_17489);
nor U18871 (N_18871,N_17517,N_16958);
xor U18872 (N_18872,N_17219,N_16879);
and U18873 (N_18873,N_17006,N_16267);
nand U18874 (N_18874,N_17994,N_16633);
xor U18875 (N_18875,N_16989,N_17989);
and U18876 (N_18876,N_17877,N_17039);
nor U18877 (N_18877,N_17725,N_16862);
or U18878 (N_18878,N_16910,N_16808);
and U18879 (N_18879,N_17124,N_17954);
nand U18880 (N_18880,N_16834,N_16666);
nand U18881 (N_18881,N_17639,N_16412);
and U18882 (N_18882,N_16471,N_17440);
or U18883 (N_18883,N_16507,N_16277);
and U18884 (N_18884,N_17218,N_16131);
nand U18885 (N_18885,N_16980,N_17450);
nand U18886 (N_18886,N_16171,N_17238);
nor U18887 (N_18887,N_17418,N_17483);
nor U18888 (N_18888,N_16368,N_17817);
or U18889 (N_18889,N_17432,N_16536);
and U18890 (N_18890,N_16732,N_17311);
and U18891 (N_18891,N_17556,N_16643);
xnor U18892 (N_18892,N_17270,N_16446);
or U18893 (N_18893,N_16226,N_17553);
nand U18894 (N_18894,N_16219,N_16870);
or U18895 (N_18895,N_16563,N_17406);
and U18896 (N_18896,N_16358,N_17999);
xnor U18897 (N_18897,N_16040,N_17963);
xor U18898 (N_18898,N_17766,N_17737);
nor U18899 (N_18899,N_16818,N_17436);
nand U18900 (N_18900,N_16281,N_17340);
nand U18901 (N_18901,N_16707,N_17015);
nor U18902 (N_18902,N_17120,N_17780);
xnor U18903 (N_18903,N_17007,N_17470);
xor U18904 (N_18904,N_17946,N_16154);
xor U18905 (N_18905,N_17559,N_17557);
and U18906 (N_18906,N_16964,N_17128);
nand U18907 (N_18907,N_16889,N_17722);
xor U18908 (N_18908,N_17000,N_16854);
or U18909 (N_18909,N_16907,N_16052);
or U18910 (N_18910,N_16564,N_16529);
nor U18911 (N_18911,N_16740,N_17624);
and U18912 (N_18912,N_17542,N_16120);
xor U18913 (N_18913,N_17433,N_17240);
xor U18914 (N_18914,N_16552,N_16135);
and U18915 (N_18915,N_16768,N_17814);
nor U18916 (N_18916,N_16797,N_16184);
or U18917 (N_18917,N_17632,N_17888);
and U18918 (N_18918,N_16962,N_16343);
xnor U18919 (N_18919,N_17893,N_17732);
and U18920 (N_18920,N_16215,N_16428);
nand U18921 (N_18921,N_16248,N_17012);
xnor U18922 (N_18922,N_16146,N_17132);
nor U18923 (N_18923,N_17769,N_17499);
or U18924 (N_18924,N_17506,N_17667);
xnor U18925 (N_18925,N_17390,N_16961);
nor U18926 (N_18926,N_16678,N_16805);
nor U18927 (N_18927,N_16493,N_17318);
or U18928 (N_18928,N_16223,N_17558);
xnor U18929 (N_18929,N_17085,N_17214);
nand U18930 (N_18930,N_17168,N_17988);
xnor U18931 (N_18931,N_16675,N_17283);
nand U18932 (N_18932,N_17970,N_17693);
nand U18933 (N_18933,N_16132,N_17655);
and U18934 (N_18934,N_16258,N_16070);
nor U18935 (N_18935,N_16155,N_17953);
nand U18936 (N_18936,N_17162,N_17603);
nor U18937 (N_18937,N_16777,N_16645);
nor U18938 (N_18938,N_16692,N_16271);
and U18939 (N_18939,N_16683,N_17560);
nand U18940 (N_18940,N_16094,N_16795);
xnor U18941 (N_18941,N_16260,N_16056);
and U18942 (N_18942,N_17577,N_17700);
nor U18943 (N_18943,N_17193,N_17735);
nand U18944 (N_18944,N_16787,N_17254);
nand U18945 (N_18945,N_16404,N_17866);
and U18946 (N_18946,N_17495,N_17545);
or U18947 (N_18947,N_17978,N_16826);
and U18948 (N_18948,N_17121,N_17840);
or U18949 (N_18949,N_16058,N_16216);
nand U18950 (N_18950,N_17448,N_16432);
xnor U18951 (N_18951,N_17612,N_16366);
nand U18952 (N_18952,N_16395,N_16356);
nand U18953 (N_18953,N_16301,N_17316);
nand U18954 (N_18954,N_16157,N_17500);
or U18955 (N_18955,N_16949,N_17758);
and U18956 (N_18956,N_16704,N_17263);
nand U18957 (N_18957,N_16824,N_16516);
xor U18958 (N_18958,N_16217,N_17373);
and U18959 (N_18959,N_17845,N_16623);
xnor U18960 (N_18960,N_17324,N_16460);
nor U18961 (N_18961,N_16371,N_16496);
xnor U18962 (N_18962,N_17252,N_16569);
and U18963 (N_18963,N_17393,N_17341);
nor U18964 (N_18964,N_16321,N_17772);
nand U18965 (N_18965,N_17801,N_17445);
and U18966 (N_18966,N_16313,N_16954);
nor U18967 (N_18967,N_17391,N_16396);
nand U18968 (N_18968,N_17699,N_17368);
nor U18969 (N_18969,N_17480,N_17635);
xnor U18970 (N_18970,N_16594,N_16762);
or U18971 (N_18971,N_16022,N_17022);
nor U18972 (N_18972,N_17264,N_16360);
nor U18973 (N_18973,N_16598,N_17578);
nand U18974 (N_18974,N_17253,N_16169);
and U18975 (N_18975,N_16174,N_16197);
or U18976 (N_18976,N_17248,N_17800);
or U18977 (N_18977,N_16543,N_16812);
nand U18978 (N_18978,N_16813,N_17879);
or U18979 (N_18979,N_17002,N_17873);
xor U18980 (N_18980,N_16067,N_16005);
nor U18981 (N_18981,N_16440,N_16246);
and U18982 (N_18982,N_17152,N_16115);
nor U18983 (N_18983,N_16068,N_17838);
and U18984 (N_18984,N_16744,N_16714);
xor U18985 (N_18985,N_16210,N_16415);
or U18986 (N_18986,N_16176,N_17806);
nor U18987 (N_18987,N_17188,N_16133);
nor U18988 (N_18988,N_16069,N_17587);
nand U18989 (N_18989,N_16606,N_16800);
xnor U18990 (N_18990,N_17665,N_16774);
nor U18991 (N_18991,N_16189,N_17381);
xor U18992 (N_18992,N_16526,N_17519);
xnor U18993 (N_18993,N_16622,N_16071);
and U18994 (N_18994,N_17108,N_17849);
and U18995 (N_18995,N_16295,N_16628);
nor U18996 (N_18996,N_17662,N_16031);
xor U18997 (N_18997,N_16880,N_16691);
xor U18998 (N_18998,N_16991,N_16595);
xnor U18999 (N_18999,N_17938,N_16480);
or U19000 (N_19000,N_16595,N_16558);
nand U19001 (N_19001,N_17844,N_16138);
nand U19002 (N_19002,N_17920,N_17494);
or U19003 (N_19003,N_17256,N_17824);
nor U19004 (N_19004,N_17712,N_17142);
nand U19005 (N_19005,N_17703,N_16870);
nor U19006 (N_19006,N_17063,N_17823);
and U19007 (N_19007,N_17764,N_17272);
nor U19008 (N_19008,N_16689,N_17465);
nand U19009 (N_19009,N_17685,N_17967);
or U19010 (N_19010,N_16720,N_16523);
and U19011 (N_19011,N_16071,N_16328);
nor U19012 (N_19012,N_16706,N_16063);
nor U19013 (N_19013,N_17109,N_17466);
or U19014 (N_19014,N_17227,N_17664);
nor U19015 (N_19015,N_17006,N_17117);
or U19016 (N_19016,N_16677,N_16626);
and U19017 (N_19017,N_16085,N_17990);
xnor U19018 (N_19018,N_16610,N_16620);
nor U19019 (N_19019,N_16831,N_17041);
or U19020 (N_19020,N_16642,N_17517);
nand U19021 (N_19021,N_17070,N_16609);
xor U19022 (N_19022,N_16695,N_16203);
or U19023 (N_19023,N_17014,N_16841);
and U19024 (N_19024,N_17184,N_16617);
and U19025 (N_19025,N_17759,N_16979);
nor U19026 (N_19026,N_17626,N_17931);
xor U19027 (N_19027,N_16444,N_16636);
nor U19028 (N_19028,N_16267,N_17078);
xor U19029 (N_19029,N_17754,N_17905);
xor U19030 (N_19030,N_17094,N_16201);
nand U19031 (N_19031,N_17280,N_16820);
or U19032 (N_19032,N_17651,N_16016);
nor U19033 (N_19033,N_17751,N_16950);
xor U19034 (N_19034,N_17098,N_17173);
or U19035 (N_19035,N_17221,N_16319);
or U19036 (N_19036,N_16903,N_17918);
or U19037 (N_19037,N_16384,N_17317);
and U19038 (N_19038,N_16845,N_16288);
xor U19039 (N_19039,N_16292,N_17708);
or U19040 (N_19040,N_17548,N_16471);
and U19041 (N_19041,N_17815,N_17086);
xnor U19042 (N_19042,N_17877,N_17646);
and U19043 (N_19043,N_17533,N_17486);
nor U19044 (N_19044,N_17528,N_16394);
and U19045 (N_19045,N_17207,N_17248);
or U19046 (N_19046,N_16180,N_17282);
or U19047 (N_19047,N_16567,N_17200);
nor U19048 (N_19048,N_17233,N_17698);
and U19049 (N_19049,N_17965,N_16501);
nor U19050 (N_19050,N_16319,N_17693);
nand U19051 (N_19051,N_17730,N_17722);
nor U19052 (N_19052,N_16360,N_17069);
and U19053 (N_19053,N_16339,N_17073);
nor U19054 (N_19054,N_16470,N_16636);
and U19055 (N_19055,N_17054,N_17776);
nor U19056 (N_19056,N_17390,N_16952);
nor U19057 (N_19057,N_17552,N_16233);
and U19058 (N_19058,N_16735,N_16783);
nor U19059 (N_19059,N_16412,N_16871);
or U19060 (N_19060,N_16628,N_16468);
nand U19061 (N_19061,N_16459,N_17730);
nand U19062 (N_19062,N_17388,N_16235);
and U19063 (N_19063,N_16585,N_16522);
and U19064 (N_19064,N_16445,N_17060);
nor U19065 (N_19065,N_17241,N_17154);
nor U19066 (N_19066,N_16623,N_17611);
nand U19067 (N_19067,N_17902,N_17733);
nor U19068 (N_19068,N_16557,N_16675);
xnor U19069 (N_19069,N_17234,N_16669);
nor U19070 (N_19070,N_16530,N_17466);
or U19071 (N_19071,N_16787,N_16138);
nand U19072 (N_19072,N_16935,N_17904);
or U19073 (N_19073,N_16002,N_17786);
xnor U19074 (N_19074,N_16972,N_17740);
xnor U19075 (N_19075,N_17078,N_16177);
xor U19076 (N_19076,N_16400,N_17403);
xor U19077 (N_19077,N_16429,N_17364);
and U19078 (N_19078,N_17970,N_16818);
nor U19079 (N_19079,N_17474,N_16707);
and U19080 (N_19080,N_17932,N_17787);
nor U19081 (N_19081,N_17405,N_17509);
nand U19082 (N_19082,N_16881,N_17931);
or U19083 (N_19083,N_17969,N_17246);
or U19084 (N_19084,N_16761,N_17798);
or U19085 (N_19085,N_16619,N_17314);
nand U19086 (N_19086,N_17272,N_17707);
and U19087 (N_19087,N_16864,N_16141);
or U19088 (N_19088,N_17159,N_17537);
and U19089 (N_19089,N_17703,N_17565);
xnor U19090 (N_19090,N_16411,N_17181);
and U19091 (N_19091,N_17050,N_16824);
nand U19092 (N_19092,N_16046,N_17158);
nor U19093 (N_19093,N_17755,N_17057);
nor U19094 (N_19094,N_17245,N_16972);
nand U19095 (N_19095,N_17148,N_16250);
nand U19096 (N_19096,N_16823,N_17541);
xnor U19097 (N_19097,N_16403,N_17914);
nor U19098 (N_19098,N_16890,N_16531);
nor U19099 (N_19099,N_16863,N_17239);
nor U19100 (N_19100,N_16007,N_17743);
and U19101 (N_19101,N_17890,N_16218);
nor U19102 (N_19102,N_16481,N_16129);
nand U19103 (N_19103,N_16849,N_16288);
or U19104 (N_19104,N_17116,N_17051);
nor U19105 (N_19105,N_16956,N_17579);
nand U19106 (N_19106,N_17487,N_17947);
and U19107 (N_19107,N_17589,N_16073);
and U19108 (N_19108,N_17323,N_16467);
nor U19109 (N_19109,N_16099,N_16296);
nand U19110 (N_19110,N_17764,N_17836);
nor U19111 (N_19111,N_16652,N_17049);
xnor U19112 (N_19112,N_17337,N_17743);
or U19113 (N_19113,N_17363,N_17055);
nor U19114 (N_19114,N_17774,N_16268);
nor U19115 (N_19115,N_16671,N_16387);
nand U19116 (N_19116,N_16342,N_16473);
nand U19117 (N_19117,N_16629,N_16739);
or U19118 (N_19118,N_17940,N_17047);
or U19119 (N_19119,N_17029,N_17445);
or U19120 (N_19120,N_16308,N_16480);
and U19121 (N_19121,N_16214,N_16626);
nor U19122 (N_19122,N_17091,N_17301);
and U19123 (N_19123,N_17679,N_16944);
xor U19124 (N_19124,N_16342,N_16535);
and U19125 (N_19125,N_16790,N_16812);
nor U19126 (N_19126,N_17563,N_16101);
nand U19127 (N_19127,N_16635,N_16705);
nand U19128 (N_19128,N_16319,N_16143);
and U19129 (N_19129,N_16480,N_17607);
nand U19130 (N_19130,N_17107,N_17528);
nor U19131 (N_19131,N_17622,N_16009);
and U19132 (N_19132,N_17967,N_17341);
or U19133 (N_19133,N_16157,N_17616);
and U19134 (N_19134,N_17976,N_17519);
and U19135 (N_19135,N_16309,N_16362);
xnor U19136 (N_19136,N_17912,N_17455);
or U19137 (N_19137,N_16384,N_16427);
or U19138 (N_19138,N_16791,N_16732);
nand U19139 (N_19139,N_16029,N_17661);
nor U19140 (N_19140,N_17793,N_16333);
or U19141 (N_19141,N_17834,N_16270);
or U19142 (N_19142,N_17930,N_16748);
nor U19143 (N_19143,N_17054,N_16533);
or U19144 (N_19144,N_17094,N_17635);
xor U19145 (N_19145,N_17324,N_16237);
nand U19146 (N_19146,N_16350,N_17740);
and U19147 (N_19147,N_16332,N_17652);
xor U19148 (N_19148,N_17986,N_17310);
nor U19149 (N_19149,N_17965,N_17094);
nand U19150 (N_19150,N_16826,N_16977);
and U19151 (N_19151,N_16000,N_17716);
or U19152 (N_19152,N_17387,N_16418);
and U19153 (N_19153,N_16891,N_17293);
nand U19154 (N_19154,N_16870,N_16340);
nor U19155 (N_19155,N_17319,N_17904);
or U19156 (N_19156,N_17836,N_16957);
and U19157 (N_19157,N_17561,N_16592);
and U19158 (N_19158,N_16196,N_17615);
xor U19159 (N_19159,N_16144,N_16568);
and U19160 (N_19160,N_16202,N_16428);
nand U19161 (N_19161,N_16040,N_16624);
and U19162 (N_19162,N_17663,N_16671);
xor U19163 (N_19163,N_17749,N_17773);
and U19164 (N_19164,N_17895,N_17665);
nand U19165 (N_19165,N_16137,N_16487);
nor U19166 (N_19166,N_17454,N_17987);
nor U19167 (N_19167,N_17757,N_16788);
nand U19168 (N_19168,N_16534,N_16667);
and U19169 (N_19169,N_16113,N_17006);
xor U19170 (N_19170,N_17526,N_17365);
nand U19171 (N_19171,N_17243,N_17272);
and U19172 (N_19172,N_17434,N_17189);
and U19173 (N_19173,N_17775,N_16568);
or U19174 (N_19174,N_16022,N_16057);
nor U19175 (N_19175,N_17714,N_17393);
nand U19176 (N_19176,N_16917,N_17871);
and U19177 (N_19177,N_16559,N_17036);
and U19178 (N_19178,N_17141,N_16365);
nand U19179 (N_19179,N_17782,N_16198);
and U19180 (N_19180,N_16500,N_17685);
nand U19181 (N_19181,N_16048,N_16114);
and U19182 (N_19182,N_16189,N_16684);
or U19183 (N_19183,N_17823,N_17944);
and U19184 (N_19184,N_16219,N_17995);
nor U19185 (N_19185,N_17482,N_16492);
xnor U19186 (N_19186,N_16848,N_16775);
and U19187 (N_19187,N_17187,N_17726);
or U19188 (N_19188,N_17578,N_16352);
nand U19189 (N_19189,N_17080,N_17360);
and U19190 (N_19190,N_17703,N_17224);
nor U19191 (N_19191,N_16330,N_17632);
xor U19192 (N_19192,N_17433,N_16139);
xnor U19193 (N_19193,N_17383,N_17543);
xor U19194 (N_19194,N_16586,N_17128);
or U19195 (N_19195,N_17440,N_16730);
nor U19196 (N_19196,N_17282,N_17517);
xor U19197 (N_19197,N_16396,N_17052);
nor U19198 (N_19198,N_17385,N_17729);
or U19199 (N_19199,N_16161,N_16678);
and U19200 (N_19200,N_16393,N_17386);
xor U19201 (N_19201,N_17483,N_17270);
nand U19202 (N_19202,N_17886,N_17206);
nor U19203 (N_19203,N_16854,N_16346);
nand U19204 (N_19204,N_16577,N_16716);
or U19205 (N_19205,N_17752,N_16959);
nor U19206 (N_19206,N_17776,N_16352);
nor U19207 (N_19207,N_16060,N_16151);
or U19208 (N_19208,N_16339,N_17136);
and U19209 (N_19209,N_16340,N_16172);
xnor U19210 (N_19210,N_17533,N_17130);
or U19211 (N_19211,N_16488,N_16126);
nor U19212 (N_19212,N_17099,N_16578);
nand U19213 (N_19213,N_16352,N_16769);
xor U19214 (N_19214,N_17154,N_17745);
nor U19215 (N_19215,N_17616,N_16375);
nor U19216 (N_19216,N_16340,N_16328);
and U19217 (N_19217,N_16691,N_17111);
nand U19218 (N_19218,N_17765,N_17317);
or U19219 (N_19219,N_17388,N_16214);
or U19220 (N_19220,N_16631,N_16718);
xor U19221 (N_19221,N_16187,N_17407);
or U19222 (N_19222,N_16259,N_16369);
nor U19223 (N_19223,N_17339,N_17006);
and U19224 (N_19224,N_16629,N_17148);
nor U19225 (N_19225,N_16800,N_17614);
nor U19226 (N_19226,N_16437,N_17127);
nor U19227 (N_19227,N_17958,N_16105);
nand U19228 (N_19228,N_17920,N_16035);
nand U19229 (N_19229,N_17015,N_16663);
nand U19230 (N_19230,N_17804,N_17369);
nand U19231 (N_19231,N_16142,N_16213);
xor U19232 (N_19232,N_16774,N_16173);
and U19233 (N_19233,N_17255,N_17247);
and U19234 (N_19234,N_16220,N_16714);
xor U19235 (N_19235,N_17336,N_17830);
or U19236 (N_19236,N_17537,N_16737);
nor U19237 (N_19237,N_17601,N_16987);
and U19238 (N_19238,N_16106,N_16999);
nor U19239 (N_19239,N_16592,N_17317);
xor U19240 (N_19240,N_16520,N_16475);
and U19241 (N_19241,N_16590,N_17086);
nand U19242 (N_19242,N_17297,N_17072);
or U19243 (N_19243,N_17626,N_16662);
nor U19244 (N_19244,N_17681,N_17844);
xnor U19245 (N_19245,N_17636,N_17208);
nor U19246 (N_19246,N_17508,N_17956);
xnor U19247 (N_19247,N_17804,N_16716);
xnor U19248 (N_19248,N_16430,N_17558);
nand U19249 (N_19249,N_17453,N_17753);
xor U19250 (N_19250,N_16523,N_17169);
xnor U19251 (N_19251,N_17246,N_17728);
or U19252 (N_19252,N_16169,N_16907);
or U19253 (N_19253,N_16746,N_16173);
nor U19254 (N_19254,N_16275,N_16675);
nand U19255 (N_19255,N_17448,N_17370);
nor U19256 (N_19256,N_16630,N_16358);
nand U19257 (N_19257,N_16778,N_16193);
nand U19258 (N_19258,N_16412,N_17943);
nand U19259 (N_19259,N_16773,N_16251);
and U19260 (N_19260,N_17467,N_17980);
and U19261 (N_19261,N_16520,N_17960);
or U19262 (N_19262,N_16924,N_17033);
and U19263 (N_19263,N_17517,N_17798);
nand U19264 (N_19264,N_16608,N_16305);
or U19265 (N_19265,N_16788,N_16406);
or U19266 (N_19266,N_16675,N_16366);
or U19267 (N_19267,N_17016,N_17487);
nor U19268 (N_19268,N_16869,N_17472);
and U19269 (N_19269,N_17778,N_16048);
or U19270 (N_19270,N_16419,N_16763);
nand U19271 (N_19271,N_16322,N_17165);
or U19272 (N_19272,N_16777,N_17044);
nand U19273 (N_19273,N_16404,N_16255);
or U19274 (N_19274,N_17701,N_17514);
nand U19275 (N_19275,N_17721,N_16469);
nor U19276 (N_19276,N_17650,N_17504);
and U19277 (N_19277,N_16431,N_17171);
nand U19278 (N_19278,N_16154,N_17784);
nand U19279 (N_19279,N_17908,N_17488);
nand U19280 (N_19280,N_17963,N_17886);
xor U19281 (N_19281,N_16482,N_16842);
nand U19282 (N_19282,N_16681,N_17754);
xor U19283 (N_19283,N_17241,N_17925);
nor U19284 (N_19284,N_17229,N_16778);
and U19285 (N_19285,N_17345,N_17871);
or U19286 (N_19286,N_17391,N_16096);
nor U19287 (N_19287,N_16029,N_17505);
nand U19288 (N_19288,N_16218,N_17217);
xor U19289 (N_19289,N_16673,N_17891);
nor U19290 (N_19290,N_16190,N_16469);
and U19291 (N_19291,N_16176,N_17523);
or U19292 (N_19292,N_17813,N_17029);
nand U19293 (N_19293,N_17461,N_16484);
nand U19294 (N_19294,N_16746,N_16287);
or U19295 (N_19295,N_16252,N_17865);
or U19296 (N_19296,N_17293,N_16398);
nor U19297 (N_19297,N_17550,N_16981);
nor U19298 (N_19298,N_16964,N_17645);
nand U19299 (N_19299,N_16387,N_17527);
xnor U19300 (N_19300,N_16773,N_16670);
nor U19301 (N_19301,N_17976,N_16188);
xor U19302 (N_19302,N_17173,N_16930);
xnor U19303 (N_19303,N_17566,N_16955);
nand U19304 (N_19304,N_16792,N_16652);
or U19305 (N_19305,N_16614,N_16301);
nand U19306 (N_19306,N_16619,N_17270);
xor U19307 (N_19307,N_16441,N_17412);
nand U19308 (N_19308,N_16715,N_16998);
xor U19309 (N_19309,N_16234,N_17604);
nor U19310 (N_19310,N_17344,N_16863);
nor U19311 (N_19311,N_16525,N_17569);
and U19312 (N_19312,N_16152,N_16813);
nor U19313 (N_19313,N_17470,N_16372);
xnor U19314 (N_19314,N_17988,N_17480);
or U19315 (N_19315,N_16095,N_16349);
nor U19316 (N_19316,N_16406,N_17970);
or U19317 (N_19317,N_16117,N_16835);
or U19318 (N_19318,N_17881,N_17218);
xnor U19319 (N_19319,N_16943,N_17109);
and U19320 (N_19320,N_16734,N_16861);
or U19321 (N_19321,N_17274,N_16547);
xnor U19322 (N_19322,N_16582,N_17341);
nor U19323 (N_19323,N_17329,N_17447);
xor U19324 (N_19324,N_17620,N_16315);
nor U19325 (N_19325,N_16121,N_16993);
nand U19326 (N_19326,N_17573,N_17634);
and U19327 (N_19327,N_17132,N_17957);
nand U19328 (N_19328,N_16663,N_16114);
or U19329 (N_19329,N_16512,N_17706);
or U19330 (N_19330,N_17881,N_17753);
and U19331 (N_19331,N_16273,N_17139);
nor U19332 (N_19332,N_17672,N_17381);
nor U19333 (N_19333,N_17761,N_16418);
or U19334 (N_19334,N_16584,N_17826);
nand U19335 (N_19335,N_16074,N_17388);
nor U19336 (N_19336,N_17127,N_16777);
or U19337 (N_19337,N_17374,N_17658);
or U19338 (N_19338,N_16311,N_17170);
and U19339 (N_19339,N_16162,N_17893);
nor U19340 (N_19340,N_17238,N_17845);
or U19341 (N_19341,N_17815,N_16057);
nand U19342 (N_19342,N_16741,N_16893);
nand U19343 (N_19343,N_17226,N_16706);
xor U19344 (N_19344,N_17133,N_16021);
nand U19345 (N_19345,N_17554,N_16173);
and U19346 (N_19346,N_17001,N_17457);
xor U19347 (N_19347,N_17739,N_16616);
and U19348 (N_19348,N_17134,N_16358);
or U19349 (N_19349,N_17840,N_17450);
xnor U19350 (N_19350,N_16123,N_17319);
nand U19351 (N_19351,N_17635,N_17374);
nor U19352 (N_19352,N_17375,N_16738);
nand U19353 (N_19353,N_16215,N_17592);
nor U19354 (N_19354,N_17352,N_17607);
nand U19355 (N_19355,N_17444,N_16319);
nand U19356 (N_19356,N_17484,N_17687);
nand U19357 (N_19357,N_16091,N_16983);
nor U19358 (N_19358,N_16552,N_17549);
and U19359 (N_19359,N_16162,N_16909);
xnor U19360 (N_19360,N_17422,N_17741);
and U19361 (N_19361,N_16063,N_16894);
nor U19362 (N_19362,N_17489,N_16588);
nand U19363 (N_19363,N_16319,N_17629);
nor U19364 (N_19364,N_16967,N_17213);
nand U19365 (N_19365,N_16240,N_16706);
nand U19366 (N_19366,N_17691,N_16601);
xor U19367 (N_19367,N_16059,N_17707);
xnor U19368 (N_19368,N_16705,N_17461);
xor U19369 (N_19369,N_17274,N_16030);
or U19370 (N_19370,N_16542,N_17490);
nor U19371 (N_19371,N_16453,N_16741);
and U19372 (N_19372,N_17659,N_17034);
nor U19373 (N_19373,N_16775,N_17356);
or U19374 (N_19374,N_17559,N_17545);
nand U19375 (N_19375,N_16819,N_17743);
or U19376 (N_19376,N_16044,N_17787);
xor U19377 (N_19377,N_16780,N_17800);
and U19378 (N_19378,N_16752,N_16202);
or U19379 (N_19379,N_17362,N_17465);
xnor U19380 (N_19380,N_16983,N_17654);
xnor U19381 (N_19381,N_17765,N_16352);
or U19382 (N_19382,N_16656,N_17138);
nand U19383 (N_19383,N_16551,N_16033);
nand U19384 (N_19384,N_17598,N_17440);
nor U19385 (N_19385,N_17927,N_17176);
or U19386 (N_19386,N_17787,N_17009);
nor U19387 (N_19387,N_16402,N_16753);
or U19388 (N_19388,N_17338,N_17194);
nand U19389 (N_19389,N_16753,N_16959);
nor U19390 (N_19390,N_17028,N_16451);
nand U19391 (N_19391,N_16948,N_16787);
xor U19392 (N_19392,N_16995,N_16004);
nor U19393 (N_19393,N_17569,N_17115);
and U19394 (N_19394,N_16018,N_17678);
or U19395 (N_19395,N_16429,N_17288);
and U19396 (N_19396,N_17505,N_17681);
nor U19397 (N_19397,N_16925,N_17418);
nand U19398 (N_19398,N_17042,N_17505);
xor U19399 (N_19399,N_16625,N_16735);
or U19400 (N_19400,N_17238,N_16590);
nor U19401 (N_19401,N_17058,N_16254);
nand U19402 (N_19402,N_16282,N_16518);
nor U19403 (N_19403,N_17054,N_16854);
xnor U19404 (N_19404,N_16088,N_17962);
nand U19405 (N_19405,N_16965,N_17974);
or U19406 (N_19406,N_16522,N_17227);
nor U19407 (N_19407,N_16727,N_16974);
nand U19408 (N_19408,N_17887,N_17369);
xnor U19409 (N_19409,N_16261,N_17382);
or U19410 (N_19410,N_17353,N_16364);
nor U19411 (N_19411,N_16722,N_16464);
xor U19412 (N_19412,N_17547,N_17321);
nand U19413 (N_19413,N_16496,N_17809);
nor U19414 (N_19414,N_17168,N_17574);
nor U19415 (N_19415,N_16712,N_16759);
and U19416 (N_19416,N_17102,N_17026);
nor U19417 (N_19417,N_16343,N_16022);
and U19418 (N_19418,N_17489,N_16653);
xnor U19419 (N_19419,N_16477,N_17278);
or U19420 (N_19420,N_17145,N_16434);
or U19421 (N_19421,N_16028,N_17918);
nand U19422 (N_19422,N_16144,N_16649);
or U19423 (N_19423,N_16717,N_17903);
xor U19424 (N_19424,N_16554,N_17801);
or U19425 (N_19425,N_17206,N_17547);
nor U19426 (N_19426,N_16346,N_17054);
nor U19427 (N_19427,N_16497,N_16614);
or U19428 (N_19428,N_16080,N_17526);
and U19429 (N_19429,N_17469,N_16287);
xnor U19430 (N_19430,N_16489,N_17076);
nor U19431 (N_19431,N_16992,N_16338);
and U19432 (N_19432,N_17271,N_16782);
and U19433 (N_19433,N_16359,N_17198);
nor U19434 (N_19434,N_16573,N_16991);
nor U19435 (N_19435,N_17444,N_17376);
nand U19436 (N_19436,N_17946,N_16500);
nand U19437 (N_19437,N_16720,N_16939);
xnor U19438 (N_19438,N_17405,N_16155);
and U19439 (N_19439,N_16365,N_17433);
xor U19440 (N_19440,N_16965,N_17216);
nand U19441 (N_19441,N_16462,N_16414);
nor U19442 (N_19442,N_17765,N_17754);
nor U19443 (N_19443,N_17185,N_17781);
nand U19444 (N_19444,N_17267,N_16655);
nor U19445 (N_19445,N_17141,N_16588);
nand U19446 (N_19446,N_17969,N_16082);
or U19447 (N_19447,N_16289,N_16287);
and U19448 (N_19448,N_17071,N_17164);
nand U19449 (N_19449,N_17602,N_17577);
or U19450 (N_19450,N_17334,N_17681);
and U19451 (N_19451,N_16852,N_17246);
and U19452 (N_19452,N_17741,N_17617);
nor U19453 (N_19453,N_16990,N_17522);
nand U19454 (N_19454,N_17973,N_17507);
nor U19455 (N_19455,N_16252,N_17455);
or U19456 (N_19456,N_16540,N_16199);
nand U19457 (N_19457,N_16031,N_16882);
or U19458 (N_19458,N_17409,N_16728);
or U19459 (N_19459,N_17663,N_17486);
nor U19460 (N_19460,N_16194,N_17838);
xor U19461 (N_19461,N_16674,N_16951);
and U19462 (N_19462,N_16209,N_17237);
nand U19463 (N_19463,N_16100,N_17946);
xor U19464 (N_19464,N_16488,N_17523);
nand U19465 (N_19465,N_16786,N_16770);
nor U19466 (N_19466,N_17126,N_16735);
nand U19467 (N_19467,N_17183,N_16000);
nor U19468 (N_19468,N_16019,N_17287);
or U19469 (N_19469,N_17169,N_17338);
and U19470 (N_19470,N_17631,N_16030);
nand U19471 (N_19471,N_17827,N_16704);
and U19472 (N_19472,N_17832,N_16960);
xnor U19473 (N_19473,N_16076,N_17725);
xor U19474 (N_19474,N_16877,N_17771);
nor U19475 (N_19475,N_17888,N_16195);
xor U19476 (N_19476,N_17126,N_17798);
xnor U19477 (N_19477,N_17549,N_17003);
or U19478 (N_19478,N_17423,N_16115);
xnor U19479 (N_19479,N_16612,N_16885);
nand U19480 (N_19480,N_17225,N_16312);
nand U19481 (N_19481,N_16102,N_16956);
or U19482 (N_19482,N_16379,N_17604);
or U19483 (N_19483,N_17237,N_16010);
or U19484 (N_19484,N_16939,N_16100);
xor U19485 (N_19485,N_16346,N_17588);
nor U19486 (N_19486,N_17851,N_17131);
and U19487 (N_19487,N_17747,N_17370);
and U19488 (N_19488,N_16105,N_17674);
xnor U19489 (N_19489,N_17911,N_17190);
nor U19490 (N_19490,N_17510,N_17564);
xnor U19491 (N_19491,N_16110,N_16160);
xnor U19492 (N_19492,N_16356,N_17640);
and U19493 (N_19493,N_17530,N_17447);
nand U19494 (N_19494,N_17833,N_16666);
or U19495 (N_19495,N_16108,N_16997);
xnor U19496 (N_19496,N_17173,N_16090);
nor U19497 (N_19497,N_16506,N_17102);
nand U19498 (N_19498,N_17457,N_16001);
or U19499 (N_19499,N_16429,N_16571);
xnor U19500 (N_19500,N_17619,N_16970);
xor U19501 (N_19501,N_17227,N_17621);
xnor U19502 (N_19502,N_16893,N_17188);
and U19503 (N_19503,N_16404,N_16109);
nor U19504 (N_19504,N_16883,N_16071);
nand U19505 (N_19505,N_17189,N_16946);
nand U19506 (N_19506,N_16794,N_17773);
xnor U19507 (N_19507,N_17253,N_17107);
nor U19508 (N_19508,N_17197,N_17092);
or U19509 (N_19509,N_17648,N_16793);
xnor U19510 (N_19510,N_16222,N_17519);
nand U19511 (N_19511,N_16385,N_17281);
or U19512 (N_19512,N_16953,N_16887);
xor U19513 (N_19513,N_17476,N_16731);
or U19514 (N_19514,N_16179,N_17435);
xnor U19515 (N_19515,N_17091,N_16713);
nand U19516 (N_19516,N_17793,N_16296);
nand U19517 (N_19517,N_16225,N_17158);
nor U19518 (N_19518,N_16841,N_17433);
xor U19519 (N_19519,N_16463,N_17164);
nor U19520 (N_19520,N_17465,N_17919);
nor U19521 (N_19521,N_16660,N_16634);
nand U19522 (N_19522,N_17869,N_16045);
nand U19523 (N_19523,N_17197,N_16284);
and U19524 (N_19524,N_17352,N_16959);
nand U19525 (N_19525,N_17137,N_17506);
nand U19526 (N_19526,N_16153,N_17979);
or U19527 (N_19527,N_17240,N_16554);
nand U19528 (N_19528,N_17926,N_16175);
or U19529 (N_19529,N_16970,N_16363);
nor U19530 (N_19530,N_16585,N_17154);
nand U19531 (N_19531,N_16479,N_17724);
nand U19532 (N_19532,N_17746,N_16227);
and U19533 (N_19533,N_16844,N_16497);
xnor U19534 (N_19534,N_16427,N_17889);
xnor U19535 (N_19535,N_17154,N_17179);
xnor U19536 (N_19536,N_17335,N_16666);
and U19537 (N_19537,N_17347,N_17220);
and U19538 (N_19538,N_17617,N_17764);
nand U19539 (N_19539,N_17262,N_16573);
or U19540 (N_19540,N_17549,N_17742);
xnor U19541 (N_19541,N_16180,N_16453);
or U19542 (N_19542,N_17064,N_17119);
xnor U19543 (N_19543,N_16631,N_16274);
xor U19544 (N_19544,N_16186,N_16080);
nand U19545 (N_19545,N_17749,N_17215);
nand U19546 (N_19546,N_16097,N_17941);
nand U19547 (N_19547,N_17158,N_16305);
and U19548 (N_19548,N_17358,N_17905);
nand U19549 (N_19549,N_17504,N_17414);
nor U19550 (N_19550,N_16622,N_17237);
or U19551 (N_19551,N_16256,N_16904);
nor U19552 (N_19552,N_17144,N_16343);
nand U19553 (N_19553,N_16704,N_17065);
and U19554 (N_19554,N_17130,N_17830);
and U19555 (N_19555,N_17893,N_17518);
nor U19556 (N_19556,N_16291,N_16090);
nor U19557 (N_19557,N_17221,N_17219);
and U19558 (N_19558,N_17098,N_17515);
nand U19559 (N_19559,N_16410,N_16287);
nand U19560 (N_19560,N_17667,N_17508);
or U19561 (N_19561,N_17725,N_17972);
or U19562 (N_19562,N_16342,N_16394);
or U19563 (N_19563,N_17215,N_17064);
nor U19564 (N_19564,N_17778,N_17252);
or U19565 (N_19565,N_17941,N_16237);
nor U19566 (N_19566,N_16610,N_17351);
nor U19567 (N_19567,N_17425,N_16382);
or U19568 (N_19568,N_17187,N_17881);
nand U19569 (N_19569,N_16250,N_17560);
or U19570 (N_19570,N_16034,N_16414);
and U19571 (N_19571,N_17966,N_16465);
nand U19572 (N_19572,N_16352,N_17385);
xor U19573 (N_19573,N_17274,N_16863);
xor U19574 (N_19574,N_17585,N_16726);
xor U19575 (N_19575,N_17283,N_17688);
nand U19576 (N_19576,N_17450,N_17870);
and U19577 (N_19577,N_16630,N_16183);
nand U19578 (N_19578,N_16246,N_17552);
xnor U19579 (N_19579,N_16466,N_17716);
nor U19580 (N_19580,N_17669,N_16473);
or U19581 (N_19581,N_16650,N_16752);
nor U19582 (N_19582,N_16944,N_16316);
and U19583 (N_19583,N_17304,N_17546);
or U19584 (N_19584,N_17566,N_17667);
nand U19585 (N_19585,N_17842,N_17223);
and U19586 (N_19586,N_16127,N_17028);
nor U19587 (N_19587,N_17822,N_16769);
xnor U19588 (N_19588,N_16721,N_17506);
or U19589 (N_19589,N_17495,N_17255);
xor U19590 (N_19590,N_16484,N_17717);
and U19591 (N_19591,N_17253,N_16888);
nor U19592 (N_19592,N_17814,N_17632);
xor U19593 (N_19593,N_16832,N_17742);
nand U19594 (N_19594,N_16833,N_17200);
or U19595 (N_19595,N_16382,N_17301);
nor U19596 (N_19596,N_17102,N_16665);
nor U19597 (N_19597,N_17371,N_16635);
nand U19598 (N_19598,N_16527,N_17279);
or U19599 (N_19599,N_17126,N_16762);
and U19600 (N_19600,N_16065,N_17174);
nand U19601 (N_19601,N_17784,N_17279);
or U19602 (N_19602,N_17518,N_16626);
xnor U19603 (N_19603,N_17353,N_16562);
and U19604 (N_19604,N_16809,N_16114);
nor U19605 (N_19605,N_17935,N_16544);
xor U19606 (N_19606,N_17134,N_16577);
nand U19607 (N_19607,N_16168,N_16238);
or U19608 (N_19608,N_16413,N_16825);
xor U19609 (N_19609,N_16047,N_16478);
nor U19610 (N_19610,N_16943,N_17709);
xnor U19611 (N_19611,N_17372,N_17353);
nor U19612 (N_19612,N_17382,N_17157);
nand U19613 (N_19613,N_17288,N_17454);
xnor U19614 (N_19614,N_17397,N_16058);
nand U19615 (N_19615,N_16184,N_16222);
and U19616 (N_19616,N_17077,N_17813);
nand U19617 (N_19617,N_16281,N_17157);
nand U19618 (N_19618,N_17741,N_16569);
and U19619 (N_19619,N_17735,N_17272);
nand U19620 (N_19620,N_16416,N_16309);
nand U19621 (N_19621,N_17259,N_16268);
nand U19622 (N_19622,N_16833,N_17519);
and U19623 (N_19623,N_17691,N_16468);
xor U19624 (N_19624,N_17845,N_16993);
or U19625 (N_19625,N_17644,N_16790);
and U19626 (N_19626,N_16679,N_16088);
xnor U19627 (N_19627,N_17541,N_17235);
nand U19628 (N_19628,N_16659,N_16667);
nand U19629 (N_19629,N_16934,N_16577);
or U19630 (N_19630,N_17478,N_17775);
nor U19631 (N_19631,N_17810,N_16879);
or U19632 (N_19632,N_17368,N_17987);
xnor U19633 (N_19633,N_17287,N_16319);
xnor U19634 (N_19634,N_17537,N_17128);
and U19635 (N_19635,N_17921,N_17599);
xnor U19636 (N_19636,N_16996,N_16353);
and U19637 (N_19637,N_17296,N_16326);
nor U19638 (N_19638,N_17755,N_16136);
and U19639 (N_19639,N_17249,N_17279);
nand U19640 (N_19640,N_17416,N_16892);
or U19641 (N_19641,N_17436,N_17882);
or U19642 (N_19642,N_17082,N_16979);
and U19643 (N_19643,N_17889,N_16083);
nand U19644 (N_19644,N_16813,N_16650);
and U19645 (N_19645,N_17986,N_16393);
nand U19646 (N_19646,N_17363,N_17453);
nand U19647 (N_19647,N_17343,N_16229);
or U19648 (N_19648,N_17703,N_16827);
and U19649 (N_19649,N_16824,N_16687);
nor U19650 (N_19650,N_16756,N_16329);
nand U19651 (N_19651,N_16668,N_17316);
xor U19652 (N_19652,N_16901,N_17076);
nor U19653 (N_19653,N_16249,N_17106);
nor U19654 (N_19654,N_16909,N_17248);
nor U19655 (N_19655,N_17056,N_16762);
nor U19656 (N_19656,N_16896,N_17160);
nor U19657 (N_19657,N_17404,N_16105);
nand U19658 (N_19658,N_17348,N_17608);
nor U19659 (N_19659,N_16102,N_16958);
xor U19660 (N_19660,N_17062,N_17984);
and U19661 (N_19661,N_16160,N_16150);
xor U19662 (N_19662,N_16888,N_17672);
nor U19663 (N_19663,N_17144,N_16373);
nor U19664 (N_19664,N_17881,N_16492);
and U19665 (N_19665,N_17514,N_16030);
and U19666 (N_19666,N_17916,N_17807);
and U19667 (N_19667,N_16409,N_17094);
xnor U19668 (N_19668,N_17934,N_17150);
and U19669 (N_19669,N_17561,N_16776);
xnor U19670 (N_19670,N_16790,N_17000);
xnor U19671 (N_19671,N_16333,N_17508);
nand U19672 (N_19672,N_17027,N_17038);
or U19673 (N_19673,N_16106,N_17097);
nand U19674 (N_19674,N_17192,N_16943);
nor U19675 (N_19675,N_17386,N_17352);
nand U19676 (N_19676,N_17704,N_16306);
xor U19677 (N_19677,N_16140,N_17003);
nand U19678 (N_19678,N_16974,N_17081);
xnor U19679 (N_19679,N_16901,N_17537);
or U19680 (N_19680,N_17589,N_17035);
and U19681 (N_19681,N_17066,N_16669);
and U19682 (N_19682,N_17514,N_17886);
and U19683 (N_19683,N_17907,N_17333);
nor U19684 (N_19684,N_16594,N_16895);
and U19685 (N_19685,N_16072,N_16179);
or U19686 (N_19686,N_16288,N_16566);
xor U19687 (N_19687,N_17035,N_16519);
nand U19688 (N_19688,N_17888,N_17762);
or U19689 (N_19689,N_16214,N_17567);
or U19690 (N_19690,N_16125,N_17831);
xor U19691 (N_19691,N_16818,N_17720);
and U19692 (N_19692,N_17401,N_16562);
and U19693 (N_19693,N_16861,N_16330);
nor U19694 (N_19694,N_17326,N_17440);
and U19695 (N_19695,N_17220,N_16211);
or U19696 (N_19696,N_17356,N_17273);
and U19697 (N_19697,N_17347,N_16037);
nand U19698 (N_19698,N_16819,N_17821);
and U19699 (N_19699,N_17225,N_16538);
and U19700 (N_19700,N_17037,N_17503);
or U19701 (N_19701,N_17676,N_16266);
nor U19702 (N_19702,N_16685,N_17600);
and U19703 (N_19703,N_16312,N_16353);
and U19704 (N_19704,N_16235,N_16463);
xor U19705 (N_19705,N_16736,N_16438);
nand U19706 (N_19706,N_17011,N_17887);
nor U19707 (N_19707,N_17897,N_17219);
or U19708 (N_19708,N_16455,N_16693);
and U19709 (N_19709,N_17706,N_17144);
and U19710 (N_19710,N_16997,N_17950);
nand U19711 (N_19711,N_16480,N_16192);
and U19712 (N_19712,N_16383,N_16485);
xor U19713 (N_19713,N_16151,N_17384);
nor U19714 (N_19714,N_16406,N_17470);
nand U19715 (N_19715,N_16262,N_17353);
xor U19716 (N_19716,N_16261,N_16124);
nor U19717 (N_19717,N_17227,N_17861);
xnor U19718 (N_19718,N_17378,N_17449);
xnor U19719 (N_19719,N_17820,N_16374);
nand U19720 (N_19720,N_17228,N_16206);
xor U19721 (N_19721,N_17126,N_17866);
nor U19722 (N_19722,N_16357,N_16370);
and U19723 (N_19723,N_17204,N_17813);
and U19724 (N_19724,N_16265,N_16703);
xnor U19725 (N_19725,N_16074,N_16916);
xor U19726 (N_19726,N_17909,N_16989);
xor U19727 (N_19727,N_16273,N_16805);
and U19728 (N_19728,N_17717,N_16765);
xor U19729 (N_19729,N_17346,N_16677);
and U19730 (N_19730,N_17006,N_17185);
xor U19731 (N_19731,N_16477,N_16780);
nor U19732 (N_19732,N_16646,N_17926);
nor U19733 (N_19733,N_17137,N_16917);
nor U19734 (N_19734,N_16175,N_16223);
nand U19735 (N_19735,N_16330,N_17735);
nor U19736 (N_19736,N_17195,N_16871);
and U19737 (N_19737,N_16536,N_17470);
xnor U19738 (N_19738,N_17378,N_16456);
nor U19739 (N_19739,N_17316,N_16878);
and U19740 (N_19740,N_16436,N_16359);
nor U19741 (N_19741,N_17968,N_16499);
or U19742 (N_19742,N_17542,N_17697);
nand U19743 (N_19743,N_17011,N_16471);
nand U19744 (N_19744,N_16110,N_16960);
nor U19745 (N_19745,N_17272,N_17753);
and U19746 (N_19746,N_16487,N_17735);
xnor U19747 (N_19747,N_16331,N_17322);
or U19748 (N_19748,N_16838,N_17496);
nand U19749 (N_19749,N_17982,N_17344);
nand U19750 (N_19750,N_17280,N_17416);
xnor U19751 (N_19751,N_17882,N_17133);
nor U19752 (N_19752,N_17532,N_16695);
or U19753 (N_19753,N_16413,N_16250);
and U19754 (N_19754,N_16435,N_17882);
and U19755 (N_19755,N_16592,N_17337);
nand U19756 (N_19756,N_16127,N_16051);
xor U19757 (N_19757,N_17419,N_17707);
nor U19758 (N_19758,N_16879,N_17922);
xor U19759 (N_19759,N_16523,N_17973);
nand U19760 (N_19760,N_17312,N_17132);
and U19761 (N_19761,N_16388,N_16922);
and U19762 (N_19762,N_16110,N_17815);
or U19763 (N_19763,N_17603,N_17515);
or U19764 (N_19764,N_17484,N_17289);
nand U19765 (N_19765,N_17054,N_16465);
xor U19766 (N_19766,N_16160,N_16209);
nor U19767 (N_19767,N_17471,N_17609);
or U19768 (N_19768,N_17930,N_16775);
nand U19769 (N_19769,N_16854,N_16429);
or U19770 (N_19770,N_17862,N_17583);
xnor U19771 (N_19771,N_17451,N_16966);
nor U19772 (N_19772,N_17337,N_17801);
and U19773 (N_19773,N_17636,N_16820);
or U19774 (N_19774,N_17545,N_16073);
nand U19775 (N_19775,N_17904,N_16464);
nor U19776 (N_19776,N_17503,N_16718);
nand U19777 (N_19777,N_16490,N_17337);
or U19778 (N_19778,N_17451,N_16285);
xnor U19779 (N_19779,N_17442,N_16279);
or U19780 (N_19780,N_17560,N_17290);
or U19781 (N_19781,N_16207,N_17197);
or U19782 (N_19782,N_16416,N_17478);
and U19783 (N_19783,N_16912,N_16358);
or U19784 (N_19784,N_16950,N_17542);
nand U19785 (N_19785,N_17613,N_16763);
xor U19786 (N_19786,N_16937,N_16234);
nor U19787 (N_19787,N_16032,N_17254);
xnor U19788 (N_19788,N_16032,N_17330);
or U19789 (N_19789,N_16205,N_17247);
nor U19790 (N_19790,N_16339,N_17607);
nand U19791 (N_19791,N_16775,N_17317);
or U19792 (N_19792,N_16953,N_17160);
nand U19793 (N_19793,N_16692,N_17267);
or U19794 (N_19794,N_17128,N_17482);
nor U19795 (N_19795,N_16673,N_16756);
and U19796 (N_19796,N_17243,N_17381);
and U19797 (N_19797,N_16381,N_16672);
or U19798 (N_19798,N_16489,N_16935);
and U19799 (N_19799,N_17753,N_16336);
or U19800 (N_19800,N_16219,N_17807);
nor U19801 (N_19801,N_17242,N_16309);
nand U19802 (N_19802,N_17167,N_16211);
and U19803 (N_19803,N_17396,N_16346);
nand U19804 (N_19804,N_17924,N_17878);
xnor U19805 (N_19805,N_16052,N_17409);
nand U19806 (N_19806,N_17384,N_16943);
xnor U19807 (N_19807,N_17841,N_17702);
or U19808 (N_19808,N_17535,N_17700);
xnor U19809 (N_19809,N_16985,N_16128);
nor U19810 (N_19810,N_17513,N_17147);
or U19811 (N_19811,N_16276,N_16453);
xor U19812 (N_19812,N_16904,N_16409);
and U19813 (N_19813,N_16372,N_17223);
nor U19814 (N_19814,N_16738,N_16625);
and U19815 (N_19815,N_17692,N_16192);
nor U19816 (N_19816,N_16894,N_16497);
nand U19817 (N_19817,N_16102,N_16388);
nor U19818 (N_19818,N_17064,N_16796);
nand U19819 (N_19819,N_16835,N_17414);
nand U19820 (N_19820,N_16421,N_16088);
and U19821 (N_19821,N_16948,N_17331);
nor U19822 (N_19822,N_17056,N_17903);
nor U19823 (N_19823,N_17151,N_17359);
nand U19824 (N_19824,N_16241,N_16762);
xnor U19825 (N_19825,N_17533,N_16041);
nand U19826 (N_19826,N_17119,N_16915);
and U19827 (N_19827,N_16367,N_17830);
or U19828 (N_19828,N_16490,N_16037);
nand U19829 (N_19829,N_17216,N_16365);
nor U19830 (N_19830,N_16184,N_16825);
xor U19831 (N_19831,N_17833,N_17650);
or U19832 (N_19832,N_16787,N_16211);
nor U19833 (N_19833,N_16458,N_17452);
xnor U19834 (N_19834,N_16342,N_17674);
or U19835 (N_19835,N_17938,N_16931);
nor U19836 (N_19836,N_17041,N_16589);
xor U19837 (N_19837,N_16767,N_17799);
nand U19838 (N_19838,N_17353,N_16817);
nand U19839 (N_19839,N_17812,N_16861);
or U19840 (N_19840,N_17863,N_16123);
xor U19841 (N_19841,N_16279,N_17154);
nor U19842 (N_19842,N_17834,N_17213);
nand U19843 (N_19843,N_17882,N_16239);
and U19844 (N_19844,N_17623,N_16424);
nor U19845 (N_19845,N_17806,N_16479);
and U19846 (N_19846,N_16267,N_17434);
or U19847 (N_19847,N_16614,N_16183);
nand U19848 (N_19848,N_17715,N_16031);
nor U19849 (N_19849,N_16992,N_16642);
xor U19850 (N_19850,N_16424,N_16039);
or U19851 (N_19851,N_16133,N_16204);
xor U19852 (N_19852,N_17034,N_16784);
nand U19853 (N_19853,N_17113,N_17563);
nor U19854 (N_19854,N_17967,N_17228);
and U19855 (N_19855,N_16783,N_16778);
and U19856 (N_19856,N_16036,N_17306);
and U19857 (N_19857,N_17287,N_17910);
xnor U19858 (N_19858,N_16386,N_17681);
nor U19859 (N_19859,N_17554,N_17658);
nor U19860 (N_19860,N_16261,N_16903);
xnor U19861 (N_19861,N_16716,N_16121);
nor U19862 (N_19862,N_17398,N_16671);
xor U19863 (N_19863,N_17372,N_16008);
nor U19864 (N_19864,N_17777,N_17978);
and U19865 (N_19865,N_16595,N_17107);
and U19866 (N_19866,N_16955,N_16297);
xnor U19867 (N_19867,N_17970,N_16825);
and U19868 (N_19868,N_16047,N_17873);
nor U19869 (N_19869,N_16019,N_17982);
xor U19870 (N_19870,N_17794,N_16897);
xnor U19871 (N_19871,N_16373,N_17779);
xnor U19872 (N_19872,N_16684,N_17326);
or U19873 (N_19873,N_17100,N_16712);
xnor U19874 (N_19874,N_16918,N_16865);
and U19875 (N_19875,N_17740,N_16142);
and U19876 (N_19876,N_17158,N_16447);
and U19877 (N_19877,N_16024,N_16925);
and U19878 (N_19878,N_17947,N_17076);
and U19879 (N_19879,N_17543,N_16298);
or U19880 (N_19880,N_17069,N_16704);
and U19881 (N_19881,N_17020,N_17071);
or U19882 (N_19882,N_16258,N_16730);
xor U19883 (N_19883,N_16231,N_17084);
xnor U19884 (N_19884,N_17308,N_17153);
or U19885 (N_19885,N_17664,N_17849);
nand U19886 (N_19886,N_17580,N_16188);
or U19887 (N_19887,N_16378,N_17157);
or U19888 (N_19888,N_17412,N_17929);
nand U19889 (N_19889,N_16024,N_17793);
nand U19890 (N_19890,N_17776,N_17641);
or U19891 (N_19891,N_16302,N_16786);
nand U19892 (N_19892,N_16199,N_17233);
and U19893 (N_19893,N_17036,N_16147);
nor U19894 (N_19894,N_16633,N_17412);
nand U19895 (N_19895,N_17989,N_16418);
nor U19896 (N_19896,N_16991,N_16006);
or U19897 (N_19897,N_16104,N_17804);
nor U19898 (N_19898,N_17447,N_17628);
nor U19899 (N_19899,N_16167,N_17758);
and U19900 (N_19900,N_16330,N_17638);
nand U19901 (N_19901,N_17302,N_16563);
or U19902 (N_19902,N_16527,N_16983);
or U19903 (N_19903,N_17667,N_17192);
nand U19904 (N_19904,N_16092,N_16403);
nand U19905 (N_19905,N_16598,N_17453);
nand U19906 (N_19906,N_17541,N_17397);
or U19907 (N_19907,N_16642,N_16524);
or U19908 (N_19908,N_17408,N_16185);
and U19909 (N_19909,N_16173,N_17509);
or U19910 (N_19910,N_16990,N_17524);
xnor U19911 (N_19911,N_17593,N_17393);
and U19912 (N_19912,N_16142,N_16923);
and U19913 (N_19913,N_16434,N_16282);
xnor U19914 (N_19914,N_17425,N_17242);
nor U19915 (N_19915,N_17864,N_17388);
nor U19916 (N_19916,N_16332,N_16973);
nor U19917 (N_19917,N_17764,N_16446);
or U19918 (N_19918,N_17153,N_16128);
and U19919 (N_19919,N_17963,N_16310);
nand U19920 (N_19920,N_16189,N_16963);
nor U19921 (N_19921,N_16683,N_17673);
xor U19922 (N_19922,N_16515,N_16726);
nor U19923 (N_19923,N_17394,N_16164);
or U19924 (N_19924,N_17318,N_17821);
nor U19925 (N_19925,N_16785,N_17845);
nor U19926 (N_19926,N_16578,N_16340);
nor U19927 (N_19927,N_17626,N_17923);
xor U19928 (N_19928,N_16317,N_16716);
and U19929 (N_19929,N_16161,N_16625);
or U19930 (N_19930,N_17958,N_16720);
nor U19931 (N_19931,N_16157,N_16467);
or U19932 (N_19932,N_17641,N_17330);
nand U19933 (N_19933,N_16828,N_16202);
or U19934 (N_19934,N_17028,N_17495);
and U19935 (N_19935,N_17699,N_16786);
nand U19936 (N_19936,N_16481,N_17472);
nand U19937 (N_19937,N_16043,N_17100);
or U19938 (N_19938,N_17182,N_17511);
xnor U19939 (N_19939,N_16998,N_16407);
nor U19940 (N_19940,N_16800,N_17373);
or U19941 (N_19941,N_17847,N_17506);
and U19942 (N_19942,N_17028,N_16159);
nor U19943 (N_19943,N_17078,N_16709);
nand U19944 (N_19944,N_17320,N_16465);
and U19945 (N_19945,N_16823,N_17118);
or U19946 (N_19946,N_16330,N_16720);
and U19947 (N_19947,N_17322,N_17740);
nand U19948 (N_19948,N_17597,N_17641);
nand U19949 (N_19949,N_16063,N_16151);
nand U19950 (N_19950,N_17331,N_16904);
or U19951 (N_19951,N_16481,N_17404);
and U19952 (N_19952,N_16569,N_17730);
nand U19953 (N_19953,N_17475,N_17055);
nand U19954 (N_19954,N_16561,N_16339);
xnor U19955 (N_19955,N_17018,N_17154);
or U19956 (N_19956,N_16188,N_17020);
xor U19957 (N_19957,N_16582,N_17040);
nor U19958 (N_19958,N_16250,N_17771);
nand U19959 (N_19959,N_17302,N_17732);
xnor U19960 (N_19960,N_16105,N_17637);
and U19961 (N_19961,N_17106,N_16408);
nand U19962 (N_19962,N_16038,N_17937);
and U19963 (N_19963,N_17857,N_16871);
xnor U19964 (N_19964,N_17019,N_17780);
and U19965 (N_19965,N_16390,N_16859);
or U19966 (N_19966,N_16684,N_16922);
xnor U19967 (N_19967,N_16667,N_16400);
nand U19968 (N_19968,N_17149,N_17070);
and U19969 (N_19969,N_16815,N_16133);
or U19970 (N_19970,N_17803,N_17466);
nand U19971 (N_19971,N_17643,N_16371);
or U19972 (N_19972,N_16187,N_17444);
or U19973 (N_19973,N_16896,N_16514);
or U19974 (N_19974,N_17736,N_16622);
nor U19975 (N_19975,N_17545,N_17678);
nand U19976 (N_19976,N_17139,N_16446);
nand U19977 (N_19977,N_17412,N_17064);
or U19978 (N_19978,N_16643,N_17923);
or U19979 (N_19979,N_16658,N_16868);
and U19980 (N_19980,N_16707,N_17326);
or U19981 (N_19981,N_16382,N_16939);
xor U19982 (N_19982,N_17645,N_17506);
or U19983 (N_19983,N_16825,N_16633);
or U19984 (N_19984,N_17721,N_17246);
nand U19985 (N_19985,N_17406,N_17830);
and U19986 (N_19986,N_17467,N_16087);
and U19987 (N_19987,N_16626,N_16019);
nand U19988 (N_19988,N_17833,N_16602);
or U19989 (N_19989,N_16363,N_17074);
nand U19990 (N_19990,N_17098,N_17498);
nor U19991 (N_19991,N_16307,N_17487);
or U19992 (N_19992,N_16956,N_16131);
xor U19993 (N_19993,N_16168,N_17182);
nor U19994 (N_19994,N_17914,N_16323);
nand U19995 (N_19995,N_17361,N_16452);
xnor U19996 (N_19996,N_17295,N_17014);
xor U19997 (N_19997,N_16832,N_16481);
or U19998 (N_19998,N_17882,N_16461);
xor U19999 (N_19999,N_16338,N_17647);
nand U20000 (N_20000,N_19036,N_18800);
nand U20001 (N_20001,N_18062,N_19369);
nor U20002 (N_20002,N_18669,N_19724);
xor U20003 (N_20003,N_18661,N_18691);
nor U20004 (N_20004,N_18330,N_18040);
nand U20005 (N_20005,N_19461,N_19764);
or U20006 (N_20006,N_18806,N_19209);
and U20007 (N_20007,N_19677,N_18607);
nand U20008 (N_20008,N_18114,N_18585);
nor U20009 (N_20009,N_18896,N_19236);
xnor U20010 (N_20010,N_19206,N_18979);
xor U20011 (N_20011,N_19229,N_18070);
nor U20012 (N_20012,N_19927,N_18413);
and U20013 (N_20013,N_19508,N_19252);
and U20014 (N_20014,N_18558,N_18518);
or U20015 (N_20015,N_19408,N_19919);
and U20016 (N_20016,N_18653,N_18651);
or U20017 (N_20017,N_18210,N_18411);
or U20018 (N_20018,N_18901,N_19345);
nand U20019 (N_20019,N_18381,N_19616);
and U20020 (N_20020,N_18679,N_19686);
nor U20021 (N_20021,N_18064,N_19890);
and U20022 (N_20022,N_18856,N_18637);
nor U20023 (N_20023,N_19270,N_19460);
xnor U20024 (N_20024,N_18935,N_18619);
xor U20025 (N_20025,N_18030,N_19184);
and U20026 (N_20026,N_18427,N_18861);
or U20027 (N_20027,N_18057,N_19348);
xor U20028 (N_20028,N_18843,N_18147);
nor U20029 (N_20029,N_18274,N_18401);
or U20030 (N_20030,N_19715,N_18096);
or U20031 (N_20031,N_19549,N_19147);
nand U20032 (N_20032,N_18279,N_19350);
nand U20033 (N_20033,N_18605,N_19498);
xor U20034 (N_20034,N_18635,N_19231);
xor U20035 (N_20035,N_19177,N_19905);
and U20036 (N_20036,N_19099,N_18655);
and U20037 (N_20037,N_19719,N_18940);
nor U20038 (N_20038,N_19753,N_19615);
nand U20039 (N_20039,N_19876,N_19988);
nor U20040 (N_20040,N_18272,N_18287);
and U20041 (N_20041,N_19219,N_18278);
xor U20042 (N_20042,N_18270,N_18068);
and U20043 (N_20043,N_19391,N_19319);
or U20044 (N_20044,N_18601,N_18506);
xor U20045 (N_20045,N_19104,N_19928);
and U20046 (N_20046,N_19906,N_18458);
and U20047 (N_20047,N_18392,N_18160);
nor U20048 (N_20048,N_18968,N_18173);
nor U20049 (N_20049,N_18532,N_19982);
xor U20050 (N_20050,N_18474,N_18025);
xnor U20051 (N_20051,N_18337,N_18898);
nand U20052 (N_20052,N_19900,N_18350);
nor U20053 (N_20053,N_18719,N_18103);
or U20054 (N_20054,N_19773,N_19993);
xor U20055 (N_20055,N_19968,N_19422);
and U20056 (N_20056,N_19805,N_18393);
xor U20057 (N_20057,N_19664,N_18403);
nand U20058 (N_20058,N_18101,N_19353);
nor U20059 (N_20059,N_19456,N_19529);
nor U20060 (N_20060,N_19392,N_18541);
nand U20061 (N_20061,N_18342,N_19593);
and U20062 (N_20062,N_19584,N_19126);
and U20063 (N_20063,N_18600,N_19495);
or U20064 (N_20064,N_18325,N_18492);
and U20065 (N_20065,N_18684,N_18914);
or U20066 (N_20066,N_18264,N_18438);
nand U20067 (N_20067,N_19793,N_18513);
or U20068 (N_20068,N_19527,N_18406);
nand U20069 (N_20069,N_19094,N_18917);
nand U20070 (N_20070,N_18459,N_19999);
and U20071 (N_20071,N_18467,N_18072);
nor U20072 (N_20072,N_18563,N_19571);
xnor U20073 (N_20073,N_19926,N_18465);
xnor U20074 (N_20074,N_19134,N_19187);
nor U20075 (N_20075,N_19577,N_19019);
and U20076 (N_20076,N_19608,N_18457);
and U20077 (N_20077,N_19636,N_19076);
xnor U20078 (N_20078,N_18308,N_18499);
xnor U20079 (N_20079,N_18053,N_19619);
nor U20080 (N_20080,N_19056,N_19895);
nand U20081 (N_20081,N_18662,N_19908);
and U20082 (N_20082,N_19443,N_19935);
nand U20083 (N_20083,N_19781,N_19752);
or U20084 (N_20084,N_18472,N_18396);
and U20085 (N_20085,N_19127,N_19092);
nand U20086 (N_20086,N_18702,N_19075);
xnor U20087 (N_20087,N_18262,N_19264);
nor U20088 (N_20088,N_18858,N_18553);
or U20089 (N_20089,N_18715,N_18723);
or U20090 (N_20090,N_19833,N_19342);
nand U20091 (N_20091,N_18190,N_19858);
nand U20092 (N_20092,N_18243,N_18616);
and U20093 (N_20093,N_18080,N_18034);
nand U20094 (N_20094,N_18306,N_18755);
nor U20095 (N_20095,N_19417,N_19803);
xnor U20096 (N_20096,N_18181,N_18146);
and U20097 (N_20097,N_19115,N_19555);
nor U20098 (N_20098,N_18199,N_19845);
xor U20099 (N_20099,N_18893,N_18491);
xor U20100 (N_20100,N_19748,N_18771);
and U20101 (N_20101,N_19305,N_18316);
or U20102 (N_20102,N_19703,N_19638);
or U20103 (N_20103,N_18905,N_19878);
xor U20104 (N_20104,N_19655,N_19378);
or U20105 (N_20105,N_19789,N_19611);
xor U20106 (N_20106,N_19871,N_19038);
xor U20107 (N_20107,N_18753,N_19225);
xnor U20108 (N_20108,N_18874,N_18549);
nand U20109 (N_20109,N_19358,N_18725);
and U20110 (N_20110,N_18952,N_18167);
nor U20111 (N_20111,N_19405,N_18934);
nor U20112 (N_20112,N_18326,N_18271);
nor U20113 (N_20113,N_19738,N_19761);
nand U20114 (N_20114,N_18764,N_19067);
and U20115 (N_20115,N_19989,N_19612);
or U20116 (N_20116,N_18084,N_19357);
xor U20117 (N_20117,N_19554,N_18945);
and U20118 (N_20118,N_18120,N_19261);
and U20119 (N_20119,N_19532,N_19827);
xnor U20120 (N_20120,N_19644,N_18688);
nor U20121 (N_20121,N_19969,N_18408);
xnor U20122 (N_20122,N_19208,N_18632);
nand U20123 (N_20123,N_18864,N_19359);
or U20124 (N_20124,N_18223,N_19741);
nor U20125 (N_20125,N_19736,N_19367);
and U20126 (N_20126,N_18156,N_19472);
xor U20127 (N_20127,N_18335,N_18424);
xnor U20128 (N_20128,N_19477,N_19063);
nor U20129 (N_20129,N_18008,N_19662);
xor U20130 (N_20130,N_19368,N_19192);
nor U20131 (N_20131,N_18341,N_19862);
xor U20132 (N_20132,N_18672,N_19487);
or U20133 (N_20133,N_18471,N_18689);
or U20134 (N_20134,N_19308,N_18422);
and U20135 (N_20135,N_18811,N_19163);
or U20136 (N_20136,N_18803,N_19976);
or U20137 (N_20137,N_19907,N_19158);
or U20138 (N_20138,N_19297,N_19710);
nor U20139 (N_20139,N_18289,N_19573);
xnor U20140 (N_20140,N_19239,N_18899);
and U20141 (N_20141,N_18744,N_18838);
or U20142 (N_20142,N_19389,N_19627);
or U20143 (N_20143,N_18721,N_19165);
xor U20144 (N_20144,N_18907,N_18624);
or U20145 (N_20145,N_18495,N_19084);
xor U20146 (N_20146,N_18011,N_18828);
nand U20147 (N_20147,N_18583,N_19060);
or U20148 (N_20148,N_18774,N_18108);
and U20149 (N_20149,N_19037,N_18926);
nor U20150 (N_20150,N_19872,N_19784);
xnor U20151 (N_20151,N_18577,N_18452);
and U20152 (N_20152,N_19483,N_19840);
or U20153 (N_20153,N_19517,N_18884);
or U20154 (N_20154,N_19996,N_19135);
nor U20155 (N_20155,N_19977,N_18107);
xnor U20156 (N_20156,N_18165,N_18244);
nand U20157 (N_20157,N_18608,N_18185);
nor U20158 (N_20158,N_18399,N_19054);
nand U20159 (N_20159,N_19288,N_18482);
or U20160 (N_20160,N_19659,N_19551);
nand U20161 (N_20161,N_19772,N_19216);
nand U20162 (N_20162,N_18727,N_19466);
and U20163 (N_20163,N_18588,N_19865);
or U20164 (N_20164,N_18370,N_18493);
or U20165 (N_20165,N_18225,N_18111);
nor U20166 (N_20166,N_19475,N_19271);
or U20167 (N_20167,N_18923,N_19595);
or U20168 (N_20168,N_19057,N_19141);
nand U20169 (N_20169,N_18464,N_18888);
nand U20170 (N_20170,N_19296,N_18509);
nand U20171 (N_20171,N_18820,N_18109);
xor U20172 (N_20172,N_19843,N_18242);
nor U20173 (N_20173,N_19541,N_19370);
and U20174 (N_20174,N_18045,N_18310);
nand U20175 (N_20175,N_19775,N_19332);
nor U20176 (N_20176,N_19875,N_19376);
or U20177 (N_20177,N_18537,N_19959);
nand U20178 (N_20178,N_19869,N_19201);
nand U20179 (N_20179,N_18017,N_19814);
xor U20180 (N_20180,N_19637,N_18266);
and U20181 (N_20181,N_19621,N_19892);
nor U20182 (N_20182,N_19321,N_18799);
nand U20183 (N_20183,N_19688,N_19138);
nor U20184 (N_20184,N_19281,N_18136);
xor U20185 (N_20185,N_18373,N_19618);
xnor U20186 (N_20186,N_18696,N_18245);
nand U20187 (N_20187,N_18463,N_19486);
nor U20188 (N_20188,N_19128,N_18962);
xnor U20189 (N_20189,N_19779,N_19089);
nand U20190 (N_20190,N_18987,N_19471);
nor U20191 (N_20191,N_19744,N_18460);
nor U20192 (N_20192,N_19630,N_19899);
nor U20193 (N_20193,N_18250,N_19235);
nand U20194 (N_20194,N_19533,N_18860);
nor U20195 (N_20195,N_19888,N_19432);
xnor U20196 (N_20196,N_19033,N_18339);
nor U20197 (N_20197,N_19142,N_18137);
and U20198 (N_20198,N_18535,N_19952);
nand U20199 (N_20199,N_19275,N_19974);
nand U20200 (N_20200,N_18054,N_19716);
xnor U20201 (N_20201,N_18311,N_19830);
or U20202 (N_20202,N_18061,N_18561);
nand U20203 (N_20203,N_18630,N_19390);
nor U20204 (N_20204,N_18200,N_18827);
nor U20205 (N_20205,N_19220,N_19384);
or U20206 (N_20206,N_19834,N_18718);
nand U20207 (N_20207,N_18999,N_18713);
nor U20208 (N_20208,N_18612,N_18834);
nor U20209 (N_20209,N_18991,N_19717);
or U20210 (N_20210,N_18484,N_19354);
nor U20211 (N_20211,N_19193,N_19301);
and U20212 (N_20212,N_19320,N_19428);
nand U20213 (N_20213,N_19095,N_18517);
and U20214 (N_20214,N_19918,N_18757);
nand U20215 (N_20215,N_18477,N_18890);
and U20216 (N_20216,N_18487,N_19942);
xnor U20217 (N_20217,N_19566,N_19985);
xor U20218 (N_20218,N_19767,N_18177);
nand U20219 (N_20219,N_18760,N_19100);
nor U20220 (N_20220,N_19912,N_19429);
nor U20221 (N_20221,N_18134,N_19485);
nand U20222 (N_20222,N_18104,N_19480);
nor U20223 (N_20223,N_19790,N_19131);
xor U20224 (N_20224,N_18257,N_18446);
nand U20225 (N_20225,N_19874,N_18969);
and U20226 (N_20226,N_19445,N_18031);
nand U20227 (N_20227,N_18739,N_19597);
xnor U20228 (N_20228,N_18903,N_19226);
and U20229 (N_20229,N_19534,N_18423);
xor U20230 (N_20230,N_19758,N_19030);
or U20231 (N_20231,N_19312,N_18404);
or U20232 (N_20232,N_19238,N_19546);
xnor U20233 (N_20233,N_19351,N_19007);
or U20234 (N_20234,N_19340,N_18789);
and U20235 (N_20235,N_18765,N_19064);
and U20236 (N_20236,N_19409,N_18873);
xor U20237 (N_20237,N_19897,N_18228);
and U20238 (N_20238,N_18380,N_19995);
nor U20239 (N_20239,N_19279,N_18439);
and U20240 (N_20240,N_19923,N_18420);
xor U20241 (N_20241,N_18117,N_19972);
xor U20242 (N_20242,N_19511,N_19800);
and U20243 (N_20243,N_18942,N_18883);
and U20244 (N_20244,N_18816,N_19170);
nor U20245 (N_20245,N_19642,N_18386);
nand U20246 (N_20246,N_18846,N_18356);
and U20247 (N_20247,N_18009,N_18248);
nor U20248 (N_20248,N_18273,N_19787);
and U20249 (N_20249,N_19420,N_18961);
nor U20250 (N_20250,N_18286,N_19058);
nand U20251 (N_20251,N_19161,N_19633);
and U20252 (N_20252,N_18218,N_19263);
and U20253 (N_20253,N_19137,N_18870);
xnor U20254 (N_20254,N_19558,N_19087);
or U20255 (N_20255,N_19822,N_18292);
nor U20256 (N_20256,N_19499,N_19617);
xor U20257 (N_20257,N_18194,N_18402);
xnor U20258 (N_20258,N_18504,N_19808);
or U20259 (N_20259,N_19535,N_19223);
or U20260 (N_20260,N_18391,N_19887);
xor U20261 (N_20261,N_19071,N_19698);
xnor U20262 (N_20262,N_18813,N_18720);
nand U20263 (N_20263,N_19658,N_19770);
nand U20264 (N_20264,N_19439,N_19401);
nand U20265 (N_20265,N_19681,N_18043);
or U20266 (N_20266,N_18020,N_19706);
nand U20267 (N_20267,N_18299,N_19467);
nor U20268 (N_20268,N_19667,N_18805);
and U20269 (N_20269,N_19813,N_19462);
nand U20270 (N_20270,N_18140,N_19675);
and U20271 (N_20271,N_18598,N_18745);
nor U20272 (N_20272,N_18695,N_19277);
xnor U20273 (N_20273,N_19157,N_19832);
nor U20274 (N_20274,N_19241,N_19596);
xor U20275 (N_20275,N_18963,N_18018);
xor U20276 (N_20276,N_18918,N_18357);
nor U20277 (N_20277,N_19806,N_18614);
and U20278 (N_20278,N_18568,N_18562);
and U20279 (N_20279,N_19222,N_18269);
and U20280 (N_20280,N_19647,N_19860);
xnor U20281 (N_20281,N_18943,N_18466);
and U20282 (N_20282,N_19243,N_18106);
nor U20283 (N_20283,N_18510,N_18302);
nor U20284 (N_20284,N_18151,N_18355);
and U20285 (N_20285,N_19478,N_18418);
and U20286 (N_20286,N_18894,N_18232);
nor U20287 (N_20287,N_18334,N_19025);
and U20288 (N_20288,N_19078,N_18220);
nand U20289 (N_20289,N_19427,N_18013);
xnor U20290 (N_20290,N_18835,N_19930);
xnor U20291 (N_20291,N_19185,N_19403);
and U20292 (N_20292,N_18946,N_19657);
nand U20293 (N_20293,N_19425,N_18397);
or U20294 (N_20294,N_18231,N_19129);
xor U20295 (N_20295,N_18582,N_18039);
nand U20296 (N_20296,N_18176,N_18318);
xor U20297 (N_20297,N_18340,N_18808);
or U20298 (N_20298,N_19629,N_19570);
and U20299 (N_20299,N_18742,N_18768);
or U20300 (N_20300,N_19837,N_19205);
nand U20301 (N_20301,N_19091,N_19902);
xor U20302 (N_20302,N_19898,N_18889);
nor U20303 (N_20303,N_18019,N_18412);
and U20304 (N_20304,N_18312,N_18857);
xor U20305 (N_20305,N_18773,N_19237);
and U20306 (N_20306,N_19762,N_19901);
xor U20307 (N_20307,N_18960,N_19842);
xor U20308 (N_20308,N_19635,N_19397);
nor U20309 (N_20309,N_19685,N_19065);
and U20310 (N_20310,N_18970,N_19178);
nand U20311 (N_20311,N_19697,N_18836);
nor U20312 (N_20312,N_18643,N_18394);
xor U20313 (N_20313,N_18930,N_19352);
nand U20314 (N_20314,N_18258,N_18448);
and U20315 (N_20315,N_18950,N_18085);
or U20316 (N_20316,N_19451,N_18209);
nor U20317 (N_20317,N_18133,N_19413);
nand U20318 (N_20318,N_19361,N_19649);
xnor U20319 (N_20319,N_19341,N_18170);
nand U20320 (N_20320,N_18633,N_19613);
and U20321 (N_20321,N_18912,N_19868);
and U20322 (N_20322,N_19318,N_19160);
and U20323 (N_20323,N_18021,N_18938);
or U20324 (N_20324,N_19861,N_18369);
nor U20325 (N_20325,N_19956,N_19143);
or U20326 (N_20326,N_18135,N_18660);
or U20327 (N_20327,N_18468,N_19856);
or U20328 (N_20328,N_18777,N_19242);
nand U20329 (N_20329,N_18360,N_19124);
nand U20330 (N_20330,N_18145,N_18815);
nor U20331 (N_20331,N_18321,N_18158);
nor U20332 (N_20332,N_18975,N_19768);
or U20333 (N_20333,N_18824,N_19419);
nand U20334 (N_20334,N_18939,N_18155);
nor U20335 (N_20335,N_19097,N_19939);
and U20336 (N_20336,N_18620,N_18113);
or U20337 (N_20337,N_19849,N_18265);
nand U20338 (N_20338,N_19922,N_18980);
xor U20339 (N_20339,N_18840,N_19692);
nand U20340 (N_20340,N_18586,N_19622);
xor U20341 (N_20341,N_19711,N_18260);
nand U20342 (N_20342,N_18236,N_19186);
and U20343 (N_20343,N_18461,N_18164);
and U20344 (N_20344,N_18233,N_19610);
and U20345 (N_20345,N_19695,N_19568);
and U20346 (N_20346,N_19669,N_18201);
and U20347 (N_20347,N_19444,N_19245);
and U20348 (N_20348,N_18694,N_19398);
xnor U20349 (N_20349,N_19010,N_19150);
xnor U20350 (N_20350,N_19743,N_19004);
xor U20351 (N_20351,N_19481,N_19228);
nand U20352 (N_20352,N_19122,N_18812);
nand U20353 (N_20353,N_18307,N_19331);
xnor U20354 (N_20354,N_18573,N_18255);
or U20355 (N_20355,N_18527,N_18037);
or U20356 (N_20356,N_18788,N_19050);
and U20357 (N_20357,N_18035,N_18436);
or U20358 (N_20358,N_19978,N_18747);
nor U20359 (N_20359,N_19146,N_18489);
xnor U20360 (N_20360,N_18826,N_18618);
nand U20361 (N_20361,N_19624,N_18703);
and U20362 (N_20362,N_18186,N_18324);
nand U20363 (N_20363,N_18049,N_19255);
nor U20364 (N_20364,N_18162,N_19096);
and U20365 (N_20365,N_19730,N_18784);
nand U20366 (N_20366,N_18869,N_19041);
nand U20367 (N_20367,N_18794,N_18994);
and U20368 (N_20368,N_18851,N_18673);
nand U20369 (N_20369,N_19410,N_18615);
nand U20370 (N_20370,N_18783,N_19654);
and U20371 (N_20371,N_18748,N_19994);
nand U20372 (N_20372,N_19528,N_19864);
nand U20373 (N_20373,N_19981,N_18483);
or U20374 (N_20374,N_19777,N_18118);
or U20375 (N_20375,N_18511,N_18609);
and U20376 (N_20376,N_18554,N_18138);
xnor U20377 (N_20377,N_18012,N_18485);
nand U20378 (N_20378,N_18595,N_19335);
nor U20379 (N_20379,N_19268,N_19623);
nor U20380 (N_20380,N_18868,N_19034);
and U20381 (N_20381,N_19195,N_18832);
and U20382 (N_20382,N_18776,N_19678);
nand U20383 (N_20383,N_19735,N_19811);
nor U20384 (N_20384,N_19375,N_19374);
and U20385 (N_20385,N_18610,N_19931);
and U20386 (N_20386,N_19022,N_18915);
and U20387 (N_20387,N_19877,N_19921);
nor U20388 (N_20388,N_18395,N_19246);
or U20389 (N_20389,N_19029,N_18119);
nand U20390 (N_20390,N_18175,N_19924);
nor U20391 (N_20391,N_19937,N_18479);
or U20392 (N_20392,N_19267,N_19377);
and U20393 (N_20393,N_18367,N_19825);
or U20394 (N_20394,N_19166,N_18410);
xor U20395 (N_20395,N_18204,N_19660);
xor U20396 (N_20396,N_18575,N_18216);
nor U20397 (N_20397,N_19510,N_19081);
or U20398 (N_20398,N_18539,N_19882);
xor U20399 (N_20399,N_19980,N_18986);
nor U20400 (N_20400,N_18368,N_18866);
nand U20401 (N_20401,N_19380,N_19572);
and U20402 (N_20402,N_19194,N_19525);
nor U20403 (N_20403,N_19960,N_19521);
xor U20404 (N_20404,N_18705,N_19070);
nor U20405 (N_20405,N_18685,N_19932);
and U20406 (N_20406,N_18732,N_18105);
nor U20407 (N_20407,N_19017,N_19778);
nor U20408 (N_20408,N_18640,N_19372);
nand U20409 (N_20409,N_18944,N_19215);
nand U20410 (N_20410,N_19329,N_19190);
or U20411 (N_20411,N_18842,N_19285);
or U20412 (N_20412,N_19802,N_19167);
or U20413 (N_20413,N_18116,N_19737);
nor U20414 (N_20414,N_19728,N_19552);
xor U20415 (N_20415,N_18936,N_18543);
xnor U20416 (N_20416,N_18507,N_19366);
nand U20417 (N_20417,N_19574,N_19093);
xor U20418 (N_20418,N_18989,N_19411);
or U20419 (N_20419,N_18400,N_19214);
nand U20420 (N_20420,N_18726,N_18481);
xor U20421 (N_20421,N_18769,N_19991);
nor U20422 (N_20422,N_18235,N_19317);
nand U20423 (N_20423,N_18428,N_18929);
or U20424 (N_20424,N_18295,N_18627);
nor U20425 (N_20425,N_19693,N_18320);
xnor U20426 (N_20426,N_19282,N_18664);
or U20427 (N_20427,N_19149,N_19749);
or U20428 (N_20428,N_19344,N_19254);
nor U20429 (N_20429,N_19538,N_18924);
and U20430 (N_20430,N_19807,N_19426);
xnor U20431 (N_20431,N_18767,N_18736);
xnor U20432 (N_20432,N_19414,N_19745);
xnor U20433 (N_20433,N_19274,N_19273);
xnor U20434 (N_20434,N_19819,N_19292);
nor U20435 (N_20435,N_18125,N_19171);
nand U20436 (N_20436,N_18886,N_18131);
xor U20437 (N_20437,N_18006,N_18831);
nand U20438 (N_20438,N_19809,N_18480);
nand U20439 (N_20439,N_18536,N_19591);
and U20440 (N_20440,N_19381,N_19590);
or U20441 (N_20441,N_19441,N_19559);
nand U20442 (N_20442,N_19073,N_18954);
nor U20443 (N_20443,N_18547,N_18810);
nor U20444 (N_20444,N_19151,N_19757);
or U20445 (N_20445,N_18211,N_19965);
or U20446 (N_20446,N_19713,N_19132);
and U20447 (N_20447,N_18349,N_18447);
xor U20448 (N_20448,N_19652,N_19459);
xor U20449 (N_20449,N_18303,N_18599);
xor U20450 (N_20450,N_19324,N_19399);
or U20451 (N_20451,N_18964,N_19962);
and U20452 (N_20452,N_18322,N_18711);
and U20453 (N_20453,N_18453,N_18848);
nor U20454 (N_20454,N_18086,N_18128);
or U20455 (N_20455,N_18126,N_19756);
nor U20456 (N_20456,N_19018,N_18364);
or U20457 (N_20457,N_19482,N_18143);
or U20458 (N_20458,N_19614,N_19123);
or U20459 (N_20459,N_19859,N_18932);
or U20460 (N_20460,N_18763,N_18390);
nand U20461 (N_20461,N_18738,N_18171);
xor U20462 (N_20462,N_19500,N_18729);
xnor U20463 (N_20463,N_18486,N_18670);
nor U20464 (N_20464,N_19560,N_18374);
and U20465 (N_20465,N_19387,N_18862);
nand U20466 (N_20466,N_19496,N_18909);
xnor U20467 (N_20467,N_19966,N_19074);
nand U20468 (N_20468,N_19603,N_18073);
or U20469 (N_20469,N_18281,N_18026);
xor U20470 (N_20470,N_19086,N_19045);
or U20471 (N_20471,N_18920,N_18309);
or U20472 (N_20472,N_18323,N_19437);
nand U20473 (N_20473,N_19512,N_18548);
nand U20474 (N_20474,N_19250,N_18581);
nor U20475 (N_20475,N_19650,N_18530);
nor U20476 (N_20476,N_19162,N_18981);
nor U20477 (N_20477,N_19172,N_19725);
and U20478 (N_20478,N_19774,N_19103);
nor U20479 (N_20479,N_18913,N_19362);
or U20480 (N_20480,N_18567,N_19562);
nor U20481 (N_20481,N_18728,N_18100);
nor U20482 (N_20482,N_19001,N_19077);
nor U20483 (N_20483,N_19696,N_19402);
nand U20484 (N_20484,N_18591,N_19310);
and U20485 (N_20485,N_18628,N_19488);
xnor U20486 (N_20486,N_18998,N_18519);
nor U20487 (N_20487,N_19973,N_19497);
nor U20488 (N_20488,N_18593,N_19531);
nor U20489 (N_20489,N_19674,N_19913);
or U20490 (N_20490,N_18704,N_18314);
nand U20491 (N_20491,N_18239,N_18284);
nand U20492 (N_20492,N_18690,N_19083);
nand U20493 (N_20493,N_18191,N_19269);
nand U20494 (N_20494,N_19240,N_18922);
nand U20495 (N_20495,N_19303,N_19818);
or U20496 (N_20496,N_18419,N_18082);
nand U20497 (N_20497,N_18580,N_19844);
or U20498 (N_20498,N_19315,N_19516);
xnor U20499 (N_20499,N_18166,N_19431);
nand U20500 (N_20500,N_18829,N_19536);
nor U20501 (N_20501,N_19153,N_19870);
or U20502 (N_20502,N_18538,N_18512);
nor U20503 (N_20503,N_18290,N_19722);
and U20504 (N_20504,N_18152,N_19565);
nor U20505 (N_20505,N_19545,N_18189);
or U20506 (N_20506,N_18168,N_19044);
nor U20507 (N_20507,N_19780,N_18163);
or U20508 (N_20508,N_19628,N_19082);
and U20509 (N_20509,N_18383,N_18178);
and U20510 (N_20510,N_19850,N_18187);
and U20511 (N_20511,N_18090,N_18603);
xnor U20512 (N_20512,N_18904,N_18351);
xor U20513 (N_20513,N_19136,N_18735);
nand U20514 (N_20514,N_18169,N_19656);
xnor U20515 (N_20515,N_19971,N_19606);
nor U20516 (N_20516,N_18144,N_19967);
and U20517 (N_20517,N_18556,N_19569);
or U20518 (N_20518,N_19746,N_18227);
and U20519 (N_20519,N_19701,N_18148);
or U20520 (N_20520,N_19663,N_19687);
or U20521 (N_20521,N_19371,N_18707);
nand U20522 (N_20522,N_19349,N_18212);
or U20523 (N_20523,N_18855,N_18529);
and U20524 (N_20524,N_18229,N_18621);
and U20525 (N_20525,N_19544,N_19015);
xor U20526 (N_20526,N_19113,N_19325);
xor U20527 (N_20527,N_19671,N_19333);
nand U20528 (N_20528,N_19189,N_19256);
or U20529 (N_20529,N_19524,N_18029);
nor U20530 (N_20530,N_18818,N_19673);
xor U20531 (N_20531,N_19727,N_18988);
xnor U20532 (N_20532,N_19003,N_19734);
and U20533 (N_20533,N_18740,N_18546);
or U20534 (N_20534,N_19006,N_18207);
and U20535 (N_20535,N_18268,N_19415);
and U20536 (N_20536,N_18088,N_19794);
nand U20537 (N_20537,N_18746,N_19200);
nand U20538 (N_20538,N_18426,N_18371);
xor U20539 (N_20539,N_18000,N_18083);
nand U20540 (N_20540,N_19867,N_19283);
nand U20541 (N_20541,N_19119,N_19118);
nand U20542 (N_20542,N_18859,N_18636);
nor U20543 (N_20543,N_18398,N_19463);
nor U20544 (N_20544,N_18678,N_19493);
and U20545 (N_20545,N_19709,N_18058);
nor U20546 (N_20546,N_19337,N_18219);
or U20547 (N_20547,N_19284,N_19731);
and U20548 (N_20548,N_19904,N_18885);
xnor U20549 (N_20549,N_18102,N_19023);
or U20550 (N_20550,N_18217,N_19213);
nand U20551 (N_20551,N_19934,N_19385);
nor U20552 (N_20552,N_18839,N_19520);
xnor U20553 (N_20553,N_18298,N_19801);
or U20554 (N_20554,N_19114,N_19174);
nand U20555 (N_20555,N_19221,N_19330);
xnor U20556 (N_20556,N_19600,N_19651);
nor U20557 (N_20557,N_18941,N_18172);
xor U20558 (N_20558,N_18967,N_19233);
nand U20559 (N_20559,N_18161,N_18867);
nor U20560 (N_20560,N_19299,N_18450);
or U20561 (N_20561,N_18900,N_18850);
or U20562 (N_20562,N_18602,N_18644);
xnor U20563 (N_20563,N_18844,N_19008);
xnor U20564 (N_20564,N_19582,N_18022);
nor U20565 (N_20565,N_18089,N_19707);
xor U20566 (N_20566,N_19509,N_18645);
nor U20567 (N_20567,N_18362,N_18366);
xor U20568 (N_20568,N_19454,N_18074);
xnor U20569 (N_20569,N_18686,N_19438);
nand U20570 (N_20570,N_18347,N_18359);
nand U20571 (N_20571,N_18797,N_19945);
nand U20572 (N_20572,N_18213,N_18379);
nor U20573 (N_20573,N_18205,N_19207);
nor U20574 (N_20574,N_19579,N_18078);
and U20575 (N_20575,N_19997,N_18435);
nor U20576 (N_20576,N_19720,N_19383);
nor U20577 (N_20577,N_18010,N_18802);
and U20578 (N_20578,N_19682,N_19938);
or U20579 (N_20579,N_19700,N_19853);
and U20580 (N_20580,N_18692,N_19021);
or U20581 (N_20581,N_18717,N_19106);
or U20582 (N_20582,N_19314,N_18157);
nor U20583 (N_20583,N_18246,N_19048);
or U20584 (N_20584,N_19107,N_19447);
xnor U20585 (N_20585,N_19583,N_19643);
nand U20586 (N_20586,N_18793,N_18892);
xnor U20587 (N_20587,N_18522,N_18282);
nor U20588 (N_20588,N_19679,N_18253);
nor U20589 (N_20589,N_18415,N_19169);
nand U20590 (N_20590,N_18626,N_18782);
and U20591 (N_20591,N_19812,N_19829);
nor U20592 (N_20592,N_18293,N_18094);
nand U20593 (N_20593,N_18551,N_19936);
nand U20594 (N_20594,N_18437,N_19943);
or U20595 (N_20595,N_19588,N_18331);
and U20596 (N_20596,N_19838,N_19530);
nand U20597 (N_20597,N_18545,N_18154);
xor U20598 (N_20598,N_18416,N_19886);
and U20599 (N_20599,N_18123,N_18743);
xor U20600 (N_20600,N_19796,N_19576);
or U20601 (N_20601,N_19760,N_19040);
or U20602 (N_20602,N_18596,N_18675);
or U20603 (N_20603,N_18995,N_18910);
nor U20604 (N_20604,N_19750,N_18804);
or U20605 (N_20605,N_19181,N_18376);
xor U20606 (N_20606,N_18700,N_18440);
xnor U20607 (N_20607,N_19210,N_18992);
nor U20608 (N_20608,N_18077,N_19666);
and U20609 (N_20609,N_18150,N_19448);
nand U20610 (N_20610,N_18638,N_19302);
xnor U20611 (N_20611,N_18781,N_18075);
xnor U20612 (N_20612,N_19338,N_18906);
and U20613 (N_20613,N_18792,N_18196);
or U20614 (N_20614,N_18267,N_19799);
or U20615 (N_20615,N_18622,N_18139);
nand U20616 (N_20616,N_19964,N_18142);
xnor U20617 (N_20617,N_18847,N_19406);
xor U20618 (N_20618,N_19975,N_19553);
nand U20619 (N_20619,N_19815,N_19198);
and U20620 (N_20620,N_19436,N_18389);
xnor U20621 (N_20621,N_18957,N_19217);
and U20622 (N_20622,N_19061,N_19453);
or U20623 (N_20623,N_18285,N_18016);
nor U20624 (N_20624,N_18183,N_18516);
and U20625 (N_20625,N_18928,N_18587);
nand U20626 (N_20626,N_19173,N_18875);
nor U20627 (N_20627,N_19851,N_19394);
or U20628 (N_20628,N_19072,N_19043);
and U20629 (N_20629,N_19537,N_19068);
or U20630 (N_20630,N_18676,N_18226);
or U20631 (N_20631,N_19155,N_18276);
or U20632 (N_20632,N_18159,N_19130);
nand U20633 (N_20633,N_19836,N_18770);
or U20634 (N_20634,N_19708,N_19705);
and U20635 (N_20635,N_19704,N_18597);
xor U20636 (N_20636,N_18574,N_18714);
xor U20637 (N_20637,N_19592,N_19987);
xor U20638 (N_20638,N_19457,N_19028);
or U20639 (N_20639,N_18852,N_19423);
or U20640 (N_20640,N_19469,N_19053);
nand U20641 (N_20641,N_18475,N_18752);
xor U20642 (N_20642,N_19880,N_19322);
xnor U20643 (N_20643,N_19718,N_18076);
and U20644 (N_20644,N_19523,N_19291);
nand U20645 (N_20645,N_18766,N_19587);
nor U20646 (N_20646,N_18876,N_18958);
and U20647 (N_20647,N_18206,N_19465);
nor U20648 (N_20648,N_19102,N_19430);
xnor U20649 (N_20649,N_18965,N_18708);
or U20650 (N_20650,N_18762,N_19950);
xnor U20651 (N_20651,N_19782,N_18733);
and U20652 (N_20652,N_19626,N_18488);
and U20653 (N_20653,N_18821,N_19440);
or U20654 (N_20654,N_18629,N_19355);
nor U20655 (N_20655,N_19879,N_19388);
or U20656 (N_20656,N_18882,N_19797);
or U20657 (N_20657,N_18927,N_18028);
and U20658 (N_20658,N_18977,N_18916);
nor U20659 (N_20659,N_19783,N_19522);
xnor U20660 (N_20660,N_18251,N_19450);
nand U20661 (N_20661,N_18659,N_19563);
or U20662 (N_20662,N_18124,N_18683);
xor U20663 (N_20663,N_18441,N_19909);
nand U20664 (N_20664,N_18344,N_18571);
nor U20665 (N_20665,N_19393,N_19539);
or U20666 (N_20666,N_19776,N_19766);
nor U20667 (N_20667,N_18192,N_18697);
and U20668 (N_20668,N_19042,N_19259);
or U20669 (N_20669,N_18384,N_18059);
or U20670 (N_20670,N_18305,N_19948);
and U20671 (N_20671,N_19961,N_18071);
nand U20672 (N_20672,N_19505,N_18193);
xor U20673 (N_20673,N_18853,N_19641);
nand U20674 (N_20674,N_19639,N_19691);
xor U20675 (N_20675,N_18382,N_18444);
or U20676 (N_20676,N_18973,N_18849);
xor U20677 (N_20677,N_19548,N_19670);
or U20678 (N_20678,N_19847,N_19002);
nor U20679 (N_20679,N_19929,N_18710);
xnor U20680 (N_20680,N_19062,N_19826);
nor U20681 (N_20681,N_19069,N_18003);
nand U20682 (N_20682,N_18122,N_19733);
nor U20683 (N_20683,N_18091,N_18496);
or U20684 (N_20684,N_19395,N_19474);
and U20685 (N_20685,N_18202,N_19765);
and U20686 (N_20686,N_18476,N_19244);
nor U20687 (N_20687,N_19604,N_18948);
nor U20688 (N_20688,N_19176,N_18454);
or U20689 (N_20689,N_18863,N_19914);
xnor U20690 (N_20690,N_19059,N_19313);
and U20691 (N_20691,N_19920,N_18589);
nand U20692 (N_20692,N_19276,N_19648);
and U20693 (N_20693,N_18001,N_18555);
and U20694 (N_20694,N_18051,N_18056);
and U20695 (N_20695,N_19740,N_18241);
xor U20696 (N_20696,N_18550,N_19645);
nor U20697 (N_20697,N_18363,N_18951);
xnor U20698 (N_20698,N_18879,N_19894);
and U20699 (N_20699,N_18514,N_19823);
or U20700 (N_20700,N_18352,N_19164);
nor U20701 (N_20701,N_18259,N_19085);
or U20702 (N_20702,N_19012,N_19133);
nor U20703 (N_20703,N_19434,N_19446);
xnor U20704 (N_20704,N_19373,N_19817);
and U20705 (N_20705,N_18974,N_19940);
and U20706 (N_20706,N_18224,N_18634);
or U20707 (N_20707,N_19547,N_19690);
xnor U20708 (N_20708,N_18378,N_18533);
xor U20709 (N_20709,N_18817,N_18345);
and U20710 (N_20710,N_18790,N_19646);
nor U20711 (N_20711,N_18617,N_19152);
xor U20712 (N_20712,N_19526,N_19684);
nand U20713 (N_20713,N_19561,N_18772);
and U20714 (N_20714,N_18785,N_18099);
nand U20715 (N_20715,N_18354,N_19182);
xor U20716 (N_20716,N_18674,N_18984);
or U20717 (N_20717,N_18442,N_18015);
xor U20718 (N_20718,N_18275,N_18188);
and U20719 (N_20719,N_19855,N_19791);
xnor U20720 (N_20720,N_18115,N_18520);
nor U20721 (N_20721,N_19795,N_19479);
nand U20722 (N_20722,N_19218,N_19676);
nor U20723 (N_20723,N_18047,N_19507);
and U20724 (N_20724,N_18291,N_18871);
nand U20725 (N_20725,N_19672,N_19442);
xnor U20726 (N_20726,N_19140,N_18592);
or U20727 (N_20727,N_18897,N_19080);
nand U20728 (N_20728,N_18141,N_19873);
nand U20729 (N_20729,N_19575,N_19896);
xnor U20730 (N_20730,N_18297,N_18300);
xor U20731 (N_20731,N_19712,N_18754);
xnor U20732 (N_20732,N_19915,N_18044);
nor U20733 (N_20733,N_18024,N_19605);
nor U20734 (N_20734,N_19893,N_18112);
xnor U20735 (N_20735,N_18976,N_18657);
xor U20736 (N_20736,N_18872,N_18333);
and U20737 (N_20737,N_19998,N_19088);
nor U20738 (N_20738,N_19828,N_19589);
or U20739 (N_20739,N_18576,N_19202);
nor U20740 (N_20740,N_18130,N_18667);
nand U20741 (N_20741,N_19653,N_18921);
xor U20742 (N_20742,N_18731,N_19009);
nor U20743 (N_20743,N_19489,N_18296);
and U20744 (N_20744,N_18263,N_18348);
or U20745 (N_20745,N_19139,N_18375);
xnor U20746 (N_20746,N_19543,N_19024);
xnor U20747 (N_20747,N_19816,N_18822);
nor U20748 (N_20748,N_19278,N_19640);
and U20749 (N_20749,N_18572,N_19759);
or U20750 (N_20750,N_18515,N_18759);
nand U20751 (N_20751,N_19049,N_19364);
xnor U20752 (N_20752,N_18971,N_19986);
and U20753 (N_20753,N_19111,N_18067);
nand U20754 (N_20754,N_19336,N_19418);
nand U20755 (N_20755,N_19911,N_19188);
xor U20756 (N_20756,N_19286,N_18666);
and U20757 (N_20757,N_19027,N_18791);
or U20758 (N_20758,N_18877,N_19047);
nor U20759 (N_20759,N_19117,N_19556);
xor U20760 (N_20760,N_18449,N_18902);
and U20761 (N_20761,N_18247,N_18525);
or U20762 (N_20762,N_18014,N_18809);
nand U20763 (N_20763,N_18343,N_19154);
xor U20764 (N_20764,N_18221,N_18470);
and U20765 (N_20765,N_18234,N_19891);
or U20766 (N_20766,N_18949,N_18798);
and U20767 (N_20767,N_18749,N_19365);
and U20768 (N_20768,N_19699,N_19586);
nand U20769 (N_20769,N_19949,N_18240);
nor U20770 (N_20770,N_18526,N_19607);
nor U20771 (N_20771,N_19889,N_19594);
nand U20772 (N_20772,N_18966,N_18837);
and U20773 (N_20773,N_19863,N_19309);
xor U20774 (N_20774,N_19311,N_18590);
and U20775 (N_20775,N_19515,N_19145);
and U20776 (N_20776,N_19501,N_18531);
or U20777 (N_20777,N_19954,N_18566);
nor U20778 (N_20778,N_18584,N_19755);
and U20779 (N_20779,N_19983,N_18796);
nor U20780 (N_20780,N_19052,N_19804);
nor U20781 (N_20781,N_19609,N_18730);
or U20782 (N_20782,N_18825,N_18737);
nand U20783 (N_20783,N_18786,N_19356);
nand U20784 (N_20784,N_18606,N_18432);
nor U20785 (N_20785,N_18055,N_19290);
or U20786 (N_20786,N_19306,N_18578);
xor U20787 (N_20787,N_18443,N_19144);
and U20788 (N_20788,N_19476,N_18990);
nand U20789 (N_20789,N_18751,N_18494);
nand U20790 (N_20790,N_19599,N_18542);
nand U20791 (N_20791,N_19468,N_19557);
or U20792 (N_20792,N_19121,N_18756);
or U20793 (N_20793,N_19464,N_19347);
xor U20794 (N_20794,N_19620,N_18336);
nor U20795 (N_20795,N_19714,N_19326);
and U20796 (N_20796,N_19665,N_18646);
nor U20797 (N_20797,N_19820,N_18417);
and U20798 (N_20798,N_18473,N_18741);
or U20799 (N_20799,N_18652,N_19035);
or U20800 (N_20800,N_19452,N_19848);
nor U20801 (N_20801,N_18656,N_19458);
and U20802 (N_20802,N_18469,N_19786);
nand U20803 (N_20803,N_18319,N_19307);
nor U20804 (N_20804,N_18414,N_18911);
and U20805 (N_20805,N_18734,N_18405);
and U20806 (N_20806,N_18528,N_19578);
or U20807 (N_20807,N_19232,N_19726);
nor U20808 (N_20808,N_19884,N_18429);
xor U20809 (N_20809,N_18434,N_18327);
nor U20810 (N_20810,N_19112,N_19721);
and U20811 (N_20811,N_19013,N_19343);
or U20812 (N_20812,N_18611,N_19506);
or U20813 (N_20813,N_19484,N_18004);
nor U20814 (N_20814,N_18865,N_18564);
nor U20815 (N_20815,N_19196,N_19026);
or U20816 (N_20816,N_19257,N_18500);
nand U20817 (N_20817,N_19249,N_19346);
xor U20818 (N_20818,N_19841,N_19990);
nand U20819 (N_20819,N_18891,N_19944);
xor U20820 (N_20820,N_19183,N_18565);
nand U20821 (N_20821,N_19771,N_18668);
nand U20822 (N_20822,N_19433,N_19694);
or U20823 (N_20823,N_18065,N_18881);
or U20824 (N_20824,N_19265,N_19567);
or U20825 (N_20825,N_18508,N_18007);
nand U20826 (N_20826,N_18214,N_19090);
xnor U20827 (N_20827,N_19120,N_18993);
nand U20828 (N_20828,N_19491,N_19014);
and U20829 (N_20829,N_19601,N_19334);
nor U20830 (N_20830,N_18570,N_18833);
nand U20831 (N_20831,N_19839,N_18501);
or U20832 (N_20832,N_19821,N_18197);
nand U20833 (N_20833,N_18953,N_19979);
or U20834 (N_20834,N_18787,N_19046);
xor U20835 (N_20835,N_19066,N_19634);
nor U20836 (N_20836,N_18931,N_19016);
xnor U20837 (N_20837,N_19382,N_18502);
and U20838 (N_20838,N_19316,N_19101);
nand U20839 (N_20839,N_18304,N_18372);
xnor U20840 (N_20840,N_18409,N_18698);
xnor U20841 (N_20841,N_18779,N_19970);
nor U20842 (N_20842,N_19109,N_18665);
xnor U20843 (N_20843,N_18521,N_18681);
nor U20844 (N_20844,N_18121,N_18724);
xor U20845 (N_20845,N_19846,N_18407);
nor U20846 (N_20846,N_18680,N_18523);
nor U20847 (N_20847,N_19831,N_19116);
xnor U20848 (N_20848,N_18524,N_19262);
or U20849 (N_20849,N_18880,N_19933);
and U20850 (N_20850,N_18560,N_19602);
nor U20851 (N_20851,N_19293,N_18110);
xnor U20852 (N_20852,N_18198,N_18534);
xor U20853 (N_20853,N_19234,N_18552);
nor U20854 (N_20854,N_19211,N_18997);
xnor U20855 (N_20855,N_18775,N_18579);
nand U20856 (N_20856,N_18005,N_18819);
and U20857 (N_20857,N_18132,N_19963);
xnor U20858 (N_20858,N_19957,N_18544);
nor U20859 (N_20859,N_18895,N_19203);
or U20860 (N_20860,N_18716,N_18887);
nor U20861 (N_20861,N_18346,N_18153);
or U20862 (N_20862,N_18092,N_19631);
nand U20863 (N_20863,N_19289,N_18036);
and U20864 (N_20864,N_18149,N_19763);
nand U20865 (N_20865,N_18301,N_19168);
or U20866 (N_20866,N_19300,N_18283);
nor U20867 (N_20867,N_18032,N_18996);
nor U20868 (N_20868,N_19490,N_19032);
nor U20869 (N_20869,N_18184,N_18823);
or U20870 (N_20870,N_19852,N_18709);
nor U20871 (N_20871,N_18332,N_18358);
and U20872 (N_20872,N_18490,N_18097);
and U20873 (N_20873,N_19916,N_19917);
nand U20874 (N_20874,N_18983,N_19953);
xnor U20875 (N_20875,N_19739,N_18503);
and U20876 (N_20876,N_18052,N_18174);
nor U20877 (N_20877,N_18701,N_18594);
and U20878 (N_20878,N_18208,N_19339);
nor U20879 (N_20879,N_19910,N_18540);
or U20880 (N_20880,N_18277,N_18256);
xor U20881 (N_20881,N_19191,N_18222);
nand U20882 (N_20882,N_19199,N_18456);
nor U20883 (N_20883,N_19632,N_19668);
nand U20884 (N_20884,N_18937,N_19280);
or U20885 (N_20885,N_18959,N_18041);
and U20886 (N_20886,N_18127,N_19625);
or U20887 (N_20887,N_18328,N_18238);
nor U20888 (N_20888,N_18180,N_18421);
nor U20889 (N_20889,N_18478,N_19785);
and U20890 (N_20890,N_18641,N_18699);
and U20891 (N_20891,N_18081,N_19835);
xnor U20892 (N_20892,N_18388,N_18095);
nand U20893 (N_20893,N_19598,N_18377);
xnor U20894 (N_20894,N_19504,N_18317);
nor U20895 (N_20895,N_19542,N_18925);
and U20896 (N_20896,N_18195,N_18982);
nor U20897 (N_20897,N_19723,N_19494);
xor U20898 (N_20898,N_19470,N_19224);
xor U20899 (N_20899,N_19400,N_19729);
or U20900 (N_20900,N_19179,N_19788);
nand U20901 (N_20901,N_18087,N_19379);
nand U20902 (N_20902,N_18023,N_18098);
nand U20903 (N_20903,N_19421,N_19079);
nor U20904 (N_20904,N_19148,N_19295);
or U20905 (N_20905,N_18430,N_19031);
and U20906 (N_20906,N_18631,N_19824);
and U20907 (N_20907,N_18956,N_18385);
nor U20908 (N_20908,N_18682,N_19266);
xnor U20909 (N_20909,N_18093,N_19866);
or U20910 (N_20910,N_19742,N_18671);
xnor U20911 (N_20911,N_19854,N_19272);
xnor U20912 (N_20912,N_19881,N_19885);
nand U20913 (N_20913,N_18845,N_18033);
and U20914 (N_20914,N_19404,N_19396);
xnor U20915 (N_20915,N_18814,N_18079);
or U20916 (N_20916,N_19903,N_18215);
nor U20917 (N_20917,N_18060,N_18778);
or U20918 (N_20918,N_19251,N_19386);
xnor U20919 (N_20919,N_19197,N_18027);
nand U20920 (N_20920,N_19323,N_19105);
nor U20921 (N_20921,N_19492,N_19580);
and U20922 (N_20922,N_19661,N_19810);
nand U20923 (N_20923,N_18750,N_19363);
nand U20924 (N_20924,N_19110,N_18069);
and U20925 (N_20925,N_18706,N_19051);
nand U20926 (N_20926,N_19000,N_19550);
nor U20927 (N_20927,N_18780,N_18353);
or U20928 (N_20928,N_19754,N_18854);
xnor U20929 (N_20929,N_19435,N_18947);
nor U20930 (N_20930,N_19248,N_19519);
and U20931 (N_20931,N_18658,N_18046);
xor U20932 (N_20932,N_19798,N_19294);
and U20933 (N_20933,N_19941,N_19951);
nand U20934 (N_20934,N_18642,N_18451);
nand U20935 (N_20935,N_19955,N_19098);
or U20936 (N_20936,N_19581,N_18807);
nor U20937 (N_20937,N_19473,N_18203);
nor U20938 (N_20938,N_19683,N_18002);
or U20939 (N_20939,N_18933,N_19304);
xor U20940 (N_20940,N_18445,N_19540);
nand U20941 (N_20941,N_19360,N_19680);
xnor U20942 (N_20942,N_18649,N_18985);
xor U20943 (N_20943,N_19769,N_18801);
or U20944 (N_20944,N_18179,N_18919);
and U20945 (N_20945,N_19732,N_18063);
nor U20946 (N_20946,N_18249,N_18687);
nor U20947 (N_20947,N_18313,N_19514);
nand U20948 (N_20948,N_19455,N_19407);
nor U20949 (N_20949,N_18048,N_18387);
nor U20950 (N_20950,N_18038,N_19585);
xor U20951 (N_20951,N_18498,N_19247);
nand U20952 (N_20952,N_18758,N_19947);
or U20953 (N_20953,N_18654,N_18129);
or U20954 (N_20954,N_18315,N_19702);
or U20955 (N_20955,N_18830,N_19958);
and U20956 (N_20956,N_19156,N_18955);
nor U20957 (N_20957,N_18712,N_18230);
nor U20958 (N_20958,N_19125,N_18722);
xor U20959 (N_20959,N_19564,N_18455);
nand U20960 (N_20960,N_18462,N_19011);
nor U20961 (N_20961,N_19298,N_18261);
or U20962 (N_20962,N_18647,N_19984);
nor U20963 (N_20963,N_19513,N_18604);
nor U20964 (N_20964,N_19230,N_19253);
nand U20965 (N_20965,N_19005,N_18841);
or U20966 (N_20966,N_19180,N_18497);
or U20967 (N_20967,N_18237,N_19424);
and U20968 (N_20968,N_18254,N_19108);
or U20969 (N_20969,N_18294,N_18677);
xnor U20970 (N_20970,N_19416,N_18365);
and U20971 (N_20971,N_18252,N_18182);
xnor U20972 (N_20972,N_19258,N_18693);
and U20973 (N_20973,N_18639,N_18625);
nand U20974 (N_20974,N_18557,N_18978);
and U20975 (N_20975,N_18972,N_18050);
xor U20976 (N_20976,N_18066,N_19175);
nand U20977 (N_20977,N_18338,N_19992);
or U20978 (N_20978,N_19327,N_18908);
nand U20979 (N_20979,N_19212,N_19747);
nand U20980 (N_20980,N_18569,N_18431);
and U20981 (N_20981,N_19260,N_19039);
nand U20982 (N_20982,N_18559,N_18623);
xnor U20983 (N_20983,N_19792,N_18425);
nand U20984 (N_20984,N_18878,N_19925);
or U20985 (N_20985,N_19449,N_19159);
xnor U20986 (N_20986,N_18280,N_19946);
nand U20987 (N_20987,N_18648,N_18795);
xnor U20988 (N_20988,N_19518,N_19204);
and U20989 (N_20989,N_19020,N_18288);
or U20990 (N_20990,N_18433,N_18361);
or U20991 (N_20991,N_18663,N_19412);
or U20992 (N_20992,N_18505,N_18329);
nand U20993 (N_20993,N_19857,N_19287);
or U20994 (N_20994,N_18042,N_18761);
and U20995 (N_20995,N_19227,N_19328);
and U20996 (N_20996,N_19689,N_19503);
nand U20997 (N_20997,N_19751,N_19883);
xnor U20998 (N_20998,N_19055,N_18650);
and U20999 (N_20999,N_18613,N_19502);
xor U21000 (N_21000,N_19246,N_19433);
nand U21001 (N_21001,N_18876,N_19190);
nand U21002 (N_21002,N_19201,N_18486);
xnor U21003 (N_21003,N_19534,N_19095);
xnor U21004 (N_21004,N_19660,N_18492);
nand U21005 (N_21005,N_19531,N_19691);
and U21006 (N_21006,N_19778,N_18831);
or U21007 (N_21007,N_18811,N_18566);
nand U21008 (N_21008,N_19136,N_19870);
or U21009 (N_21009,N_18004,N_19750);
and U21010 (N_21010,N_19315,N_18544);
and U21011 (N_21011,N_18148,N_19621);
nand U21012 (N_21012,N_18461,N_19351);
nor U21013 (N_21013,N_19515,N_19811);
xor U21014 (N_21014,N_19616,N_19847);
and U21015 (N_21015,N_18862,N_19742);
nor U21016 (N_21016,N_19667,N_18966);
and U21017 (N_21017,N_18014,N_19613);
and U21018 (N_21018,N_19152,N_19977);
and U21019 (N_21019,N_19705,N_19584);
nor U21020 (N_21020,N_19680,N_18769);
nand U21021 (N_21021,N_18576,N_18236);
nor U21022 (N_21022,N_18518,N_18850);
or U21023 (N_21023,N_19103,N_19876);
nor U21024 (N_21024,N_18108,N_18330);
xnor U21025 (N_21025,N_18365,N_18414);
or U21026 (N_21026,N_19356,N_18527);
or U21027 (N_21027,N_18191,N_18455);
nor U21028 (N_21028,N_19710,N_18783);
nor U21029 (N_21029,N_19838,N_19974);
xnor U21030 (N_21030,N_18855,N_19551);
or U21031 (N_21031,N_19521,N_18920);
or U21032 (N_21032,N_18568,N_18037);
or U21033 (N_21033,N_18123,N_18523);
nand U21034 (N_21034,N_18123,N_19633);
or U21035 (N_21035,N_19209,N_18024);
nand U21036 (N_21036,N_19647,N_19901);
or U21037 (N_21037,N_18228,N_19545);
nor U21038 (N_21038,N_19266,N_18096);
or U21039 (N_21039,N_19704,N_18731);
nor U21040 (N_21040,N_19047,N_18058);
xnor U21041 (N_21041,N_19379,N_18753);
and U21042 (N_21042,N_18945,N_19818);
nand U21043 (N_21043,N_18761,N_18202);
nand U21044 (N_21044,N_19324,N_19923);
and U21045 (N_21045,N_18248,N_18058);
nor U21046 (N_21046,N_19189,N_18973);
and U21047 (N_21047,N_19145,N_19146);
xnor U21048 (N_21048,N_18365,N_19460);
or U21049 (N_21049,N_18254,N_19930);
xnor U21050 (N_21050,N_18579,N_18416);
xor U21051 (N_21051,N_18558,N_18863);
xor U21052 (N_21052,N_19271,N_19223);
nor U21053 (N_21053,N_18567,N_19959);
xor U21054 (N_21054,N_19681,N_18563);
nand U21055 (N_21055,N_18391,N_19886);
or U21056 (N_21056,N_18687,N_18828);
xnor U21057 (N_21057,N_18776,N_19563);
or U21058 (N_21058,N_19572,N_18209);
or U21059 (N_21059,N_19720,N_19074);
or U21060 (N_21060,N_18428,N_18502);
and U21061 (N_21061,N_18040,N_18436);
or U21062 (N_21062,N_18432,N_18552);
or U21063 (N_21063,N_19518,N_19582);
xnor U21064 (N_21064,N_18551,N_18285);
or U21065 (N_21065,N_18381,N_19950);
or U21066 (N_21066,N_18670,N_19169);
nand U21067 (N_21067,N_19738,N_19091);
nand U21068 (N_21068,N_18147,N_18372);
xnor U21069 (N_21069,N_18989,N_18828);
nor U21070 (N_21070,N_19822,N_18274);
nor U21071 (N_21071,N_19543,N_19027);
or U21072 (N_21072,N_19646,N_19671);
xor U21073 (N_21073,N_18891,N_19644);
xor U21074 (N_21074,N_19079,N_19334);
xor U21075 (N_21075,N_18038,N_19701);
or U21076 (N_21076,N_19658,N_19414);
and U21077 (N_21077,N_19795,N_18616);
xor U21078 (N_21078,N_18359,N_19484);
nand U21079 (N_21079,N_19709,N_19435);
nor U21080 (N_21080,N_19896,N_19373);
nor U21081 (N_21081,N_19860,N_19795);
and U21082 (N_21082,N_18856,N_18219);
or U21083 (N_21083,N_19787,N_19479);
or U21084 (N_21084,N_19474,N_19215);
nor U21085 (N_21085,N_19906,N_18802);
xor U21086 (N_21086,N_19822,N_19067);
nand U21087 (N_21087,N_19968,N_18931);
nand U21088 (N_21088,N_18758,N_18035);
xor U21089 (N_21089,N_19684,N_18709);
nor U21090 (N_21090,N_19557,N_19951);
nand U21091 (N_21091,N_18469,N_18969);
nand U21092 (N_21092,N_18489,N_18235);
nand U21093 (N_21093,N_18275,N_19650);
nand U21094 (N_21094,N_18883,N_19584);
or U21095 (N_21095,N_18734,N_19146);
xnor U21096 (N_21096,N_18362,N_18892);
or U21097 (N_21097,N_19729,N_19010);
or U21098 (N_21098,N_18536,N_19927);
and U21099 (N_21099,N_18125,N_18137);
xnor U21100 (N_21100,N_18849,N_19984);
nand U21101 (N_21101,N_19308,N_19953);
or U21102 (N_21102,N_18351,N_18468);
and U21103 (N_21103,N_18612,N_19413);
or U21104 (N_21104,N_18810,N_19771);
and U21105 (N_21105,N_18972,N_19671);
or U21106 (N_21106,N_19605,N_18517);
xor U21107 (N_21107,N_18582,N_19711);
nor U21108 (N_21108,N_18463,N_18720);
nand U21109 (N_21109,N_18494,N_19840);
and U21110 (N_21110,N_19274,N_18758);
nor U21111 (N_21111,N_19231,N_18467);
and U21112 (N_21112,N_19160,N_18718);
nor U21113 (N_21113,N_18479,N_18182);
nand U21114 (N_21114,N_19253,N_19371);
xor U21115 (N_21115,N_18285,N_18592);
xnor U21116 (N_21116,N_18224,N_19329);
nand U21117 (N_21117,N_18783,N_19555);
or U21118 (N_21118,N_19009,N_18415);
xor U21119 (N_21119,N_19342,N_18732);
and U21120 (N_21120,N_19086,N_18480);
nor U21121 (N_21121,N_19441,N_18332);
xor U21122 (N_21122,N_19696,N_19447);
or U21123 (N_21123,N_19288,N_19896);
or U21124 (N_21124,N_18875,N_19532);
xnor U21125 (N_21125,N_19928,N_18543);
xnor U21126 (N_21126,N_18046,N_18340);
or U21127 (N_21127,N_19454,N_18427);
and U21128 (N_21128,N_18822,N_18106);
xor U21129 (N_21129,N_18048,N_19234);
nor U21130 (N_21130,N_18038,N_18376);
and U21131 (N_21131,N_18431,N_18345);
or U21132 (N_21132,N_19662,N_19431);
or U21133 (N_21133,N_19933,N_18945);
and U21134 (N_21134,N_19304,N_19950);
nor U21135 (N_21135,N_19153,N_19137);
nand U21136 (N_21136,N_18287,N_19676);
xnor U21137 (N_21137,N_19828,N_19125);
or U21138 (N_21138,N_19612,N_18678);
or U21139 (N_21139,N_18995,N_18352);
and U21140 (N_21140,N_19057,N_18137);
and U21141 (N_21141,N_18329,N_19235);
xnor U21142 (N_21142,N_19213,N_19125);
or U21143 (N_21143,N_18824,N_19014);
xnor U21144 (N_21144,N_19506,N_19641);
nand U21145 (N_21145,N_18412,N_19119);
nand U21146 (N_21146,N_18863,N_18513);
xnor U21147 (N_21147,N_18675,N_18246);
nor U21148 (N_21148,N_19221,N_19777);
xor U21149 (N_21149,N_19753,N_18614);
nor U21150 (N_21150,N_18024,N_19109);
or U21151 (N_21151,N_19502,N_18893);
xnor U21152 (N_21152,N_18048,N_19035);
nand U21153 (N_21153,N_18242,N_19085);
nor U21154 (N_21154,N_19525,N_19840);
nor U21155 (N_21155,N_19412,N_19867);
or U21156 (N_21156,N_19886,N_19805);
nand U21157 (N_21157,N_18185,N_19358);
nand U21158 (N_21158,N_18109,N_19218);
or U21159 (N_21159,N_18386,N_19033);
or U21160 (N_21160,N_19916,N_18534);
or U21161 (N_21161,N_19766,N_18879);
xnor U21162 (N_21162,N_19524,N_18694);
and U21163 (N_21163,N_19968,N_18170);
or U21164 (N_21164,N_19391,N_18856);
nor U21165 (N_21165,N_19130,N_19115);
nand U21166 (N_21166,N_19071,N_19705);
and U21167 (N_21167,N_18340,N_18842);
nand U21168 (N_21168,N_19416,N_18030);
nand U21169 (N_21169,N_19486,N_18306);
and U21170 (N_21170,N_19264,N_18859);
xor U21171 (N_21171,N_19022,N_19023);
or U21172 (N_21172,N_18645,N_19133);
nor U21173 (N_21173,N_18648,N_18668);
nor U21174 (N_21174,N_19478,N_18842);
and U21175 (N_21175,N_18675,N_18572);
nor U21176 (N_21176,N_19393,N_18885);
xnor U21177 (N_21177,N_18212,N_18470);
nand U21178 (N_21178,N_18396,N_18638);
xor U21179 (N_21179,N_19179,N_19838);
and U21180 (N_21180,N_18089,N_18985);
or U21181 (N_21181,N_18319,N_19806);
xor U21182 (N_21182,N_19659,N_19343);
nand U21183 (N_21183,N_19176,N_19819);
and U21184 (N_21184,N_19037,N_19385);
nor U21185 (N_21185,N_18739,N_18895);
and U21186 (N_21186,N_18175,N_19966);
xor U21187 (N_21187,N_18205,N_18758);
and U21188 (N_21188,N_19377,N_19743);
nand U21189 (N_21189,N_19371,N_19784);
and U21190 (N_21190,N_19112,N_19900);
nand U21191 (N_21191,N_19904,N_18063);
and U21192 (N_21192,N_19874,N_18544);
and U21193 (N_21193,N_19680,N_19520);
or U21194 (N_21194,N_19461,N_18719);
xor U21195 (N_21195,N_18212,N_19916);
xnor U21196 (N_21196,N_18959,N_19023);
nor U21197 (N_21197,N_19768,N_19981);
xor U21198 (N_21198,N_19682,N_18425);
or U21199 (N_21199,N_19463,N_19646);
xor U21200 (N_21200,N_18601,N_18507);
xor U21201 (N_21201,N_19274,N_18527);
nand U21202 (N_21202,N_19516,N_19575);
nor U21203 (N_21203,N_19959,N_19474);
xor U21204 (N_21204,N_19618,N_18299);
nor U21205 (N_21205,N_19357,N_18693);
nor U21206 (N_21206,N_18076,N_19321);
xnor U21207 (N_21207,N_18387,N_19920);
or U21208 (N_21208,N_19861,N_19695);
nor U21209 (N_21209,N_18017,N_18121);
and U21210 (N_21210,N_18520,N_19348);
and U21211 (N_21211,N_18279,N_19034);
xnor U21212 (N_21212,N_19053,N_19118);
xnor U21213 (N_21213,N_18997,N_18154);
nor U21214 (N_21214,N_19385,N_18529);
nor U21215 (N_21215,N_19112,N_18487);
nor U21216 (N_21216,N_18154,N_19040);
xnor U21217 (N_21217,N_19180,N_19892);
nand U21218 (N_21218,N_19254,N_19276);
nand U21219 (N_21219,N_18216,N_18100);
nor U21220 (N_21220,N_18579,N_19143);
and U21221 (N_21221,N_18692,N_18412);
nand U21222 (N_21222,N_18110,N_19904);
nand U21223 (N_21223,N_19835,N_18048);
nand U21224 (N_21224,N_18043,N_18690);
nor U21225 (N_21225,N_18094,N_18047);
or U21226 (N_21226,N_19550,N_18460);
nor U21227 (N_21227,N_18489,N_18162);
nand U21228 (N_21228,N_18962,N_19144);
nand U21229 (N_21229,N_19447,N_19952);
or U21230 (N_21230,N_18946,N_18546);
nor U21231 (N_21231,N_19281,N_19610);
xnor U21232 (N_21232,N_19227,N_18354);
nand U21233 (N_21233,N_19694,N_19443);
xor U21234 (N_21234,N_18340,N_18308);
xnor U21235 (N_21235,N_19843,N_18809);
or U21236 (N_21236,N_19954,N_19815);
xor U21237 (N_21237,N_18425,N_19195);
nor U21238 (N_21238,N_18875,N_18972);
and U21239 (N_21239,N_18159,N_18061);
nand U21240 (N_21240,N_18490,N_18109);
nand U21241 (N_21241,N_19181,N_18674);
and U21242 (N_21242,N_19208,N_19201);
xnor U21243 (N_21243,N_19633,N_18542);
or U21244 (N_21244,N_18431,N_18802);
xnor U21245 (N_21245,N_18043,N_19613);
or U21246 (N_21246,N_19410,N_18020);
nor U21247 (N_21247,N_19532,N_18124);
or U21248 (N_21248,N_18119,N_18390);
and U21249 (N_21249,N_19939,N_19554);
and U21250 (N_21250,N_19533,N_19344);
xnor U21251 (N_21251,N_18891,N_19819);
xnor U21252 (N_21252,N_18724,N_19042);
nand U21253 (N_21253,N_18369,N_18915);
and U21254 (N_21254,N_18328,N_19501);
and U21255 (N_21255,N_19824,N_19447);
and U21256 (N_21256,N_18974,N_18500);
and U21257 (N_21257,N_19538,N_19733);
nor U21258 (N_21258,N_19927,N_18726);
and U21259 (N_21259,N_19872,N_19480);
nor U21260 (N_21260,N_19771,N_19766);
nor U21261 (N_21261,N_19940,N_18592);
nand U21262 (N_21262,N_19632,N_18533);
nand U21263 (N_21263,N_18272,N_19199);
nor U21264 (N_21264,N_19860,N_18781);
and U21265 (N_21265,N_18485,N_18340);
xnor U21266 (N_21266,N_19383,N_18092);
or U21267 (N_21267,N_18190,N_18612);
and U21268 (N_21268,N_18270,N_19042);
or U21269 (N_21269,N_18736,N_18460);
xnor U21270 (N_21270,N_18967,N_18885);
or U21271 (N_21271,N_18369,N_18967);
or U21272 (N_21272,N_18840,N_19899);
and U21273 (N_21273,N_19140,N_18035);
nor U21274 (N_21274,N_19912,N_19793);
xor U21275 (N_21275,N_18751,N_18514);
and U21276 (N_21276,N_18078,N_18058);
xnor U21277 (N_21277,N_19659,N_18722);
or U21278 (N_21278,N_19878,N_19957);
or U21279 (N_21279,N_18958,N_19109);
xnor U21280 (N_21280,N_18819,N_18262);
and U21281 (N_21281,N_19936,N_18102);
nand U21282 (N_21282,N_19856,N_18732);
or U21283 (N_21283,N_18452,N_18754);
nand U21284 (N_21284,N_18552,N_19226);
nand U21285 (N_21285,N_18353,N_19169);
nor U21286 (N_21286,N_18821,N_18368);
nand U21287 (N_21287,N_18439,N_19175);
xor U21288 (N_21288,N_19897,N_19949);
nand U21289 (N_21289,N_19984,N_18934);
nor U21290 (N_21290,N_18761,N_19132);
and U21291 (N_21291,N_19138,N_18902);
nor U21292 (N_21292,N_18297,N_18118);
or U21293 (N_21293,N_18836,N_19067);
nor U21294 (N_21294,N_19684,N_18433);
and U21295 (N_21295,N_18855,N_19853);
and U21296 (N_21296,N_18566,N_18561);
nand U21297 (N_21297,N_18806,N_19633);
nor U21298 (N_21298,N_19302,N_19460);
nor U21299 (N_21299,N_19998,N_19875);
nor U21300 (N_21300,N_19947,N_18823);
or U21301 (N_21301,N_19206,N_19659);
nor U21302 (N_21302,N_18280,N_19760);
or U21303 (N_21303,N_18192,N_19555);
xor U21304 (N_21304,N_19640,N_19492);
xor U21305 (N_21305,N_18578,N_19337);
nor U21306 (N_21306,N_19534,N_18427);
or U21307 (N_21307,N_19948,N_19736);
xor U21308 (N_21308,N_18933,N_18588);
xnor U21309 (N_21309,N_19940,N_19312);
nand U21310 (N_21310,N_18868,N_18049);
and U21311 (N_21311,N_18233,N_19591);
and U21312 (N_21312,N_18873,N_18216);
xor U21313 (N_21313,N_18528,N_18137);
nand U21314 (N_21314,N_19835,N_19863);
xor U21315 (N_21315,N_18371,N_18779);
xnor U21316 (N_21316,N_18780,N_19927);
or U21317 (N_21317,N_18658,N_18547);
nand U21318 (N_21318,N_19811,N_19012);
or U21319 (N_21319,N_19227,N_18848);
xnor U21320 (N_21320,N_18988,N_18514);
nor U21321 (N_21321,N_19594,N_18386);
and U21322 (N_21322,N_18247,N_18415);
and U21323 (N_21323,N_19732,N_18587);
nand U21324 (N_21324,N_19675,N_19158);
nor U21325 (N_21325,N_18723,N_19667);
and U21326 (N_21326,N_19288,N_19141);
nand U21327 (N_21327,N_18429,N_18464);
nor U21328 (N_21328,N_18554,N_18969);
xor U21329 (N_21329,N_18700,N_19390);
or U21330 (N_21330,N_19425,N_19998);
or U21331 (N_21331,N_18713,N_18065);
or U21332 (N_21332,N_18327,N_18606);
nor U21333 (N_21333,N_18058,N_18765);
and U21334 (N_21334,N_18342,N_18911);
and U21335 (N_21335,N_19387,N_18908);
nor U21336 (N_21336,N_18847,N_19414);
or U21337 (N_21337,N_19035,N_19488);
or U21338 (N_21338,N_18679,N_18270);
xor U21339 (N_21339,N_18395,N_19338);
nand U21340 (N_21340,N_18161,N_18951);
nand U21341 (N_21341,N_19404,N_18921);
nand U21342 (N_21342,N_19639,N_18218);
or U21343 (N_21343,N_19049,N_18702);
or U21344 (N_21344,N_19295,N_18525);
xor U21345 (N_21345,N_18658,N_18417);
nor U21346 (N_21346,N_19233,N_19764);
or U21347 (N_21347,N_19839,N_18936);
xor U21348 (N_21348,N_18267,N_19544);
nand U21349 (N_21349,N_18193,N_18981);
nand U21350 (N_21350,N_18222,N_19930);
xnor U21351 (N_21351,N_19472,N_18689);
or U21352 (N_21352,N_18254,N_18699);
xnor U21353 (N_21353,N_19717,N_18006);
or U21354 (N_21354,N_18585,N_18371);
or U21355 (N_21355,N_19003,N_18084);
or U21356 (N_21356,N_19926,N_18528);
nor U21357 (N_21357,N_19866,N_19241);
nor U21358 (N_21358,N_19967,N_19325);
xor U21359 (N_21359,N_18355,N_18510);
xor U21360 (N_21360,N_18446,N_19529);
xnor U21361 (N_21361,N_19069,N_19679);
and U21362 (N_21362,N_19542,N_19082);
xnor U21363 (N_21363,N_19242,N_18198);
xor U21364 (N_21364,N_18891,N_19586);
or U21365 (N_21365,N_19809,N_19425);
nor U21366 (N_21366,N_19133,N_19987);
or U21367 (N_21367,N_18978,N_19650);
and U21368 (N_21368,N_19847,N_19574);
nand U21369 (N_21369,N_19445,N_18161);
or U21370 (N_21370,N_18615,N_19903);
and U21371 (N_21371,N_19610,N_19421);
nor U21372 (N_21372,N_19946,N_19262);
nand U21373 (N_21373,N_18904,N_19546);
or U21374 (N_21374,N_18730,N_18754);
nor U21375 (N_21375,N_19209,N_19503);
nand U21376 (N_21376,N_18479,N_19926);
nand U21377 (N_21377,N_19696,N_18162);
xor U21378 (N_21378,N_18106,N_19687);
nand U21379 (N_21379,N_18264,N_19198);
and U21380 (N_21380,N_18494,N_19392);
xor U21381 (N_21381,N_18646,N_19156);
xor U21382 (N_21382,N_19016,N_18646);
xnor U21383 (N_21383,N_18822,N_18757);
or U21384 (N_21384,N_19653,N_19473);
nand U21385 (N_21385,N_18523,N_19289);
and U21386 (N_21386,N_19004,N_18095);
and U21387 (N_21387,N_18880,N_18847);
or U21388 (N_21388,N_18263,N_18999);
and U21389 (N_21389,N_18733,N_19432);
nor U21390 (N_21390,N_19857,N_19426);
nor U21391 (N_21391,N_19814,N_19456);
nor U21392 (N_21392,N_19976,N_18340);
nand U21393 (N_21393,N_19428,N_19050);
xor U21394 (N_21394,N_18650,N_19164);
or U21395 (N_21395,N_19220,N_18913);
or U21396 (N_21396,N_18684,N_18368);
nand U21397 (N_21397,N_19610,N_19828);
xor U21398 (N_21398,N_19079,N_18846);
nand U21399 (N_21399,N_18188,N_19139);
and U21400 (N_21400,N_18084,N_18983);
nor U21401 (N_21401,N_19810,N_18976);
and U21402 (N_21402,N_18980,N_19788);
or U21403 (N_21403,N_18807,N_18366);
and U21404 (N_21404,N_18908,N_19883);
xor U21405 (N_21405,N_19693,N_19072);
xnor U21406 (N_21406,N_18808,N_19102);
or U21407 (N_21407,N_19155,N_19294);
and U21408 (N_21408,N_18185,N_19546);
nor U21409 (N_21409,N_18917,N_18808);
xor U21410 (N_21410,N_19093,N_18361);
and U21411 (N_21411,N_19348,N_19956);
and U21412 (N_21412,N_19518,N_19756);
nand U21413 (N_21413,N_19190,N_19293);
nand U21414 (N_21414,N_19828,N_18477);
or U21415 (N_21415,N_18448,N_18678);
or U21416 (N_21416,N_18172,N_19588);
nor U21417 (N_21417,N_18823,N_19045);
nand U21418 (N_21418,N_18620,N_19701);
nand U21419 (N_21419,N_19210,N_19435);
or U21420 (N_21420,N_19203,N_18371);
xor U21421 (N_21421,N_18748,N_18754);
and U21422 (N_21422,N_18927,N_18347);
or U21423 (N_21423,N_19601,N_19289);
or U21424 (N_21424,N_18046,N_19901);
nand U21425 (N_21425,N_18468,N_19576);
nand U21426 (N_21426,N_18726,N_18465);
xnor U21427 (N_21427,N_19364,N_19509);
xor U21428 (N_21428,N_19464,N_18187);
xor U21429 (N_21429,N_19346,N_18831);
or U21430 (N_21430,N_18663,N_18566);
or U21431 (N_21431,N_19694,N_19876);
and U21432 (N_21432,N_19411,N_18403);
nor U21433 (N_21433,N_18570,N_18794);
and U21434 (N_21434,N_18657,N_18705);
or U21435 (N_21435,N_19761,N_18299);
nand U21436 (N_21436,N_19401,N_19710);
and U21437 (N_21437,N_18199,N_19678);
nor U21438 (N_21438,N_18596,N_18794);
nor U21439 (N_21439,N_18226,N_19324);
or U21440 (N_21440,N_19733,N_18612);
nor U21441 (N_21441,N_18355,N_19417);
xnor U21442 (N_21442,N_18176,N_19247);
xnor U21443 (N_21443,N_19673,N_18099);
xnor U21444 (N_21444,N_18699,N_18098);
or U21445 (N_21445,N_18650,N_18798);
and U21446 (N_21446,N_18202,N_19950);
and U21447 (N_21447,N_19797,N_18557);
and U21448 (N_21448,N_19971,N_19862);
or U21449 (N_21449,N_18341,N_19750);
xnor U21450 (N_21450,N_18723,N_18359);
xnor U21451 (N_21451,N_18276,N_18467);
and U21452 (N_21452,N_19582,N_18936);
nand U21453 (N_21453,N_18371,N_19397);
nor U21454 (N_21454,N_19563,N_18899);
nor U21455 (N_21455,N_19905,N_19605);
or U21456 (N_21456,N_19530,N_18693);
or U21457 (N_21457,N_19940,N_18295);
and U21458 (N_21458,N_18315,N_18351);
and U21459 (N_21459,N_19793,N_19867);
and U21460 (N_21460,N_19085,N_18026);
or U21461 (N_21461,N_18541,N_18646);
xnor U21462 (N_21462,N_19509,N_19010);
nand U21463 (N_21463,N_18617,N_18814);
nand U21464 (N_21464,N_18647,N_18421);
or U21465 (N_21465,N_19625,N_19109);
xor U21466 (N_21466,N_18681,N_18694);
and U21467 (N_21467,N_19167,N_18852);
xnor U21468 (N_21468,N_18208,N_19166);
xnor U21469 (N_21469,N_18843,N_18507);
nand U21470 (N_21470,N_18552,N_18705);
xor U21471 (N_21471,N_18240,N_18795);
nand U21472 (N_21472,N_18698,N_19404);
nand U21473 (N_21473,N_18300,N_18866);
nor U21474 (N_21474,N_18916,N_18741);
or U21475 (N_21475,N_18190,N_18930);
nand U21476 (N_21476,N_19602,N_18194);
and U21477 (N_21477,N_18450,N_18986);
nand U21478 (N_21478,N_19708,N_18416);
nand U21479 (N_21479,N_18968,N_19913);
nor U21480 (N_21480,N_19379,N_19516);
or U21481 (N_21481,N_19007,N_19332);
and U21482 (N_21482,N_18160,N_19147);
nand U21483 (N_21483,N_19094,N_19724);
xnor U21484 (N_21484,N_18582,N_18137);
nor U21485 (N_21485,N_19265,N_18110);
nand U21486 (N_21486,N_18669,N_19825);
nand U21487 (N_21487,N_18683,N_18728);
or U21488 (N_21488,N_18307,N_18830);
or U21489 (N_21489,N_19572,N_18004);
and U21490 (N_21490,N_19965,N_18139);
or U21491 (N_21491,N_19355,N_19049);
nor U21492 (N_21492,N_18613,N_18836);
and U21493 (N_21493,N_19619,N_19189);
and U21494 (N_21494,N_18524,N_19964);
and U21495 (N_21495,N_19486,N_18904);
nor U21496 (N_21496,N_18056,N_19569);
and U21497 (N_21497,N_18771,N_19511);
nand U21498 (N_21498,N_19749,N_18223);
or U21499 (N_21499,N_19432,N_19213);
or U21500 (N_21500,N_19231,N_18026);
nor U21501 (N_21501,N_18769,N_19005);
nor U21502 (N_21502,N_19983,N_18095);
and U21503 (N_21503,N_19348,N_19285);
nand U21504 (N_21504,N_19170,N_19959);
and U21505 (N_21505,N_19856,N_19811);
nor U21506 (N_21506,N_18715,N_19974);
and U21507 (N_21507,N_19734,N_18132);
xor U21508 (N_21508,N_18313,N_18302);
and U21509 (N_21509,N_19511,N_19412);
xnor U21510 (N_21510,N_19677,N_19914);
xor U21511 (N_21511,N_19474,N_19450);
nor U21512 (N_21512,N_18765,N_18998);
and U21513 (N_21513,N_19797,N_18831);
nand U21514 (N_21514,N_19636,N_18641);
nor U21515 (N_21515,N_18320,N_19717);
nor U21516 (N_21516,N_19260,N_19949);
nand U21517 (N_21517,N_19577,N_18335);
nor U21518 (N_21518,N_19668,N_18365);
nor U21519 (N_21519,N_18230,N_18542);
and U21520 (N_21520,N_19082,N_19367);
or U21521 (N_21521,N_18793,N_19054);
and U21522 (N_21522,N_18531,N_19654);
or U21523 (N_21523,N_19735,N_19631);
and U21524 (N_21524,N_19156,N_19708);
nor U21525 (N_21525,N_19497,N_19832);
or U21526 (N_21526,N_18733,N_19813);
nand U21527 (N_21527,N_18636,N_19289);
nand U21528 (N_21528,N_18608,N_18209);
xor U21529 (N_21529,N_19780,N_19892);
nor U21530 (N_21530,N_19792,N_19806);
nor U21531 (N_21531,N_18439,N_19216);
nand U21532 (N_21532,N_18606,N_18317);
or U21533 (N_21533,N_18590,N_18592);
nand U21534 (N_21534,N_18721,N_18327);
nand U21535 (N_21535,N_19706,N_18863);
or U21536 (N_21536,N_19197,N_19320);
nor U21537 (N_21537,N_18050,N_19731);
nand U21538 (N_21538,N_18065,N_18718);
and U21539 (N_21539,N_18553,N_18885);
xor U21540 (N_21540,N_18575,N_18188);
and U21541 (N_21541,N_19728,N_19823);
and U21542 (N_21542,N_18815,N_18241);
nor U21543 (N_21543,N_18305,N_18823);
nor U21544 (N_21544,N_19287,N_18998);
nor U21545 (N_21545,N_19320,N_19347);
or U21546 (N_21546,N_19106,N_19457);
and U21547 (N_21547,N_19549,N_19732);
and U21548 (N_21548,N_19639,N_19919);
and U21549 (N_21549,N_18794,N_19473);
nand U21550 (N_21550,N_18209,N_19618);
or U21551 (N_21551,N_19060,N_19452);
nor U21552 (N_21552,N_18289,N_18364);
nand U21553 (N_21553,N_18847,N_18434);
nand U21554 (N_21554,N_19304,N_19456);
or U21555 (N_21555,N_18056,N_19473);
xnor U21556 (N_21556,N_18809,N_18617);
nand U21557 (N_21557,N_18954,N_18751);
or U21558 (N_21558,N_19562,N_18745);
or U21559 (N_21559,N_19299,N_18843);
xor U21560 (N_21560,N_18194,N_19841);
or U21561 (N_21561,N_19285,N_19913);
and U21562 (N_21562,N_19084,N_18991);
nor U21563 (N_21563,N_18054,N_19987);
nand U21564 (N_21564,N_18577,N_19059);
xor U21565 (N_21565,N_18673,N_18772);
or U21566 (N_21566,N_19057,N_19688);
or U21567 (N_21567,N_18797,N_18548);
nor U21568 (N_21568,N_18659,N_19964);
nand U21569 (N_21569,N_18744,N_18767);
xnor U21570 (N_21570,N_18209,N_18670);
or U21571 (N_21571,N_19597,N_18329);
xor U21572 (N_21572,N_18112,N_19258);
nand U21573 (N_21573,N_18191,N_18142);
nor U21574 (N_21574,N_19093,N_18970);
nor U21575 (N_21575,N_19193,N_18091);
nand U21576 (N_21576,N_19347,N_19276);
and U21577 (N_21577,N_19205,N_18382);
xnor U21578 (N_21578,N_19502,N_19898);
or U21579 (N_21579,N_19771,N_19292);
nand U21580 (N_21580,N_19499,N_18838);
nor U21581 (N_21581,N_19530,N_18312);
and U21582 (N_21582,N_18258,N_18120);
xnor U21583 (N_21583,N_18084,N_18553);
nand U21584 (N_21584,N_18629,N_18531);
and U21585 (N_21585,N_19371,N_18786);
or U21586 (N_21586,N_18551,N_18035);
xor U21587 (N_21587,N_19712,N_19177);
or U21588 (N_21588,N_18674,N_18312);
nand U21589 (N_21589,N_18203,N_19190);
nor U21590 (N_21590,N_18605,N_18729);
xnor U21591 (N_21591,N_18319,N_18542);
xor U21592 (N_21592,N_19152,N_19407);
or U21593 (N_21593,N_18275,N_19845);
and U21594 (N_21594,N_19859,N_19351);
xnor U21595 (N_21595,N_18071,N_18580);
and U21596 (N_21596,N_18617,N_18006);
xnor U21597 (N_21597,N_19865,N_18608);
nand U21598 (N_21598,N_19320,N_19896);
and U21599 (N_21599,N_18264,N_19290);
nor U21600 (N_21600,N_18899,N_18240);
and U21601 (N_21601,N_19543,N_19401);
and U21602 (N_21602,N_18588,N_18790);
nor U21603 (N_21603,N_19533,N_18144);
or U21604 (N_21604,N_18046,N_19522);
nor U21605 (N_21605,N_18969,N_19257);
nand U21606 (N_21606,N_18901,N_19521);
xnor U21607 (N_21607,N_19083,N_19884);
and U21608 (N_21608,N_18582,N_19355);
xor U21609 (N_21609,N_18651,N_19397);
and U21610 (N_21610,N_19079,N_18147);
and U21611 (N_21611,N_18187,N_18244);
nand U21612 (N_21612,N_18622,N_18384);
nand U21613 (N_21613,N_18820,N_18652);
and U21614 (N_21614,N_19929,N_19055);
or U21615 (N_21615,N_19327,N_19953);
and U21616 (N_21616,N_18286,N_18546);
or U21617 (N_21617,N_18286,N_19857);
nand U21618 (N_21618,N_18229,N_18304);
or U21619 (N_21619,N_19473,N_18197);
nand U21620 (N_21620,N_18792,N_19622);
and U21621 (N_21621,N_19172,N_18207);
and U21622 (N_21622,N_19495,N_18675);
and U21623 (N_21623,N_18585,N_18081);
nor U21624 (N_21624,N_18949,N_19925);
nand U21625 (N_21625,N_18574,N_18744);
nor U21626 (N_21626,N_19757,N_19164);
or U21627 (N_21627,N_19188,N_19122);
nor U21628 (N_21628,N_18197,N_19461);
or U21629 (N_21629,N_19724,N_18431);
nor U21630 (N_21630,N_18989,N_18518);
nand U21631 (N_21631,N_19934,N_18788);
or U21632 (N_21632,N_19480,N_19591);
or U21633 (N_21633,N_18863,N_18877);
nand U21634 (N_21634,N_19405,N_18479);
and U21635 (N_21635,N_19267,N_18064);
xnor U21636 (N_21636,N_19657,N_19846);
or U21637 (N_21637,N_18400,N_18371);
xnor U21638 (N_21638,N_18126,N_19675);
xnor U21639 (N_21639,N_19412,N_19658);
or U21640 (N_21640,N_19937,N_19486);
or U21641 (N_21641,N_18898,N_18161);
nand U21642 (N_21642,N_19724,N_18533);
and U21643 (N_21643,N_19109,N_19952);
and U21644 (N_21644,N_19318,N_18627);
and U21645 (N_21645,N_18284,N_19203);
nand U21646 (N_21646,N_19248,N_18525);
xnor U21647 (N_21647,N_18660,N_18408);
nor U21648 (N_21648,N_19822,N_19495);
nand U21649 (N_21649,N_19615,N_18804);
nor U21650 (N_21650,N_18771,N_19575);
and U21651 (N_21651,N_19948,N_19995);
nor U21652 (N_21652,N_19261,N_18009);
nand U21653 (N_21653,N_18033,N_19987);
xor U21654 (N_21654,N_18842,N_19390);
xnor U21655 (N_21655,N_19114,N_19635);
xor U21656 (N_21656,N_18089,N_18229);
or U21657 (N_21657,N_19506,N_18103);
nand U21658 (N_21658,N_18882,N_18577);
nand U21659 (N_21659,N_19980,N_18619);
nor U21660 (N_21660,N_19956,N_19662);
and U21661 (N_21661,N_19382,N_19573);
nand U21662 (N_21662,N_19811,N_18707);
and U21663 (N_21663,N_19391,N_18704);
nor U21664 (N_21664,N_19532,N_19984);
xnor U21665 (N_21665,N_19980,N_18256);
or U21666 (N_21666,N_19400,N_18366);
and U21667 (N_21667,N_19497,N_19159);
and U21668 (N_21668,N_18144,N_19991);
or U21669 (N_21669,N_19695,N_18076);
nor U21670 (N_21670,N_18891,N_19440);
xor U21671 (N_21671,N_19204,N_18759);
and U21672 (N_21672,N_19199,N_18424);
and U21673 (N_21673,N_18159,N_19196);
xnor U21674 (N_21674,N_18852,N_19177);
xnor U21675 (N_21675,N_19349,N_19543);
xor U21676 (N_21676,N_18233,N_18299);
and U21677 (N_21677,N_19325,N_19117);
xnor U21678 (N_21678,N_18112,N_19036);
and U21679 (N_21679,N_19455,N_19944);
nor U21680 (N_21680,N_18002,N_19789);
or U21681 (N_21681,N_18480,N_19766);
xor U21682 (N_21682,N_18488,N_18303);
xnor U21683 (N_21683,N_18258,N_18621);
nor U21684 (N_21684,N_18751,N_18691);
nor U21685 (N_21685,N_19341,N_19464);
and U21686 (N_21686,N_18254,N_19256);
and U21687 (N_21687,N_18567,N_19977);
and U21688 (N_21688,N_19904,N_18625);
xnor U21689 (N_21689,N_19263,N_18273);
nand U21690 (N_21690,N_18759,N_18148);
or U21691 (N_21691,N_19557,N_18144);
or U21692 (N_21692,N_18272,N_19968);
nand U21693 (N_21693,N_19701,N_19784);
nand U21694 (N_21694,N_18040,N_19157);
and U21695 (N_21695,N_19982,N_19920);
or U21696 (N_21696,N_18890,N_19216);
xor U21697 (N_21697,N_19574,N_19322);
nand U21698 (N_21698,N_19768,N_18845);
or U21699 (N_21699,N_18196,N_19027);
and U21700 (N_21700,N_18046,N_18222);
nor U21701 (N_21701,N_19632,N_18219);
xor U21702 (N_21702,N_18371,N_18384);
nor U21703 (N_21703,N_18833,N_19508);
nand U21704 (N_21704,N_18552,N_18791);
and U21705 (N_21705,N_19162,N_18671);
nand U21706 (N_21706,N_19710,N_19069);
xnor U21707 (N_21707,N_18769,N_19555);
nor U21708 (N_21708,N_19838,N_18715);
xnor U21709 (N_21709,N_18347,N_18557);
or U21710 (N_21710,N_18142,N_18385);
xnor U21711 (N_21711,N_18960,N_19499);
nand U21712 (N_21712,N_19848,N_18901);
xnor U21713 (N_21713,N_19775,N_18633);
xor U21714 (N_21714,N_19946,N_19222);
nor U21715 (N_21715,N_18302,N_19474);
and U21716 (N_21716,N_18552,N_19908);
nand U21717 (N_21717,N_19623,N_19338);
xor U21718 (N_21718,N_19119,N_19681);
nor U21719 (N_21719,N_19777,N_18905);
nand U21720 (N_21720,N_18988,N_18573);
nand U21721 (N_21721,N_18819,N_18153);
and U21722 (N_21722,N_19693,N_18999);
or U21723 (N_21723,N_19542,N_19137);
nor U21724 (N_21724,N_18570,N_19056);
xnor U21725 (N_21725,N_18102,N_19083);
xor U21726 (N_21726,N_18349,N_19343);
or U21727 (N_21727,N_18559,N_18122);
nand U21728 (N_21728,N_19244,N_19543);
and U21729 (N_21729,N_18576,N_19654);
xnor U21730 (N_21730,N_19569,N_19586);
xor U21731 (N_21731,N_19385,N_18661);
nand U21732 (N_21732,N_18741,N_19628);
xnor U21733 (N_21733,N_19857,N_18568);
nand U21734 (N_21734,N_18509,N_18123);
and U21735 (N_21735,N_19201,N_18459);
nand U21736 (N_21736,N_18025,N_18269);
xor U21737 (N_21737,N_18591,N_18390);
nor U21738 (N_21738,N_18221,N_18939);
nand U21739 (N_21739,N_19747,N_19668);
nor U21740 (N_21740,N_18579,N_18938);
xor U21741 (N_21741,N_19905,N_19978);
nand U21742 (N_21742,N_18155,N_18456);
and U21743 (N_21743,N_19396,N_18054);
or U21744 (N_21744,N_19552,N_19247);
nor U21745 (N_21745,N_19855,N_19406);
nand U21746 (N_21746,N_19423,N_18013);
and U21747 (N_21747,N_18381,N_19656);
nor U21748 (N_21748,N_19320,N_19111);
nor U21749 (N_21749,N_18916,N_19313);
xnor U21750 (N_21750,N_18215,N_19446);
nor U21751 (N_21751,N_18349,N_18391);
xnor U21752 (N_21752,N_18928,N_19601);
xnor U21753 (N_21753,N_18608,N_19925);
xor U21754 (N_21754,N_18098,N_19805);
nand U21755 (N_21755,N_19890,N_18401);
and U21756 (N_21756,N_19309,N_19769);
or U21757 (N_21757,N_18544,N_19923);
or U21758 (N_21758,N_18179,N_19064);
and U21759 (N_21759,N_19266,N_19638);
nand U21760 (N_21760,N_18084,N_18185);
and U21761 (N_21761,N_19104,N_19983);
or U21762 (N_21762,N_18073,N_19064);
or U21763 (N_21763,N_19842,N_18407);
nand U21764 (N_21764,N_19135,N_18142);
and U21765 (N_21765,N_18227,N_18771);
xnor U21766 (N_21766,N_18017,N_18142);
and U21767 (N_21767,N_19595,N_18550);
or U21768 (N_21768,N_18227,N_19982);
and U21769 (N_21769,N_19049,N_18212);
xor U21770 (N_21770,N_18663,N_18879);
and U21771 (N_21771,N_18319,N_19023);
nor U21772 (N_21772,N_19594,N_19076);
nor U21773 (N_21773,N_18149,N_18960);
or U21774 (N_21774,N_19513,N_19924);
or U21775 (N_21775,N_19695,N_19776);
or U21776 (N_21776,N_19817,N_19497);
nand U21777 (N_21777,N_19490,N_18036);
xnor U21778 (N_21778,N_18121,N_18775);
nor U21779 (N_21779,N_18929,N_18586);
and U21780 (N_21780,N_19631,N_18267);
xor U21781 (N_21781,N_19155,N_18088);
nand U21782 (N_21782,N_18800,N_19773);
or U21783 (N_21783,N_19290,N_18644);
nor U21784 (N_21784,N_19789,N_19037);
or U21785 (N_21785,N_18180,N_18444);
xnor U21786 (N_21786,N_18802,N_18941);
nor U21787 (N_21787,N_18305,N_18400);
or U21788 (N_21788,N_19036,N_19889);
xor U21789 (N_21789,N_19086,N_19528);
nand U21790 (N_21790,N_19605,N_18727);
xor U21791 (N_21791,N_19511,N_18129);
or U21792 (N_21792,N_19585,N_18045);
nand U21793 (N_21793,N_18326,N_18455);
nand U21794 (N_21794,N_19218,N_19848);
nor U21795 (N_21795,N_18884,N_18357);
nand U21796 (N_21796,N_18313,N_18753);
nand U21797 (N_21797,N_19535,N_18204);
nor U21798 (N_21798,N_18190,N_18742);
and U21799 (N_21799,N_19611,N_18787);
xnor U21800 (N_21800,N_18705,N_19651);
or U21801 (N_21801,N_18552,N_19644);
or U21802 (N_21802,N_18477,N_19209);
and U21803 (N_21803,N_18987,N_19278);
nand U21804 (N_21804,N_19969,N_19845);
nor U21805 (N_21805,N_19203,N_18660);
xnor U21806 (N_21806,N_19066,N_19479);
or U21807 (N_21807,N_18142,N_18411);
xor U21808 (N_21808,N_18542,N_18137);
nor U21809 (N_21809,N_19403,N_18617);
xor U21810 (N_21810,N_19952,N_19740);
nor U21811 (N_21811,N_19528,N_18136);
nand U21812 (N_21812,N_19326,N_19163);
or U21813 (N_21813,N_19361,N_19798);
xnor U21814 (N_21814,N_19357,N_18383);
or U21815 (N_21815,N_19752,N_18621);
nand U21816 (N_21816,N_18772,N_19702);
or U21817 (N_21817,N_19090,N_19940);
or U21818 (N_21818,N_19616,N_18992);
xnor U21819 (N_21819,N_18731,N_18287);
nor U21820 (N_21820,N_18778,N_19217);
nand U21821 (N_21821,N_18408,N_18738);
nor U21822 (N_21822,N_19709,N_19162);
and U21823 (N_21823,N_18703,N_19998);
xor U21824 (N_21824,N_18174,N_19670);
and U21825 (N_21825,N_19038,N_18165);
nand U21826 (N_21826,N_18355,N_19277);
and U21827 (N_21827,N_19821,N_18062);
or U21828 (N_21828,N_19907,N_18156);
and U21829 (N_21829,N_18562,N_19660);
xnor U21830 (N_21830,N_18229,N_18269);
xor U21831 (N_21831,N_19695,N_18772);
nand U21832 (N_21832,N_19631,N_18686);
or U21833 (N_21833,N_18498,N_18920);
nor U21834 (N_21834,N_19157,N_19880);
nand U21835 (N_21835,N_18753,N_19331);
and U21836 (N_21836,N_19971,N_19707);
or U21837 (N_21837,N_18644,N_18372);
or U21838 (N_21838,N_19716,N_19602);
nor U21839 (N_21839,N_18653,N_19322);
or U21840 (N_21840,N_18133,N_19488);
xor U21841 (N_21841,N_19631,N_18804);
and U21842 (N_21842,N_19989,N_19263);
or U21843 (N_21843,N_18865,N_19670);
nand U21844 (N_21844,N_18897,N_19748);
nor U21845 (N_21845,N_18078,N_18635);
xor U21846 (N_21846,N_18476,N_19693);
nand U21847 (N_21847,N_19752,N_19317);
or U21848 (N_21848,N_19022,N_19679);
and U21849 (N_21849,N_18761,N_19963);
nor U21850 (N_21850,N_18555,N_19756);
nor U21851 (N_21851,N_19133,N_19732);
xnor U21852 (N_21852,N_18583,N_18772);
nor U21853 (N_21853,N_19875,N_19667);
or U21854 (N_21854,N_19704,N_19329);
nor U21855 (N_21855,N_18976,N_19068);
nand U21856 (N_21856,N_18397,N_19103);
or U21857 (N_21857,N_19171,N_18863);
xnor U21858 (N_21858,N_19473,N_19288);
or U21859 (N_21859,N_18722,N_19396);
nor U21860 (N_21860,N_18430,N_18840);
nand U21861 (N_21861,N_18358,N_18916);
nor U21862 (N_21862,N_19686,N_19187);
or U21863 (N_21863,N_19609,N_18865);
xor U21864 (N_21864,N_18422,N_18250);
and U21865 (N_21865,N_18430,N_18154);
and U21866 (N_21866,N_19152,N_18740);
or U21867 (N_21867,N_18394,N_18260);
nor U21868 (N_21868,N_19898,N_18948);
nor U21869 (N_21869,N_19317,N_19451);
or U21870 (N_21870,N_18772,N_18955);
and U21871 (N_21871,N_19069,N_18371);
nand U21872 (N_21872,N_19684,N_18658);
and U21873 (N_21873,N_19432,N_19407);
xor U21874 (N_21874,N_18159,N_18329);
or U21875 (N_21875,N_18431,N_19938);
nor U21876 (N_21876,N_19004,N_19201);
xor U21877 (N_21877,N_19404,N_19410);
and U21878 (N_21878,N_19931,N_19466);
nand U21879 (N_21879,N_19054,N_19035);
or U21880 (N_21880,N_18526,N_18603);
xnor U21881 (N_21881,N_19203,N_19073);
and U21882 (N_21882,N_19117,N_19572);
or U21883 (N_21883,N_19500,N_19481);
or U21884 (N_21884,N_19436,N_18284);
xnor U21885 (N_21885,N_18074,N_19752);
or U21886 (N_21886,N_19578,N_19101);
or U21887 (N_21887,N_18686,N_18898);
nand U21888 (N_21888,N_18749,N_18622);
or U21889 (N_21889,N_19916,N_19417);
nor U21890 (N_21890,N_19917,N_18753);
nand U21891 (N_21891,N_19713,N_19415);
xnor U21892 (N_21892,N_18436,N_19471);
nand U21893 (N_21893,N_18236,N_19863);
and U21894 (N_21894,N_19587,N_18579);
xnor U21895 (N_21895,N_18239,N_19716);
and U21896 (N_21896,N_19665,N_19051);
or U21897 (N_21897,N_19558,N_18426);
xnor U21898 (N_21898,N_18778,N_18682);
and U21899 (N_21899,N_18366,N_18388);
xor U21900 (N_21900,N_19549,N_19104);
nor U21901 (N_21901,N_19865,N_18070);
nor U21902 (N_21902,N_19742,N_19836);
nand U21903 (N_21903,N_19496,N_19167);
nor U21904 (N_21904,N_18440,N_18068);
or U21905 (N_21905,N_19168,N_19937);
xnor U21906 (N_21906,N_18510,N_18547);
nor U21907 (N_21907,N_19472,N_19930);
and U21908 (N_21908,N_18855,N_19333);
nand U21909 (N_21909,N_18858,N_18668);
nand U21910 (N_21910,N_18157,N_19684);
xnor U21911 (N_21911,N_18029,N_18208);
or U21912 (N_21912,N_18195,N_19942);
nand U21913 (N_21913,N_19753,N_18747);
nand U21914 (N_21914,N_18577,N_19091);
xnor U21915 (N_21915,N_18920,N_18404);
and U21916 (N_21916,N_18537,N_19690);
or U21917 (N_21917,N_18153,N_18745);
xor U21918 (N_21918,N_19554,N_19577);
xnor U21919 (N_21919,N_18120,N_19479);
nor U21920 (N_21920,N_19218,N_19208);
xor U21921 (N_21921,N_19946,N_19535);
nand U21922 (N_21922,N_19487,N_18245);
nand U21923 (N_21923,N_19417,N_18140);
xor U21924 (N_21924,N_18725,N_18771);
nand U21925 (N_21925,N_18631,N_18381);
xnor U21926 (N_21926,N_18500,N_18632);
nor U21927 (N_21927,N_19673,N_18608);
and U21928 (N_21928,N_18790,N_19416);
nor U21929 (N_21929,N_19286,N_18309);
or U21930 (N_21930,N_18642,N_18705);
nand U21931 (N_21931,N_19378,N_18573);
xor U21932 (N_21932,N_18350,N_18002);
xnor U21933 (N_21933,N_19811,N_19180);
nor U21934 (N_21934,N_18770,N_19366);
or U21935 (N_21935,N_18122,N_19214);
or U21936 (N_21936,N_18697,N_19171);
xor U21937 (N_21937,N_18961,N_18970);
nand U21938 (N_21938,N_19833,N_19773);
nor U21939 (N_21939,N_19829,N_19749);
nand U21940 (N_21940,N_19896,N_18198);
or U21941 (N_21941,N_18971,N_18828);
nand U21942 (N_21942,N_18591,N_18885);
and U21943 (N_21943,N_19293,N_19159);
nor U21944 (N_21944,N_19788,N_18663);
xor U21945 (N_21945,N_19743,N_18036);
nand U21946 (N_21946,N_18177,N_18632);
or U21947 (N_21947,N_19510,N_19433);
or U21948 (N_21948,N_18370,N_19048);
nand U21949 (N_21949,N_19627,N_19964);
nor U21950 (N_21950,N_18893,N_18396);
xor U21951 (N_21951,N_19938,N_18706);
or U21952 (N_21952,N_19989,N_19696);
and U21953 (N_21953,N_19792,N_19351);
and U21954 (N_21954,N_18993,N_18766);
xnor U21955 (N_21955,N_19633,N_19825);
xnor U21956 (N_21956,N_18385,N_18311);
and U21957 (N_21957,N_18169,N_18095);
and U21958 (N_21958,N_18383,N_19000);
xor U21959 (N_21959,N_18523,N_19740);
nor U21960 (N_21960,N_19035,N_18219);
xnor U21961 (N_21961,N_19283,N_19608);
or U21962 (N_21962,N_19008,N_19683);
xnor U21963 (N_21963,N_18164,N_19929);
nor U21964 (N_21964,N_19820,N_19010);
and U21965 (N_21965,N_18974,N_19396);
nor U21966 (N_21966,N_18470,N_19486);
nor U21967 (N_21967,N_18285,N_19939);
and U21968 (N_21968,N_19103,N_19298);
nor U21969 (N_21969,N_18447,N_19698);
xor U21970 (N_21970,N_19910,N_18926);
nor U21971 (N_21971,N_18158,N_18297);
nor U21972 (N_21972,N_19301,N_18664);
and U21973 (N_21973,N_18805,N_19115);
or U21974 (N_21974,N_18569,N_18468);
xor U21975 (N_21975,N_19763,N_18182);
and U21976 (N_21976,N_18010,N_19148);
nor U21977 (N_21977,N_18418,N_19062);
nor U21978 (N_21978,N_19765,N_19100);
xor U21979 (N_21979,N_18633,N_19307);
nor U21980 (N_21980,N_19928,N_19285);
nor U21981 (N_21981,N_18335,N_19611);
xor U21982 (N_21982,N_18661,N_18848);
and U21983 (N_21983,N_19700,N_18824);
or U21984 (N_21984,N_19286,N_19125);
nand U21985 (N_21985,N_18822,N_19490);
nor U21986 (N_21986,N_19305,N_19196);
or U21987 (N_21987,N_19453,N_18065);
nand U21988 (N_21988,N_19592,N_18610);
xor U21989 (N_21989,N_19800,N_18558);
nand U21990 (N_21990,N_18873,N_18030);
nand U21991 (N_21991,N_19859,N_19010);
nor U21992 (N_21992,N_18530,N_19534);
nor U21993 (N_21993,N_19429,N_18242);
nor U21994 (N_21994,N_18463,N_18692);
and U21995 (N_21995,N_19364,N_18783);
or U21996 (N_21996,N_19339,N_19933);
xnor U21997 (N_21997,N_19924,N_19553);
xnor U21998 (N_21998,N_19051,N_19141);
nand U21999 (N_21999,N_18213,N_19257);
xnor U22000 (N_22000,N_21033,N_21315);
xor U22001 (N_22001,N_20209,N_20949);
and U22002 (N_22002,N_21590,N_21109);
xnor U22003 (N_22003,N_20329,N_20187);
or U22004 (N_22004,N_21909,N_21709);
or U22005 (N_22005,N_20514,N_20610);
nor U22006 (N_22006,N_21297,N_20399);
nor U22007 (N_22007,N_21387,N_20350);
nand U22008 (N_22008,N_20821,N_21232);
and U22009 (N_22009,N_20696,N_21536);
or U22010 (N_22010,N_21056,N_21507);
xor U22011 (N_22011,N_21410,N_21365);
xor U22012 (N_22012,N_20150,N_20737);
nand U22013 (N_22013,N_21135,N_21293);
xnor U22014 (N_22014,N_20781,N_21695);
xnor U22015 (N_22015,N_20380,N_21597);
xnor U22016 (N_22016,N_20709,N_20438);
or U22017 (N_22017,N_20025,N_21389);
nor U22018 (N_22018,N_21133,N_21376);
or U22019 (N_22019,N_20365,N_21867);
nand U22020 (N_22020,N_20988,N_20048);
or U22021 (N_22021,N_21339,N_21999);
and U22022 (N_22022,N_20413,N_21492);
xor U22023 (N_22023,N_21242,N_20138);
nor U22024 (N_22024,N_20481,N_21101);
or U22025 (N_22025,N_20944,N_21271);
nand U22026 (N_22026,N_21490,N_21355);
xnor U22027 (N_22027,N_21829,N_20152);
nor U22028 (N_22028,N_21878,N_20328);
nand U22029 (N_22029,N_20089,N_21579);
xnor U22030 (N_22030,N_20278,N_20050);
xnor U22031 (N_22031,N_21209,N_21923);
and U22032 (N_22032,N_21324,N_21766);
nand U22033 (N_22033,N_21151,N_20607);
nor U22034 (N_22034,N_20293,N_20546);
or U22035 (N_22035,N_21066,N_21500);
xor U22036 (N_22036,N_20796,N_21247);
nor U22037 (N_22037,N_21152,N_21683);
and U22038 (N_22038,N_21237,N_20721);
nand U22039 (N_22039,N_21021,N_20450);
xnor U22040 (N_22040,N_20368,N_20661);
xor U22041 (N_22041,N_21974,N_21664);
nor U22042 (N_22042,N_21108,N_21004);
or U22043 (N_22043,N_20398,N_20954);
nor U22044 (N_22044,N_20464,N_20057);
nor U22045 (N_22045,N_21042,N_21982);
nor U22046 (N_22046,N_21868,N_21599);
nand U22047 (N_22047,N_20947,N_21091);
or U22048 (N_22048,N_21116,N_21710);
nand U22049 (N_22049,N_20909,N_21892);
or U22050 (N_22050,N_21431,N_20680);
and U22051 (N_22051,N_20857,N_21910);
and U22052 (N_22052,N_21094,N_21268);
nand U22053 (N_22053,N_20609,N_20600);
and U22054 (N_22054,N_20297,N_21498);
nand U22055 (N_22055,N_20778,N_21142);
or U22056 (N_22056,N_20810,N_21074);
nor U22057 (N_22057,N_21262,N_20316);
xnor U22058 (N_22058,N_20096,N_20714);
and U22059 (N_22059,N_21501,N_21838);
nor U22060 (N_22060,N_20026,N_21306);
xnor U22061 (N_22061,N_20597,N_20237);
and U22062 (N_22062,N_20518,N_20121);
and U22063 (N_22063,N_21001,N_21913);
and U22064 (N_22064,N_21699,N_21880);
nand U22065 (N_22065,N_20162,N_21055);
and U22066 (N_22066,N_20492,N_21893);
or U22067 (N_22067,N_20034,N_21879);
xnor U22068 (N_22068,N_21534,N_21456);
or U22069 (N_22069,N_21491,N_21092);
nand U22070 (N_22070,N_20912,N_20357);
nand U22071 (N_22071,N_21052,N_20540);
nor U22072 (N_22072,N_20344,N_20155);
or U22073 (N_22073,N_20407,N_21029);
nand U22074 (N_22074,N_21162,N_20184);
nand U22075 (N_22075,N_21251,N_20531);
or U22076 (N_22076,N_21650,N_21429);
and U22077 (N_22077,N_21637,N_21062);
and U22078 (N_22078,N_21160,N_20405);
xnor U22079 (N_22079,N_21214,N_20488);
and U22080 (N_22080,N_20742,N_20654);
xnor U22081 (N_22081,N_20467,N_20123);
nor U22082 (N_22082,N_20345,N_20183);
nand U22083 (N_22083,N_21844,N_21150);
xor U22084 (N_22084,N_20151,N_21640);
nand U22085 (N_22085,N_20740,N_20364);
nand U22086 (N_22086,N_21728,N_20157);
or U22087 (N_22087,N_21316,N_21856);
nand U22088 (N_22088,N_21660,N_20422);
and U22089 (N_22089,N_21243,N_21426);
and U22090 (N_22090,N_20074,N_21937);
xor U22091 (N_22091,N_20462,N_21864);
nor U22092 (N_22092,N_20880,N_20700);
nor U22093 (N_22093,N_20430,N_20071);
nand U22094 (N_22094,N_20159,N_20541);
nor U22095 (N_22095,N_20894,N_21677);
and U22096 (N_22096,N_20629,N_20707);
nor U22097 (N_22097,N_21964,N_21745);
nor U22098 (N_22098,N_20308,N_20489);
and U22099 (N_22099,N_20594,N_20750);
or U22100 (N_22100,N_20861,N_20961);
and U22101 (N_22101,N_20994,N_20687);
and U22102 (N_22102,N_20606,N_20186);
nand U22103 (N_22103,N_21520,N_20190);
xnor U22104 (N_22104,N_21208,N_20993);
nor U22105 (N_22105,N_20019,N_21628);
nor U22106 (N_22106,N_20896,N_21960);
nor U22107 (N_22107,N_21447,N_20615);
nor U22108 (N_22108,N_21687,N_20480);
and U22109 (N_22109,N_21577,N_21851);
or U22110 (N_22110,N_20276,N_21379);
or U22111 (N_22111,N_20161,N_21360);
nor U22112 (N_22112,N_20567,N_21043);
and U22113 (N_22113,N_20081,N_20082);
and U22114 (N_22114,N_20979,N_20213);
xor U22115 (N_22115,N_20200,N_21485);
or U22116 (N_22116,N_21886,N_20148);
or U22117 (N_22117,N_21825,N_20746);
nor U22118 (N_22118,N_21286,N_21702);
and U22119 (N_22119,N_20999,N_20494);
and U22120 (N_22120,N_21285,N_20106);
and U22121 (N_22121,N_21646,N_20719);
xor U22122 (N_22122,N_21688,N_21516);
or U22123 (N_22123,N_21971,N_21873);
and U22124 (N_22124,N_20473,N_20094);
and U22125 (N_22125,N_20469,N_20599);
xnor U22126 (N_22126,N_21483,N_20290);
or U22127 (N_22127,N_20243,N_21141);
nand U22128 (N_22128,N_20315,N_21434);
nand U22129 (N_22129,N_21013,N_20419);
nor U22130 (N_22130,N_20093,N_21254);
and U22131 (N_22131,N_21918,N_20589);
nor U22132 (N_22132,N_20616,N_21450);
nor U22133 (N_22133,N_20353,N_20114);
nor U22134 (N_22134,N_20614,N_20620);
or U22135 (N_22135,N_20374,N_21802);
or U22136 (N_22136,N_21994,N_20028);
or U22137 (N_22137,N_20506,N_20976);
nor U22138 (N_22138,N_20053,N_21951);
or U22139 (N_22139,N_21822,N_20671);
nand U22140 (N_22140,N_20009,N_20261);
and U22141 (N_22141,N_20327,N_21096);
nand U22142 (N_22142,N_20824,N_20173);
or U22143 (N_22143,N_21678,N_20250);
or U22144 (N_22144,N_21063,N_21192);
xnor U22145 (N_22145,N_20545,N_20475);
xnor U22146 (N_22146,N_21437,N_20558);
xnor U22147 (N_22147,N_21352,N_21428);
nor U22148 (N_22148,N_20453,N_21138);
or U22149 (N_22149,N_20552,N_21415);
or U22150 (N_22150,N_20710,N_20998);
nand U22151 (N_22151,N_20128,N_20142);
nand U22152 (N_22152,N_21551,N_21464);
xor U22153 (N_22153,N_21302,N_21606);
nor U22154 (N_22154,N_20834,N_20694);
nand U22155 (N_22155,N_21676,N_20883);
xor U22156 (N_22156,N_20641,N_20015);
nand U22157 (N_22157,N_21082,N_20387);
and U22158 (N_22158,N_20655,N_20862);
and U22159 (N_22159,N_20022,N_21290);
nand U22160 (N_22160,N_20853,N_20577);
nor U22161 (N_22161,N_20692,N_21222);
and U22162 (N_22162,N_20252,N_20685);
or U22163 (N_22163,N_21540,N_20215);
nand U22164 (N_22164,N_20145,N_20601);
and U22165 (N_22165,N_20512,N_21778);
or U22166 (N_22166,N_21479,N_21050);
nor U22167 (N_22167,N_20633,N_21330);
nor U22168 (N_22168,N_21451,N_21189);
and U22169 (N_22169,N_20131,N_21201);
nand U22170 (N_22170,N_20588,N_20231);
nand U22171 (N_22171,N_21182,N_21395);
and U22172 (N_22172,N_20660,N_21115);
nor U22173 (N_22173,N_20177,N_20455);
or U22174 (N_22174,N_21539,N_21146);
or U22175 (N_22175,N_21611,N_21436);
and U22176 (N_22176,N_21735,N_20471);
or U22177 (N_22177,N_21872,N_21835);
nand U22178 (N_22178,N_20220,N_21724);
or U22179 (N_22179,N_20521,N_21184);
and U22180 (N_22180,N_21481,N_21968);
xor U22181 (N_22181,N_21154,N_21284);
nand U22182 (N_22182,N_20491,N_20332);
xnor U22183 (N_22183,N_21080,N_21430);
xor U22184 (N_22184,N_21403,N_21327);
nor U22185 (N_22185,N_20156,N_21391);
nand U22186 (N_22186,N_21995,N_21409);
or U22187 (N_22187,N_20664,N_21468);
and U22188 (N_22188,N_20990,N_20669);
and U22189 (N_22189,N_21973,N_20608);
xnor U22190 (N_22190,N_21341,N_21503);
nand U22191 (N_22191,N_21629,N_21535);
xnor U22192 (N_22192,N_20920,N_21553);
nor U22193 (N_22193,N_21946,N_21039);
and U22194 (N_22194,N_20561,N_20593);
and U22195 (N_22195,N_21380,N_21749);
and U22196 (N_22196,N_20864,N_20100);
nor U22197 (N_22197,N_20795,N_21773);
xnor U22198 (N_22198,N_21077,N_20535);
nor U22199 (N_22199,N_21976,N_21943);
or U22200 (N_22200,N_20216,N_21600);
nor U22201 (N_22201,N_20466,N_20264);
nor U22202 (N_22202,N_21333,N_20638);
nor U22203 (N_22203,N_20863,N_20951);
and U22204 (N_22204,N_20806,N_20507);
xnor U22205 (N_22205,N_21236,N_21986);
nand U22206 (N_22206,N_21731,N_20956);
xor U22207 (N_22207,N_20902,N_20066);
or U22208 (N_22208,N_21642,N_21616);
or U22209 (N_22209,N_20943,N_20679);
nor U22210 (N_22210,N_20431,N_20918);
nor U22211 (N_22211,N_21439,N_21719);
nor U22212 (N_22212,N_20921,N_20051);
xor U22213 (N_22213,N_21213,N_20634);
xnor U22214 (N_22214,N_20741,N_21518);
nand U22215 (N_22215,N_20367,N_20748);
xor U22216 (N_22216,N_20612,N_21848);
or U22217 (N_22217,N_21343,N_21031);
nor U22218 (N_22218,N_21662,N_21028);
or U22219 (N_22219,N_20559,N_20371);
nor U22220 (N_22220,N_21764,N_21277);
nor U22221 (N_22221,N_21340,N_20309);
nor U22222 (N_22222,N_21040,N_20408);
or U22223 (N_22223,N_21947,N_20557);
xnor U22224 (N_22224,N_21163,N_20139);
xor U22225 (N_22225,N_21014,N_21705);
xnor U22226 (N_22226,N_21344,N_20170);
or U22227 (N_22227,N_20836,N_20112);
nand U22228 (N_22228,N_20706,N_21275);
xor U22229 (N_22229,N_20060,N_20504);
nor U22230 (N_22230,N_21147,N_21882);
xor U22231 (N_22231,N_21930,N_21808);
xor U22232 (N_22232,N_20233,N_20321);
nor U22233 (N_22233,N_21278,N_20505);
and U22234 (N_22234,N_20705,N_20105);
or U22235 (N_22235,N_21252,N_20087);
nor U22236 (N_22236,N_21668,N_20726);
or U22237 (N_22237,N_21026,N_20965);
nor U22238 (N_22238,N_21244,N_21682);
nand U22239 (N_22239,N_21124,N_21800);
nand U22240 (N_22240,N_20622,N_21128);
and U22241 (N_22241,N_20793,N_21538);
xor U22242 (N_22242,N_20851,N_20765);
nand U22243 (N_22243,N_21895,N_20476);
xor U22244 (N_22244,N_20985,N_21005);
and U22245 (N_22245,N_21165,N_21461);
nand U22246 (N_22246,N_20639,N_21003);
and U22247 (N_22247,N_20485,N_20032);
and U22248 (N_22248,N_20715,N_20772);
nand U22249 (N_22249,N_20977,N_21168);
nand U22250 (N_22250,N_21148,N_21854);
and U22251 (N_22251,N_20194,N_20981);
nand U22252 (N_22252,N_20938,N_21321);
nand U22253 (N_22253,N_21963,N_21367);
nor U22254 (N_22254,N_20447,N_20412);
nand U22255 (N_22255,N_20141,N_21506);
and U22256 (N_22256,N_21693,N_20570);
xor U22257 (N_22257,N_21869,N_21090);
xnor U22258 (N_22258,N_21644,N_21624);
nand U22259 (N_22259,N_21940,N_20035);
nand U22260 (N_22260,N_20320,N_20067);
or U22261 (N_22261,N_20298,N_21980);
nor U22262 (N_22262,N_21898,N_21266);
and U22263 (N_22263,N_21070,N_21794);
nor U22264 (N_22264,N_20259,N_21670);
xnor U22265 (N_22265,N_21806,N_20360);
nor U22266 (N_22266,N_20826,N_21020);
and U22267 (N_22267,N_20611,N_21862);
and U22268 (N_22268,N_21310,N_21299);
nand U22269 (N_22269,N_21566,N_21350);
nand U22270 (N_22270,N_20953,N_21186);
and U22271 (N_22271,N_20940,N_20925);
or U22272 (N_22272,N_20247,N_21657);
and U22273 (N_22273,N_20381,N_20840);
xnor U22274 (N_22274,N_20236,N_21753);
nor U22275 (N_22275,N_20586,N_21024);
or U22276 (N_22276,N_21348,N_21852);
or U22277 (N_22277,N_20666,N_21075);
and U22278 (N_22278,N_20792,N_20547);
and U22279 (N_22279,N_21009,N_21790);
nor U22280 (N_22280,N_21261,N_20870);
nor U22281 (N_22281,N_21057,N_20333);
or U22282 (N_22282,N_21765,N_20759);
nand U22283 (N_22283,N_21193,N_21296);
nor U22284 (N_22284,N_21499,N_20269);
and U22285 (N_22285,N_21820,N_20901);
or U22286 (N_22286,N_20527,N_20662);
and U22287 (N_22287,N_21086,N_21661);
xnor U22288 (N_22288,N_20133,N_20738);
nand U22289 (N_22289,N_20126,N_20650);
nor U22290 (N_22290,N_21533,N_21480);
nand U22291 (N_22291,N_21458,N_20487);
xnor U22292 (N_22292,N_21061,N_20744);
nor U22293 (N_22293,N_21972,N_21030);
nor U22294 (N_22294,N_21459,N_21239);
nor U22295 (N_22295,N_20343,N_20084);
or U22296 (N_22296,N_20798,N_20887);
or U22297 (N_22297,N_21076,N_21767);
nand U22298 (N_22298,N_20083,N_20299);
or U22299 (N_22299,N_20513,N_20733);
or U22300 (N_22300,N_20347,N_21981);
or U22301 (N_22301,N_20871,N_21233);
xnor U22302 (N_22302,N_21552,N_21174);
nand U22303 (N_22303,N_20843,N_21925);
nor U22304 (N_22304,N_21839,N_20681);
and U22305 (N_22305,N_21861,N_20058);
and U22306 (N_22306,N_21545,N_21761);
xor U22307 (N_22307,N_20076,N_20065);
xnor U22308 (N_22308,N_20045,N_21358);
nand U22309 (N_22309,N_21206,N_21750);
nor U22310 (N_22310,N_20199,N_20850);
and U22311 (N_22311,N_21441,N_21807);
and U22312 (N_22312,N_20673,N_20869);
and U22313 (N_22313,N_21303,N_21402);
or U22314 (N_22314,N_21388,N_20510);
nor U22315 (N_22315,N_20910,N_20052);
xor U22316 (N_22316,N_21068,N_20509);
nor U22317 (N_22317,N_20534,N_20049);
nand U22318 (N_22318,N_20149,N_20820);
or U22319 (N_22319,N_20273,N_21627);
nand U22320 (N_22320,N_21489,N_20729);
and U22321 (N_22321,N_20339,N_21263);
nor U22322 (N_22322,N_20361,N_20479);
and U22323 (N_22323,N_20785,N_20144);
nand U22324 (N_22324,N_21161,N_21989);
xor U22325 (N_22325,N_21811,N_20424);
or U22326 (N_22326,N_20542,N_20691);
nor U22327 (N_22327,N_21037,N_21405);
nand U22328 (N_22328,N_20036,N_21957);
nor U22329 (N_22329,N_20303,N_20454);
xor U22330 (N_22330,N_21706,N_20153);
nand U22331 (N_22331,N_20246,N_20932);
xnor U22332 (N_22332,N_20584,N_21801);
xnor U22333 (N_22333,N_21435,N_21111);
and U22334 (N_22334,N_20583,N_20446);
and U22335 (N_22335,N_21818,N_20042);
and U22336 (N_22336,N_21051,N_21667);
nor U22337 (N_22337,N_21809,N_20794);
and U22338 (N_22338,N_20369,N_20749);
nand U22339 (N_22339,N_20286,N_21855);
xnor U22340 (N_22340,N_21651,N_21685);
nand U22341 (N_22341,N_21928,N_21328);
xnor U22342 (N_22342,N_20027,N_21496);
and U22343 (N_22343,N_20970,N_20493);
nor U22344 (N_22344,N_21572,N_20693);
nor U22345 (N_22345,N_20031,N_21784);
nor U22346 (N_22346,N_20728,N_21530);
and U22347 (N_22347,N_21203,N_21543);
and U22348 (N_22348,N_21527,N_20301);
or U22349 (N_22349,N_20665,N_20352);
and U22350 (N_22350,N_21273,N_20948);
and U22351 (N_22351,N_21860,N_20288);
nand U22352 (N_22352,N_20676,N_21058);
or U22353 (N_22353,N_20336,N_21272);
and U22354 (N_22354,N_20983,N_21265);
xnor U22355 (N_22355,N_21532,N_20804);
nand U22356 (N_22356,N_20179,N_20078);
nand U22357 (N_22357,N_21803,N_20569);
nor U22358 (N_22358,N_20978,N_20030);
nand U22359 (N_22359,N_21849,N_21698);
nor U22360 (N_22360,N_20683,N_20926);
or U22361 (N_22361,N_21961,N_20415);
or U22362 (N_22362,N_20244,N_21122);
nand U22363 (N_22363,N_20585,N_20182);
xor U22364 (N_22364,N_20950,N_20827);
and U22365 (N_22365,N_20091,N_20059);
nor U22366 (N_22366,N_20385,N_20704);
nor U22367 (N_22367,N_21674,N_21763);
nand U22368 (N_22368,N_21639,N_20136);
xnor U22369 (N_22369,N_20118,N_20193);
or U22370 (N_22370,N_20474,N_21605);
and U22371 (N_22371,N_20115,N_21176);
nor U22372 (N_22372,N_21965,N_20224);
or U22373 (N_22373,N_20029,N_21181);
xnor U22374 (N_22374,N_21465,N_21411);
nand U22375 (N_22375,N_20952,N_21319);
nand U22376 (N_22376,N_20735,N_21656);
nor U22377 (N_22377,N_20571,N_20204);
and U22378 (N_22378,N_21497,N_20241);
nor U22379 (N_22379,N_21777,N_21899);
or U22380 (N_22380,N_20260,N_20900);
or U22381 (N_22381,N_20211,N_20079);
nand U22382 (N_22382,N_20372,N_20354);
nand U22383 (N_22383,N_21159,N_21522);
and U22384 (N_22384,N_21023,N_20110);
xnor U22385 (N_22385,N_21412,N_21812);
nand U22386 (N_22386,N_20645,N_21515);
nor U22387 (N_22387,N_21107,N_21783);
nand U22388 (N_22388,N_20109,N_21308);
and U22389 (N_22389,N_20291,N_21495);
and U22390 (N_22390,N_20515,N_21269);
nand U22391 (N_22391,N_20443,N_21555);
or U22392 (N_22392,N_20086,N_21137);
xor U22393 (N_22393,N_20168,N_20366);
xnor U22394 (N_22394,N_20120,N_21593);
xnor U22395 (N_22395,N_21740,N_21573);
xnor U22396 (N_22396,N_21198,N_20695);
and U22397 (N_22397,N_20143,N_20452);
and U22398 (N_22398,N_21334,N_21183);
nor U22399 (N_22399,N_20482,N_20124);
nor U22400 (N_22400,N_20922,N_20005);
xor U22401 (N_22401,N_20957,N_20495);
nor U22402 (N_22402,N_20538,N_20682);
or U22403 (N_22403,N_21591,N_20971);
xor U22404 (N_22404,N_21889,N_21104);
nor U22405 (N_22405,N_21920,N_20562);
xor U22406 (N_22406,N_21235,N_20217);
and U22407 (N_22407,N_21118,N_20272);
or U22408 (N_22408,N_21787,N_21721);
nor U22409 (N_22409,N_20623,N_21905);
xnor U22410 (N_22410,N_21774,N_21145);
and U22411 (N_22411,N_20295,N_20739);
nor U22412 (N_22412,N_21796,N_21840);
xor U22413 (N_22413,N_21114,N_21433);
xor U22414 (N_22414,N_20876,N_20038);
nand U22415 (N_22415,N_20899,N_20502);
xor U22416 (N_22416,N_21167,N_20905);
or U22417 (N_22417,N_20519,N_21392);
and U22418 (N_22418,N_20960,N_20478);
nand U22419 (N_22419,N_20396,N_21228);
nor U22420 (N_22420,N_21647,N_20718);
or U22421 (N_22421,N_20849,N_20451);
xnor U22422 (N_22422,N_21155,N_21249);
and U22423 (N_22423,N_20873,N_20814);
nor U22424 (N_22424,N_20459,N_20219);
or U22425 (N_22425,N_20539,N_20055);
and U22426 (N_22426,N_20812,N_21103);
nor U22427 (N_22427,N_20470,N_20537);
nor U22428 (N_22428,N_20668,N_20874);
xnor U22429 (N_22429,N_20439,N_21220);
or U22430 (N_22430,N_21488,N_20757);
and U22431 (N_22431,N_21173,N_21353);
and U22432 (N_22432,N_20310,N_20117);
nor U22433 (N_22433,N_21313,N_21875);
nand U22434 (N_22434,N_21841,N_21821);
nor U22435 (N_22435,N_21325,N_20214);
nand U22436 (N_22436,N_21797,N_20931);
and U22437 (N_22437,N_21569,N_21751);
nand U22438 (N_22438,N_21900,N_21514);
nand U22439 (N_22439,N_21099,N_20391);
and U22440 (N_22440,N_20958,N_21472);
and U22441 (N_22441,N_20014,N_20490);
xor U22442 (N_22442,N_21517,N_20575);
or U22443 (N_22443,N_20617,N_20690);
or U22444 (N_22444,N_20348,N_20674);
and U22445 (N_22445,N_21748,N_21666);
and U22446 (N_22446,N_20181,N_20727);
xnor U22447 (N_22447,N_21658,N_20895);
nor U22448 (N_22448,N_21136,N_20382);
or U22449 (N_22449,N_20158,N_20147);
nor U22450 (N_22450,N_21127,N_21032);
or U22451 (N_22451,N_20725,N_21362);
or U22452 (N_22452,N_21356,N_20845);
xor U22453 (N_22453,N_20764,N_20460);
nor U22454 (N_22454,N_21322,N_21883);
and U22455 (N_22455,N_20279,N_21393);
xor U22456 (N_22456,N_20730,N_21939);
nand U22457 (N_22457,N_21788,N_21396);
or U22458 (N_22458,N_21385,N_21166);
and U22459 (N_22459,N_21349,N_20881);
nand U22460 (N_22460,N_21563,N_20113);
xnor U22461 (N_22461,N_21487,N_20206);
and U22462 (N_22462,N_21992,N_21072);
xnor U22463 (N_22463,N_21255,N_20913);
or U22464 (N_22464,N_20813,N_21716);
or U22465 (N_22465,N_20776,N_21817);
and U22466 (N_22466,N_21419,N_20678);
nand U22467 (N_22467,N_21226,N_21291);
xnor U22468 (N_22468,N_20501,N_21620);
and U22469 (N_22469,N_20020,N_21320);
xor U22470 (N_22470,N_20986,N_20132);
nand U22471 (N_22471,N_20859,N_20628);
or U22472 (N_22472,N_20817,N_21592);
or U22473 (N_22473,N_20061,N_20822);
nand U22474 (N_22474,N_21589,N_21416);
nor U22475 (N_22475,N_21842,N_21945);
nor U22476 (N_22476,N_20867,N_21603);
xnor U22477 (N_22477,N_20805,N_20257);
xor U22478 (N_22478,N_21541,N_20389);
xor U22479 (N_22479,N_21125,N_21065);
and U22480 (N_22480,N_20090,N_20780);
or U22481 (N_22481,N_20442,N_21594);
nand U22482 (N_22482,N_21399,N_21635);
and U22483 (N_22483,N_20911,N_20072);
nor U22484 (N_22484,N_21703,N_20189);
xnor U22485 (N_22485,N_21510,N_20621);
nand U22486 (N_22486,N_21301,N_20356);
nand U22487 (N_22487,N_21554,N_20300);
or U22488 (N_22488,N_21314,N_20722);
and U22489 (N_22489,N_21229,N_21954);
xnor U22490 (N_22490,N_21460,N_20929);
xor U22491 (N_22491,N_20903,N_20923);
nand U22492 (N_22492,N_20208,N_20831);
xnor U22493 (N_22493,N_20974,N_20982);
xor U22494 (N_22494,N_21830,N_21420);
or U22495 (N_22495,N_20024,N_21558);
and U22496 (N_22496,N_20543,N_21007);
xnor U22497 (N_22497,N_21386,N_20317);
and U22498 (N_22498,N_20790,N_20004);
nor U22499 (N_22499,N_21587,N_21614);
or U22500 (N_22500,N_20167,N_20283);
and U22501 (N_22501,N_20003,N_21281);
xor U22502 (N_22502,N_21218,N_20355);
xnor U22503 (N_22503,N_21565,N_20379);
nor U22504 (N_22504,N_21338,N_20285);
xor U22505 (N_22505,N_21512,N_20165);
and U22506 (N_22506,N_20769,N_20263);
nor U22507 (N_22507,N_21401,N_21288);
or U22508 (N_22508,N_21734,N_21576);
and U22509 (N_22509,N_20330,N_21095);
xnor U22510 (N_22510,N_21083,N_20016);
nor U22511 (N_22511,N_20774,N_21826);
nand U22512 (N_22512,N_21054,N_21571);
nand U22513 (N_22513,N_20331,N_20946);
xnor U22514 (N_22514,N_21078,N_21726);
and U22515 (N_22515,N_20815,N_21071);
or U22516 (N_22516,N_20255,N_20897);
or U22517 (N_22517,N_21914,N_21225);
nor U22518 (N_22518,N_20636,N_20833);
nor U22519 (N_22519,N_20941,N_21016);
xnor U22520 (N_22520,N_21106,N_20229);
nor U22521 (N_22521,N_20129,N_20865);
xnor U22522 (N_22522,N_20630,N_21513);
nand U22523 (N_22523,N_21962,N_21736);
and U22524 (N_22524,N_21126,N_21169);
or U22525 (N_22525,N_20403,N_20797);
and U22526 (N_22526,N_20670,N_21445);
and U22527 (N_22527,N_21250,N_21977);
and U22528 (N_22528,N_20743,N_20936);
nor U22529 (N_22529,N_20251,N_20618);
or U22530 (N_22530,N_21549,N_21623);
nand U22531 (N_22531,N_21701,N_20969);
and U22532 (N_22532,N_20172,N_21630);
nand U22533 (N_22533,N_21351,N_20659);
nand U22534 (N_22534,N_20370,N_20777);
nand U22535 (N_22535,N_20893,N_20075);
xor U22536 (N_22536,N_21596,N_21729);
nand U22537 (N_22537,N_21318,N_20847);
and U22538 (N_22538,N_20335,N_21890);
or U22539 (N_22539,N_20054,N_21793);
or U22540 (N_22540,N_21267,N_20846);
xor U22541 (N_22541,N_20713,N_20322);
nand U22542 (N_22542,N_20752,N_20281);
nor U22543 (N_22543,N_20578,N_21584);
and U22544 (N_22544,N_21443,N_20287);
and U22545 (N_22545,N_20717,N_20313);
or U22546 (N_22546,N_20296,N_20312);
xor U22547 (N_22547,N_20756,N_21309);
and U22548 (N_22548,N_21582,N_21292);
nand U22549 (N_22549,N_20898,N_20334);
nand U22550 (N_22550,N_20525,N_21824);
and U22551 (N_22551,N_20107,N_20647);
or U22552 (N_22552,N_21632,N_21924);
or U22553 (N_22553,N_21727,N_21874);
nand U22554 (N_22554,N_21347,N_21175);
or U22555 (N_22555,N_21739,N_20294);
nand U22556 (N_22556,N_20458,N_21470);
xnor U22557 (N_22557,N_21248,N_20642);
nor U22558 (N_22558,N_21955,N_21471);
xor U22559 (N_22559,N_20522,N_20520);
nor U22560 (N_22560,N_20195,N_21626);
xor U22561 (N_22561,N_20548,N_21941);
xnor U22562 (N_22562,N_21368,N_21217);
nor U22563 (N_22563,N_20788,N_21486);
or U22564 (N_22564,N_20503,N_21345);
or U22565 (N_22565,N_20463,N_21234);
or U22566 (N_22566,N_20390,N_20001);
or U22567 (N_22567,N_20854,N_21179);
and U22568 (N_22568,N_21689,N_21567);
nand U22569 (N_22569,N_20013,N_21827);
nor U22570 (N_22570,N_21547,N_21178);
nand U22571 (N_22571,N_21548,N_21475);
nor U22572 (N_22572,N_20037,N_21531);
nand U22573 (N_22573,N_20268,N_21329);
nor U22574 (N_22574,N_20169,N_21164);
nor U22575 (N_22575,N_20763,N_20755);
xor U22576 (N_22576,N_20837,N_21190);
and U22577 (N_22577,N_20282,N_20425);
xor U22578 (N_22578,N_21690,N_21649);
xnor U22579 (N_22579,N_20337,N_21612);
nor U22580 (N_22580,N_20423,N_20825);
or U22581 (N_22581,N_20500,N_20377);
or U22582 (N_22582,N_21929,N_20119);
nand U22583 (N_22583,N_21884,N_21828);
or U22584 (N_22584,N_21770,N_20908);
or U22585 (N_22585,N_21073,N_21438);
and U22586 (N_22586,N_21559,N_21942);
nor U22587 (N_22587,N_20362,N_20675);
or U22588 (N_22588,N_20884,N_20040);
nand U22589 (N_22589,N_21756,N_20207);
xnor U22590 (N_22590,N_21737,N_20404);
xnor U22591 (N_22591,N_21585,N_21509);
xor U22592 (N_22592,N_21158,N_21449);
or U22593 (N_22593,N_20305,N_21085);
or U22594 (N_22594,N_21197,N_21130);
and U22595 (N_22595,N_21885,N_21832);
nor U22596 (N_22596,N_20202,N_20731);
or U22597 (N_22597,N_20565,N_21795);
nand U22598 (N_22598,N_20656,N_21455);
nor U22599 (N_22599,N_21686,N_21400);
nand U22600 (N_22600,N_20205,N_20761);
nand U22601 (N_22601,N_20324,N_20484);
xor U22602 (N_22602,N_21786,N_20819);
nor U22603 (N_22603,N_21768,N_21454);
or U22604 (N_22604,N_21245,N_21967);
nand U22605 (N_22605,N_21833,N_21215);
and U22606 (N_22606,N_21363,N_20689);
nand U22607 (N_22607,N_21110,N_20566);
nand U22608 (N_22608,N_20346,N_21779);
nand U22609 (N_22609,N_20603,N_21908);
or U22610 (N_22610,N_20457,N_20564);
nor U22611 (N_22611,N_21300,N_21949);
nand U22612 (N_22612,N_20635,N_20592);
and U22613 (N_22613,N_21525,N_20409);
xnor U22614 (N_22614,N_21953,N_21210);
or U22615 (N_22615,N_20046,N_21397);
and U22616 (N_22616,N_20393,N_21732);
and U22617 (N_22617,N_20358,N_21870);
and U22618 (N_22618,N_20176,N_21508);
xor U22619 (N_22619,N_20553,N_20766);
nor U22620 (N_22620,N_20904,N_21969);
nand U22621 (N_22621,N_21238,N_20935);
and U22622 (N_22622,N_20576,N_20980);
nand U22623 (N_22623,N_21815,N_20627);
or U22624 (N_22624,N_20852,N_21258);
xor U22625 (N_22625,N_21781,N_20916);
nor U22626 (N_22626,N_21588,N_20582);
nand U22627 (N_22627,N_20417,N_21084);
nand U22628 (N_22628,N_20832,N_21669);
nand U22629 (N_22629,N_21195,N_21523);
nor U22630 (N_22630,N_21093,N_21199);
xor U22631 (N_22631,N_20551,N_21715);
or U22632 (N_22632,N_21816,N_21601);
xor U22633 (N_22633,N_20445,N_21782);
nor U22634 (N_22634,N_21187,N_20631);
xnor U22635 (N_22635,N_20858,N_20497);
xnor U22636 (N_22636,N_21185,N_21866);
nor U22637 (N_22637,N_20939,N_20047);
nor U22638 (N_22638,N_20311,N_21602);
xor U22639 (N_22639,N_21615,N_21132);
xor U22640 (N_22640,N_21744,N_21776);
nand U22641 (N_22641,N_20441,N_21041);
nor U22642 (N_22642,N_21700,N_20373);
or U22643 (N_22643,N_20127,N_21194);
nand U22644 (N_22644,N_21000,N_20021);
and U22645 (N_22645,N_21791,N_20686);
or U22646 (N_22646,N_20652,N_20275);
and U22647 (N_22647,N_20188,N_20137);
or U22648 (N_22648,N_20196,N_20754);
and U22649 (N_22649,N_20420,N_20434);
or U22650 (N_22650,N_21157,N_21718);
nand U22651 (N_22651,N_20720,N_20803);
nand U22652 (N_22652,N_21891,N_20070);
xor U22653 (N_22653,N_21448,N_21469);
xor U22654 (N_22654,N_20800,N_20449);
nand U22655 (N_22655,N_20580,N_21926);
and U22656 (N_22656,N_20964,N_21047);
nor U22657 (N_22657,N_21717,N_20770);
nor U22658 (N_22658,N_21894,N_20018);
nand U22659 (N_22659,N_20240,N_21204);
or U22660 (N_22660,N_20302,N_21636);
nand U22661 (N_22661,N_21607,N_21283);
nand U22662 (N_22662,N_21048,N_21311);
and U22663 (N_22663,N_21224,N_20400);
or U22664 (N_22664,N_20536,N_20767);
or U22665 (N_22665,N_20508,N_20529);
nor U22666 (N_22666,N_21335,N_21634);
xor U22667 (N_22667,N_20791,N_21304);
xnor U22668 (N_22668,N_20062,N_20962);
nor U22669 (N_22669,N_21814,N_20008);
nand U22670 (N_22670,N_20292,N_20444);
nor U22671 (N_22671,N_20802,N_21406);
and U22672 (N_22672,N_21568,N_21526);
and U22673 (N_22673,N_20418,N_21743);
nand U22674 (N_22674,N_21414,N_21711);
xnor U22675 (N_22675,N_20017,N_21257);
xor U22676 (N_22676,N_20421,N_21177);
nor U22677 (N_22677,N_20928,N_21064);
nor U22678 (N_22678,N_21733,N_21556);
and U22679 (N_22679,N_20598,N_21102);
xor U22680 (N_22680,N_21046,N_21097);
or U22681 (N_22681,N_21357,N_21741);
nor U22682 (N_22682,N_20891,N_21704);
nor U22683 (N_22683,N_21053,N_21991);
nor U22684 (N_22684,N_21772,N_21679);
xnor U22685 (N_22685,N_21675,N_20440);
nor U22686 (N_22686,N_20550,N_20012);
and U22687 (N_22687,N_20745,N_21067);
nor U22688 (N_22688,N_21671,N_21998);
and U22689 (N_22689,N_21100,N_21044);
nand U22690 (N_22690,N_21069,N_20555);
or U22691 (N_22691,N_20221,N_21887);
xnor U22692 (N_22692,N_20697,N_21673);
and U22693 (N_22693,N_20888,N_21006);
xor U22694 (N_22694,N_20688,N_21253);
or U22695 (N_22695,N_21404,N_21241);
xor U22696 (N_22696,N_21935,N_20258);
and U22697 (N_22697,N_21876,N_21696);
nor U22698 (N_22698,N_20266,N_21332);
and U22699 (N_22699,N_21810,N_20319);
nor U22700 (N_22700,N_21625,N_21354);
and U22701 (N_22701,N_21474,N_20351);
nor U22702 (N_22702,N_21139,N_21931);
xnor U22703 (N_22703,N_21342,N_20924);
or U22704 (N_22704,N_20375,N_20712);
nor U22705 (N_22705,N_21759,N_20056);
xor U22706 (N_22706,N_20885,N_20427);
nor U22707 (N_22707,N_21002,N_21714);
nand U22708 (N_22708,N_21457,N_20996);
or U22709 (N_22709,N_20359,N_21871);
nand U22710 (N_22710,N_20006,N_21117);
nor U22711 (N_22711,N_21985,N_21785);
and U22712 (N_22712,N_20829,N_21697);
xnor U22713 (N_22713,N_20587,N_21098);
and U22714 (N_22714,N_20043,N_21384);
xor U22715 (N_22715,N_21877,N_21202);
nand U22716 (N_22716,N_20069,N_21652);
xnor U22717 (N_22717,N_21619,N_21578);
xnor U22718 (N_22718,N_20426,N_21746);
nor U22719 (N_22719,N_20643,N_21713);
and U22720 (N_22720,N_20579,N_21618);
and U22721 (N_22721,N_21912,N_20937);
xor U22722 (N_22722,N_20875,N_20625);
or U22723 (N_22723,N_21595,N_21149);
nand U22724 (N_22724,N_20968,N_21442);
xnor U22725 (N_22725,N_20613,N_21346);
xor U22726 (N_22726,N_20108,N_21035);
xor U22727 (N_22727,N_20995,N_21398);
nand U22728 (N_22728,N_21888,N_20146);
or U22729 (N_22729,N_20383,N_20632);
nor U22730 (N_22730,N_21231,N_20274);
and U22731 (N_22731,N_21916,N_20228);
and U22732 (N_22732,N_20872,N_21659);
nor U22733 (N_22733,N_20416,N_21617);
and U22734 (N_22734,N_20429,N_21608);
xor U22735 (N_22735,N_20125,N_20363);
and U22736 (N_22736,N_21843,N_20245);
nor U22737 (N_22737,N_21246,N_21294);
nand U22738 (N_22738,N_20855,N_21654);
nor U22739 (N_22739,N_21792,N_21478);
nand U22740 (N_22740,N_20103,N_21983);
or U22741 (N_22741,N_20435,N_21823);
nand U22742 (N_22742,N_21425,N_21494);
nand U22743 (N_22743,N_20838,N_21769);
xor U22744 (N_22744,N_21274,N_21570);
xor U22745 (N_22745,N_21361,N_21804);
or U22746 (N_22746,N_21493,N_21859);
or U22747 (N_22747,N_21089,N_20860);
nor U22748 (N_22748,N_20092,N_21948);
nor U22749 (N_22749,N_20163,N_21663);
xor U22750 (N_22750,N_20342,N_21979);
nand U22751 (N_22751,N_20392,N_20198);
and U22752 (N_22752,N_21371,N_21264);
nand U22753 (N_22753,N_21413,N_21337);
nand U22754 (N_22754,N_21762,N_21105);
and U22755 (N_22755,N_20684,N_21813);
and U22756 (N_22756,N_21907,N_21427);
nand U22757 (N_22757,N_21707,N_20959);
nor U22758 (N_22758,N_20992,N_21915);
or U22759 (N_22759,N_21336,N_20604);
nor U22760 (N_22760,N_21011,N_21129);
or U22761 (N_22761,N_20180,N_20828);
and U22762 (N_22762,N_21672,N_20602);
xor U22763 (N_22763,N_20104,N_20984);
nor U22764 (N_22764,N_21240,N_21079);
or U22765 (N_22765,N_20323,N_21837);
or U22766 (N_22766,N_21484,N_21452);
nor U22767 (N_22767,N_21665,N_21546);
and U22768 (N_22768,N_20699,N_20915);
nor U22769 (N_22769,N_20758,N_20626);
nor U22770 (N_22770,N_21374,N_21902);
xnor U22771 (N_22771,N_21938,N_20549);
xor U22772 (N_22772,N_20972,N_20063);
and U22773 (N_22773,N_21780,N_21289);
nor U22774 (N_22774,N_21956,N_21988);
nor U22775 (N_22775,N_21934,N_21256);
nand U22776 (N_22776,N_21799,N_20201);
or U22777 (N_22777,N_20945,N_21641);
xnor U22778 (N_22778,N_21896,N_20325);
or U22779 (N_22779,N_20753,N_20657);
xor U22780 (N_22780,N_21120,N_20134);
or U22781 (N_22781,N_20786,N_20573);
or U22782 (N_22782,N_21708,N_21171);
xor U22783 (N_22783,N_20716,N_20927);
nand U22784 (N_22784,N_20848,N_20011);
xor U22785 (N_22785,N_20218,N_21408);
nand U22786 (N_22786,N_21381,N_21958);
nand U22787 (N_22787,N_21648,N_21188);
or U22788 (N_22788,N_20101,N_20222);
nand U22789 (N_22789,N_20002,N_21692);
or U22790 (N_22790,N_21446,N_20523);
and U22791 (N_22791,N_20338,N_21524);
or U22792 (N_22792,N_20768,N_20809);
xnor U22793 (N_22793,N_21557,N_21730);
and U22794 (N_22794,N_21805,N_20563);
nor U22795 (N_22795,N_20239,N_20242);
and U22796 (N_22796,N_21372,N_20433);
and U22797 (N_22797,N_20064,N_20437);
xnor U22798 (N_22798,N_21259,N_21010);
and U22799 (N_22799,N_21144,N_21112);
nand U22800 (N_22800,N_20039,N_21153);
xor U22801 (N_22801,N_20468,N_21422);
nor U22802 (N_22802,N_21580,N_20963);
and U22803 (N_22803,N_20967,N_21119);
and U22804 (N_22804,N_20192,N_20856);
nand U22805 (N_22805,N_21407,N_20388);
nor U22806 (N_22806,N_20164,N_20701);
xnor U22807 (N_22807,N_20111,N_20517);
or U22808 (N_22808,N_20212,N_21287);
or U22809 (N_22809,N_21466,N_21113);
nand U22810 (N_22810,N_21383,N_20267);
and U22811 (N_22811,N_21561,N_20000);
nor U22812 (N_22812,N_20154,N_20378);
and U22813 (N_22813,N_21901,N_20789);
and U22814 (N_22814,N_20526,N_20185);
or U22815 (N_22815,N_21680,N_20116);
nor U22816 (N_22816,N_21919,N_20653);
or U22817 (N_22817,N_20340,N_20226);
nand U22818 (N_22818,N_21906,N_21537);
and U22819 (N_22819,N_20088,N_21087);
and U22820 (N_22820,N_21691,N_20174);
xnor U22821 (N_22821,N_20289,N_20210);
or U22822 (N_22822,N_20818,N_21984);
and U22823 (N_22823,N_21834,N_21476);
xor U22824 (N_22824,N_21544,N_21681);
or U22825 (N_22825,N_21172,N_20483);
nand U22826 (N_22826,N_20782,N_21712);
nand U22827 (N_22827,N_20530,N_21738);
nand U22828 (N_22828,N_20677,N_20667);
nor U22829 (N_22829,N_20942,N_20197);
xnor U22830 (N_22830,N_20277,N_21140);
xor U22831 (N_22831,N_20099,N_20917);
nor U22832 (N_22832,N_20987,N_20544);
or U22833 (N_22833,N_20306,N_21212);
or U22834 (N_22834,N_21847,N_21850);
nor U22835 (N_22835,N_21223,N_21643);
nor U22836 (N_22836,N_21081,N_20401);
or U22837 (N_22837,N_21655,N_20256);
and U22838 (N_22838,N_21375,N_20318);
and U22839 (N_22839,N_20033,N_20658);
or U22840 (N_22840,N_21858,N_20711);
and U22841 (N_22841,N_21684,N_20394);
and U22842 (N_22842,N_21424,N_21959);
and U22843 (N_22843,N_20747,N_20595);
xor U22844 (N_22844,N_20077,N_20866);
or U22845 (N_22845,N_20304,N_20648);
nand U22846 (N_22846,N_20835,N_20879);
or U22847 (N_22847,N_21583,N_20775);
nor U22848 (N_22848,N_20326,N_21609);
nand U22849 (N_22849,N_20498,N_20411);
nand U22850 (N_22850,N_20225,N_20762);
xor U22851 (N_22851,N_20010,N_20160);
nand U22852 (N_22852,N_21836,N_20314);
nand U22853 (N_22853,N_21230,N_20989);
nor U22854 (N_22854,N_20080,N_20823);
or U22855 (N_22855,N_21542,N_21022);
and U22856 (N_22856,N_21211,N_20830);
and U22857 (N_22857,N_21221,N_20892);
nand U22858 (N_22858,N_21017,N_20262);
nand U22859 (N_22859,N_21562,N_20068);
nor U22860 (N_22860,N_21143,N_20889);
nand U22861 (N_22861,N_20532,N_20732);
xor U22862 (N_22862,N_21723,N_21694);
nor U22863 (N_22863,N_21505,N_20973);
nor U22864 (N_22864,N_21156,N_21504);
or U22865 (N_22865,N_20672,N_20839);
nor U22866 (N_22866,N_21462,N_20140);
nor U22867 (N_22867,N_20724,N_21725);
nor U22868 (N_22868,N_21134,N_21018);
xnor U22869 (N_22869,N_21560,N_21180);
xnor U22870 (N_22870,N_21917,N_21045);
nand U22871 (N_22871,N_21921,N_21604);
xnor U22872 (N_22872,N_20175,N_20882);
nor U22873 (N_22873,N_21049,N_20097);
nor U22874 (N_22874,N_21312,N_20472);
nor U22875 (N_22875,N_21897,N_20166);
nor U22876 (N_22876,N_21276,N_20702);
nand U22877 (N_22877,N_20736,N_20171);
nand U22878 (N_22878,N_20930,N_21382);
and U22879 (N_22879,N_21207,N_21390);
and U22880 (N_22880,N_21200,N_20619);
nand U22881 (N_22881,N_20811,N_20799);
xor U22882 (N_22882,N_21903,N_21377);
xor U22883 (N_22883,N_20461,N_21366);
or U22884 (N_22884,N_21519,N_20223);
xnor U22885 (N_22885,N_20556,N_20386);
and U22886 (N_22886,N_21359,N_21440);
or U22887 (N_22887,N_21034,N_21760);
xnor U22888 (N_22888,N_21088,N_21911);
nor U22889 (N_22889,N_21323,N_20384);
xnor U22890 (N_22890,N_20486,N_20238);
or U22891 (N_22891,N_20397,N_21993);
xnor U22892 (N_22892,N_21758,N_20044);
xor U22893 (N_22893,N_21432,N_20271);
nand U22894 (N_22894,N_21845,N_21798);
or U22895 (N_22895,N_21012,N_21027);
nand U22896 (N_22896,N_21019,N_20644);
xnor U22897 (N_22897,N_21881,N_20465);
or U22898 (N_22898,N_20414,N_20428);
nand U22899 (N_22899,N_20230,N_21933);
and U22900 (N_22900,N_21936,N_20102);
or U22901 (N_22901,N_20248,N_20130);
and U22902 (N_22902,N_21423,N_20410);
nor U22903 (N_22903,N_20760,N_20007);
nand U22904 (N_22904,N_21008,N_20877);
or U22905 (N_22905,N_21990,N_20436);
or U22906 (N_22906,N_20402,N_21378);
and U22907 (N_22907,N_20787,N_20649);
and U22908 (N_22908,N_20591,N_21757);
nor U22909 (N_22909,N_21564,N_21613);
nand U22910 (N_22910,N_21966,N_20624);
nand U22911 (N_22911,N_20249,N_20807);
nand U22912 (N_22912,N_20234,N_21369);
and U22913 (N_22913,N_21633,N_20997);
or U22914 (N_22914,N_21819,N_20933);
and U22915 (N_22915,N_20708,N_21904);
xnor U22916 (N_22916,N_21123,N_20783);
xor U22917 (N_22917,N_21846,N_20265);
xor U22918 (N_22918,N_21922,N_20073);
nand U22919 (N_22919,N_21550,N_20955);
xor U22920 (N_22920,N_21219,N_21927);
nand U22921 (N_22921,N_20698,N_20890);
nand U22922 (N_22922,N_21326,N_21638);
or U22923 (N_22923,N_21060,N_21038);
nand U22924 (N_22924,N_21978,N_21987);
and U22925 (N_22925,N_21453,N_20253);
or U22926 (N_22926,N_20568,N_20934);
nand U22927 (N_22927,N_21755,N_21586);
and U22928 (N_22928,N_20605,N_20023);
nand U22929 (N_22929,N_21853,N_20284);
and U22930 (N_22930,N_20041,N_21298);
or U22931 (N_22931,N_21521,N_21529);
nand U22932 (N_22932,N_21015,N_20456);
xnor U22933 (N_22933,N_21581,N_20907);
or U22934 (N_22934,N_20496,N_21421);
nand U22935 (N_22935,N_21305,N_21511);
nor U22936 (N_22936,N_21025,N_21131);
or U22937 (N_22937,N_20280,N_20906);
nor U22938 (N_22938,N_20801,N_21950);
nor U22939 (N_22939,N_21477,N_21932);
nor U22940 (N_22940,N_20349,N_21279);
nor U22941 (N_22941,N_21747,N_20554);
and U22942 (N_22942,N_21610,N_20640);
and U22943 (N_22943,N_20477,N_21857);
and U22944 (N_22944,N_20178,N_20516);
and U22945 (N_22945,N_20376,N_20703);
and U22946 (N_22946,N_20406,N_20341);
xor U22947 (N_22947,N_21216,N_20596);
xnor U22948 (N_22948,N_21752,N_21370);
nor U22949 (N_22949,N_21598,N_21467);
xor U22950 (N_22950,N_20227,N_21502);
and U22951 (N_22951,N_21418,N_20878);
or U22952 (N_22952,N_20095,N_20868);
xor U22953 (N_22953,N_20723,N_21996);
nor U22954 (N_22954,N_20886,N_21975);
nand U22955 (N_22955,N_21364,N_21574);
nor U22956 (N_22956,N_20574,N_20734);
and U22957 (N_22957,N_21653,N_21170);
nor U22958 (N_22958,N_21754,N_20395);
nand U22959 (N_22959,N_21944,N_20771);
and U22960 (N_22960,N_21282,N_21720);
and U22961 (N_22961,N_20135,N_21865);
xor U22962 (N_22962,N_20203,N_20914);
nor U22963 (N_22963,N_20646,N_21863);
xnor U22964 (N_22964,N_21394,N_21331);
or U22965 (N_22965,N_20779,N_21191);
xnor U22966 (N_22966,N_20511,N_20499);
or U22967 (N_22967,N_20590,N_20191);
xor U22968 (N_22968,N_20572,N_21621);
nand U22969 (N_22969,N_21260,N_21295);
nor U22970 (N_22970,N_20560,N_21280);
nor U22971 (N_22971,N_20808,N_21205);
xor U22972 (N_22972,N_20524,N_21482);
nand U22973 (N_22973,N_20844,N_20751);
nor U22974 (N_22974,N_20991,N_21307);
or U22975 (N_22975,N_21952,N_21789);
and U22976 (N_22976,N_20533,N_21831);
nand U22977 (N_22977,N_21742,N_20307);
nor U22978 (N_22978,N_20966,N_20919);
nor U22979 (N_22979,N_21059,N_21036);
xor U22980 (N_22980,N_21631,N_21473);
nor U22981 (N_22981,N_21444,N_21270);
and U22982 (N_22982,N_20637,N_20841);
and U22983 (N_22983,N_21722,N_21196);
and U22984 (N_22984,N_20651,N_20773);
nand U22985 (N_22985,N_21622,N_20270);
nor U22986 (N_22986,N_20098,N_20122);
and U22987 (N_22987,N_20085,N_21575);
and U22988 (N_22988,N_20232,N_20581);
xor U22989 (N_22989,N_20816,N_21771);
nand U22990 (N_22990,N_20842,N_21528);
or U22991 (N_22991,N_21970,N_21373);
nand U22992 (N_22992,N_21775,N_20528);
nand U22993 (N_22993,N_20663,N_21121);
nand U22994 (N_22994,N_21463,N_21317);
and U22995 (N_22995,N_21645,N_20448);
or U22996 (N_22996,N_21417,N_21997);
xor U22997 (N_22997,N_21227,N_20254);
nor U22998 (N_22998,N_20975,N_20235);
or U22999 (N_22999,N_20784,N_20432);
xnor U23000 (N_23000,N_21473,N_21011);
and U23001 (N_23001,N_21969,N_20208);
nor U23002 (N_23002,N_21078,N_20866);
and U23003 (N_23003,N_21096,N_21457);
nor U23004 (N_23004,N_20709,N_20233);
nand U23005 (N_23005,N_21666,N_21121);
nor U23006 (N_23006,N_21003,N_21111);
xnor U23007 (N_23007,N_20376,N_20331);
xor U23008 (N_23008,N_21544,N_20439);
and U23009 (N_23009,N_21236,N_21615);
nand U23010 (N_23010,N_20241,N_21126);
xor U23011 (N_23011,N_21498,N_20522);
and U23012 (N_23012,N_20031,N_21606);
nand U23013 (N_23013,N_20872,N_20081);
xor U23014 (N_23014,N_20657,N_20581);
or U23015 (N_23015,N_20585,N_20483);
xnor U23016 (N_23016,N_20168,N_20064);
xnor U23017 (N_23017,N_20825,N_20231);
xnor U23018 (N_23018,N_20329,N_21900);
nand U23019 (N_23019,N_20261,N_21860);
nor U23020 (N_23020,N_21629,N_20423);
nor U23021 (N_23021,N_21066,N_21363);
xnor U23022 (N_23022,N_21724,N_21391);
and U23023 (N_23023,N_21456,N_20103);
nor U23024 (N_23024,N_20098,N_21675);
or U23025 (N_23025,N_20986,N_20047);
nor U23026 (N_23026,N_20315,N_20629);
nor U23027 (N_23027,N_20717,N_20750);
xor U23028 (N_23028,N_21610,N_21231);
and U23029 (N_23029,N_21373,N_21944);
nor U23030 (N_23030,N_20762,N_20823);
xnor U23031 (N_23031,N_21948,N_21251);
or U23032 (N_23032,N_21354,N_20816);
nand U23033 (N_23033,N_21987,N_20679);
or U23034 (N_23034,N_20047,N_21284);
and U23035 (N_23035,N_21421,N_21289);
or U23036 (N_23036,N_20656,N_20488);
or U23037 (N_23037,N_20845,N_21603);
nor U23038 (N_23038,N_20031,N_20663);
and U23039 (N_23039,N_20709,N_21618);
nand U23040 (N_23040,N_21836,N_20891);
xor U23041 (N_23041,N_21557,N_21469);
nand U23042 (N_23042,N_20786,N_20444);
or U23043 (N_23043,N_20100,N_21181);
xor U23044 (N_23044,N_20434,N_20700);
and U23045 (N_23045,N_21971,N_20836);
and U23046 (N_23046,N_20539,N_20795);
or U23047 (N_23047,N_20708,N_21314);
and U23048 (N_23048,N_20748,N_20426);
and U23049 (N_23049,N_20342,N_20951);
or U23050 (N_23050,N_20084,N_20218);
xnor U23051 (N_23051,N_20241,N_21270);
xor U23052 (N_23052,N_20663,N_20389);
or U23053 (N_23053,N_21731,N_21887);
nand U23054 (N_23054,N_21942,N_21613);
nor U23055 (N_23055,N_21566,N_21339);
xnor U23056 (N_23056,N_20565,N_21925);
and U23057 (N_23057,N_20893,N_20354);
nor U23058 (N_23058,N_21519,N_21385);
and U23059 (N_23059,N_20623,N_20709);
and U23060 (N_23060,N_20751,N_21568);
or U23061 (N_23061,N_21292,N_21744);
or U23062 (N_23062,N_21219,N_21102);
nor U23063 (N_23063,N_20302,N_21031);
nand U23064 (N_23064,N_20392,N_20310);
or U23065 (N_23065,N_20109,N_21654);
nor U23066 (N_23066,N_20034,N_21801);
and U23067 (N_23067,N_20412,N_21308);
nand U23068 (N_23068,N_21785,N_21852);
xor U23069 (N_23069,N_21326,N_20520);
or U23070 (N_23070,N_21549,N_21916);
and U23071 (N_23071,N_21223,N_20282);
xor U23072 (N_23072,N_21335,N_21667);
nand U23073 (N_23073,N_20664,N_20805);
and U23074 (N_23074,N_21023,N_20127);
and U23075 (N_23075,N_20042,N_21430);
nor U23076 (N_23076,N_20586,N_21226);
or U23077 (N_23077,N_21588,N_21906);
and U23078 (N_23078,N_21894,N_21930);
or U23079 (N_23079,N_20422,N_20011);
nor U23080 (N_23080,N_20787,N_21606);
or U23081 (N_23081,N_20484,N_20179);
or U23082 (N_23082,N_20900,N_20162);
or U23083 (N_23083,N_21030,N_21047);
nand U23084 (N_23084,N_20681,N_21764);
xnor U23085 (N_23085,N_21782,N_21072);
and U23086 (N_23086,N_20548,N_21580);
nand U23087 (N_23087,N_21555,N_21349);
and U23088 (N_23088,N_21248,N_21986);
xnor U23089 (N_23089,N_21186,N_21363);
xor U23090 (N_23090,N_21996,N_20288);
nand U23091 (N_23091,N_21915,N_21354);
xnor U23092 (N_23092,N_20112,N_20071);
xnor U23093 (N_23093,N_21047,N_20481);
nor U23094 (N_23094,N_21449,N_21808);
or U23095 (N_23095,N_21481,N_20768);
nand U23096 (N_23096,N_21745,N_21622);
xor U23097 (N_23097,N_20359,N_21782);
and U23098 (N_23098,N_21686,N_20523);
nand U23099 (N_23099,N_21059,N_21106);
nand U23100 (N_23100,N_20363,N_21206);
nor U23101 (N_23101,N_21398,N_21693);
or U23102 (N_23102,N_20680,N_20322);
nand U23103 (N_23103,N_20324,N_20563);
nand U23104 (N_23104,N_21895,N_21620);
and U23105 (N_23105,N_21747,N_20024);
xnor U23106 (N_23106,N_20078,N_21150);
nand U23107 (N_23107,N_21529,N_20143);
or U23108 (N_23108,N_20653,N_20802);
xnor U23109 (N_23109,N_21278,N_20468);
and U23110 (N_23110,N_21708,N_20611);
and U23111 (N_23111,N_21041,N_20544);
xnor U23112 (N_23112,N_20563,N_20220);
and U23113 (N_23113,N_20579,N_21633);
and U23114 (N_23114,N_21304,N_21915);
nor U23115 (N_23115,N_20111,N_20751);
xor U23116 (N_23116,N_21244,N_20317);
or U23117 (N_23117,N_20978,N_21418);
or U23118 (N_23118,N_21434,N_20872);
or U23119 (N_23119,N_21064,N_20650);
nand U23120 (N_23120,N_21935,N_20242);
nand U23121 (N_23121,N_20360,N_21417);
nor U23122 (N_23122,N_21267,N_21164);
and U23123 (N_23123,N_21310,N_20378);
nand U23124 (N_23124,N_21543,N_21285);
nor U23125 (N_23125,N_21146,N_21055);
nor U23126 (N_23126,N_21597,N_21122);
nand U23127 (N_23127,N_21313,N_20650);
nand U23128 (N_23128,N_20564,N_21603);
nor U23129 (N_23129,N_20172,N_21115);
and U23130 (N_23130,N_21295,N_20380);
xnor U23131 (N_23131,N_21924,N_21407);
xnor U23132 (N_23132,N_20097,N_20039);
nand U23133 (N_23133,N_21301,N_20863);
or U23134 (N_23134,N_20659,N_20866);
nand U23135 (N_23135,N_20865,N_21026);
xor U23136 (N_23136,N_21495,N_21773);
nand U23137 (N_23137,N_20111,N_21129);
xor U23138 (N_23138,N_21798,N_21405);
and U23139 (N_23139,N_21535,N_20262);
or U23140 (N_23140,N_20390,N_20616);
or U23141 (N_23141,N_20921,N_21868);
nand U23142 (N_23142,N_20606,N_20637);
nor U23143 (N_23143,N_20727,N_20972);
xnor U23144 (N_23144,N_21047,N_20259);
and U23145 (N_23145,N_20460,N_21169);
xor U23146 (N_23146,N_20291,N_21664);
nand U23147 (N_23147,N_21111,N_20611);
and U23148 (N_23148,N_21164,N_21109);
or U23149 (N_23149,N_20135,N_21898);
nor U23150 (N_23150,N_20803,N_21997);
xor U23151 (N_23151,N_21973,N_20441);
nor U23152 (N_23152,N_21591,N_21384);
nand U23153 (N_23153,N_21037,N_20226);
nand U23154 (N_23154,N_20397,N_20074);
or U23155 (N_23155,N_21775,N_21302);
or U23156 (N_23156,N_20956,N_21358);
xnor U23157 (N_23157,N_20144,N_21495);
nor U23158 (N_23158,N_20210,N_20129);
nand U23159 (N_23159,N_20441,N_21103);
or U23160 (N_23160,N_21832,N_21544);
or U23161 (N_23161,N_20682,N_21268);
or U23162 (N_23162,N_21450,N_21275);
nand U23163 (N_23163,N_20694,N_21134);
nand U23164 (N_23164,N_20890,N_20116);
and U23165 (N_23165,N_20343,N_21825);
nand U23166 (N_23166,N_21585,N_20110);
or U23167 (N_23167,N_20383,N_21072);
nand U23168 (N_23168,N_20350,N_21118);
and U23169 (N_23169,N_21468,N_21079);
or U23170 (N_23170,N_20125,N_20565);
nand U23171 (N_23171,N_20840,N_20907);
and U23172 (N_23172,N_20514,N_20580);
nor U23173 (N_23173,N_21290,N_20708);
and U23174 (N_23174,N_20487,N_21286);
nand U23175 (N_23175,N_21082,N_21095);
nand U23176 (N_23176,N_21473,N_20821);
nand U23177 (N_23177,N_20331,N_21367);
and U23178 (N_23178,N_20851,N_20383);
nor U23179 (N_23179,N_20939,N_21564);
xnor U23180 (N_23180,N_21000,N_21462);
nand U23181 (N_23181,N_20505,N_21046);
nor U23182 (N_23182,N_20904,N_21150);
nand U23183 (N_23183,N_20746,N_21354);
nand U23184 (N_23184,N_21218,N_21786);
xor U23185 (N_23185,N_20167,N_20711);
nand U23186 (N_23186,N_20278,N_20816);
or U23187 (N_23187,N_21989,N_21101);
nor U23188 (N_23188,N_21892,N_21296);
xnor U23189 (N_23189,N_20622,N_21854);
xor U23190 (N_23190,N_20160,N_20673);
nor U23191 (N_23191,N_21345,N_20122);
and U23192 (N_23192,N_20983,N_21908);
or U23193 (N_23193,N_20708,N_20379);
nor U23194 (N_23194,N_21663,N_21725);
nand U23195 (N_23195,N_21818,N_20580);
and U23196 (N_23196,N_20441,N_21356);
or U23197 (N_23197,N_20494,N_21883);
and U23198 (N_23198,N_21675,N_21990);
or U23199 (N_23199,N_21740,N_21539);
or U23200 (N_23200,N_20366,N_20151);
nand U23201 (N_23201,N_20622,N_20234);
or U23202 (N_23202,N_21426,N_20750);
xnor U23203 (N_23203,N_21747,N_21044);
nor U23204 (N_23204,N_21347,N_20171);
or U23205 (N_23205,N_21745,N_20026);
nand U23206 (N_23206,N_21152,N_21358);
or U23207 (N_23207,N_20873,N_20458);
nor U23208 (N_23208,N_20918,N_20593);
or U23209 (N_23209,N_21542,N_21444);
nand U23210 (N_23210,N_21509,N_20535);
nor U23211 (N_23211,N_20293,N_20717);
nor U23212 (N_23212,N_21067,N_20515);
xor U23213 (N_23213,N_20262,N_21372);
or U23214 (N_23214,N_21969,N_21622);
or U23215 (N_23215,N_20173,N_20735);
and U23216 (N_23216,N_21966,N_20217);
nor U23217 (N_23217,N_21698,N_21099);
and U23218 (N_23218,N_21768,N_20110);
or U23219 (N_23219,N_20674,N_20732);
xor U23220 (N_23220,N_21091,N_21893);
or U23221 (N_23221,N_20040,N_21145);
and U23222 (N_23222,N_20437,N_21676);
or U23223 (N_23223,N_20737,N_20119);
or U23224 (N_23224,N_20940,N_20204);
and U23225 (N_23225,N_21446,N_20114);
or U23226 (N_23226,N_21994,N_21757);
nor U23227 (N_23227,N_20014,N_21280);
nand U23228 (N_23228,N_20285,N_21907);
nand U23229 (N_23229,N_21730,N_21802);
nand U23230 (N_23230,N_20417,N_20198);
nand U23231 (N_23231,N_21128,N_21865);
xnor U23232 (N_23232,N_21725,N_20456);
nor U23233 (N_23233,N_21063,N_20571);
nand U23234 (N_23234,N_21366,N_20284);
xor U23235 (N_23235,N_20572,N_20635);
nand U23236 (N_23236,N_20026,N_20060);
nand U23237 (N_23237,N_21564,N_21145);
and U23238 (N_23238,N_20522,N_21381);
and U23239 (N_23239,N_21435,N_20371);
nand U23240 (N_23240,N_20544,N_21335);
nand U23241 (N_23241,N_21144,N_20168);
and U23242 (N_23242,N_20324,N_21757);
xor U23243 (N_23243,N_20977,N_21933);
nor U23244 (N_23244,N_20371,N_20400);
nor U23245 (N_23245,N_20114,N_21679);
or U23246 (N_23246,N_21093,N_21640);
nand U23247 (N_23247,N_21143,N_20372);
or U23248 (N_23248,N_21166,N_20343);
xor U23249 (N_23249,N_20739,N_20964);
or U23250 (N_23250,N_20612,N_21137);
xnor U23251 (N_23251,N_21582,N_20651);
nand U23252 (N_23252,N_20190,N_21917);
xnor U23253 (N_23253,N_21099,N_21276);
and U23254 (N_23254,N_21661,N_21081);
and U23255 (N_23255,N_21039,N_20296);
or U23256 (N_23256,N_20086,N_20413);
and U23257 (N_23257,N_21634,N_21629);
and U23258 (N_23258,N_20365,N_20441);
nand U23259 (N_23259,N_20139,N_20661);
nand U23260 (N_23260,N_20922,N_21261);
nor U23261 (N_23261,N_20238,N_20132);
or U23262 (N_23262,N_21990,N_20085);
xor U23263 (N_23263,N_20369,N_21800);
xnor U23264 (N_23264,N_21495,N_21799);
xor U23265 (N_23265,N_21795,N_21275);
and U23266 (N_23266,N_20869,N_21936);
xor U23267 (N_23267,N_21859,N_21142);
nor U23268 (N_23268,N_21728,N_20690);
and U23269 (N_23269,N_20169,N_20534);
or U23270 (N_23270,N_20403,N_20788);
or U23271 (N_23271,N_21085,N_20660);
nand U23272 (N_23272,N_20160,N_20943);
nor U23273 (N_23273,N_20210,N_20836);
and U23274 (N_23274,N_20298,N_20702);
xnor U23275 (N_23275,N_20401,N_20721);
or U23276 (N_23276,N_20075,N_20489);
nor U23277 (N_23277,N_20251,N_21293);
or U23278 (N_23278,N_21328,N_20995);
and U23279 (N_23279,N_21939,N_21562);
and U23280 (N_23280,N_21582,N_20318);
nand U23281 (N_23281,N_21344,N_21724);
nand U23282 (N_23282,N_20997,N_21544);
nand U23283 (N_23283,N_20200,N_20910);
or U23284 (N_23284,N_21641,N_21866);
or U23285 (N_23285,N_21561,N_21997);
nor U23286 (N_23286,N_21542,N_20261);
and U23287 (N_23287,N_20547,N_21902);
or U23288 (N_23288,N_21626,N_21091);
and U23289 (N_23289,N_20397,N_21758);
nor U23290 (N_23290,N_21831,N_21611);
nand U23291 (N_23291,N_21801,N_20938);
nor U23292 (N_23292,N_21151,N_20602);
nor U23293 (N_23293,N_20146,N_21365);
nor U23294 (N_23294,N_21018,N_21244);
or U23295 (N_23295,N_20682,N_21164);
and U23296 (N_23296,N_20058,N_21511);
nor U23297 (N_23297,N_20077,N_20173);
nand U23298 (N_23298,N_20895,N_20929);
and U23299 (N_23299,N_20976,N_21597);
nand U23300 (N_23300,N_21573,N_21216);
nand U23301 (N_23301,N_20756,N_20930);
xnor U23302 (N_23302,N_21234,N_21540);
nand U23303 (N_23303,N_21803,N_20945);
nand U23304 (N_23304,N_20937,N_20561);
nor U23305 (N_23305,N_21934,N_20512);
and U23306 (N_23306,N_21619,N_21932);
nand U23307 (N_23307,N_21395,N_21708);
xor U23308 (N_23308,N_20698,N_21707);
and U23309 (N_23309,N_21648,N_20580);
nand U23310 (N_23310,N_20624,N_20639);
nor U23311 (N_23311,N_20086,N_21761);
or U23312 (N_23312,N_21391,N_20914);
and U23313 (N_23313,N_21750,N_21443);
nand U23314 (N_23314,N_21308,N_21149);
xor U23315 (N_23315,N_20916,N_20550);
nand U23316 (N_23316,N_21506,N_20955);
nand U23317 (N_23317,N_21086,N_21012);
xor U23318 (N_23318,N_21710,N_21611);
or U23319 (N_23319,N_21209,N_20240);
and U23320 (N_23320,N_21625,N_21656);
nand U23321 (N_23321,N_20977,N_20727);
nand U23322 (N_23322,N_20010,N_20827);
xnor U23323 (N_23323,N_20972,N_20476);
xnor U23324 (N_23324,N_21152,N_20745);
or U23325 (N_23325,N_21575,N_20896);
xor U23326 (N_23326,N_20548,N_21994);
nor U23327 (N_23327,N_21091,N_21504);
nand U23328 (N_23328,N_20130,N_20291);
xor U23329 (N_23329,N_21098,N_21864);
xor U23330 (N_23330,N_20355,N_20524);
and U23331 (N_23331,N_21217,N_20818);
xnor U23332 (N_23332,N_21028,N_20894);
nand U23333 (N_23333,N_21334,N_21775);
nand U23334 (N_23334,N_21815,N_21012);
and U23335 (N_23335,N_21283,N_21078);
and U23336 (N_23336,N_20855,N_20725);
and U23337 (N_23337,N_20446,N_21764);
and U23338 (N_23338,N_20517,N_20453);
nor U23339 (N_23339,N_21292,N_21036);
nor U23340 (N_23340,N_20239,N_20552);
and U23341 (N_23341,N_21808,N_21289);
or U23342 (N_23342,N_20735,N_21890);
and U23343 (N_23343,N_20465,N_21335);
xor U23344 (N_23344,N_20817,N_21752);
or U23345 (N_23345,N_20864,N_21530);
and U23346 (N_23346,N_21888,N_20265);
nand U23347 (N_23347,N_21948,N_20230);
nand U23348 (N_23348,N_20836,N_20777);
xnor U23349 (N_23349,N_20936,N_21872);
xnor U23350 (N_23350,N_21982,N_21588);
or U23351 (N_23351,N_21028,N_21537);
or U23352 (N_23352,N_20958,N_20101);
and U23353 (N_23353,N_21973,N_21412);
nand U23354 (N_23354,N_21964,N_20625);
and U23355 (N_23355,N_21269,N_21932);
nor U23356 (N_23356,N_21727,N_20877);
nor U23357 (N_23357,N_20335,N_21069);
xnor U23358 (N_23358,N_20682,N_21616);
xnor U23359 (N_23359,N_21934,N_20396);
or U23360 (N_23360,N_20379,N_20000);
or U23361 (N_23361,N_20109,N_21033);
nand U23362 (N_23362,N_20912,N_21030);
nand U23363 (N_23363,N_20111,N_20368);
or U23364 (N_23364,N_20357,N_20506);
and U23365 (N_23365,N_20243,N_21450);
and U23366 (N_23366,N_20186,N_21183);
xnor U23367 (N_23367,N_20332,N_21728);
and U23368 (N_23368,N_21067,N_21852);
and U23369 (N_23369,N_20179,N_21735);
nor U23370 (N_23370,N_21894,N_20140);
xnor U23371 (N_23371,N_21594,N_20609);
and U23372 (N_23372,N_21805,N_21257);
nand U23373 (N_23373,N_21169,N_21132);
xnor U23374 (N_23374,N_21472,N_21528);
nand U23375 (N_23375,N_20781,N_21583);
or U23376 (N_23376,N_21020,N_20049);
xnor U23377 (N_23377,N_20444,N_21698);
nor U23378 (N_23378,N_20627,N_21640);
or U23379 (N_23379,N_20962,N_20598);
xor U23380 (N_23380,N_20925,N_21686);
nor U23381 (N_23381,N_20825,N_21028);
nor U23382 (N_23382,N_21947,N_20414);
nand U23383 (N_23383,N_20945,N_20979);
nand U23384 (N_23384,N_21448,N_20887);
nor U23385 (N_23385,N_20079,N_20297);
and U23386 (N_23386,N_20167,N_20950);
and U23387 (N_23387,N_21583,N_21727);
xor U23388 (N_23388,N_21110,N_20313);
xor U23389 (N_23389,N_20832,N_21083);
nand U23390 (N_23390,N_20558,N_20769);
or U23391 (N_23391,N_21137,N_21228);
or U23392 (N_23392,N_21519,N_21722);
xnor U23393 (N_23393,N_21589,N_21305);
nand U23394 (N_23394,N_21477,N_21723);
nand U23395 (N_23395,N_21795,N_20216);
xor U23396 (N_23396,N_21839,N_21762);
or U23397 (N_23397,N_20984,N_21660);
and U23398 (N_23398,N_21881,N_20573);
nand U23399 (N_23399,N_21689,N_21153);
nand U23400 (N_23400,N_21842,N_20322);
or U23401 (N_23401,N_20539,N_20520);
and U23402 (N_23402,N_20680,N_21240);
nand U23403 (N_23403,N_21567,N_21804);
and U23404 (N_23404,N_20164,N_20771);
nand U23405 (N_23405,N_20443,N_20065);
nand U23406 (N_23406,N_20686,N_21451);
xnor U23407 (N_23407,N_21723,N_21143);
xnor U23408 (N_23408,N_21630,N_21331);
or U23409 (N_23409,N_20521,N_20425);
and U23410 (N_23410,N_20281,N_21819);
xnor U23411 (N_23411,N_20024,N_20448);
and U23412 (N_23412,N_20798,N_21771);
and U23413 (N_23413,N_20373,N_20774);
and U23414 (N_23414,N_20959,N_20829);
or U23415 (N_23415,N_21484,N_20623);
xor U23416 (N_23416,N_20449,N_21159);
or U23417 (N_23417,N_21113,N_21462);
xnor U23418 (N_23418,N_20293,N_20777);
or U23419 (N_23419,N_20028,N_21529);
nor U23420 (N_23420,N_20033,N_20369);
nor U23421 (N_23421,N_20384,N_20052);
nor U23422 (N_23422,N_20413,N_20883);
nand U23423 (N_23423,N_20003,N_21423);
or U23424 (N_23424,N_21203,N_21652);
and U23425 (N_23425,N_21587,N_21651);
and U23426 (N_23426,N_20999,N_20955);
nor U23427 (N_23427,N_20316,N_20928);
and U23428 (N_23428,N_21056,N_21589);
xor U23429 (N_23429,N_21693,N_21390);
and U23430 (N_23430,N_20283,N_21750);
and U23431 (N_23431,N_21998,N_21080);
xor U23432 (N_23432,N_21297,N_20908);
and U23433 (N_23433,N_21258,N_20442);
xor U23434 (N_23434,N_20307,N_21998);
or U23435 (N_23435,N_21578,N_20771);
nor U23436 (N_23436,N_20342,N_21616);
nor U23437 (N_23437,N_21378,N_20549);
or U23438 (N_23438,N_21013,N_20014);
xor U23439 (N_23439,N_20643,N_20467);
nand U23440 (N_23440,N_21684,N_21609);
nor U23441 (N_23441,N_21727,N_21173);
and U23442 (N_23442,N_21823,N_21943);
nand U23443 (N_23443,N_20796,N_20576);
or U23444 (N_23444,N_20677,N_20302);
and U23445 (N_23445,N_21149,N_21072);
xor U23446 (N_23446,N_20944,N_20204);
and U23447 (N_23447,N_21983,N_21785);
xnor U23448 (N_23448,N_20622,N_21366);
and U23449 (N_23449,N_20337,N_20649);
xnor U23450 (N_23450,N_20040,N_20012);
and U23451 (N_23451,N_20758,N_20916);
and U23452 (N_23452,N_21552,N_20700);
nor U23453 (N_23453,N_20564,N_21465);
nor U23454 (N_23454,N_20758,N_20433);
nand U23455 (N_23455,N_21946,N_20982);
nand U23456 (N_23456,N_20748,N_21567);
nand U23457 (N_23457,N_20287,N_20757);
or U23458 (N_23458,N_20925,N_20259);
nor U23459 (N_23459,N_20330,N_20630);
nand U23460 (N_23460,N_21394,N_21007);
xor U23461 (N_23461,N_21290,N_21249);
and U23462 (N_23462,N_20237,N_21328);
and U23463 (N_23463,N_21762,N_20390);
nor U23464 (N_23464,N_20571,N_20388);
or U23465 (N_23465,N_20013,N_21933);
and U23466 (N_23466,N_20131,N_21858);
nand U23467 (N_23467,N_20304,N_21337);
nor U23468 (N_23468,N_21433,N_20655);
and U23469 (N_23469,N_20694,N_20583);
nand U23470 (N_23470,N_20113,N_20929);
xnor U23471 (N_23471,N_21551,N_21983);
nor U23472 (N_23472,N_20991,N_21748);
or U23473 (N_23473,N_20285,N_20823);
nor U23474 (N_23474,N_20971,N_20217);
nor U23475 (N_23475,N_20997,N_21062);
or U23476 (N_23476,N_21849,N_20321);
or U23477 (N_23477,N_21661,N_21772);
or U23478 (N_23478,N_21067,N_20721);
xor U23479 (N_23479,N_21493,N_20006);
nor U23480 (N_23480,N_21980,N_21889);
nor U23481 (N_23481,N_21439,N_20349);
xnor U23482 (N_23482,N_20757,N_21672);
nand U23483 (N_23483,N_21863,N_21876);
nor U23484 (N_23484,N_21416,N_20397);
nor U23485 (N_23485,N_20563,N_20048);
nor U23486 (N_23486,N_21565,N_21039);
or U23487 (N_23487,N_21499,N_21061);
xor U23488 (N_23488,N_21728,N_21286);
nor U23489 (N_23489,N_20982,N_20817);
and U23490 (N_23490,N_21395,N_20159);
xor U23491 (N_23491,N_21585,N_20045);
or U23492 (N_23492,N_20962,N_21548);
and U23493 (N_23493,N_21645,N_20027);
xnor U23494 (N_23494,N_20072,N_21069);
xor U23495 (N_23495,N_20500,N_21640);
nand U23496 (N_23496,N_21350,N_20219);
xor U23497 (N_23497,N_21355,N_21818);
nor U23498 (N_23498,N_20657,N_20534);
nor U23499 (N_23499,N_20689,N_21064);
nor U23500 (N_23500,N_20652,N_20768);
nor U23501 (N_23501,N_20099,N_21054);
or U23502 (N_23502,N_20084,N_20645);
xor U23503 (N_23503,N_21450,N_20108);
or U23504 (N_23504,N_20573,N_20967);
or U23505 (N_23505,N_20938,N_21981);
and U23506 (N_23506,N_20526,N_21834);
nand U23507 (N_23507,N_21302,N_20191);
nor U23508 (N_23508,N_21975,N_20308);
nand U23509 (N_23509,N_21111,N_21329);
nand U23510 (N_23510,N_20356,N_20263);
xor U23511 (N_23511,N_21490,N_20083);
xnor U23512 (N_23512,N_20869,N_20823);
nor U23513 (N_23513,N_21216,N_20845);
xnor U23514 (N_23514,N_21678,N_20715);
nor U23515 (N_23515,N_20590,N_21293);
nand U23516 (N_23516,N_20298,N_20334);
and U23517 (N_23517,N_20823,N_21096);
nor U23518 (N_23518,N_21309,N_21434);
or U23519 (N_23519,N_20850,N_20714);
nand U23520 (N_23520,N_21925,N_20556);
nand U23521 (N_23521,N_20101,N_20519);
xnor U23522 (N_23522,N_20975,N_21275);
nor U23523 (N_23523,N_20727,N_20103);
xnor U23524 (N_23524,N_21460,N_20808);
or U23525 (N_23525,N_20545,N_20770);
nand U23526 (N_23526,N_21048,N_20330);
nor U23527 (N_23527,N_21663,N_20748);
nor U23528 (N_23528,N_20879,N_20358);
nor U23529 (N_23529,N_20783,N_21011);
or U23530 (N_23530,N_20885,N_20452);
nand U23531 (N_23531,N_20935,N_21455);
or U23532 (N_23532,N_21817,N_20002);
or U23533 (N_23533,N_21720,N_20735);
xor U23534 (N_23534,N_21889,N_20014);
or U23535 (N_23535,N_21750,N_21015);
nand U23536 (N_23536,N_21330,N_20414);
and U23537 (N_23537,N_21648,N_21570);
or U23538 (N_23538,N_20679,N_20470);
nand U23539 (N_23539,N_20063,N_21143);
or U23540 (N_23540,N_20755,N_21147);
and U23541 (N_23541,N_20329,N_20497);
xor U23542 (N_23542,N_20493,N_20379);
or U23543 (N_23543,N_20569,N_21944);
nor U23544 (N_23544,N_21020,N_20172);
or U23545 (N_23545,N_20803,N_21465);
and U23546 (N_23546,N_21831,N_20083);
or U23547 (N_23547,N_21722,N_21744);
xnor U23548 (N_23548,N_21123,N_21614);
and U23549 (N_23549,N_21669,N_21147);
or U23550 (N_23550,N_20649,N_21319);
xor U23551 (N_23551,N_20798,N_20777);
or U23552 (N_23552,N_21007,N_20552);
nor U23553 (N_23553,N_21234,N_20228);
and U23554 (N_23554,N_20497,N_21498);
and U23555 (N_23555,N_21194,N_21331);
or U23556 (N_23556,N_20409,N_20556);
nand U23557 (N_23557,N_21316,N_21709);
and U23558 (N_23558,N_20758,N_21741);
nand U23559 (N_23559,N_20996,N_21608);
xnor U23560 (N_23560,N_20828,N_21957);
and U23561 (N_23561,N_20780,N_21305);
xnor U23562 (N_23562,N_20369,N_21566);
nand U23563 (N_23563,N_21811,N_21516);
or U23564 (N_23564,N_20323,N_20804);
xor U23565 (N_23565,N_21168,N_21396);
xnor U23566 (N_23566,N_20231,N_21946);
or U23567 (N_23567,N_21362,N_21167);
nand U23568 (N_23568,N_20202,N_20458);
xor U23569 (N_23569,N_21036,N_20148);
and U23570 (N_23570,N_20162,N_20888);
xnor U23571 (N_23571,N_21856,N_20470);
and U23572 (N_23572,N_20709,N_20796);
nor U23573 (N_23573,N_21883,N_20151);
xor U23574 (N_23574,N_20395,N_20127);
and U23575 (N_23575,N_21402,N_21093);
xnor U23576 (N_23576,N_20481,N_21236);
xnor U23577 (N_23577,N_21241,N_21296);
and U23578 (N_23578,N_20523,N_21342);
xnor U23579 (N_23579,N_20629,N_20193);
xnor U23580 (N_23580,N_20236,N_21040);
xnor U23581 (N_23581,N_21038,N_20123);
or U23582 (N_23582,N_21398,N_20333);
and U23583 (N_23583,N_20359,N_20811);
nor U23584 (N_23584,N_20164,N_20253);
xor U23585 (N_23585,N_21033,N_21877);
and U23586 (N_23586,N_20786,N_21981);
xor U23587 (N_23587,N_20308,N_21421);
or U23588 (N_23588,N_21616,N_20010);
nor U23589 (N_23589,N_20539,N_20038);
or U23590 (N_23590,N_20945,N_20106);
or U23591 (N_23591,N_20206,N_20470);
or U23592 (N_23592,N_20910,N_20062);
and U23593 (N_23593,N_20616,N_21430);
nor U23594 (N_23594,N_21221,N_20330);
xnor U23595 (N_23595,N_20961,N_21150);
xor U23596 (N_23596,N_20777,N_20530);
or U23597 (N_23597,N_21251,N_21479);
or U23598 (N_23598,N_20734,N_21737);
nor U23599 (N_23599,N_20797,N_20436);
nand U23600 (N_23600,N_20082,N_21104);
nand U23601 (N_23601,N_21497,N_20639);
xor U23602 (N_23602,N_20293,N_21001);
or U23603 (N_23603,N_21784,N_21378);
or U23604 (N_23604,N_21042,N_20555);
and U23605 (N_23605,N_21098,N_21262);
or U23606 (N_23606,N_20454,N_21406);
nand U23607 (N_23607,N_21816,N_21079);
xnor U23608 (N_23608,N_21655,N_21635);
xnor U23609 (N_23609,N_21030,N_21049);
nor U23610 (N_23610,N_20593,N_20910);
and U23611 (N_23611,N_21866,N_21002);
nand U23612 (N_23612,N_20476,N_21885);
xnor U23613 (N_23613,N_20407,N_20775);
nand U23614 (N_23614,N_20525,N_20235);
or U23615 (N_23615,N_21108,N_21731);
nand U23616 (N_23616,N_21718,N_21439);
and U23617 (N_23617,N_21165,N_21536);
nand U23618 (N_23618,N_20126,N_20368);
or U23619 (N_23619,N_20570,N_20173);
or U23620 (N_23620,N_21542,N_21963);
nor U23621 (N_23621,N_20365,N_21234);
nand U23622 (N_23622,N_20668,N_20272);
and U23623 (N_23623,N_20637,N_21468);
and U23624 (N_23624,N_20059,N_21725);
nand U23625 (N_23625,N_20540,N_20512);
xnor U23626 (N_23626,N_21453,N_20921);
xor U23627 (N_23627,N_20798,N_20497);
xnor U23628 (N_23628,N_21528,N_20059);
xnor U23629 (N_23629,N_21882,N_21288);
or U23630 (N_23630,N_20403,N_21850);
and U23631 (N_23631,N_21535,N_21755);
xor U23632 (N_23632,N_21062,N_21483);
nor U23633 (N_23633,N_21493,N_21084);
nand U23634 (N_23634,N_21788,N_21956);
xnor U23635 (N_23635,N_20980,N_21899);
xor U23636 (N_23636,N_20869,N_20609);
nand U23637 (N_23637,N_21498,N_20379);
and U23638 (N_23638,N_21857,N_20097);
or U23639 (N_23639,N_20116,N_21809);
and U23640 (N_23640,N_20210,N_20952);
or U23641 (N_23641,N_21598,N_21054);
xor U23642 (N_23642,N_21007,N_20528);
nor U23643 (N_23643,N_20765,N_20953);
xnor U23644 (N_23644,N_21883,N_21071);
and U23645 (N_23645,N_20293,N_20300);
nand U23646 (N_23646,N_21349,N_21692);
and U23647 (N_23647,N_20257,N_21941);
xnor U23648 (N_23648,N_21387,N_21205);
xor U23649 (N_23649,N_20103,N_20479);
nor U23650 (N_23650,N_21390,N_20590);
and U23651 (N_23651,N_21885,N_20607);
nor U23652 (N_23652,N_20733,N_20904);
nand U23653 (N_23653,N_20043,N_21650);
and U23654 (N_23654,N_20146,N_20847);
and U23655 (N_23655,N_20312,N_20957);
xnor U23656 (N_23656,N_21537,N_21650);
nand U23657 (N_23657,N_21231,N_20959);
nor U23658 (N_23658,N_20301,N_21697);
xnor U23659 (N_23659,N_21280,N_20008);
or U23660 (N_23660,N_21671,N_20330);
nand U23661 (N_23661,N_21906,N_20724);
and U23662 (N_23662,N_21692,N_21654);
nor U23663 (N_23663,N_20298,N_20601);
nor U23664 (N_23664,N_21970,N_20235);
or U23665 (N_23665,N_21710,N_21449);
xor U23666 (N_23666,N_21630,N_21067);
and U23667 (N_23667,N_20187,N_20934);
nand U23668 (N_23668,N_21971,N_20239);
and U23669 (N_23669,N_20550,N_21690);
and U23670 (N_23670,N_20815,N_20923);
or U23671 (N_23671,N_20772,N_20838);
xor U23672 (N_23672,N_21212,N_21826);
and U23673 (N_23673,N_21429,N_20880);
nor U23674 (N_23674,N_21749,N_21672);
and U23675 (N_23675,N_20226,N_20764);
xor U23676 (N_23676,N_21737,N_21246);
nand U23677 (N_23677,N_20576,N_21168);
or U23678 (N_23678,N_20529,N_21564);
xnor U23679 (N_23679,N_20367,N_21447);
or U23680 (N_23680,N_20250,N_21072);
or U23681 (N_23681,N_20692,N_20478);
xor U23682 (N_23682,N_20107,N_20879);
xor U23683 (N_23683,N_21444,N_21229);
and U23684 (N_23684,N_21035,N_21463);
nor U23685 (N_23685,N_21528,N_21812);
nor U23686 (N_23686,N_21141,N_20119);
nor U23687 (N_23687,N_21719,N_20062);
xor U23688 (N_23688,N_21250,N_21168);
nor U23689 (N_23689,N_20136,N_20852);
nand U23690 (N_23690,N_21895,N_20243);
nor U23691 (N_23691,N_20241,N_20581);
xnor U23692 (N_23692,N_20618,N_20080);
xor U23693 (N_23693,N_20612,N_20374);
or U23694 (N_23694,N_21686,N_20861);
nor U23695 (N_23695,N_21350,N_21226);
and U23696 (N_23696,N_20782,N_20590);
xnor U23697 (N_23697,N_20536,N_21397);
nor U23698 (N_23698,N_20243,N_20129);
nand U23699 (N_23699,N_21856,N_21772);
nand U23700 (N_23700,N_20655,N_21278);
xor U23701 (N_23701,N_21393,N_20206);
xor U23702 (N_23702,N_20211,N_20773);
nor U23703 (N_23703,N_21958,N_20843);
nand U23704 (N_23704,N_21590,N_21582);
and U23705 (N_23705,N_21711,N_20078);
nand U23706 (N_23706,N_20925,N_20652);
nand U23707 (N_23707,N_21713,N_20296);
or U23708 (N_23708,N_20161,N_21318);
nor U23709 (N_23709,N_21171,N_21208);
nor U23710 (N_23710,N_20837,N_20169);
and U23711 (N_23711,N_20798,N_21236);
or U23712 (N_23712,N_21957,N_20301);
and U23713 (N_23713,N_20529,N_21587);
nand U23714 (N_23714,N_21622,N_20425);
or U23715 (N_23715,N_20099,N_20274);
nand U23716 (N_23716,N_20134,N_21321);
xnor U23717 (N_23717,N_20223,N_21617);
or U23718 (N_23718,N_20873,N_21534);
and U23719 (N_23719,N_21417,N_21391);
and U23720 (N_23720,N_20906,N_21828);
nand U23721 (N_23721,N_21181,N_21402);
nor U23722 (N_23722,N_20867,N_20174);
nand U23723 (N_23723,N_21598,N_21602);
or U23724 (N_23724,N_21882,N_21260);
and U23725 (N_23725,N_20476,N_21407);
nor U23726 (N_23726,N_20540,N_20626);
xnor U23727 (N_23727,N_21453,N_20663);
xnor U23728 (N_23728,N_21902,N_21860);
or U23729 (N_23729,N_21335,N_20327);
xor U23730 (N_23730,N_20837,N_20456);
or U23731 (N_23731,N_21009,N_21238);
or U23732 (N_23732,N_20635,N_21368);
nand U23733 (N_23733,N_20452,N_20935);
nor U23734 (N_23734,N_20382,N_20778);
xnor U23735 (N_23735,N_21532,N_20061);
or U23736 (N_23736,N_21518,N_21271);
or U23737 (N_23737,N_21913,N_21862);
nor U23738 (N_23738,N_20556,N_21051);
or U23739 (N_23739,N_20459,N_20115);
or U23740 (N_23740,N_20427,N_21638);
nor U23741 (N_23741,N_21708,N_20432);
nor U23742 (N_23742,N_20003,N_21444);
nor U23743 (N_23743,N_21335,N_20181);
or U23744 (N_23744,N_21457,N_20396);
and U23745 (N_23745,N_21127,N_20285);
xnor U23746 (N_23746,N_21741,N_20279);
or U23747 (N_23747,N_21363,N_20761);
nand U23748 (N_23748,N_20831,N_21018);
nand U23749 (N_23749,N_20549,N_20859);
nand U23750 (N_23750,N_20246,N_21507);
or U23751 (N_23751,N_20169,N_20142);
nor U23752 (N_23752,N_21050,N_20370);
nand U23753 (N_23753,N_21617,N_20123);
xnor U23754 (N_23754,N_20086,N_21155);
xnor U23755 (N_23755,N_21116,N_20612);
nor U23756 (N_23756,N_20347,N_21910);
or U23757 (N_23757,N_21180,N_20676);
nor U23758 (N_23758,N_20619,N_21226);
or U23759 (N_23759,N_20058,N_20014);
nand U23760 (N_23760,N_20268,N_20343);
nand U23761 (N_23761,N_20796,N_21457);
and U23762 (N_23762,N_20909,N_21226);
xor U23763 (N_23763,N_21374,N_20026);
or U23764 (N_23764,N_21870,N_20208);
or U23765 (N_23765,N_20199,N_21250);
nand U23766 (N_23766,N_20118,N_20453);
xnor U23767 (N_23767,N_21524,N_20007);
xor U23768 (N_23768,N_21369,N_21576);
and U23769 (N_23769,N_21025,N_20940);
nand U23770 (N_23770,N_21969,N_20357);
and U23771 (N_23771,N_21653,N_20365);
nor U23772 (N_23772,N_21321,N_21339);
xor U23773 (N_23773,N_21182,N_21279);
nand U23774 (N_23774,N_20012,N_20366);
or U23775 (N_23775,N_21767,N_20826);
or U23776 (N_23776,N_21013,N_21939);
nor U23777 (N_23777,N_20211,N_20069);
nand U23778 (N_23778,N_20317,N_21298);
or U23779 (N_23779,N_20259,N_21076);
and U23780 (N_23780,N_20185,N_20092);
nor U23781 (N_23781,N_21915,N_20899);
or U23782 (N_23782,N_20270,N_20430);
nand U23783 (N_23783,N_21214,N_20281);
xnor U23784 (N_23784,N_20946,N_20741);
and U23785 (N_23785,N_20250,N_21835);
xor U23786 (N_23786,N_20269,N_20940);
xor U23787 (N_23787,N_21312,N_20274);
xor U23788 (N_23788,N_20893,N_20892);
or U23789 (N_23789,N_21930,N_20159);
nor U23790 (N_23790,N_21159,N_21557);
or U23791 (N_23791,N_20399,N_20190);
or U23792 (N_23792,N_21882,N_21953);
or U23793 (N_23793,N_21850,N_21716);
xor U23794 (N_23794,N_21713,N_20264);
nand U23795 (N_23795,N_20027,N_21330);
xnor U23796 (N_23796,N_21024,N_21092);
nor U23797 (N_23797,N_20946,N_20215);
or U23798 (N_23798,N_20393,N_20208);
nor U23799 (N_23799,N_21388,N_20307);
or U23800 (N_23800,N_21473,N_21711);
nand U23801 (N_23801,N_20989,N_21772);
nor U23802 (N_23802,N_20134,N_20770);
xor U23803 (N_23803,N_20181,N_20328);
and U23804 (N_23804,N_21980,N_20563);
xnor U23805 (N_23805,N_20215,N_21008);
nor U23806 (N_23806,N_21036,N_21214);
xnor U23807 (N_23807,N_21742,N_20796);
or U23808 (N_23808,N_21334,N_20130);
nand U23809 (N_23809,N_20242,N_20438);
or U23810 (N_23810,N_21482,N_20345);
nor U23811 (N_23811,N_20733,N_21745);
xnor U23812 (N_23812,N_21675,N_21567);
nand U23813 (N_23813,N_21243,N_21804);
nand U23814 (N_23814,N_20917,N_20209);
xor U23815 (N_23815,N_20111,N_20031);
and U23816 (N_23816,N_20556,N_21954);
and U23817 (N_23817,N_20215,N_20464);
or U23818 (N_23818,N_20227,N_20221);
and U23819 (N_23819,N_21985,N_21319);
and U23820 (N_23820,N_21971,N_20663);
xor U23821 (N_23821,N_20683,N_21204);
xnor U23822 (N_23822,N_20151,N_20710);
and U23823 (N_23823,N_20034,N_20728);
nand U23824 (N_23824,N_21825,N_20834);
nand U23825 (N_23825,N_20241,N_21732);
xnor U23826 (N_23826,N_21742,N_20489);
nand U23827 (N_23827,N_21257,N_21322);
and U23828 (N_23828,N_20450,N_21585);
xnor U23829 (N_23829,N_20732,N_20079);
xnor U23830 (N_23830,N_21536,N_20389);
nor U23831 (N_23831,N_21101,N_20383);
nand U23832 (N_23832,N_21664,N_20013);
or U23833 (N_23833,N_20207,N_20846);
and U23834 (N_23834,N_21409,N_21804);
nor U23835 (N_23835,N_20036,N_20796);
nor U23836 (N_23836,N_21902,N_20320);
nor U23837 (N_23837,N_21198,N_21325);
nor U23838 (N_23838,N_20705,N_20047);
and U23839 (N_23839,N_21894,N_20628);
xor U23840 (N_23840,N_20361,N_20366);
xor U23841 (N_23841,N_20985,N_20528);
nor U23842 (N_23842,N_21916,N_20210);
or U23843 (N_23843,N_20753,N_20312);
nand U23844 (N_23844,N_20508,N_21220);
and U23845 (N_23845,N_20922,N_21207);
and U23846 (N_23846,N_20266,N_21124);
nor U23847 (N_23847,N_21303,N_21389);
or U23848 (N_23848,N_21952,N_21980);
and U23849 (N_23849,N_20803,N_21228);
nor U23850 (N_23850,N_20388,N_21806);
and U23851 (N_23851,N_20966,N_20842);
and U23852 (N_23852,N_21443,N_21862);
nor U23853 (N_23853,N_21782,N_21588);
nor U23854 (N_23854,N_20456,N_21708);
nor U23855 (N_23855,N_20362,N_20940);
and U23856 (N_23856,N_20938,N_21065);
nand U23857 (N_23857,N_20727,N_20109);
and U23858 (N_23858,N_21936,N_21773);
and U23859 (N_23859,N_21812,N_21340);
nor U23860 (N_23860,N_20945,N_20978);
or U23861 (N_23861,N_21302,N_20421);
and U23862 (N_23862,N_21456,N_21250);
nor U23863 (N_23863,N_20063,N_21592);
and U23864 (N_23864,N_21912,N_20211);
and U23865 (N_23865,N_21405,N_21546);
nand U23866 (N_23866,N_20802,N_20556);
and U23867 (N_23867,N_20555,N_20142);
nand U23868 (N_23868,N_20958,N_21849);
xor U23869 (N_23869,N_21841,N_20197);
nand U23870 (N_23870,N_20381,N_20804);
nand U23871 (N_23871,N_21692,N_21856);
nor U23872 (N_23872,N_21496,N_20137);
xor U23873 (N_23873,N_21515,N_21500);
nor U23874 (N_23874,N_21317,N_20453);
xor U23875 (N_23875,N_20747,N_20200);
and U23876 (N_23876,N_20244,N_21823);
xnor U23877 (N_23877,N_21777,N_21516);
or U23878 (N_23878,N_20458,N_20493);
or U23879 (N_23879,N_20894,N_20720);
nand U23880 (N_23880,N_20485,N_20428);
and U23881 (N_23881,N_20330,N_21318);
or U23882 (N_23882,N_20782,N_21882);
or U23883 (N_23883,N_21573,N_21387);
and U23884 (N_23884,N_21051,N_20669);
nand U23885 (N_23885,N_21198,N_21469);
xor U23886 (N_23886,N_21753,N_20947);
nand U23887 (N_23887,N_21027,N_21461);
or U23888 (N_23888,N_20710,N_21734);
xnor U23889 (N_23889,N_21938,N_21865);
nor U23890 (N_23890,N_20577,N_20627);
nand U23891 (N_23891,N_20487,N_20376);
or U23892 (N_23892,N_20297,N_21083);
or U23893 (N_23893,N_20263,N_20454);
and U23894 (N_23894,N_21369,N_20942);
and U23895 (N_23895,N_20778,N_20091);
and U23896 (N_23896,N_20510,N_21394);
nand U23897 (N_23897,N_20514,N_20887);
nand U23898 (N_23898,N_20504,N_21388);
and U23899 (N_23899,N_21372,N_21884);
nand U23900 (N_23900,N_20941,N_21309);
xnor U23901 (N_23901,N_20963,N_20666);
nand U23902 (N_23902,N_21681,N_20924);
nor U23903 (N_23903,N_20580,N_20901);
and U23904 (N_23904,N_20898,N_21589);
xor U23905 (N_23905,N_20920,N_20298);
nor U23906 (N_23906,N_21786,N_21257);
nand U23907 (N_23907,N_20740,N_21420);
and U23908 (N_23908,N_21437,N_21820);
nor U23909 (N_23909,N_21022,N_20742);
nor U23910 (N_23910,N_21385,N_21613);
nor U23911 (N_23911,N_21162,N_21894);
or U23912 (N_23912,N_21000,N_21333);
xor U23913 (N_23913,N_20970,N_20147);
nor U23914 (N_23914,N_21978,N_20675);
xor U23915 (N_23915,N_21726,N_21357);
xor U23916 (N_23916,N_20815,N_21634);
and U23917 (N_23917,N_21596,N_20613);
and U23918 (N_23918,N_21386,N_21410);
nand U23919 (N_23919,N_21389,N_20887);
or U23920 (N_23920,N_21519,N_20833);
nor U23921 (N_23921,N_20406,N_21469);
nor U23922 (N_23922,N_21578,N_21627);
nor U23923 (N_23923,N_20267,N_21839);
or U23924 (N_23924,N_20501,N_21645);
nor U23925 (N_23925,N_21013,N_21780);
and U23926 (N_23926,N_20912,N_20766);
nor U23927 (N_23927,N_21091,N_20685);
or U23928 (N_23928,N_20421,N_20720);
and U23929 (N_23929,N_20531,N_21689);
xnor U23930 (N_23930,N_21800,N_20997);
and U23931 (N_23931,N_20170,N_21259);
nor U23932 (N_23932,N_21973,N_21063);
xor U23933 (N_23933,N_20901,N_20482);
nor U23934 (N_23934,N_21820,N_21897);
and U23935 (N_23935,N_21219,N_21172);
or U23936 (N_23936,N_20695,N_20587);
nor U23937 (N_23937,N_21318,N_20955);
xor U23938 (N_23938,N_21165,N_20688);
nor U23939 (N_23939,N_20860,N_20504);
nor U23940 (N_23940,N_21807,N_20258);
and U23941 (N_23941,N_21492,N_21354);
nand U23942 (N_23942,N_21194,N_20340);
nor U23943 (N_23943,N_21227,N_21354);
and U23944 (N_23944,N_21509,N_20216);
xor U23945 (N_23945,N_20395,N_21318);
and U23946 (N_23946,N_21135,N_21336);
nand U23947 (N_23947,N_21820,N_20430);
nor U23948 (N_23948,N_20758,N_21679);
and U23949 (N_23949,N_20417,N_20415);
nor U23950 (N_23950,N_20276,N_21892);
and U23951 (N_23951,N_21145,N_20329);
and U23952 (N_23952,N_21494,N_21191);
nor U23953 (N_23953,N_21746,N_21572);
and U23954 (N_23954,N_20249,N_20221);
nor U23955 (N_23955,N_21987,N_21099);
or U23956 (N_23956,N_20181,N_20172);
nor U23957 (N_23957,N_21512,N_21812);
nand U23958 (N_23958,N_20690,N_20423);
nand U23959 (N_23959,N_21219,N_21002);
xor U23960 (N_23960,N_20079,N_20543);
nand U23961 (N_23961,N_20593,N_20396);
nand U23962 (N_23962,N_21023,N_21790);
and U23963 (N_23963,N_20510,N_21447);
and U23964 (N_23964,N_21778,N_20698);
or U23965 (N_23965,N_20349,N_20474);
nand U23966 (N_23966,N_20226,N_20757);
and U23967 (N_23967,N_21486,N_21655);
and U23968 (N_23968,N_21266,N_20617);
nor U23969 (N_23969,N_20859,N_21273);
nand U23970 (N_23970,N_21631,N_21288);
and U23971 (N_23971,N_21865,N_20983);
or U23972 (N_23972,N_20624,N_21859);
xor U23973 (N_23973,N_21330,N_21856);
nor U23974 (N_23974,N_21098,N_20953);
xor U23975 (N_23975,N_20208,N_20833);
nor U23976 (N_23976,N_21610,N_21324);
xnor U23977 (N_23977,N_20333,N_20421);
nor U23978 (N_23978,N_21464,N_20103);
xnor U23979 (N_23979,N_21189,N_21966);
nor U23980 (N_23980,N_20899,N_20496);
nor U23981 (N_23981,N_20125,N_20649);
or U23982 (N_23982,N_21133,N_21544);
xor U23983 (N_23983,N_20840,N_21771);
nor U23984 (N_23984,N_21939,N_21540);
nand U23985 (N_23985,N_21742,N_20300);
xor U23986 (N_23986,N_20900,N_20580);
and U23987 (N_23987,N_21420,N_21030);
xor U23988 (N_23988,N_21825,N_20732);
and U23989 (N_23989,N_20324,N_21463);
or U23990 (N_23990,N_20038,N_20436);
and U23991 (N_23991,N_20831,N_20810);
nor U23992 (N_23992,N_20842,N_20868);
or U23993 (N_23993,N_20874,N_20166);
or U23994 (N_23994,N_21412,N_20574);
xnor U23995 (N_23995,N_21138,N_21408);
nor U23996 (N_23996,N_21132,N_21989);
nor U23997 (N_23997,N_20959,N_21061);
or U23998 (N_23998,N_21102,N_21960);
nand U23999 (N_23999,N_20523,N_20950);
xor U24000 (N_24000,N_22985,N_22130);
nor U24001 (N_24001,N_22378,N_22305);
nand U24002 (N_24002,N_22835,N_22541);
xnor U24003 (N_24003,N_22781,N_23852);
nand U24004 (N_24004,N_22940,N_23017);
nor U24005 (N_24005,N_22685,N_23492);
or U24006 (N_24006,N_23599,N_22884);
xnor U24007 (N_24007,N_22692,N_22244);
nand U24008 (N_24008,N_22280,N_22261);
nand U24009 (N_24009,N_23483,N_23983);
or U24010 (N_24010,N_22028,N_23523);
and U24011 (N_24011,N_22135,N_22599);
xor U24012 (N_24012,N_22777,N_22732);
or U24013 (N_24013,N_23952,N_23662);
or U24014 (N_24014,N_23358,N_23682);
nor U24015 (N_24015,N_22089,N_22990);
xnor U24016 (N_24016,N_22441,N_23762);
nand U24017 (N_24017,N_23761,N_23420);
nor U24018 (N_24018,N_22399,N_22639);
and U24019 (N_24019,N_23873,N_22537);
xor U24020 (N_24020,N_23688,N_22375);
and U24021 (N_24021,N_23512,N_22314);
or U24022 (N_24022,N_23959,N_22512);
or U24023 (N_24023,N_22726,N_22859);
and U24024 (N_24024,N_23602,N_23767);
xor U24025 (N_24025,N_23713,N_22741);
nand U24026 (N_24026,N_23985,N_22914);
nand U24027 (N_24027,N_23047,N_23435);
and U24028 (N_24028,N_23151,N_23223);
xnor U24029 (N_24029,N_22418,N_22501);
nor U24030 (N_24030,N_22307,N_23920);
xnor U24031 (N_24031,N_22576,N_23575);
or U24032 (N_24032,N_22191,N_22768);
nand U24033 (N_24033,N_23166,N_23617);
nor U24034 (N_24034,N_22572,N_22344);
nor U24035 (N_24035,N_22707,N_23993);
and U24036 (N_24036,N_22054,N_23621);
nor U24037 (N_24037,N_22025,N_23604);
or U24038 (N_24038,N_22247,N_22640);
xnor U24039 (N_24039,N_22225,N_23659);
and U24040 (N_24040,N_22531,N_22704);
nor U24041 (N_24041,N_22604,N_22571);
or U24042 (N_24042,N_23708,N_22747);
xnor U24043 (N_24043,N_23600,N_22624);
or U24044 (N_24044,N_22535,N_23516);
nand U24045 (N_24045,N_23109,N_22429);
and U24046 (N_24046,N_22632,N_23350);
or U24047 (N_24047,N_23697,N_22578);
and U24048 (N_24048,N_22878,N_23215);
and U24049 (N_24049,N_23302,N_23172);
nor U24050 (N_24050,N_23861,N_23637);
xnor U24051 (N_24051,N_23149,N_22478);
nand U24052 (N_24052,N_22053,N_23179);
nor U24053 (N_24053,N_22434,N_22162);
nand U24054 (N_24054,N_23609,N_22829);
or U24055 (N_24055,N_22543,N_22310);
and U24056 (N_24056,N_22118,N_22839);
nand U24057 (N_24057,N_22352,N_22950);
xnor U24058 (N_24058,N_23676,N_22547);
nor U24059 (N_24059,N_22407,N_23209);
or U24060 (N_24060,N_23954,N_22754);
or U24061 (N_24061,N_23967,N_22023);
nor U24062 (N_24062,N_22350,N_23772);
xnor U24063 (N_24063,N_23913,N_22369);
xor U24064 (N_24064,N_22461,N_22855);
and U24065 (N_24065,N_22708,N_22973);
nor U24066 (N_24066,N_23564,N_23860);
nor U24067 (N_24067,N_23737,N_22979);
nand U24068 (N_24068,N_23468,N_22984);
nand U24069 (N_24069,N_23125,N_23670);
nand U24070 (N_24070,N_23187,N_22511);
nor U24071 (N_24071,N_23042,N_23392);
nor U24072 (N_24072,N_22267,N_22913);
nor U24073 (N_24073,N_23606,N_22619);
xor U24074 (N_24074,N_23283,N_23155);
and U24075 (N_24075,N_23494,N_23411);
nand U24076 (N_24076,N_22390,N_23982);
and U24077 (N_24077,N_23856,N_22893);
nand U24078 (N_24078,N_23890,N_22313);
and U24079 (N_24079,N_23072,N_22200);
nor U24080 (N_24080,N_23243,N_22129);
and U24081 (N_24081,N_22076,N_23196);
or U24082 (N_24082,N_22532,N_22816);
xnor U24083 (N_24083,N_22966,N_23778);
nor U24084 (N_24084,N_22096,N_23629);
nor U24085 (N_24085,N_22733,N_23165);
nand U24086 (N_24086,N_22084,N_23934);
xor U24087 (N_24087,N_22909,N_22231);
nor U24088 (N_24088,N_23539,N_23971);
xnor U24089 (N_24089,N_23990,N_23603);
or U24090 (N_24090,N_23769,N_22046);
nand U24091 (N_24091,N_22370,N_23784);
and U24092 (N_24092,N_23807,N_22981);
nand U24093 (N_24093,N_22653,N_23069);
or U24094 (N_24094,N_22018,N_22479);
or U24095 (N_24095,N_22103,N_23693);
or U24096 (N_24096,N_22204,N_23672);
nor U24097 (N_24097,N_23324,N_23396);
nor U24098 (N_24098,N_22301,N_22083);
and U24099 (N_24099,N_23686,N_22652);
and U24100 (N_24100,N_23844,N_22651);
nor U24101 (N_24101,N_22097,N_22294);
xor U24102 (N_24102,N_22682,N_23050);
and U24103 (N_24103,N_23244,N_22368);
and U24104 (N_24104,N_22505,N_23889);
nand U24105 (N_24105,N_23063,N_22365);
or U24106 (N_24106,N_23865,N_22110);
nor U24107 (N_24107,N_22630,N_22615);
and U24108 (N_24108,N_22686,N_22299);
nor U24109 (N_24109,N_22150,N_22935);
or U24110 (N_24110,N_22568,N_23286);
xor U24111 (N_24111,N_23430,N_22376);
nor U24112 (N_24112,N_23595,N_23882);
or U24113 (N_24113,N_22219,N_23938);
xor U24114 (N_24114,N_23416,N_23156);
or U24115 (N_24115,N_23611,N_23111);
xor U24116 (N_24116,N_22464,N_22320);
nand U24117 (N_24117,N_22991,N_22870);
nor U24118 (N_24118,N_22166,N_22793);
or U24119 (N_24119,N_23378,N_23267);
and U24120 (N_24120,N_23221,N_22485);
xor U24121 (N_24121,N_23351,N_23858);
or U24122 (N_24122,N_22269,N_22058);
or U24123 (N_24123,N_23746,N_23666);
nand U24124 (N_24124,N_22782,N_23463);
nand U24125 (N_24125,N_22513,N_22260);
and U24126 (N_24126,N_23367,N_22425);
or U24127 (N_24127,N_23946,N_22300);
xor U24128 (N_24128,N_23277,N_22761);
and U24129 (N_24129,N_23241,N_23372);
and U24130 (N_24130,N_23674,N_23306);
nand U24131 (N_24131,N_22798,N_22721);
or U24132 (N_24132,N_23450,N_22493);
or U24133 (N_24133,N_22924,N_23944);
or U24134 (N_24134,N_23871,N_22713);
xor U24135 (N_24135,N_23195,N_23102);
and U24136 (N_24136,N_22032,N_22149);
nand U24137 (N_24137,N_23817,N_23357);
nand U24138 (N_24138,N_22833,N_22767);
nand U24139 (N_24139,N_22437,N_23353);
nor U24140 (N_24140,N_22169,N_22740);
and U24141 (N_24141,N_23783,N_22759);
nand U24142 (N_24142,N_22308,N_23320);
nand U24143 (N_24143,N_22748,N_23691);
and U24144 (N_24144,N_23835,N_22538);
or U24145 (N_24145,N_22549,N_23004);
nor U24146 (N_24146,N_23189,N_22391);
nor U24147 (N_24147,N_23054,N_22820);
and U24148 (N_24148,N_22115,N_22766);
nand U24149 (N_24149,N_23466,N_22423);
xnor U24150 (N_24150,N_22958,N_23660);
nor U24151 (N_24151,N_23768,N_22551);
nor U24152 (N_24152,N_23003,N_22936);
or U24153 (N_24153,N_23675,N_22185);
and U24154 (N_24154,N_22928,N_22451);
or U24155 (N_24155,N_23775,N_22889);
or U24156 (N_24156,N_23405,N_23633);
nor U24157 (N_24157,N_23608,N_22815);
xor U24158 (N_24158,N_23104,N_22021);
xor U24159 (N_24159,N_23044,N_22542);
xnor U24160 (N_24160,N_22736,N_22163);
nor U24161 (N_24161,N_23265,N_22447);
nor U24162 (N_24162,N_22142,N_23936);
xor U24163 (N_24163,N_23082,N_22837);
and U24164 (N_24164,N_23643,N_22643);
nor U24165 (N_24165,N_22003,N_22047);
xor U24166 (N_24166,N_22265,N_22373);
or U24167 (N_24167,N_22845,N_22088);
xor U24168 (N_24168,N_22232,N_23118);
nand U24169 (N_24169,N_23458,N_22670);
and U24170 (N_24170,N_22005,N_22172);
nor U24171 (N_24171,N_22976,N_23425);
and U24172 (N_24172,N_23041,N_23878);
xor U24173 (N_24173,N_23526,N_23587);
nor U24174 (N_24174,N_22016,N_23549);
xor U24175 (N_24175,N_22916,N_22671);
nor U24176 (N_24176,N_22211,N_22540);
nand U24177 (N_24177,N_23665,N_23016);
xor U24178 (N_24178,N_23544,N_23311);
nor U24179 (N_24179,N_23089,N_22738);
and U24180 (N_24180,N_23304,N_23412);
nor U24181 (N_24181,N_22846,N_22679);
and U24182 (N_24182,N_23780,N_23798);
and U24183 (N_24183,N_22031,N_23057);
nand U24184 (N_24184,N_23359,N_22421);
nor U24185 (N_24185,N_22044,N_23777);
or U24186 (N_24186,N_22156,N_23476);
and U24187 (N_24187,N_23825,N_23640);
nand U24188 (N_24188,N_22729,N_23730);
or U24189 (N_24189,N_23487,N_22459);
xnor U24190 (N_24190,N_22108,N_22949);
nand U24191 (N_24191,N_22631,N_23218);
nand U24192 (N_24192,N_22330,N_22471);
and U24193 (N_24193,N_23256,N_22710);
nand U24194 (N_24194,N_23178,N_22903);
or U24195 (N_24195,N_22959,N_23510);
and U24196 (N_24196,N_23576,N_22457);
xnor U24197 (N_24197,N_23153,N_22298);
and U24198 (N_24198,N_22011,N_22687);
nand U24199 (N_24199,N_23143,N_23380);
xnor U24200 (N_24200,N_23441,N_23885);
and U24201 (N_24201,N_22050,N_23011);
nand U24202 (N_24202,N_22151,N_22943);
and U24203 (N_24203,N_23554,N_22817);
nor U24204 (N_24204,N_22797,N_22220);
nand U24205 (N_24205,N_22205,N_22324);
and U24206 (N_24206,N_22545,N_23075);
nor U24207 (N_24207,N_22109,N_23655);
and U24208 (N_24208,N_22414,N_22771);
and U24209 (N_24209,N_22024,N_22270);
nor U24210 (N_24210,N_22987,N_22450);
or U24211 (N_24211,N_23915,N_22198);
or U24212 (N_24212,N_22873,N_22483);
xnor U24213 (N_24213,N_22069,N_22379);
and U24214 (N_24214,N_22992,N_23532);
or U24215 (N_24215,N_22847,N_23386);
xnor U24216 (N_24216,N_23091,N_23584);
nand U24217 (N_24217,N_23771,N_22051);
xor U24218 (N_24218,N_22467,N_22562);
nor U24219 (N_24219,N_23354,N_22802);
nor U24220 (N_24220,N_23800,N_23360);
nand U24221 (N_24221,N_23428,N_23826);
xor U24222 (N_24222,N_23446,N_22408);
and U24223 (N_24223,N_22811,N_22867);
nand U24224 (N_24224,N_23028,N_22857);
and U24225 (N_24225,N_23181,N_22625);
or U24226 (N_24226,N_22393,N_23384);
nand U24227 (N_24227,N_22674,N_23269);
and U24228 (N_24228,N_22287,N_23725);
xor U24229 (N_24229,N_22203,N_22402);
or U24230 (N_24230,N_22794,N_23126);
xnor U24231 (N_24231,N_22406,N_22477);
or U24232 (N_24232,N_22645,N_22312);
or U24233 (N_24233,N_22090,N_22251);
nand U24234 (N_24234,N_23872,N_22720);
nor U24235 (N_24235,N_22361,N_23830);
xnor U24236 (N_24236,N_22932,N_23094);
nand U24237 (N_24237,N_22500,N_22877);
nand U24238 (N_24238,N_23619,N_23315);
nor U24239 (N_24239,N_23741,N_22711);
or U24240 (N_24240,N_22607,N_22977);
nand U24241 (N_24241,N_22502,N_23563);
or U24242 (N_24242,N_22519,N_23188);
xnor U24243 (N_24243,N_22061,N_23142);
and U24244 (N_24244,N_23081,N_23454);
and U24245 (N_24245,N_22623,N_23939);
nand U24246 (N_24246,N_22947,N_22929);
and U24247 (N_24247,N_23432,N_23793);
and U24248 (N_24248,N_22481,N_23170);
xnor U24249 (N_24249,N_23719,N_22286);
nor U24250 (N_24250,N_23711,N_23689);
and U24251 (N_24251,N_22799,N_22517);
and U24252 (N_24252,N_22552,N_23018);
and U24253 (N_24253,N_22331,N_23912);
or U24254 (N_24254,N_22642,N_23698);
and U24255 (N_24255,N_23816,N_23369);
nor U24256 (N_24256,N_23052,N_23314);
or U24257 (N_24257,N_22066,N_22259);
nor U24258 (N_24258,N_23438,N_23226);
or U24259 (N_24259,N_22161,N_23524);
xnor U24260 (N_24260,N_23298,N_22258);
nor U24261 (N_24261,N_22875,N_22214);
nor U24262 (N_24262,N_23064,N_23870);
or U24263 (N_24263,N_23043,N_23339);
and U24264 (N_24264,N_23904,N_22941);
nand U24265 (N_24265,N_22480,N_23853);
or U24266 (N_24266,N_22342,N_23199);
or U24267 (N_24267,N_23007,N_23884);
xnor U24268 (N_24268,N_22667,N_23429);
nor U24269 (N_24269,N_22444,N_22760);
xnor U24270 (N_24270,N_23121,N_23914);
nor U24271 (N_24271,N_23289,N_22460);
nand U24272 (N_24272,N_23085,N_23998);
nand U24273 (N_24273,N_22487,N_23203);
nand U24274 (N_24274,N_22114,N_23514);
nor U24275 (N_24275,N_23397,N_22275);
nand U24276 (N_24276,N_23424,N_23841);
nand U24277 (N_24277,N_23467,N_22001);
or U24278 (N_24278,N_22188,N_22174);
nor U24279 (N_24279,N_22718,N_22957);
xor U24280 (N_24280,N_23211,N_22473);
and U24281 (N_24281,N_23900,N_23902);
and U24282 (N_24282,N_23293,N_23399);
or U24283 (N_24283,N_22779,N_22919);
nand U24284 (N_24284,N_22888,N_23377);
xor U24285 (N_24285,N_23418,N_23035);
or U24286 (N_24286,N_22605,N_23832);
or U24287 (N_24287,N_23796,N_23403);
nor U24288 (N_24288,N_23908,N_23667);
nor U24289 (N_24289,N_23930,N_22019);
nor U24290 (N_24290,N_23183,N_23374);
nand U24291 (N_24291,N_23079,N_23076);
and U24292 (N_24292,N_23947,N_23477);
xnor U24293 (N_24293,N_22579,N_23225);
or U24294 (N_24294,N_23319,N_22925);
and U24295 (N_24295,N_23417,N_23144);
or U24296 (N_24296,N_23014,N_23005);
xnor U24297 (N_24297,N_22222,N_23994);
and U24298 (N_24298,N_23543,N_23597);
and U24299 (N_24299,N_22693,N_22567);
xor U24300 (N_24300,N_22548,N_22911);
xnor U24301 (N_24301,N_23250,N_22073);
nand U24302 (N_24302,N_22918,N_23519);
xnor U24303 (N_24303,N_23799,N_23231);
xor U24304 (N_24304,N_22117,N_23536);
or U24305 (N_24305,N_23823,N_22577);
xnor U24306 (N_24306,N_22742,N_22327);
xor U24307 (N_24307,N_22648,N_23127);
and U24308 (N_24308,N_23864,N_22183);
xor U24309 (N_24309,N_22785,N_23336);
or U24310 (N_24310,N_22250,N_23831);
nand U24311 (N_24311,N_23677,N_22539);
or U24312 (N_24312,N_22589,N_23220);
and U24313 (N_24313,N_23026,N_22297);
or U24314 (N_24314,N_23452,N_23135);
nor U24315 (N_24315,N_22601,N_23961);
and U24316 (N_24316,N_23055,N_22049);
nor U24317 (N_24317,N_23486,N_22676);
nand U24318 (N_24318,N_23238,N_22696);
xnor U24319 (N_24319,N_23820,N_23132);
nor U24320 (N_24320,N_23586,N_23918);
nand U24321 (N_24321,N_22237,N_23605);
xnor U24322 (N_24322,N_23625,N_23517);
nand U24323 (N_24323,N_22059,N_22284);
and U24324 (N_24324,N_22336,N_22248);
and U24325 (N_24325,N_23006,N_22787);
nand U24326 (N_24326,N_22659,N_22836);
nand U24327 (N_24327,N_23210,N_23242);
nand U24328 (N_24328,N_23090,N_23812);
or U24329 (N_24329,N_22014,N_23036);
xnor U24330 (N_24330,N_22510,N_22585);
xor U24331 (N_24331,N_22806,N_22405);
nor U24332 (N_24332,N_22555,N_22334);
or U24333 (N_24333,N_23236,N_22852);
or U24334 (N_24334,N_23992,N_23909);
xor U24335 (N_24335,N_22348,N_23995);
nand U24336 (N_24336,N_22661,N_23855);
nand U24337 (N_24337,N_23493,N_22784);
nand U24338 (N_24338,N_22235,N_22316);
nor U24339 (N_24339,N_22600,N_23765);
and U24340 (N_24340,N_23426,N_23390);
nand U24341 (N_24341,N_23582,N_23529);
nor U24342 (N_24342,N_22553,N_22234);
and U24343 (N_24343,N_22626,N_23634);
or U24344 (N_24344,N_23099,N_23547);
and U24345 (N_24345,N_23579,N_22879);
nor U24346 (N_24346,N_23347,N_23702);
nor U24347 (N_24347,N_23325,N_23222);
and U24348 (N_24348,N_22930,N_22168);
xnor U24349 (N_24349,N_23182,N_22896);
xnor U24350 (N_24350,N_23840,N_23572);
xnor U24351 (N_24351,N_23837,N_23818);
xor U24352 (N_24352,N_23888,N_23364);
and U24353 (N_24353,N_23124,N_23434);
xnor U24354 (N_24354,N_22106,N_22080);
nand U24355 (N_24355,N_22134,N_22840);
or U24356 (N_24356,N_23001,N_23522);
and U24357 (N_24357,N_23518,N_23177);
xnor U24358 (N_24358,N_22319,N_22484);
nor U24359 (N_24359,N_22524,N_23128);
nor U24360 (N_24360,N_22063,N_23262);
nor U24361 (N_24361,N_22786,N_23112);
nand U24362 (N_24362,N_23999,N_23919);
xor U24363 (N_24363,N_22170,N_22085);
nor U24364 (N_24364,N_22574,N_23440);
xor U24365 (N_24365,N_23048,N_23834);
or U24366 (N_24366,N_22603,N_23857);
and U24367 (N_24367,N_23484,N_22194);
or U24368 (N_24368,N_22999,N_23671);
xnor U24369 (N_24369,N_23694,N_23437);
xnor U24370 (N_24370,N_23246,N_23049);
and U24371 (N_24371,N_23530,N_22560);
and U24372 (N_24372,N_22395,N_22616);
nor U24373 (N_24373,N_22119,N_22566);
and U24374 (N_24374,N_22669,N_23789);
xnor U24375 (N_24375,N_23059,N_22881);
nand U24376 (N_24376,N_22594,N_22431);
and U24377 (N_24377,N_23721,N_22665);
or U24378 (N_24378,N_22443,N_23387);
and U24379 (N_24379,N_22716,N_22008);
xor U24380 (N_24380,N_23577,N_22905);
or U24381 (N_24381,N_23764,N_22995);
or U24382 (N_24382,N_22629,N_23540);
xnor U24383 (N_24383,N_22960,N_23490);
xnor U24384 (N_24384,N_22148,N_22355);
nand U24385 (N_24385,N_23776,N_22303);
nor U24386 (N_24386,N_23457,N_23015);
xor U24387 (N_24387,N_23436,N_22394);
nand U24388 (N_24388,N_23107,N_23239);
nand U24389 (N_24389,N_22217,N_22010);
nor U24390 (N_24390,N_22180,N_23464);
and U24391 (N_24391,N_23804,N_22666);
nor U24392 (N_24392,N_22554,N_22392);
nand U24393 (N_24393,N_22776,N_23080);
nor U24394 (N_24394,N_23453,N_22243);
nor U24395 (N_24395,N_22637,N_23010);
xnor U24396 (N_24396,N_22094,N_22187);
nor U24397 (N_24397,N_23201,N_22963);
xnor U24398 (N_24398,N_22563,N_22725);
xnor U24399 (N_24399,N_23758,N_23976);
xor U24400 (N_24400,N_23499,N_23419);
and U24401 (N_24401,N_23866,N_22606);
nor U24402 (N_24402,N_23025,N_22812);
and U24403 (N_24403,N_23191,N_23652);
xor U24404 (N_24404,N_22831,N_23383);
nor U24405 (N_24405,N_23683,N_23162);
nand U24406 (N_24406,N_23284,N_23021);
or U24407 (N_24407,N_22278,N_22207);
and U24408 (N_24408,N_23555,N_23160);
and U24409 (N_24409,N_22264,N_23973);
xor U24410 (N_24410,N_22842,N_22856);
nand U24411 (N_24411,N_22143,N_22986);
xnor U24412 (N_24412,N_22321,N_22948);
nand U24413 (N_24413,N_23867,N_22364);
or U24414 (N_24414,N_23552,N_22874);
or U24415 (N_24415,N_23363,N_22961);
xor U24416 (N_24416,N_23876,N_23726);
nand U24417 (N_24417,N_23809,N_23745);
and U24418 (N_24418,N_22819,N_22683);
and U24419 (N_24419,N_22416,N_22105);
nand U24420 (N_24420,N_22463,N_22075);
nand U24421 (N_24421,N_23729,N_22614);
and U24422 (N_24422,N_23479,N_22899);
and U24423 (N_24423,N_23657,N_22534);
nor U24424 (N_24424,N_23557,N_22388);
or U24425 (N_24425,N_23471,N_23299);
nand U24426 (N_24426,N_23842,N_23168);
and U24427 (N_24427,N_23718,N_22453);
nor U24428 (N_24428,N_22969,N_23815);
and U24429 (N_24429,N_22681,N_22843);
nand U24430 (N_24430,N_23422,N_23527);
nor U24431 (N_24431,N_22422,N_22801);
xor U24432 (N_24432,N_22848,N_23949);
nand U24433 (N_24433,N_22971,N_22598);
and U24434 (N_24434,N_23092,N_23561);
and U24435 (N_24435,N_23313,N_22488);
nand U24436 (N_24436,N_22673,N_22882);
and U24437 (N_24437,N_22112,N_23098);
xnor U24438 (N_24438,N_23644,N_22951);
and U24439 (N_24439,N_22660,N_22057);
or U24440 (N_24440,N_22609,N_23274);
and U24441 (N_24441,N_22827,N_23271);
xnor U24442 (N_24442,N_23895,N_23308);
xnor U24443 (N_24443,N_23296,N_23774);
or U24444 (N_24444,N_23593,N_23309);
nand U24445 (N_24445,N_22684,N_22730);
nor U24446 (N_24446,N_23559,N_23850);
or U24447 (N_24447,N_23366,N_22347);
or U24448 (N_24448,N_23344,N_23773);
nor U24449 (N_24449,N_22098,N_22153);
and U24450 (N_24450,N_23122,N_22650);
or U24451 (N_24451,N_23445,N_23355);
nand U24452 (N_24452,N_22157,N_23056);
xnor U24453 (N_24453,N_23280,N_23747);
nor U24454 (N_24454,N_23147,N_22055);
xnor U24455 (N_24455,N_22739,N_23491);
and U24456 (N_24456,N_23537,N_23828);
or U24457 (N_24457,N_22077,N_22384);
nand U24458 (N_24458,N_23504,N_22184);
and U24459 (N_24459,N_22082,N_23395);
and U24460 (N_24460,N_22454,N_22672);
and U24461 (N_24461,N_23376,N_22141);
and U24462 (N_24462,N_22715,N_22608);
or U24463 (N_24463,N_22403,N_23928);
xor U24464 (N_24464,N_22830,N_23610);
and U24465 (N_24465,N_22036,N_22382);
and U24466 (N_24466,N_22723,N_23679);
and U24467 (N_24467,N_22689,N_22041);
xor U24468 (N_24468,N_23590,N_22257);
nor U24469 (N_24469,N_22854,N_22868);
and U24470 (N_24470,N_23568,N_23558);
nand U24471 (N_24471,N_23573,N_23008);
nand U24472 (N_24472,N_23779,N_23734);
xor U24473 (N_24473,N_22927,N_22256);
and U24474 (N_24474,N_22807,N_23760);
xnor U24475 (N_24475,N_22751,N_23978);
nand U24476 (N_24476,N_23965,N_22295);
nor U24477 (N_24477,N_23272,N_23507);
nor U24478 (N_24478,N_22351,N_22561);
or U24479 (N_24479,N_23935,N_22952);
and U24480 (N_24480,N_23110,N_22862);
nand U24481 (N_24481,N_22814,N_23498);
xnor U24482 (N_24482,N_22302,N_23839);
or U24483 (N_24483,N_22850,N_23500);
or U24484 (N_24484,N_23788,N_23031);
or U24485 (N_24485,N_22591,N_22937);
and U24486 (N_24486,N_22805,N_23171);
and U24487 (N_24487,N_23233,N_23029);
and U24488 (N_24488,N_23365,N_23120);
nor U24489 (N_24489,N_22292,N_23136);
or U24490 (N_24490,N_22946,N_23700);
nand U24491 (N_24491,N_22417,N_22749);
or U24492 (N_24492,N_22864,N_23381);
or U24493 (N_24493,N_23312,N_22904);
or U24494 (N_24494,N_23455,N_22213);
xor U24495 (N_24495,N_23157,N_23303);
nand U24496 (N_24496,N_22705,N_22627);
nor U24497 (N_24497,N_23066,N_23097);
nand U24498 (N_24498,N_22516,N_22033);
nor U24499 (N_24499,N_22136,N_23343);
nand U24500 (N_24500,N_23404,N_22397);
nand U24501 (N_24501,N_22430,N_22998);
or U24502 (N_24502,N_23134,N_22559);
xor U24503 (N_24503,N_23969,N_22190);
nor U24504 (N_24504,N_23371,N_22332);
or U24505 (N_24505,N_22346,N_23391);
or U24506 (N_24506,N_22590,N_23581);
nor U24507 (N_24507,N_23161,N_23770);
nand U24508 (N_24508,N_22452,N_23329);
and U24509 (N_24509,N_23415,N_23802);
and U24510 (N_24510,N_22289,N_22506);
nor U24511 (N_24511,N_22068,N_22954);
and U24512 (N_24512,N_23742,N_23086);
and U24513 (N_24513,N_22360,N_22769);
nor U24514 (N_24514,N_23032,N_22039);
xnor U24515 (N_24515,N_22339,N_23334);
and U24516 (N_24516,N_23520,N_22849);
nor U24517 (N_24517,N_23521,N_23207);
and U24518 (N_24518,N_22887,N_23923);
nand U24519 (N_24519,N_23307,N_23740);
xor U24520 (N_24520,N_23528,N_23724);
and U24521 (N_24521,N_23687,N_22086);
and U24522 (N_24522,N_23862,N_22714);
and U24523 (N_24523,N_22341,N_22448);
or U24524 (N_24524,N_23950,N_23000);
and U24525 (N_24525,N_23562,N_23270);
nand U24526 (N_24526,N_23851,N_23279);
xnor U24527 (N_24527,N_22030,N_22617);
and U24528 (N_24528,N_22530,N_22139);
nand U24529 (N_24529,N_23553,N_23658);
nand U24530 (N_24530,N_22910,N_22528);
nor U24531 (N_24531,N_22756,N_22886);
or U24532 (N_24532,N_23940,N_22592);
xnor U24533 (N_24533,N_22206,N_22029);
nor U24534 (N_24534,N_22311,N_23907);
xnor U24535 (N_24535,N_22246,N_22872);
nor U24536 (N_24536,N_23893,N_22263);
nand U24537 (N_24537,N_22201,N_22866);
nand U24538 (N_24538,N_22727,N_22853);
xor U24539 (N_24539,N_22268,N_22962);
nand U24540 (N_24540,N_23955,N_23039);
nor U24541 (N_24541,N_23574,N_22439);
or U24542 (N_24542,N_23546,N_23656);
or U24543 (N_24543,N_23316,N_23988);
and U24544 (N_24544,N_22792,N_23152);
xnor U24545 (N_24545,N_22374,N_22424);
nor U24546 (N_24546,N_22009,N_22102);
nor U24547 (N_24547,N_23560,N_22618);
nand U24548 (N_24548,N_23037,N_22389);
and U24549 (N_24549,N_22834,N_23488);
nand U24550 (N_24550,N_22596,N_22647);
nor U24551 (N_24551,N_22508,N_23249);
nor U24552 (N_24552,N_22249,N_23881);
or U24553 (N_24553,N_22492,N_22221);
and U24554 (N_24554,N_22942,N_23409);
and U24555 (N_24555,N_22658,N_23905);
and U24556 (N_24556,N_22209,N_22354);
xnor U24557 (N_24557,N_23827,N_22004);
xor U24558 (N_24558,N_23202,N_23465);
xor U24559 (N_24559,N_23838,N_22012);
nor U24560 (N_24560,N_22610,N_23548);
xnor U24561 (N_24561,N_23744,N_22093);
nand U24562 (N_24562,N_23692,N_22015);
xnor U24563 (N_24563,N_23295,N_23863);
nor U24564 (N_24564,N_22147,N_22433);
nand U24565 (N_24565,N_23154,N_22900);
or U24566 (N_24566,N_23180,N_23074);
xor U24567 (N_24567,N_23328,N_22345);
nand U24568 (N_24568,N_23212,N_23623);
nor U24569 (N_24569,N_23062,N_22734);
and U24570 (N_24570,N_23953,N_23368);
and U24571 (N_24571,N_23894,N_22982);
xor U24572 (N_24572,N_22385,N_23925);
nand U24573 (N_24573,N_22178,N_23123);
or U24574 (N_24574,N_23116,N_23794);
and U24575 (N_24575,N_23846,N_23732);
nor U24576 (N_24576,N_22233,N_22790);
nand U24577 (N_24577,N_22800,N_23093);
xor U24578 (N_24578,N_22173,N_22335);
nor U24579 (N_24579,N_22656,N_22514);
or U24580 (N_24580,N_22271,N_22722);
nor U24581 (N_24581,N_22613,N_22272);
nor U24582 (N_24582,N_23848,N_23264);
nor U24583 (N_24583,N_22529,N_22491);
and U24584 (N_24584,N_23618,N_23073);
and U24585 (N_24585,N_23186,N_23023);
nand U24586 (N_24586,N_22074,N_22367);
xnor U24587 (N_24587,N_22822,N_22703);
nor U24588 (N_24588,N_23245,N_23051);
xor U24589 (N_24589,N_22876,N_23503);
xor U24590 (N_24590,N_22458,N_23591);
nand U24591 (N_24591,N_23678,N_22894);
or U24592 (N_24592,N_23795,N_23485);
nor U24593 (N_24593,N_23991,N_23981);
and U24594 (N_24594,N_22775,N_23663);
and U24595 (N_24595,N_22724,N_22890);
nor U24596 (N_24596,N_23755,N_23892);
or U24597 (N_24597,N_23394,N_22750);
xor U24598 (N_24598,N_22636,N_23184);
nand U24599 (N_24599,N_22757,N_22804);
xnor U24600 (N_24600,N_23506,N_22752);
xnor U24601 (N_24601,N_22241,N_23030);
nand U24602 (N_24602,N_22466,N_23330);
xnor U24603 (N_24603,N_22956,N_22920);
nor U24604 (N_24604,N_23481,N_23261);
nand U24605 (N_24605,N_23717,N_22690);
nor U24606 (N_24606,N_23087,N_22698);
or U24607 (N_24607,N_23903,N_22880);
nor U24608 (N_24608,N_23792,N_22343);
nand U24609 (N_24609,N_23578,N_23534);
or U24610 (N_24610,N_23146,N_23787);
nor U24611 (N_24611,N_23836,N_23647);
xnor U24612 (N_24612,N_22100,N_23766);
nor U24613 (N_24613,N_23948,N_23736);
nand U24614 (N_24614,N_23198,N_22239);
nand U24615 (N_24615,N_22079,N_23664);
nand U24616 (N_24616,N_22586,N_23478);
nor U24617 (N_24617,N_22719,N_22017);
or U24618 (N_24618,N_22527,N_22140);
and U24619 (N_24619,N_22283,N_22953);
and U24620 (N_24620,N_22737,N_23921);
nor U24621 (N_24621,N_22182,N_22897);
and U24622 (N_24622,N_23012,N_22809);
or U24623 (N_24623,N_23106,N_22791);
or U24624 (N_24624,N_23045,N_22497);
xnor U24625 (N_24625,N_23237,N_22869);
or U24626 (N_24626,N_22902,N_22228);
and U24627 (N_24627,N_22037,N_23260);
nand U24628 (N_24628,N_22828,N_22885);
nor U24629 (N_24629,N_23980,N_22359);
xnor U24630 (N_24630,N_23797,N_23868);
or U24631 (N_24631,N_22818,N_22381);
xnor U24632 (N_24632,N_23845,N_22357);
and U24633 (N_24633,N_22580,N_23252);
nand U24634 (N_24634,N_22780,N_23345);
nor U24635 (N_24635,N_23922,N_23349);
xor U24636 (N_24636,N_22242,N_23801);
or U24637 (N_24637,N_22042,N_22199);
or U24638 (N_24638,N_22997,N_23607);
or U24639 (N_24639,N_23984,N_23291);
or U24640 (N_24640,N_22922,N_22620);
nor U24641 (N_24641,N_23701,N_23723);
or U24642 (N_24642,N_22974,N_22588);
nor U24643 (N_24643,N_22655,N_23974);
nand U24644 (N_24644,N_22668,N_22515);
nand U24645 (N_24645,N_23727,N_23373);
or U24646 (N_24646,N_23958,N_23346);
and U24647 (N_24647,N_22821,N_22582);
xnor U24648 (N_24648,N_22764,N_23601);
nor U24649 (N_24649,N_23690,N_22366);
nor U24650 (N_24650,N_23247,N_23630);
or U24651 (N_24651,N_22428,N_23414);
nand U24652 (N_24652,N_23810,N_23635);
or U24653 (N_24653,N_23649,N_23100);
nor U24654 (N_24654,N_22223,N_23943);
nor U24655 (N_24655,N_23615,N_22116);
nor U24656 (N_24656,N_23214,N_22372);
xor U24657 (N_24657,N_22907,N_22641);
nor U24658 (N_24658,N_23229,N_22475);
nor U24659 (N_24659,N_22123,N_22412);
and U24660 (N_24660,N_23883,N_23305);
xnor U24661 (N_24661,N_23388,N_23105);
nor U24662 (N_24662,N_23645,N_22838);
and U24663 (N_24663,N_22013,N_23444);
xor U24664 (N_24664,N_22763,N_22575);
or U24665 (N_24665,N_23987,N_22731);
nand U24666 (N_24666,N_22279,N_22230);
nand U24667 (N_24667,N_23235,N_23714);
nand U24668 (N_24668,N_22933,N_23019);
nor U24669 (N_24669,N_23756,N_22349);
nand U24670 (N_24670,N_23297,N_23133);
and U24671 (N_24671,N_22550,N_23627);
or U24672 (N_24672,N_23164,N_22411);
or U24673 (N_24673,N_23996,N_23699);
or U24674 (N_24674,N_23113,N_23898);
or U24675 (N_24675,N_23227,N_22525);
or U24676 (N_24676,N_23083,N_23096);
nor U24677 (N_24677,N_22062,N_23899);
nor U24678 (N_24678,N_23880,N_23550);
or U24679 (N_24679,N_22197,N_22772);
nor U24680 (N_24680,N_23673,N_22858);
nand U24681 (N_24681,N_22564,N_23803);
or U24682 (N_24682,N_22646,N_23957);
nand U24683 (N_24683,N_23385,N_22121);
or U24684 (N_24684,N_22983,N_23167);
and U24685 (N_24685,N_22252,N_23684);
and U24686 (N_24686,N_23791,N_23977);
or U24687 (N_24687,N_22773,N_22468);
or U24688 (N_24688,N_22810,N_22131);
or U24689 (N_24689,N_23585,N_23200);
or U24690 (N_24690,N_23333,N_23937);
or U24691 (N_24691,N_22254,N_23129);
xor U24692 (N_24692,N_23859,N_22557);
or U24693 (N_24693,N_22544,N_23459);
nand U24694 (N_24694,N_22965,N_23058);
or U24695 (N_24695,N_23034,N_22934);
nand U24696 (N_24696,N_22065,N_22099);
nand U24697 (N_24697,N_22917,N_23781);
xnor U24698 (N_24698,N_23139,N_23228);
xnor U24699 (N_24699,N_23910,N_22224);
or U24700 (N_24700,N_23847,N_23715);
nand U24701 (N_24701,N_23217,N_22165);
and U24702 (N_24702,N_22216,N_22474);
and U24703 (N_24703,N_23703,N_23728);
and U24704 (N_24704,N_23400,N_23638);
xnor U24705 (N_24705,N_23790,N_22276);
nor U24706 (N_24706,N_22227,N_23782);
nand U24707 (N_24707,N_22813,N_22113);
and U24708 (N_24708,N_23230,N_22420);
and U24709 (N_24709,N_22398,N_22509);
nor U24710 (N_24710,N_23456,N_22362);
or U24711 (N_24711,N_22789,N_22104);
or U24712 (N_24712,N_23997,N_23282);
nand U24713 (N_24713,N_22644,N_22634);
and U24714 (N_24714,N_22363,N_22315);
and U24715 (N_24715,N_23989,N_23754);
xor U24716 (N_24716,N_22132,N_22070);
nor U24717 (N_24717,N_22144,N_23067);
xor U24718 (N_24718,N_23566,N_22002);
nand U24719 (N_24719,N_23401,N_23427);
xnor U24720 (N_24720,N_22306,N_23322);
nor U24721 (N_24721,N_23077,N_23716);
nor U24722 (N_24722,N_23323,N_23733);
and U24723 (N_24723,N_23805,N_23495);
xor U24724 (N_24724,N_22520,N_22353);
and U24725 (N_24725,N_22915,N_22449);
or U24726 (N_24726,N_22432,N_23808);
and U24727 (N_24727,N_22126,N_23342);
xnor U24728 (N_24728,N_22383,N_23749);
and U24729 (N_24729,N_22770,N_23194);
or U24730 (N_24730,N_22597,N_22706);
xor U24731 (N_24731,N_22489,N_22462);
nand U24732 (N_24732,N_23275,N_22435);
or U24733 (N_24733,N_22164,N_23571);
nand U24734 (N_24734,N_23046,N_23193);
xnor U24735 (N_24735,N_22583,N_22000);
nand U24736 (N_24736,N_23750,N_22824);
or U24737 (N_24737,N_22633,N_23956);
and U24738 (N_24738,N_23705,N_22883);
and U24739 (N_24739,N_22803,N_23622);
and U24740 (N_24740,N_23174,N_22410);
xor U24741 (N_24741,N_23024,N_23362);
xor U24742 (N_24742,N_23751,N_22240);
or U24743 (N_24743,N_23696,N_22318);
and U24744 (N_24744,N_23158,N_23525);
and U24745 (N_24745,N_22158,N_22753);
and U24746 (N_24746,N_22317,N_22503);
xnor U24747 (N_24747,N_23616,N_22700);
xnor U24748 (N_24748,N_22326,N_22912);
xor U24749 (N_24749,N_22923,N_22052);
or U24750 (N_24750,N_23294,N_23317);
nor U24751 (N_24751,N_22095,N_22413);
and U24752 (N_24752,N_23695,N_22387);
nor U24753 (N_24753,N_22469,N_22678);
nand U24754 (N_24754,N_22701,N_23916);
or U24755 (N_24755,N_23421,N_23874);
or U24756 (N_24756,N_23192,N_23060);
xor U24757 (N_24757,N_22159,N_22386);
or U24758 (N_24758,N_22565,N_23108);
or U24759 (N_24759,N_23541,N_22908);
and U24760 (N_24760,N_23119,N_23763);
nor U24761 (N_24761,N_23743,N_23103);
or U24762 (N_24762,N_22906,N_23101);
nor U24763 (N_24763,N_22944,N_23451);
xor U24764 (N_24764,N_22056,N_22657);
xor U24765 (N_24765,N_23213,N_23931);
nor U24766 (N_24766,N_22419,N_22861);
nor U24767 (N_24767,N_23375,N_22795);
or U24768 (N_24768,N_23963,N_23443);
nand U24769 (N_24769,N_22825,N_23138);
xnor U24770 (N_24770,N_22060,N_23759);
and U24771 (N_24771,N_22891,N_23535);
and U24772 (N_24772,N_22496,N_23497);
xnor U24773 (N_24773,N_23318,N_23786);
or U24774 (N_24774,N_22325,N_23439);
nor U24775 (N_24775,N_23614,N_22978);
or U24776 (N_24776,N_22495,N_23511);
xor U24777 (N_24777,N_22446,N_23009);
xnor U24778 (N_24778,N_23141,N_23542);
or U24779 (N_24779,N_23114,N_23628);
and U24780 (N_24780,N_23338,N_22455);
and U24781 (N_24781,N_22533,N_23070);
or U24782 (N_24782,N_23470,N_23406);
and U24783 (N_24783,N_23588,N_22006);
xor U24784 (N_24784,N_23442,N_22628);
xor U24785 (N_24785,N_22138,N_22111);
and U24786 (N_24786,N_23472,N_22296);
nor U24787 (N_24787,N_23356,N_23824);
nor U24788 (N_24788,N_23653,N_23130);
xnor U24789 (N_24789,N_23408,N_22664);
xor U24790 (N_24790,N_22744,N_22507);
or U24791 (N_24791,N_22975,N_22081);
nor U24792 (N_24792,N_22709,N_22034);
and U24793 (N_24793,N_22155,N_22020);
or U24794 (N_24794,N_23084,N_22035);
and U24795 (N_24795,N_22067,N_23173);
xor U24796 (N_24796,N_22680,N_22078);
xnor U24797 (N_24797,N_23567,N_23869);
xnor U24798 (N_24798,N_22072,N_22593);
and U24799 (N_24799,N_23137,N_22137);
and U24800 (N_24800,N_23620,N_22133);
and U24801 (N_24801,N_23460,N_23505);
nor U24802 (N_24802,N_23911,N_23821);
or U24803 (N_24803,N_22377,N_23206);
nor U24804 (N_24804,N_23720,N_22445);
or U24805 (N_24805,N_22796,N_22175);
or U24806 (N_24806,N_23340,N_23276);
nor U24807 (N_24807,N_22146,N_22765);
and U24808 (N_24808,N_22892,N_23654);
nand U24809 (N_24809,N_22189,N_22945);
or U24810 (N_24810,N_23447,N_23022);
xor U24811 (N_24811,N_23061,N_23583);
xnor U24812 (N_24812,N_22273,N_22573);
xnor U24813 (N_24813,N_22470,N_22436);
or U24814 (N_24814,N_23942,N_23975);
nor U24815 (N_24815,N_22823,N_22027);
or U24816 (N_24816,N_22167,N_22285);
and U24817 (N_24817,N_23475,N_22931);
nand U24818 (N_24818,N_23473,N_22304);
and U24819 (N_24819,N_22404,N_22048);
nand U24820 (N_24820,N_22970,N_23204);
nand U24821 (N_24821,N_22465,N_23945);
and U24822 (N_24822,N_23580,N_22778);
and U24823 (N_24823,N_22196,N_23268);
and U24824 (N_24824,N_23854,N_22699);
or U24825 (N_24825,N_22309,N_22442);
and U24826 (N_24826,N_23932,N_22863);
or U24827 (N_24827,N_23515,N_22415);
or U24828 (N_24828,N_22171,N_23285);
nor U24829 (N_24829,N_23669,N_22808);
xor U24830 (N_24830,N_22176,N_22329);
and U24831 (N_24831,N_23814,N_22556);
and U24832 (N_24832,N_22755,N_22358);
nand U24833 (N_24833,N_23216,N_23962);
nor U24834 (N_24834,N_23175,N_22865);
nand U24835 (N_24835,N_23819,N_23901);
and U24836 (N_24836,N_22939,N_22844);
nand U24837 (N_24837,N_23361,N_22526);
or U24838 (N_24838,N_23020,N_23402);
or U24839 (N_24839,N_23002,N_22340);
or U24840 (N_24840,N_22371,N_22635);
and U24841 (N_24841,N_23917,N_23053);
or U24842 (N_24842,N_23502,N_23288);
and U24843 (N_24843,N_23879,N_22125);
and U24844 (N_24844,N_23639,N_22181);
nand U24845 (N_24845,N_22546,N_23407);
or U24846 (N_24846,N_23169,N_23509);
nor U24847 (N_24847,N_22322,N_22282);
nor U24848 (N_24848,N_23829,N_23849);
nor U24849 (N_24849,N_22026,N_23533);
xor U24850 (N_24850,N_23027,N_22409);
or U24851 (N_24851,N_22145,N_23972);
nor U24852 (N_24852,N_22695,N_23651);
and U24853 (N_24853,N_23331,N_23843);
xor U24854 (N_24854,N_22426,N_23300);
and U24855 (N_24855,N_23941,N_23341);
nor U24856 (N_24856,N_22728,N_23352);
or U24857 (N_24857,N_22602,N_22281);
xor U24858 (N_24858,N_23722,N_22536);
xnor U24859 (N_24859,N_22654,N_23219);
xnor U24860 (N_24860,N_22266,N_22895);
or U24861 (N_24861,N_23624,N_22186);
and U24862 (N_24862,N_23205,N_23327);
or U24863 (N_24863,N_22964,N_22064);
or U24864 (N_24864,N_23140,N_23266);
or U24865 (N_24865,N_22611,N_23661);
xnor U24866 (N_24866,N_22697,N_22456);
xnor U24867 (N_24867,N_23551,N_23569);
nand U24868 (N_24868,N_23731,N_23301);
xor U24869 (N_24869,N_23710,N_22274);
nand U24870 (N_24870,N_22128,N_22482);
xor U24871 (N_24871,N_23190,N_22218);
or U24872 (N_24872,N_23811,N_22955);
nor U24873 (N_24873,N_23641,N_22745);
nand U24874 (N_24874,N_22972,N_22486);
xnor U24875 (N_24875,N_23565,N_23078);
and U24876 (N_24876,N_22774,N_23709);
nand U24877 (N_24877,N_23145,N_22179);
xor U24878 (N_24878,N_23706,N_23933);
and U24879 (N_24879,N_23538,N_22675);
nand U24880 (N_24880,N_23712,N_23248);
nand U24881 (N_24881,N_22255,N_22212);
or U24882 (N_24882,N_22122,N_23095);
and U24883 (N_24883,N_23646,N_22202);
xnor U24884 (N_24884,N_23240,N_23208);
or U24885 (N_24885,N_22622,N_22401);
nor U24886 (N_24886,N_23979,N_23224);
nor U24887 (N_24887,N_23822,N_23513);
nor U24888 (N_24888,N_22226,N_23088);
and U24889 (N_24889,N_23556,N_23273);
nand U24890 (N_24890,N_23813,N_22440);
and U24891 (N_24891,N_23897,N_23642);
nand U24892 (N_24892,N_23065,N_22584);
xor U24893 (N_24893,N_22735,N_22154);
nand U24894 (N_24894,N_22523,N_22438);
nor U24895 (N_24895,N_22968,N_23482);
or U24896 (N_24896,N_22677,N_22788);
and U24897 (N_24897,N_23785,N_22851);
or U24898 (N_24898,N_23148,N_23545);
and U24899 (N_24899,N_23748,N_23176);
nand U24900 (N_24900,N_22262,N_23926);
nor U24901 (N_24901,N_23287,N_23960);
nor U24902 (N_24902,N_22860,N_23806);
and U24903 (N_24903,N_23681,N_22518);
or U24904 (N_24904,N_23131,N_22921);
xnor U24905 (N_24905,N_23480,N_23251);
nand U24906 (N_24906,N_22177,N_22994);
and U24907 (N_24907,N_23163,N_22038);
or U24908 (N_24908,N_23348,N_22688);
and U24909 (N_24909,N_23159,N_22427);
xnor U24910 (N_24910,N_22277,N_22293);
nand U24911 (N_24911,N_23332,N_22236);
nand U24912 (N_24912,N_22253,N_22338);
and U24913 (N_24913,N_22193,N_22087);
xnor U24914 (N_24914,N_23254,N_23068);
nand U24915 (N_24915,N_22926,N_22967);
or U24916 (N_24916,N_23685,N_22522);
xor U24917 (N_24917,N_22356,N_22581);
or U24918 (N_24918,N_23389,N_23197);
and U24919 (N_24919,N_23986,N_22472);
or U24920 (N_24920,N_23924,N_22127);
nand U24921 (N_24921,N_22612,N_23431);
xnor U24922 (N_24922,N_23281,N_22717);
xnor U24923 (N_24923,N_23648,N_23951);
and U24924 (N_24924,N_22621,N_23757);
nor U24925 (N_24925,N_23234,N_23253);
nand U24926 (N_24926,N_22476,N_23496);
nor U24927 (N_24927,N_22091,N_23589);
and U24928 (N_24928,N_23379,N_22980);
and U24929 (N_24929,N_23598,N_23257);
and U24930 (N_24930,N_23150,N_23594);
nand U24931 (N_24931,N_22988,N_22712);
or U24932 (N_24932,N_23335,N_23596);
and U24933 (N_24933,N_22758,N_22662);
nor U24934 (N_24934,N_23321,N_23448);
or U24935 (N_24935,N_22107,N_23469);
and U24936 (N_24936,N_22558,N_22989);
nor U24937 (N_24937,N_23461,N_23337);
xnor U24938 (N_24938,N_22071,N_22871);
nand U24939 (N_24939,N_23013,N_22898);
or U24940 (N_24940,N_22043,N_23612);
nand U24941 (N_24941,N_23508,N_23185);
or U24942 (N_24942,N_23449,N_23877);
and U24943 (N_24943,N_23290,N_22746);
nor U24944 (N_24944,N_23680,N_22826);
xor U24945 (N_24945,N_23739,N_22521);
or U24946 (N_24946,N_22663,N_22195);
nor U24947 (N_24947,N_23636,N_22245);
nor U24948 (N_24948,N_22229,N_23891);
nand U24949 (N_24949,N_23531,N_22498);
nor U24950 (N_24950,N_22993,N_23613);
or U24951 (N_24951,N_22160,N_22045);
nor U24952 (N_24952,N_22649,N_23232);
nand U24953 (N_24953,N_22702,N_23263);
xnor U24954 (N_24954,N_22290,N_22337);
or U24955 (N_24955,N_22490,N_23489);
or U24956 (N_24956,N_23326,N_23929);
and U24957 (N_24957,N_23735,N_23398);
and U24958 (N_24958,N_23632,N_22494);
and U24959 (N_24959,N_22208,N_23752);
and U24960 (N_24960,N_22901,N_23370);
and U24961 (N_24961,N_22215,N_23259);
or U24962 (N_24962,N_22504,N_22938);
nand U24963 (N_24963,N_23033,N_23278);
and U24964 (N_24964,N_23393,N_22288);
nor U24965 (N_24965,N_23115,N_22210);
nand U24966 (N_24966,N_22570,N_23117);
or U24967 (N_24967,N_23833,N_22120);
and U24968 (N_24968,N_23258,N_22092);
or U24969 (N_24969,N_22007,N_23707);
xnor U24970 (N_24970,N_22333,N_23906);
xor U24971 (N_24971,N_23927,N_22323);
nand U24972 (N_24972,N_23474,N_22396);
nand U24973 (N_24973,N_22587,N_23704);
nor U24974 (N_24974,N_22691,N_23738);
nand U24975 (N_24975,N_23886,N_23501);
or U24976 (N_24976,N_23038,N_23570);
or U24977 (N_24977,N_22595,N_22499);
nand U24978 (N_24978,N_23423,N_23875);
nor U24979 (N_24979,N_23650,N_23970);
or U24980 (N_24980,N_22152,N_22743);
or U24981 (N_24981,N_23631,N_23462);
and U24982 (N_24982,N_23753,N_23413);
and U24983 (N_24983,N_23382,N_23433);
nand U24984 (N_24984,N_23310,N_22291);
and U24985 (N_24985,N_22124,N_22638);
xnor U24986 (N_24986,N_23626,N_23968);
nor U24987 (N_24987,N_22380,N_23040);
and U24988 (N_24988,N_22040,N_23887);
and U24989 (N_24989,N_22328,N_22569);
and U24990 (N_24990,N_23410,N_22101);
or U24991 (N_24991,N_22022,N_22762);
nand U24992 (N_24992,N_23071,N_22783);
xor U24993 (N_24993,N_23896,N_22841);
and U24994 (N_24994,N_23592,N_23964);
and U24995 (N_24995,N_23966,N_22694);
nor U24996 (N_24996,N_22238,N_22192);
and U24997 (N_24997,N_22996,N_23292);
nor U24998 (N_24998,N_22400,N_23255);
nor U24999 (N_24999,N_23668,N_22832);
xnor U25000 (N_25000,N_23372,N_23079);
nor U25001 (N_25001,N_23208,N_23701);
and U25002 (N_25002,N_22200,N_22429);
nand U25003 (N_25003,N_22438,N_23296);
nor U25004 (N_25004,N_22182,N_23816);
or U25005 (N_25005,N_23837,N_23170);
nor U25006 (N_25006,N_22667,N_23881);
or U25007 (N_25007,N_22368,N_22985);
xor U25008 (N_25008,N_22398,N_23620);
or U25009 (N_25009,N_22513,N_22523);
or U25010 (N_25010,N_22171,N_23384);
or U25011 (N_25011,N_22473,N_23587);
nand U25012 (N_25012,N_22942,N_22081);
or U25013 (N_25013,N_23081,N_23293);
nand U25014 (N_25014,N_22334,N_23541);
and U25015 (N_25015,N_23177,N_22493);
nand U25016 (N_25016,N_22199,N_22520);
or U25017 (N_25017,N_22373,N_22472);
or U25018 (N_25018,N_22434,N_23223);
and U25019 (N_25019,N_23323,N_23342);
nand U25020 (N_25020,N_22623,N_23063);
nand U25021 (N_25021,N_22437,N_22849);
or U25022 (N_25022,N_23748,N_23213);
xnor U25023 (N_25023,N_22009,N_22907);
nor U25024 (N_25024,N_22903,N_23566);
or U25025 (N_25025,N_22729,N_23781);
and U25026 (N_25026,N_23367,N_22524);
or U25027 (N_25027,N_22422,N_23869);
nand U25028 (N_25028,N_22569,N_22358);
and U25029 (N_25029,N_23444,N_22452);
nand U25030 (N_25030,N_22762,N_22457);
nand U25031 (N_25031,N_22351,N_22792);
xor U25032 (N_25032,N_23355,N_23363);
or U25033 (N_25033,N_23985,N_23657);
or U25034 (N_25034,N_23152,N_23250);
nor U25035 (N_25035,N_23666,N_22156);
and U25036 (N_25036,N_22477,N_22482);
xor U25037 (N_25037,N_22711,N_22134);
nor U25038 (N_25038,N_22777,N_23607);
nand U25039 (N_25039,N_23020,N_23994);
nor U25040 (N_25040,N_22646,N_23460);
nand U25041 (N_25041,N_23171,N_22801);
and U25042 (N_25042,N_23414,N_23649);
xor U25043 (N_25043,N_23870,N_22405);
or U25044 (N_25044,N_23670,N_22883);
and U25045 (N_25045,N_23664,N_22264);
xnor U25046 (N_25046,N_23986,N_23480);
xnor U25047 (N_25047,N_22306,N_22804);
and U25048 (N_25048,N_22303,N_22458);
xnor U25049 (N_25049,N_22157,N_23544);
and U25050 (N_25050,N_23448,N_23536);
nand U25051 (N_25051,N_23620,N_23288);
nor U25052 (N_25052,N_22120,N_22694);
xor U25053 (N_25053,N_22435,N_22657);
or U25054 (N_25054,N_22831,N_23830);
or U25055 (N_25055,N_23625,N_22475);
nor U25056 (N_25056,N_23196,N_22414);
or U25057 (N_25057,N_22954,N_22420);
or U25058 (N_25058,N_23208,N_22028);
nand U25059 (N_25059,N_23584,N_23620);
or U25060 (N_25060,N_23082,N_23173);
nand U25061 (N_25061,N_22238,N_22064);
and U25062 (N_25062,N_23830,N_23959);
or U25063 (N_25063,N_22408,N_22543);
nand U25064 (N_25064,N_22337,N_23882);
nor U25065 (N_25065,N_22093,N_22481);
or U25066 (N_25066,N_22557,N_22984);
and U25067 (N_25067,N_23354,N_23738);
and U25068 (N_25068,N_22899,N_22339);
nand U25069 (N_25069,N_22945,N_23370);
or U25070 (N_25070,N_23162,N_22570);
or U25071 (N_25071,N_23691,N_22999);
and U25072 (N_25072,N_22687,N_23705);
nor U25073 (N_25073,N_22774,N_22596);
nand U25074 (N_25074,N_23790,N_22678);
or U25075 (N_25075,N_22297,N_22347);
nand U25076 (N_25076,N_23382,N_23223);
nor U25077 (N_25077,N_22298,N_23638);
or U25078 (N_25078,N_22802,N_22000);
nor U25079 (N_25079,N_23735,N_22632);
xor U25080 (N_25080,N_22363,N_22372);
and U25081 (N_25081,N_23352,N_23419);
nor U25082 (N_25082,N_22878,N_22237);
nand U25083 (N_25083,N_23980,N_22512);
and U25084 (N_25084,N_23158,N_23973);
or U25085 (N_25085,N_23995,N_22235);
and U25086 (N_25086,N_22308,N_22484);
nor U25087 (N_25087,N_22781,N_23326);
nand U25088 (N_25088,N_22301,N_23830);
xnor U25089 (N_25089,N_22638,N_22969);
or U25090 (N_25090,N_23224,N_22370);
xnor U25091 (N_25091,N_22264,N_22366);
nand U25092 (N_25092,N_23881,N_23268);
and U25093 (N_25093,N_23578,N_23296);
or U25094 (N_25094,N_22306,N_22998);
nand U25095 (N_25095,N_23044,N_23201);
nor U25096 (N_25096,N_23540,N_22253);
and U25097 (N_25097,N_23854,N_22489);
nor U25098 (N_25098,N_22638,N_22951);
nand U25099 (N_25099,N_22567,N_22842);
and U25100 (N_25100,N_23674,N_22575);
or U25101 (N_25101,N_22493,N_23830);
xnor U25102 (N_25102,N_23643,N_23614);
and U25103 (N_25103,N_22334,N_23928);
or U25104 (N_25104,N_22313,N_22134);
nor U25105 (N_25105,N_22822,N_23957);
and U25106 (N_25106,N_22238,N_22081);
nor U25107 (N_25107,N_22987,N_23105);
nor U25108 (N_25108,N_22335,N_23436);
nor U25109 (N_25109,N_23443,N_23142);
nor U25110 (N_25110,N_22782,N_22544);
or U25111 (N_25111,N_23876,N_22331);
xnor U25112 (N_25112,N_23282,N_22152);
nand U25113 (N_25113,N_23098,N_22135);
xor U25114 (N_25114,N_22099,N_23043);
xnor U25115 (N_25115,N_23719,N_23164);
nor U25116 (N_25116,N_22988,N_22234);
nor U25117 (N_25117,N_22745,N_23925);
nor U25118 (N_25118,N_22121,N_23821);
or U25119 (N_25119,N_22288,N_23606);
nor U25120 (N_25120,N_22714,N_23914);
xor U25121 (N_25121,N_23241,N_22386);
nor U25122 (N_25122,N_22075,N_22741);
nand U25123 (N_25123,N_23854,N_23997);
or U25124 (N_25124,N_23825,N_23693);
nand U25125 (N_25125,N_22820,N_23053);
nor U25126 (N_25126,N_23420,N_22865);
and U25127 (N_25127,N_23887,N_23089);
xnor U25128 (N_25128,N_23854,N_23911);
nor U25129 (N_25129,N_22498,N_22223);
nand U25130 (N_25130,N_23871,N_23227);
or U25131 (N_25131,N_23417,N_23420);
nor U25132 (N_25132,N_23801,N_22833);
nor U25133 (N_25133,N_23924,N_22233);
nand U25134 (N_25134,N_23920,N_23897);
nor U25135 (N_25135,N_22408,N_23665);
and U25136 (N_25136,N_23405,N_23472);
nor U25137 (N_25137,N_22085,N_23529);
and U25138 (N_25138,N_22112,N_22924);
and U25139 (N_25139,N_22814,N_22011);
and U25140 (N_25140,N_23975,N_23126);
and U25141 (N_25141,N_22368,N_22389);
and U25142 (N_25142,N_23297,N_22452);
or U25143 (N_25143,N_22334,N_23687);
nand U25144 (N_25144,N_22191,N_22222);
and U25145 (N_25145,N_23855,N_22559);
xnor U25146 (N_25146,N_23227,N_22629);
or U25147 (N_25147,N_23528,N_23295);
nand U25148 (N_25148,N_22363,N_23855);
nor U25149 (N_25149,N_22773,N_22586);
xor U25150 (N_25150,N_23502,N_23138);
nor U25151 (N_25151,N_22845,N_22529);
nand U25152 (N_25152,N_22578,N_22401);
and U25153 (N_25153,N_23261,N_23366);
and U25154 (N_25154,N_23728,N_23262);
or U25155 (N_25155,N_23780,N_23883);
or U25156 (N_25156,N_23145,N_23758);
xnor U25157 (N_25157,N_22231,N_23302);
or U25158 (N_25158,N_23115,N_23684);
or U25159 (N_25159,N_23796,N_22021);
nand U25160 (N_25160,N_23804,N_22400);
nand U25161 (N_25161,N_22994,N_23998);
and U25162 (N_25162,N_23101,N_23754);
nand U25163 (N_25163,N_23198,N_22340);
xnor U25164 (N_25164,N_23881,N_23328);
nor U25165 (N_25165,N_22144,N_23759);
nor U25166 (N_25166,N_22354,N_22018);
xor U25167 (N_25167,N_22926,N_23145);
nor U25168 (N_25168,N_23740,N_23874);
nand U25169 (N_25169,N_22403,N_22716);
xor U25170 (N_25170,N_22405,N_23124);
xnor U25171 (N_25171,N_23635,N_22853);
and U25172 (N_25172,N_22284,N_23712);
nand U25173 (N_25173,N_22867,N_23764);
or U25174 (N_25174,N_22562,N_23991);
or U25175 (N_25175,N_22727,N_23970);
and U25176 (N_25176,N_22275,N_23005);
xor U25177 (N_25177,N_23003,N_23173);
nor U25178 (N_25178,N_22719,N_23129);
xor U25179 (N_25179,N_23507,N_23870);
nand U25180 (N_25180,N_22049,N_22112);
or U25181 (N_25181,N_22509,N_22797);
nor U25182 (N_25182,N_22991,N_23157);
or U25183 (N_25183,N_23776,N_22667);
xor U25184 (N_25184,N_22218,N_22349);
nor U25185 (N_25185,N_22444,N_23025);
xor U25186 (N_25186,N_22308,N_23921);
or U25187 (N_25187,N_22934,N_22541);
nor U25188 (N_25188,N_23075,N_23558);
xor U25189 (N_25189,N_22865,N_22056);
nor U25190 (N_25190,N_23239,N_23460);
nand U25191 (N_25191,N_22489,N_22414);
or U25192 (N_25192,N_22987,N_23640);
xnor U25193 (N_25193,N_22301,N_22522);
and U25194 (N_25194,N_23570,N_23439);
nand U25195 (N_25195,N_22825,N_23761);
and U25196 (N_25196,N_23321,N_22332);
nand U25197 (N_25197,N_22759,N_23459);
nor U25198 (N_25198,N_22094,N_22530);
xor U25199 (N_25199,N_22265,N_22931);
nand U25200 (N_25200,N_22930,N_22944);
and U25201 (N_25201,N_23622,N_22992);
xnor U25202 (N_25202,N_22634,N_22470);
or U25203 (N_25203,N_23341,N_23873);
xnor U25204 (N_25204,N_22348,N_23917);
nand U25205 (N_25205,N_23734,N_22013);
or U25206 (N_25206,N_23955,N_22304);
or U25207 (N_25207,N_22117,N_23759);
and U25208 (N_25208,N_23469,N_23610);
nand U25209 (N_25209,N_23000,N_22337);
or U25210 (N_25210,N_22644,N_23154);
nor U25211 (N_25211,N_22986,N_22359);
or U25212 (N_25212,N_23141,N_22189);
nor U25213 (N_25213,N_23803,N_22751);
and U25214 (N_25214,N_23307,N_23334);
nand U25215 (N_25215,N_22851,N_23693);
nor U25216 (N_25216,N_23781,N_23975);
xor U25217 (N_25217,N_23334,N_22516);
nand U25218 (N_25218,N_22504,N_22913);
xnor U25219 (N_25219,N_23799,N_23763);
xor U25220 (N_25220,N_23952,N_23375);
xor U25221 (N_25221,N_22695,N_22948);
nor U25222 (N_25222,N_23203,N_23553);
nand U25223 (N_25223,N_22422,N_22783);
nand U25224 (N_25224,N_22458,N_23933);
nor U25225 (N_25225,N_22496,N_23480);
xor U25226 (N_25226,N_22044,N_22411);
xor U25227 (N_25227,N_22135,N_22281);
nand U25228 (N_25228,N_23441,N_23797);
nand U25229 (N_25229,N_22069,N_22019);
nand U25230 (N_25230,N_23764,N_23349);
or U25231 (N_25231,N_22045,N_22038);
nand U25232 (N_25232,N_23501,N_23386);
or U25233 (N_25233,N_23001,N_23385);
nand U25234 (N_25234,N_23666,N_23194);
and U25235 (N_25235,N_23616,N_23266);
or U25236 (N_25236,N_22647,N_23778);
or U25237 (N_25237,N_23468,N_23312);
nor U25238 (N_25238,N_23227,N_22134);
xnor U25239 (N_25239,N_23870,N_23389);
or U25240 (N_25240,N_22607,N_23911);
nor U25241 (N_25241,N_22854,N_22922);
nor U25242 (N_25242,N_22137,N_23688);
and U25243 (N_25243,N_22585,N_22774);
xnor U25244 (N_25244,N_22171,N_22862);
xor U25245 (N_25245,N_23793,N_23941);
or U25246 (N_25246,N_23626,N_23706);
xnor U25247 (N_25247,N_23577,N_22770);
xnor U25248 (N_25248,N_22120,N_22515);
and U25249 (N_25249,N_22696,N_22303);
and U25250 (N_25250,N_22658,N_22490);
or U25251 (N_25251,N_22809,N_22742);
nor U25252 (N_25252,N_22658,N_22739);
nor U25253 (N_25253,N_23055,N_22462);
nor U25254 (N_25254,N_23911,N_23061);
nor U25255 (N_25255,N_22317,N_22672);
and U25256 (N_25256,N_23321,N_23994);
nor U25257 (N_25257,N_22242,N_22698);
nand U25258 (N_25258,N_22833,N_23969);
and U25259 (N_25259,N_22963,N_22313);
and U25260 (N_25260,N_22984,N_23064);
xor U25261 (N_25261,N_23567,N_22819);
and U25262 (N_25262,N_22179,N_23954);
nor U25263 (N_25263,N_22315,N_22188);
and U25264 (N_25264,N_22532,N_22370);
nor U25265 (N_25265,N_22695,N_23485);
and U25266 (N_25266,N_22322,N_23206);
nand U25267 (N_25267,N_22331,N_22350);
or U25268 (N_25268,N_22277,N_23106);
nor U25269 (N_25269,N_22287,N_22368);
nand U25270 (N_25270,N_23480,N_23786);
nand U25271 (N_25271,N_22160,N_22515);
xor U25272 (N_25272,N_22209,N_23847);
or U25273 (N_25273,N_23872,N_23423);
nor U25274 (N_25274,N_23950,N_23467);
nor U25275 (N_25275,N_22736,N_22958);
xor U25276 (N_25276,N_22124,N_22882);
xnor U25277 (N_25277,N_23054,N_22181);
or U25278 (N_25278,N_23253,N_22840);
or U25279 (N_25279,N_22842,N_23662);
or U25280 (N_25280,N_22549,N_22823);
xor U25281 (N_25281,N_23298,N_23054);
or U25282 (N_25282,N_22163,N_23736);
and U25283 (N_25283,N_22754,N_22941);
nor U25284 (N_25284,N_22011,N_22727);
and U25285 (N_25285,N_23095,N_22135);
nor U25286 (N_25286,N_23766,N_22513);
and U25287 (N_25287,N_22249,N_23724);
xnor U25288 (N_25288,N_22636,N_23583);
xor U25289 (N_25289,N_22910,N_22111);
or U25290 (N_25290,N_23200,N_22808);
nand U25291 (N_25291,N_23453,N_23025);
or U25292 (N_25292,N_23808,N_22091);
and U25293 (N_25293,N_23539,N_23687);
nor U25294 (N_25294,N_23022,N_23777);
or U25295 (N_25295,N_23877,N_22072);
xnor U25296 (N_25296,N_22680,N_22076);
xnor U25297 (N_25297,N_23151,N_22934);
and U25298 (N_25298,N_22011,N_23748);
nor U25299 (N_25299,N_23437,N_22917);
and U25300 (N_25300,N_23160,N_22526);
nand U25301 (N_25301,N_22015,N_23024);
xor U25302 (N_25302,N_23622,N_22547);
or U25303 (N_25303,N_22404,N_22750);
nor U25304 (N_25304,N_22349,N_22933);
nor U25305 (N_25305,N_23992,N_22543);
nor U25306 (N_25306,N_23522,N_23453);
nor U25307 (N_25307,N_22429,N_23549);
nor U25308 (N_25308,N_23421,N_23976);
xor U25309 (N_25309,N_22510,N_22151);
xor U25310 (N_25310,N_22829,N_23631);
nor U25311 (N_25311,N_22974,N_23704);
xnor U25312 (N_25312,N_22772,N_23497);
or U25313 (N_25313,N_22374,N_23377);
nand U25314 (N_25314,N_22093,N_22692);
nand U25315 (N_25315,N_23756,N_22405);
and U25316 (N_25316,N_23747,N_22681);
nand U25317 (N_25317,N_23265,N_22083);
xor U25318 (N_25318,N_22404,N_23276);
nor U25319 (N_25319,N_22389,N_23831);
nand U25320 (N_25320,N_23855,N_22054);
xor U25321 (N_25321,N_23845,N_23876);
xnor U25322 (N_25322,N_23124,N_23114);
or U25323 (N_25323,N_22383,N_22591);
nor U25324 (N_25324,N_23163,N_22567);
or U25325 (N_25325,N_23962,N_22205);
or U25326 (N_25326,N_22543,N_22634);
nor U25327 (N_25327,N_23844,N_23722);
or U25328 (N_25328,N_22874,N_23009);
nand U25329 (N_25329,N_22678,N_23265);
nand U25330 (N_25330,N_23882,N_23165);
nand U25331 (N_25331,N_23629,N_23264);
nand U25332 (N_25332,N_22039,N_23728);
nand U25333 (N_25333,N_22554,N_22956);
nand U25334 (N_25334,N_23425,N_23670);
and U25335 (N_25335,N_23393,N_22105);
and U25336 (N_25336,N_22892,N_23438);
nor U25337 (N_25337,N_23543,N_22705);
and U25338 (N_25338,N_23007,N_23993);
nand U25339 (N_25339,N_22786,N_23709);
nor U25340 (N_25340,N_22745,N_23232);
nand U25341 (N_25341,N_22842,N_23645);
nor U25342 (N_25342,N_23088,N_23405);
nor U25343 (N_25343,N_23211,N_22828);
xnor U25344 (N_25344,N_22648,N_22516);
nor U25345 (N_25345,N_23985,N_22396);
nand U25346 (N_25346,N_23438,N_22003);
nor U25347 (N_25347,N_22342,N_22412);
and U25348 (N_25348,N_22680,N_23447);
nand U25349 (N_25349,N_22998,N_22130);
and U25350 (N_25350,N_22103,N_22904);
and U25351 (N_25351,N_22029,N_22237);
or U25352 (N_25352,N_22357,N_22485);
or U25353 (N_25353,N_22480,N_23232);
xor U25354 (N_25354,N_22903,N_23015);
nand U25355 (N_25355,N_23572,N_22423);
or U25356 (N_25356,N_23764,N_22915);
or U25357 (N_25357,N_23781,N_22586);
nor U25358 (N_25358,N_22022,N_23331);
or U25359 (N_25359,N_22566,N_22467);
xnor U25360 (N_25360,N_22420,N_23631);
and U25361 (N_25361,N_23130,N_23244);
xnor U25362 (N_25362,N_22677,N_22442);
and U25363 (N_25363,N_22612,N_23462);
xnor U25364 (N_25364,N_22821,N_23683);
nand U25365 (N_25365,N_23204,N_22781);
nand U25366 (N_25366,N_22604,N_22274);
nor U25367 (N_25367,N_23546,N_22174);
xor U25368 (N_25368,N_22687,N_23420);
and U25369 (N_25369,N_22861,N_23564);
nand U25370 (N_25370,N_22331,N_22081);
or U25371 (N_25371,N_22245,N_23112);
and U25372 (N_25372,N_23272,N_22030);
and U25373 (N_25373,N_22043,N_22734);
nand U25374 (N_25374,N_22928,N_22514);
xor U25375 (N_25375,N_22243,N_23951);
and U25376 (N_25376,N_23678,N_22405);
xnor U25377 (N_25377,N_22970,N_22776);
or U25378 (N_25378,N_22129,N_23546);
nand U25379 (N_25379,N_23704,N_23122);
xor U25380 (N_25380,N_23864,N_23052);
nand U25381 (N_25381,N_22483,N_22878);
nor U25382 (N_25382,N_23714,N_22410);
nor U25383 (N_25383,N_23855,N_23322);
and U25384 (N_25384,N_23285,N_23044);
and U25385 (N_25385,N_23011,N_22155);
xor U25386 (N_25386,N_23103,N_23971);
xor U25387 (N_25387,N_23014,N_22606);
or U25388 (N_25388,N_23154,N_22852);
or U25389 (N_25389,N_23726,N_23530);
nor U25390 (N_25390,N_23197,N_23324);
xnor U25391 (N_25391,N_23915,N_23994);
xor U25392 (N_25392,N_22471,N_23993);
xor U25393 (N_25393,N_22467,N_23849);
nand U25394 (N_25394,N_23030,N_23997);
and U25395 (N_25395,N_22462,N_23964);
or U25396 (N_25396,N_23637,N_22422);
xor U25397 (N_25397,N_22656,N_23544);
nand U25398 (N_25398,N_22947,N_22085);
and U25399 (N_25399,N_23559,N_22489);
xor U25400 (N_25400,N_22550,N_23301);
nand U25401 (N_25401,N_22851,N_22719);
nor U25402 (N_25402,N_23352,N_23433);
nand U25403 (N_25403,N_22814,N_23972);
xnor U25404 (N_25404,N_23394,N_23177);
xnor U25405 (N_25405,N_23150,N_22239);
nand U25406 (N_25406,N_23987,N_23552);
xor U25407 (N_25407,N_22307,N_23751);
nor U25408 (N_25408,N_23012,N_22297);
nor U25409 (N_25409,N_23766,N_22278);
nor U25410 (N_25410,N_23517,N_22140);
or U25411 (N_25411,N_22534,N_22971);
and U25412 (N_25412,N_23163,N_22656);
and U25413 (N_25413,N_22493,N_22841);
and U25414 (N_25414,N_22044,N_23104);
and U25415 (N_25415,N_22023,N_23917);
and U25416 (N_25416,N_23483,N_23777);
or U25417 (N_25417,N_22355,N_23419);
nor U25418 (N_25418,N_23382,N_22826);
or U25419 (N_25419,N_22814,N_22612);
nand U25420 (N_25420,N_22805,N_23919);
nand U25421 (N_25421,N_23796,N_22244);
xor U25422 (N_25422,N_22736,N_22415);
nor U25423 (N_25423,N_23437,N_23705);
nand U25424 (N_25424,N_22277,N_22142);
xnor U25425 (N_25425,N_23306,N_22440);
and U25426 (N_25426,N_22458,N_22842);
or U25427 (N_25427,N_22001,N_22870);
and U25428 (N_25428,N_23971,N_23989);
and U25429 (N_25429,N_22135,N_22964);
xor U25430 (N_25430,N_22215,N_23558);
nand U25431 (N_25431,N_22673,N_22160);
or U25432 (N_25432,N_22591,N_23813);
nand U25433 (N_25433,N_23101,N_23696);
nor U25434 (N_25434,N_23423,N_23033);
xnor U25435 (N_25435,N_23421,N_23284);
nand U25436 (N_25436,N_22988,N_23972);
nand U25437 (N_25437,N_23400,N_22307);
xor U25438 (N_25438,N_22586,N_23124);
and U25439 (N_25439,N_23154,N_22266);
nand U25440 (N_25440,N_23342,N_22129);
and U25441 (N_25441,N_23848,N_23321);
or U25442 (N_25442,N_23115,N_23670);
nor U25443 (N_25443,N_22783,N_23392);
nand U25444 (N_25444,N_22403,N_23295);
or U25445 (N_25445,N_22432,N_22727);
nand U25446 (N_25446,N_22341,N_22926);
nand U25447 (N_25447,N_22346,N_23624);
or U25448 (N_25448,N_23706,N_22633);
nor U25449 (N_25449,N_22743,N_22714);
nand U25450 (N_25450,N_22108,N_23058);
nand U25451 (N_25451,N_22965,N_22280);
xnor U25452 (N_25452,N_22806,N_22848);
xnor U25453 (N_25453,N_23875,N_22486);
and U25454 (N_25454,N_23347,N_23534);
or U25455 (N_25455,N_22712,N_22577);
nor U25456 (N_25456,N_23223,N_22277);
or U25457 (N_25457,N_23930,N_22552);
or U25458 (N_25458,N_23508,N_22518);
nor U25459 (N_25459,N_23131,N_22720);
nor U25460 (N_25460,N_23157,N_22655);
or U25461 (N_25461,N_23710,N_22812);
nor U25462 (N_25462,N_23241,N_22399);
nand U25463 (N_25463,N_22577,N_22238);
and U25464 (N_25464,N_22278,N_22245);
and U25465 (N_25465,N_22303,N_23120);
nand U25466 (N_25466,N_23889,N_23167);
nor U25467 (N_25467,N_22186,N_22452);
or U25468 (N_25468,N_22451,N_22933);
nand U25469 (N_25469,N_23684,N_22952);
nor U25470 (N_25470,N_22991,N_23833);
nor U25471 (N_25471,N_23064,N_23138);
and U25472 (N_25472,N_22497,N_23298);
xor U25473 (N_25473,N_22368,N_22355);
or U25474 (N_25474,N_23996,N_22819);
or U25475 (N_25475,N_23316,N_22776);
or U25476 (N_25476,N_23591,N_23087);
and U25477 (N_25477,N_22324,N_22270);
xor U25478 (N_25478,N_23770,N_23528);
or U25479 (N_25479,N_22065,N_22546);
or U25480 (N_25480,N_23923,N_22995);
nand U25481 (N_25481,N_23380,N_23968);
nor U25482 (N_25482,N_22169,N_23355);
nand U25483 (N_25483,N_23305,N_23115);
or U25484 (N_25484,N_22238,N_22540);
nand U25485 (N_25485,N_23708,N_22259);
nand U25486 (N_25486,N_22134,N_23533);
xnor U25487 (N_25487,N_22254,N_22166);
nor U25488 (N_25488,N_23506,N_23233);
or U25489 (N_25489,N_22052,N_23024);
nand U25490 (N_25490,N_23793,N_23556);
and U25491 (N_25491,N_22757,N_23336);
and U25492 (N_25492,N_23138,N_23036);
nor U25493 (N_25493,N_23504,N_22388);
nor U25494 (N_25494,N_22117,N_23379);
xor U25495 (N_25495,N_22779,N_23683);
nand U25496 (N_25496,N_22426,N_23364);
nor U25497 (N_25497,N_22130,N_22294);
nor U25498 (N_25498,N_23393,N_23680);
xnor U25499 (N_25499,N_23445,N_23496);
xor U25500 (N_25500,N_22370,N_23926);
or U25501 (N_25501,N_22720,N_23010);
or U25502 (N_25502,N_23451,N_22861);
or U25503 (N_25503,N_22511,N_22361);
nor U25504 (N_25504,N_23405,N_22717);
or U25505 (N_25505,N_22980,N_23423);
nand U25506 (N_25506,N_23670,N_23820);
and U25507 (N_25507,N_22192,N_23519);
xnor U25508 (N_25508,N_23780,N_23714);
or U25509 (N_25509,N_22848,N_22743);
nand U25510 (N_25510,N_22255,N_23191);
nor U25511 (N_25511,N_22807,N_23964);
and U25512 (N_25512,N_23434,N_22952);
or U25513 (N_25513,N_22930,N_22079);
xnor U25514 (N_25514,N_22467,N_22542);
and U25515 (N_25515,N_22435,N_23404);
nor U25516 (N_25516,N_23149,N_23102);
and U25517 (N_25517,N_22219,N_23611);
or U25518 (N_25518,N_23495,N_22714);
nand U25519 (N_25519,N_22035,N_22684);
nand U25520 (N_25520,N_23741,N_22343);
or U25521 (N_25521,N_22173,N_23987);
nand U25522 (N_25522,N_23736,N_22500);
nor U25523 (N_25523,N_22908,N_22000);
xor U25524 (N_25524,N_22174,N_23739);
nor U25525 (N_25525,N_22179,N_23548);
or U25526 (N_25526,N_23133,N_23822);
and U25527 (N_25527,N_23356,N_23370);
or U25528 (N_25528,N_23420,N_23508);
nand U25529 (N_25529,N_23042,N_22549);
nand U25530 (N_25530,N_23418,N_23491);
nor U25531 (N_25531,N_23182,N_23672);
or U25532 (N_25532,N_23772,N_23542);
or U25533 (N_25533,N_22500,N_22473);
nor U25534 (N_25534,N_23795,N_22271);
and U25535 (N_25535,N_22943,N_23861);
and U25536 (N_25536,N_22099,N_23689);
xnor U25537 (N_25537,N_23118,N_23484);
and U25538 (N_25538,N_22056,N_22047);
nand U25539 (N_25539,N_22138,N_23402);
or U25540 (N_25540,N_23539,N_23448);
nor U25541 (N_25541,N_22019,N_23080);
nor U25542 (N_25542,N_23709,N_23032);
and U25543 (N_25543,N_22696,N_22318);
xor U25544 (N_25544,N_23679,N_23445);
xnor U25545 (N_25545,N_23699,N_23371);
xor U25546 (N_25546,N_23950,N_22360);
or U25547 (N_25547,N_23735,N_23203);
and U25548 (N_25548,N_23765,N_23994);
xor U25549 (N_25549,N_23581,N_23121);
nand U25550 (N_25550,N_23879,N_22466);
nor U25551 (N_25551,N_23064,N_23593);
and U25552 (N_25552,N_22985,N_23279);
and U25553 (N_25553,N_22737,N_22570);
nand U25554 (N_25554,N_23237,N_23269);
or U25555 (N_25555,N_22379,N_23237);
nand U25556 (N_25556,N_23289,N_23839);
and U25557 (N_25557,N_22342,N_22445);
or U25558 (N_25558,N_22294,N_22286);
nor U25559 (N_25559,N_23951,N_23784);
xnor U25560 (N_25560,N_22576,N_22604);
and U25561 (N_25561,N_23097,N_23536);
xnor U25562 (N_25562,N_22194,N_22745);
or U25563 (N_25563,N_22348,N_22134);
and U25564 (N_25564,N_22263,N_23348);
or U25565 (N_25565,N_22837,N_23495);
nor U25566 (N_25566,N_22141,N_22565);
nor U25567 (N_25567,N_22672,N_23425);
and U25568 (N_25568,N_23713,N_23656);
nand U25569 (N_25569,N_23887,N_22654);
or U25570 (N_25570,N_23307,N_23153);
xor U25571 (N_25571,N_22641,N_23361);
or U25572 (N_25572,N_23947,N_23750);
nand U25573 (N_25573,N_23428,N_23676);
xnor U25574 (N_25574,N_23487,N_23481);
nor U25575 (N_25575,N_23116,N_23137);
and U25576 (N_25576,N_23245,N_22826);
and U25577 (N_25577,N_22704,N_23861);
nor U25578 (N_25578,N_23530,N_23588);
nor U25579 (N_25579,N_23174,N_23014);
xnor U25580 (N_25580,N_23824,N_22271);
and U25581 (N_25581,N_22062,N_23448);
and U25582 (N_25582,N_23901,N_22575);
nand U25583 (N_25583,N_22846,N_22377);
or U25584 (N_25584,N_22492,N_23088);
and U25585 (N_25585,N_22530,N_23500);
and U25586 (N_25586,N_22838,N_22212);
and U25587 (N_25587,N_23340,N_23429);
nor U25588 (N_25588,N_23373,N_22030);
xor U25589 (N_25589,N_23584,N_22994);
or U25590 (N_25590,N_23860,N_22060);
xnor U25591 (N_25591,N_23123,N_22127);
and U25592 (N_25592,N_22606,N_23500);
or U25593 (N_25593,N_22481,N_23513);
and U25594 (N_25594,N_23560,N_22168);
nand U25595 (N_25595,N_23861,N_23475);
nand U25596 (N_25596,N_22195,N_22643);
or U25597 (N_25597,N_22310,N_23365);
nor U25598 (N_25598,N_22970,N_22313);
nor U25599 (N_25599,N_23274,N_22978);
nand U25600 (N_25600,N_22266,N_22428);
and U25601 (N_25601,N_23726,N_23443);
and U25602 (N_25602,N_23661,N_22275);
xnor U25603 (N_25603,N_23930,N_23191);
nand U25604 (N_25604,N_23307,N_23494);
xor U25605 (N_25605,N_22843,N_23697);
xor U25606 (N_25606,N_22653,N_22540);
nand U25607 (N_25607,N_23416,N_23342);
or U25608 (N_25608,N_23154,N_23358);
and U25609 (N_25609,N_22522,N_22761);
and U25610 (N_25610,N_23337,N_22239);
and U25611 (N_25611,N_23137,N_23524);
nor U25612 (N_25612,N_23146,N_23460);
xor U25613 (N_25613,N_23978,N_22973);
and U25614 (N_25614,N_23891,N_23407);
or U25615 (N_25615,N_23596,N_23785);
or U25616 (N_25616,N_22420,N_22904);
nor U25617 (N_25617,N_23578,N_23393);
nor U25618 (N_25618,N_23390,N_23559);
or U25619 (N_25619,N_23833,N_22836);
or U25620 (N_25620,N_22709,N_23901);
nor U25621 (N_25621,N_23527,N_23539);
nand U25622 (N_25622,N_23638,N_23648);
and U25623 (N_25623,N_22477,N_23045);
nor U25624 (N_25624,N_22598,N_22802);
nand U25625 (N_25625,N_23833,N_22682);
and U25626 (N_25626,N_23178,N_22080);
nor U25627 (N_25627,N_23796,N_22841);
and U25628 (N_25628,N_23870,N_22934);
nand U25629 (N_25629,N_23800,N_22066);
nor U25630 (N_25630,N_23960,N_23606);
nor U25631 (N_25631,N_23108,N_22147);
nor U25632 (N_25632,N_22043,N_22423);
or U25633 (N_25633,N_22161,N_23012);
and U25634 (N_25634,N_23055,N_23744);
or U25635 (N_25635,N_23815,N_23433);
or U25636 (N_25636,N_22190,N_23985);
nand U25637 (N_25637,N_23420,N_22793);
xnor U25638 (N_25638,N_23368,N_22726);
and U25639 (N_25639,N_23114,N_22236);
and U25640 (N_25640,N_22854,N_22660);
nor U25641 (N_25641,N_23587,N_23842);
nand U25642 (N_25642,N_23925,N_22263);
nand U25643 (N_25643,N_23596,N_23966);
xnor U25644 (N_25644,N_22103,N_22176);
nor U25645 (N_25645,N_23885,N_22249);
nand U25646 (N_25646,N_23050,N_23026);
xnor U25647 (N_25647,N_22117,N_22714);
nand U25648 (N_25648,N_23158,N_22931);
nor U25649 (N_25649,N_22482,N_22167);
nand U25650 (N_25650,N_23183,N_22136);
nand U25651 (N_25651,N_23229,N_22045);
nor U25652 (N_25652,N_23290,N_22917);
nor U25653 (N_25653,N_23414,N_23291);
nor U25654 (N_25654,N_23443,N_22029);
nor U25655 (N_25655,N_23628,N_23291);
and U25656 (N_25656,N_23219,N_22605);
or U25657 (N_25657,N_23756,N_22982);
or U25658 (N_25658,N_22816,N_22071);
or U25659 (N_25659,N_23876,N_23540);
nand U25660 (N_25660,N_22738,N_22136);
nand U25661 (N_25661,N_23492,N_22199);
nor U25662 (N_25662,N_23605,N_23008);
or U25663 (N_25663,N_23575,N_23608);
xor U25664 (N_25664,N_22820,N_22263);
nand U25665 (N_25665,N_22954,N_23594);
or U25666 (N_25666,N_22661,N_22364);
xor U25667 (N_25667,N_22486,N_23669);
nor U25668 (N_25668,N_22235,N_22409);
and U25669 (N_25669,N_23574,N_22625);
nor U25670 (N_25670,N_23478,N_23605);
or U25671 (N_25671,N_23976,N_23821);
xor U25672 (N_25672,N_22178,N_22367);
and U25673 (N_25673,N_23483,N_23523);
xor U25674 (N_25674,N_22918,N_23158);
nand U25675 (N_25675,N_23297,N_22087);
and U25676 (N_25676,N_23723,N_23078);
or U25677 (N_25677,N_22596,N_23399);
and U25678 (N_25678,N_22526,N_23140);
nor U25679 (N_25679,N_22395,N_22169);
nand U25680 (N_25680,N_23917,N_22195);
nand U25681 (N_25681,N_22505,N_22835);
nand U25682 (N_25682,N_22125,N_22792);
xor U25683 (N_25683,N_22365,N_22349);
or U25684 (N_25684,N_23980,N_22315);
or U25685 (N_25685,N_22561,N_22554);
or U25686 (N_25686,N_23817,N_23989);
xnor U25687 (N_25687,N_22953,N_22470);
and U25688 (N_25688,N_23936,N_23998);
xor U25689 (N_25689,N_23836,N_23026);
or U25690 (N_25690,N_23957,N_23637);
or U25691 (N_25691,N_23770,N_22067);
and U25692 (N_25692,N_22906,N_23803);
xnor U25693 (N_25693,N_23972,N_23780);
and U25694 (N_25694,N_22859,N_22763);
nand U25695 (N_25695,N_22355,N_22960);
nor U25696 (N_25696,N_23088,N_22713);
nor U25697 (N_25697,N_22276,N_23248);
xnor U25698 (N_25698,N_23128,N_22904);
or U25699 (N_25699,N_22774,N_22112);
or U25700 (N_25700,N_23278,N_22583);
or U25701 (N_25701,N_22927,N_22744);
nand U25702 (N_25702,N_23439,N_23753);
or U25703 (N_25703,N_22724,N_23784);
or U25704 (N_25704,N_23801,N_22121);
nand U25705 (N_25705,N_23170,N_22600);
nor U25706 (N_25706,N_23401,N_23436);
and U25707 (N_25707,N_23376,N_23856);
nand U25708 (N_25708,N_22095,N_23053);
nand U25709 (N_25709,N_23030,N_23647);
xor U25710 (N_25710,N_23065,N_23850);
nor U25711 (N_25711,N_22593,N_23502);
xnor U25712 (N_25712,N_22206,N_22976);
xor U25713 (N_25713,N_22746,N_22713);
nor U25714 (N_25714,N_23178,N_22503);
nor U25715 (N_25715,N_22704,N_23555);
nand U25716 (N_25716,N_22901,N_22899);
xnor U25717 (N_25717,N_23100,N_22906);
and U25718 (N_25718,N_22896,N_23988);
or U25719 (N_25719,N_23811,N_23644);
or U25720 (N_25720,N_22237,N_23744);
and U25721 (N_25721,N_23698,N_22602);
nand U25722 (N_25722,N_23942,N_23160);
nand U25723 (N_25723,N_23555,N_22194);
nor U25724 (N_25724,N_22750,N_23326);
or U25725 (N_25725,N_23707,N_23497);
and U25726 (N_25726,N_23112,N_22952);
xnor U25727 (N_25727,N_22942,N_23721);
nor U25728 (N_25728,N_22454,N_22116);
or U25729 (N_25729,N_23633,N_22560);
and U25730 (N_25730,N_23245,N_22437);
and U25731 (N_25731,N_22777,N_23828);
or U25732 (N_25732,N_23511,N_23487);
or U25733 (N_25733,N_23302,N_23126);
nor U25734 (N_25734,N_23365,N_23219);
xor U25735 (N_25735,N_22217,N_23748);
and U25736 (N_25736,N_22877,N_23154);
nor U25737 (N_25737,N_23880,N_22343);
and U25738 (N_25738,N_22172,N_23240);
or U25739 (N_25739,N_22642,N_23070);
nor U25740 (N_25740,N_23588,N_22712);
xor U25741 (N_25741,N_22751,N_22816);
nor U25742 (N_25742,N_23282,N_22202);
nor U25743 (N_25743,N_23144,N_22003);
xor U25744 (N_25744,N_23747,N_23442);
and U25745 (N_25745,N_23541,N_23728);
nand U25746 (N_25746,N_23317,N_23612);
and U25747 (N_25747,N_23633,N_22237);
and U25748 (N_25748,N_23081,N_22102);
or U25749 (N_25749,N_23482,N_23984);
or U25750 (N_25750,N_23794,N_22840);
and U25751 (N_25751,N_22846,N_22710);
xnor U25752 (N_25752,N_23191,N_22384);
or U25753 (N_25753,N_23171,N_22325);
or U25754 (N_25754,N_22796,N_22502);
or U25755 (N_25755,N_23073,N_23417);
nand U25756 (N_25756,N_22474,N_23576);
and U25757 (N_25757,N_23730,N_23036);
nand U25758 (N_25758,N_22902,N_23069);
xor U25759 (N_25759,N_23711,N_23570);
and U25760 (N_25760,N_22175,N_22436);
nor U25761 (N_25761,N_23244,N_23455);
nand U25762 (N_25762,N_23554,N_23783);
or U25763 (N_25763,N_23664,N_23230);
or U25764 (N_25764,N_23254,N_22486);
xor U25765 (N_25765,N_22667,N_22039);
nor U25766 (N_25766,N_22673,N_23332);
and U25767 (N_25767,N_22505,N_23210);
xnor U25768 (N_25768,N_22780,N_22172);
nand U25769 (N_25769,N_23260,N_22714);
nand U25770 (N_25770,N_22705,N_22941);
and U25771 (N_25771,N_23409,N_23592);
and U25772 (N_25772,N_22444,N_22856);
and U25773 (N_25773,N_23124,N_22540);
and U25774 (N_25774,N_22833,N_23555);
or U25775 (N_25775,N_22220,N_22669);
xnor U25776 (N_25776,N_22751,N_23573);
xor U25777 (N_25777,N_23452,N_23251);
or U25778 (N_25778,N_22980,N_22036);
xor U25779 (N_25779,N_23071,N_22940);
xor U25780 (N_25780,N_22916,N_23903);
nor U25781 (N_25781,N_23194,N_23748);
nand U25782 (N_25782,N_22171,N_23286);
nor U25783 (N_25783,N_23677,N_23416);
nand U25784 (N_25784,N_22308,N_23035);
nand U25785 (N_25785,N_22712,N_22127);
nand U25786 (N_25786,N_23023,N_23681);
nor U25787 (N_25787,N_22176,N_22111);
or U25788 (N_25788,N_22538,N_22153);
and U25789 (N_25789,N_23180,N_22777);
and U25790 (N_25790,N_22037,N_22456);
nor U25791 (N_25791,N_23340,N_23927);
nor U25792 (N_25792,N_23211,N_22231);
nand U25793 (N_25793,N_23424,N_22522);
or U25794 (N_25794,N_23041,N_22968);
xnor U25795 (N_25795,N_23400,N_22741);
xor U25796 (N_25796,N_23085,N_22426);
nand U25797 (N_25797,N_22637,N_23467);
or U25798 (N_25798,N_22029,N_23813);
or U25799 (N_25799,N_22003,N_22339);
and U25800 (N_25800,N_23163,N_23439);
or U25801 (N_25801,N_23127,N_22868);
nor U25802 (N_25802,N_23669,N_23007);
or U25803 (N_25803,N_22478,N_23998);
and U25804 (N_25804,N_23584,N_23595);
and U25805 (N_25805,N_22489,N_23178);
and U25806 (N_25806,N_22132,N_22481);
xnor U25807 (N_25807,N_22999,N_23142);
or U25808 (N_25808,N_23591,N_22120);
and U25809 (N_25809,N_23012,N_22330);
nor U25810 (N_25810,N_22617,N_22697);
and U25811 (N_25811,N_22735,N_22043);
nor U25812 (N_25812,N_22441,N_23876);
or U25813 (N_25813,N_23767,N_23462);
xnor U25814 (N_25814,N_22350,N_22413);
and U25815 (N_25815,N_23676,N_22109);
nand U25816 (N_25816,N_22445,N_23322);
or U25817 (N_25817,N_23137,N_23600);
xnor U25818 (N_25818,N_23671,N_22943);
xnor U25819 (N_25819,N_22355,N_22566);
nor U25820 (N_25820,N_22271,N_22442);
nor U25821 (N_25821,N_22475,N_23260);
nand U25822 (N_25822,N_23770,N_23669);
nand U25823 (N_25823,N_22927,N_23052);
and U25824 (N_25824,N_22205,N_22716);
and U25825 (N_25825,N_22456,N_23254);
nand U25826 (N_25826,N_23625,N_23220);
and U25827 (N_25827,N_22143,N_22503);
or U25828 (N_25828,N_23417,N_22106);
nand U25829 (N_25829,N_23137,N_23038);
xor U25830 (N_25830,N_23976,N_23215);
nand U25831 (N_25831,N_23977,N_23388);
and U25832 (N_25832,N_22187,N_23152);
xnor U25833 (N_25833,N_23381,N_23127);
xor U25834 (N_25834,N_23339,N_22591);
xor U25835 (N_25835,N_22224,N_22063);
or U25836 (N_25836,N_22182,N_23547);
xnor U25837 (N_25837,N_22380,N_22560);
nand U25838 (N_25838,N_23451,N_22139);
or U25839 (N_25839,N_23364,N_22652);
nand U25840 (N_25840,N_23480,N_23622);
or U25841 (N_25841,N_22811,N_22926);
nor U25842 (N_25842,N_22350,N_22336);
xor U25843 (N_25843,N_22153,N_22049);
nand U25844 (N_25844,N_22035,N_22052);
nand U25845 (N_25845,N_23777,N_22787);
or U25846 (N_25846,N_23659,N_22358);
nor U25847 (N_25847,N_23658,N_22315);
xor U25848 (N_25848,N_23039,N_23705);
xnor U25849 (N_25849,N_23078,N_22476);
nor U25850 (N_25850,N_23335,N_22673);
nand U25851 (N_25851,N_23586,N_23145);
nand U25852 (N_25852,N_23161,N_23790);
nor U25853 (N_25853,N_23842,N_22403);
nor U25854 (N_25854,N_22467,N_22671);
xor U25855 (N_25855,N_23646,N_23379);
nor U25856 (N_25856,N_22753,N_22341);
nor U25857 (N_25857,N_23876,N_22165);
or U25858 (N_25858,N_22779,N_23006);
and U25859 (N_25859,N_23492,N_23170);
nor U25860 (N_25860,N_23021,N_23936);
and U25861 (N_25861,N_22473,N_23553);
nand U25862 (N_25862,N_23791,N_22950);
xnor U25863 (N_25863,N_23389,N_23477);
xnor U25864 (N_25864,N_22065,N_23858);
nand U25865 (N_25865,N_23486,N_23063);
or U25866 (N_25866,N_23461,N_23063);
xnor U25867 (N_25867,N_22897,N_22987);
or U25868 (N_25868,N_23943,N_22721);
xor U25869 (N_25869,N_23288,N_23627);
nand U25870 (N_25870,N_22465,N_22320);
nor U25871 (N_25871,N_23495,N_22874);
nand U25872 (N_25872,N_23050,N_23096);
or U25873 (N_25873,N_22180,N_23566);
or U25874 (N_25874,N_23773,N_23421);
nor U25875 (N_25875,N_22333,N_22221);
or U25876 (N_25876,N_23146,N_22903);
nor U25877 (N_25877,N_22562,N_22612);
xnor U25878 (N_25878,N_23533,N_23011);
and U25879 (N_25879,N_22415,N_22625);
and U25880 (N_25880,N_22815,N_23157);
or U25881 (N_25881,N_23765,N_22094);
nand U25882 (N_25882,N_23900,N_22362);
nand U25883 (N_25883,N_23553,N_23058);
and U25884 (N_25884,N_22275,N_22497);
xnor U25885 (N_25885,N_23526,N_23585);
or U25886 (N_25886,N_23489,N_23510);
nand U25887 (N_25887,N_23891,N_23611);
and U25888 (N_25888,N_23544,N_22204);
or U25889 (N_25889,N_23124,N_22956);
nand U25890 (N_25890,N_23573,N_22654);
nor U25891 (N_25891,N_23448,N_23788);
and U25892 (N_25892,N_23648,N_22142);
and U25893 (N_25893,N_22623,N_22109);
nor U25894 (N_25894,N_22019,N_23532);
nand U25895 (N_25895,N_23960,N_22035);
nand U25896 (N_25896,N_23897,N_23921);
and U25897 (N_25897,N_22184,N_22533);
nor U25898 (N_25898,N_22232,N_22501);
or U25899 (N_25899,N_22998,N_23863);
xor U25900 (N_25900,N_23748,N_22840);
nand U25901 (N_25901,N_22964,N_22096);
or U25902 (N_25902,N_23248,N_22365);
or U25903 (N_25903,N_23391,N_22622);
nand U25904 (N_25904,N_23119,N_22288);
and U25905 (N_25905,N_22681,N_22830);
nor U25906 (N_25906,N_22489,N_22709);
nand U25907 (N_25907,N_22491,N_23992);
nand U25908 (N_25908,N_22527,N_23351);
or U25909 (N_25909,N_22955,N_22170);
or U25910 (N_25910,N_23173,N_22108);
and U25911 (N_25911,N_23821,N_22657);
and U25912 (N_25912,N_23691,N_23190);
and U25913 (N_25913,N_23469,N_22685);
or U25914 (N_25914,N_22675,N_23450);
nand U25915 (N_25915,N_23716,N_22704);
and U25916 (N_25916,N_23624,N_23712);
and U25917 (N_25917,N_23213,N_23453);
and U25918 (N_25918,N_23131,N_23178);
xor U25919 (N_25919,N_23993,N_23082);
nand U25920 (N_25920,N_23725,N_23451);
nor U25921 (N_25921,N_22700,N_23699);
nor U25922 (N_25922,N_22517,N_22163);
and U25923 (N_25923,N_23784,N_23855);
and U25924 (N_25924,N_22108,N_22189);
or U25925 (N_25925,N_23732,N_22216);
and U25926 (N_25926,N_22908,N_22293);
and U25927 (N_25927,N_23620,N_22490);
and U25928 (N_25928,N_22150,N_23679);
or U25929 (N_25929,N_23379,N_23974);
nand U25930 (N_25930,N_22230,N_22414);
or U25931 (N_25931,N_22302,N_23592);
and U25932 (N_25932,N_22702,N_23441);
or U25933 (N_25933,N_22665,N_23051);
xnor U25934 (N_25934,N_22595,N_23661);
or U25935 (N_25935,N_23153,N_23785);
nand U25936 (N_25936,N_22864,N_23205);
xnor U25937 (N_25937,N_23112,N_22014);
xor U25938 (N_25938,N_23818,N_22128);
xnor U25939 (N_25939,N_23984,N_23980);
and U25940 (N_25940,N_23948,N_22051);
and U25941 (N_25941,N_22425,N_23380);
or U25942 (N_25942,N_22100,N_23246);
and U25943 (N_25943,N_23089,N_23070);
nor U25944 (N_25944,N_22056,N_23438);
nor U25945 (N_25945,N_23999,N_23717);
xor U25946 (N_25946,N_22908,N_23765);
and U25947 (N_25947,N_22891,N_22196);
nand U25948 (N_25948,N_23365,N_22305);
nand U25949 (N_25949,N_22196,N_23975);
and U25950 (N_25950,N_23240,N_23429);
and U25951 (N_25951,N_23068,N_22837);
nor U25952 (N_25952,N_23014,N_23242);
or U25953 (N_25953,N_23980,N_22185);
and U25954 (N_25954,N_23800,N_22497);
nand U25955 (N_25955,N_23354,N_23752);
or U25956 (N_25956,N_23867,N_23439);
xor U25957 (N_25957,N_23928,N_23895);
and U25958 (N_25958,N_22383,N_23119);
xnor U25959 (N_25959,N_23226,N_23194);
xnor U25960 (N_25960,N_22794,N_22117);
nand U25961 (N_25961,N_22138,N_22189);
nor U25962 (N_25962,N_22424,N_22502);
xnor U25963 (N_25963,N_23109,N_22738);
or U25964 (N_25964,N_22363,N_22405);
or U25965 (N_25965,N_23371,N_23909);
or U25966 (N_25966,N_22503,N_22717);
or U25967 (N_25967,N_23137,N_23590);
and U25968 (N_25968,N_23460,N_22527);
nor U25969 (N_25969,N_23984,N_23971);
nand U25970 (N_25970,N_23682,N_22987);
and U25971 (N_25971,N_22681,N_23024);
nand U25972 (N_25972,N_22965,N_23495);
nand U25973 (N_25973,N_23530,N_23442);
nor U25974 (N_25974,N_23127,N_23376);
nand U25975 (N_25975,N_22916,N_22008);
nand U25976 (N_25976,N_23115,N_23938);
nand U25977 (N_25977,N_23274,N_22486);
nor U25978 (N_25978,N_23660,N_22652);
and U25979 (N_25979,N_23698,N_22192);
or U25980 (N_25980,N_23527,N_22630);
or U25981 (N_25981,N_23654,N_22067);
or U25982 (N_25982,N_22661,N_23249);
nand U25983 (N_25983,N_22892,N_23029);
nand U25984 (N_25984,N_23734,N_22330);
nor U25985 (N_25985,N_23387,N_22370);
and U25986 (N_25986,N_22539,N_22381);
xor U25987 (N_25987,N_22647,N_23039);
nor U25988 (N_25988,N_23297,N_23530);
and U25989 (N_25989,N_22804,N_23663);
xnor U25990 (N_25990,N_22748,N_23161);
and U25991 (N_25991,N_22769,N_22301);
nand U25992 (N_25992,N_23362,N_22872);
nor U25993 (N_25993,N_22079,N_23539);
xor U25994 (N_25994,N_22357,N_23607);
xor U25995 (N_25995,N_22877,N_22255);
and U25996 (N_25996,N_23197,N_23969);
nor U25997 (N_25997,N_23896,N_23984);
xnor U25998 (N_25998,N_23398,N_22722);
nand U25999 (N_25999,N_22872,N_22142);
xnor U26000 (N_26000,N_24776,N_25770);
and U26001 (N_26001,N_24556,N_25460);
or U26002 (N_26002,N_25294,N_25323);
xnor U26003 (N_26003,N_24346,N_24859);
nand U26004 (N_26004,N_24136,N_25258);
xor U26005 (N_26005,N_25873,N_24258);
and U26006 (N_26006,N_25473,N_24297);
and U26007 (N_26007,N_24237,N_25621);
or U26008 (N_26008,N_24707,N_24806);
and U26009 (N_26009,N_24722,N_25774);
nor U26010 (N_26010,N_24303,N_25634);
nand U26011 (N_26011,N_24882,N_24466);
and U26012 (N_26012,N_24240,N_25681);
and U26013 (N_26013,N_25646,N_25185);
xnor U26014 (N_26014,N_24100,N_25654);
xor U26015 (N_26015,N_25914,N_25936);
nor U26016 (N_26016,N_25406,N_25313);
nand U26017 (N_26017,N_24811,N_25735);
nor U26018 (N_26018,N_25483,N_24044);
or U26019 (N_26019,N_24443,N_24078);
and U26020 (N_26020,N_25949,N_25499);
or U26021 (N_26021,N_25943,N_24016);
xor U26022 (N_26022,N_24642,N_25251);
nor U26023 (N_26023,N_24692,N_24116);
xnor U26024 (N_26024,N_25032,N_25158);
nand U26025 (N_26025,N_25363,N_24274);
nand U26026 (N_26026,N_25026,N_25801);
nor U26027 (N_26027,N_25910,N_25782);
nand U26028 (N_26028,N_24641,N_25769);
or U26029 (N_26029,N_24082,N_25933);
xnor U26030 (N_26030,N_25418,N_25245);
and U26031 (N_26031,N_25331,N_25624);
nor U26032 (N_26032,N_25340,N_24400);
xor U26033 (N_26033,N_24038,N_24096);
nor U26034 (N_26034,N_25558,N_25538);
and U26035 (N_26035,N_24706,N_25237);
or U26036 (N_26036,N_25713,N_24747);
or U26037 (N_26037,N_25253,N_25966);
and U26038 (N_26038,N_24936,N_24890);
and U26039 (N_26039,N_24305,N_24661);
or U26040 (N_26040,N_25560,N_24061);
and U26041 (N_26041,N_24479,N_25484);
or U26042 (N_26042,N_24458,N_25069);
or U26043 (N_26043,N_24517,N_25934);
nor U26044 (N_26044,N_24500,N_25061);
xnor U26045 (N_26045,N_25403,N_25030);
xnor U26046 (N_26046,N_25886,N_24716);
nand U26047 (N_26047,N_24204,N_25053);
or U26048 (N_26048,N_24165,N_24293);
or U26049 (N_26049,N_25375,N_25194);
or U26050 (N_26050,N_24126,N_24771);
xor U26051 (N_26051,N_24732,N_24537);
xnor U26052 (N_26052,N_24087,N_25764);
xnor U26053 (N_26053,N_24306,N_24298);
nand U26054 (N_26054,N_24627,N_25271);
nand U26055 (N_26055,N_25120,N_25391);
nand U26056 (N_26056,N_24526,N_24975);
xor U26057 (N_26057,N_24964,N_24769);
or U26058 (N_26058,N_24270,N_24825);
xnor U26059 (N_26059,N_25401,N_24555);
nand U26060 (N_26060,N_25448,N_24155);
or U26061 (N_26061,N_24621,N_25159);
and U26062 (N_26062,N_24327,N_25344);
nor U26063 (N_26063,N_25579,N_24688);
xnor U26064 (N_26064,N_25348,N_24362);
and U26065 (N_26065,N_24307,N_24893);
or U26066 (N_26066,N_24587,N_24591);
nor U26067 (N_26067,N_25687,N_24075);
and U26068 (N_26068,N_24501,N_25626);
nor U26069 (N_26069,N_25817,N_25037);
nand U26070 (N_26070,N_24956,N_25367);
nor U26071 (N_26071,N_24002,N_24674);
nor U26072 (N_26072,N_24328,N_25711);
nand U26073 (N_26073,N_25786,N_25419);
nor U26074 (N_26074,N_25077,N_25150);
or U26075 (N_26075,N_25939,N_25458);
nor U26076 (N_26076,N_25749,N_25369);
and U26077 (N_26077,N_25585,N_24276);
nand U26078 (N_26078,N_24915,N_24084);
nand U26079 (N_26079,N_25320,N_24213);
xor U26080 (N_26080,N_24224,N_24329);
and U26081 (N_26081,N_24903,N_24753);
nand U26082 (N_26082,N_25227,N_24310);
nand U26083 (N_26083,N_25364,N_24389);
nor U26084 (N_26084,N_25426,N_25005);
nor U26085 (N_26085,N_25924,N_25928);
or U26086 (N_26086,N_25075,N_25855);
xnor U26087 (N_26087,N_25311,N_24000);
xnor U26088 (N_26088,N_25112,N_25953);
or U26089 (N_26089,N_25976,N_25880);
nor U26090 (N_26090,N_25704,N_25605);
and U26091 (N_26091,N_24390,N_24239);
or U26092 (N_26092,N_24251,N_25049);
nor U26093 (N_26093,N_24348,N_24145);
nand U26094 (N_26094,N_24595,N_24432);
nor U26095 (N_26095,N_25034,N_25494);
xnor U26096 (N_26096,N_24447,N_25950);
xnor U26097 (N_26097,N_25969,N_24992);
and U26098 (N_26098,N_24812,N_25087);
nand U26099 (N_26099,N_24892,N_24386);
and U26100 (N_26100,N_24634,N_24906);
and U26101 (N_26101,N_25368,N_24871);
xnor U26102 (N_26102,N_24436,N_25612);
nand U26103 (N_26103,N_24832,N_24995);
or U26104 (N_26104,N_25440,N_24754);
xnor U26105 (N_26105,N_24062,N_24993);
xor U26106 (N_26106,N_24454,N_25705);
nor U26107 (N_26107,N_25822,N_24219);
nor U26108 (N_26108,N_25507,N_25894);
xor U26109 (N_26109,N_25652,N_24847);
nor U26110 (N_26110,N_25213,N_24865);
and U26111 (N_26111,N_24336,N_24668);
nand U26112 (N_26112,N_25768,N_24648);
nor U26113 (N_26113,N_24569,N_25386);
xnor U26114 (N_26114,N_25312,N_25398);
and U26115 (N_26115,N_25290,N_25022);
xnor U26116 (N_26116,N_24201,N_25777);
and U26117 (N_26117,N_24824,N_25610);
nand U26118 (N_26118,N_25490,N_25909);
nand U26119 (N_26119,N_24394,N_24001);
xnor U26120 (N_26120,N_24818,N_24218);
xnor U26121 (N_26121,N_24367,N_25736);
and U26122 (N_26122,N_25619,N_25962);
or U26123 (N_26123,N_25200,N_24843);
nor U26124 (N_26124,N_24004,N_25385);
nor U26125 (N_26125,N_24081,N_25356);
nand U26126 (N_26126,N_24283,N_25668);
xor U26127 (N_26127,N_25964,N_24299);
nor U26128 (N_26128,N_25593,N_24281);
and U26129 (N_26129,N_24817,N_25677);
nand U26130 (N_26130,N_24854,N_24808);
and U26131 (N_26131,N_25671,N_25230);
nor U26132 (N_26132,N_25043,N_24863);
and U26133 (N_26133,N_24068,N_24007);
xnor U26134 (N_26134,N_25887,N_24941);
xor U26135 (N_26135,N_25932,N_24534);
and U26136 (N_26136,N_24042,N_24114);
xnor U26137 (N_26137,N_25196,N_25137);
or U26138 (N_26138,N_24459,N_24066);
or U26139 (N_26139,N_25653,N_25173);
or U26140 (N_26140,N_24259,N_25211);
nor U26141 (N_26141,N_25465,N_25732);
xnor U26142 (N_26142,N_24723,N_24037);
and U26143 (N_26143,N_25149,N_24907);
and U26144 (N_26144,N_25788,N_24577);
or U26145 (N_26145,N_25812,N_24523);
or U26146 (N_26146,N_25374,N_25999);
xnor U26147 (N_26147,N_24045,N_25620);
xor U26148 (N_26148,N_25903,N_25338);
nor U26149 (N_26149,N_25319,N_25337);
xor U26150 (N_26150,N_24131,N_24831);
and U26151 (N_26151,N_24530,N_25779);
nand U26152 (N_26152,N_24809,N_24758);
and U26153 (N_26153,N_25411,N_24491);
xnor U26154 (N_26154,N_24997,N_24564);
or U26155 (N_26155,N_25335,N_25154);
xnor U26156 (N_26156,N_25508,N_25202);
and U26157 (N_26157,N_25658,N_25265);
nor U26158 (N_26158,N_24088,N_24406);
and U26159 (N_26159,N_25901,N_24381);
nor U26160 (N_26160,N_25918,N_24550);
or U26161 (N_26161,N_24885,N_25378);
xor U26162 (N_26162,N_25189,N_25274);
or U26163 (N_26163,N_25577,N_25463);
and U26164 (N_26164,N_24380,N_25461);
nor U26165 (N_26165,N_25804,N_25689);
and U26166 (N_26166,N_25633,N_25045);
xor U26167 (N_26167,N_25618,N_24989);
and U26168 (N_26168,N_24428,N_25091);
nand U26169 (N_26169,N_25707,N_25446);
nor U26170 (N_26170,N_25772,N_24969);
and U26171 (N_26171,N_25815,N_24884);
or U26172 (N_26172,N_24122,N_24424);
and U26173 (N_26173,N_25882,N_24146);
or U26174 (N_26174,N_25803,N_25183);
and U26175 (N_26175,N_25156,N_25958);
or U26176 (N_26176,N_25896,N_25500);
or U26177 (N_26177,N_25225,N_24946);
xor U26178 (N_26178,N_25549,N_25082);
xnor U26179 (N_26179,N_25751,N_25868);
or U26180 (N_26180,N_25818,N_24408);
nor U26181 (N_26181,N_25414,N_25197);
and U26182 (N_26182,N_24541,N_25728);
nor U26183 (N_26183,N_25016,N_24911);
nor U26184 (N_26184,N_25683,N_24981);
nor U26185 (N_26185,N_25963,N_24069);
or U26186 (N_26186,N_25951,N_24023);
xnor U26187 (N_26187,N_24721,N_24469);
or U26188 (N_26188,N_25642,N_25790);
xor U26189 (N_26189,N_25545,N_24645);
nand U26190 (N_26190,N_25512,N_24192);
and U26191 (N_26191,N_24495,N_25645);
or U26192 (N_26192,N_25306,N_25478);
xor U26193 (N_26193,N_25021,N_25761);
or U26194 (N_26194,N_24195,N_24301);
nand U26195 (N_26195,N_25935,N_24411);
xnor U26196 (N_26196,N_24783,N_24904);
or U26197 (N_26197,N_25404,N_25063);
and U26198 (N_26198,N_24777,N_25036);
and U26199 (N_26199,N_25365,N_25255);
xor U26200 (N_26200,N_25810,N_25572);
and U26201 (N_26201,N_25002,N_24717);
and U26202 (N_26202,N_24363,N_25960);
or U26203 (N_26203,N_25254,N_25979);
or U26204 (N_26204,N_25808,N_24853);
xnor U26205 (N_26205,N_24954,N_25003);
and U26206 (N_26206,N_25064,N_24790);
nor U26207 (N_26207,N_24942,N_24644);
or U26208 (N_26208,N_24697,N_25423);
and U26209 (N_26209,N_24193,N_24639);
and U26210 (N_26210,N_24349,N_24848);
nor U26211 (N_26211,N_24172,N_24143);
and U26212 (N_26212,N_25542,N_24515);
nand U26213 (N_26213,N_25302,N_25783);
nor U26214 (N_26214,N_25522,N_24091);
xnor U26215 (N_26215,N_25724,N_24664);
nand U26216 (N_26216,N_24482,N_24319);
or U26217 (N_26217,N_25941,N_25971);
or U26218 (N_26218,N_24288,N_25123);
nor U26219 (N_26219,N_24191,N_25206);
nor U26220 (N_26220,N_24130,N_25675);
and U26221 (N_26221,N_24207,N_24080);
nor U26222 (N_26222,N_24908,N_24189);
or U26223 (N_26223,N_25346,N_25826);
nand U26224 (N_26224,N_24633,N_24508);
nor U26225 (N_26225,N_24382,N_24905);
nand U26226 (N_26226,N_25480,N_24573);
or U26227 (N_26227,N_25252,N_25472);
nor U26228 (N_26228,N_24222,N_25929);
or U26229 (N_26229,N_24181,N_25118);
xor U26230 (N_26230,N_24142,N_25526);
xor U26231 (N_26231,N_25760,N_25190);
xor U26232 (N_26232,N_24286,N_24860);
nor U26233 (N_26233,N_25470,N_25144);
nand U26234 (N_26234,N_24967,N_25131);
xnor U26235 (N_26235,N_25372,N_25991);
nand U26236 (N_26236,N_25959,N_24008);
and U26237 (N_26237,N_25492,N_25574);
nand U26238 (N_26238,N_25543,N_24211);
or U26239 (N_26239,N_25066,N_24687);
or U26240 (N_26240,N_25359,N_25433);
and U26241 (N_26241,N_24450,N_24830);
nor U26242 (N_26242,N_24881,N_24140);
and U26243 (N_26243,N_25065,N_24779);
nand U26244 (N_26244,N_25553,N_24617);
and U26245 (N_26245,N_25048,N_25357);
nor U26246 (N_26246,N_25347,N_25521);
nand U26247 (N_26247,N_25682,N_24602);
and U26248 (N_26248,N_24353,N_24528);
and U26249 (N_26249,N_25600,N_24356);
xor U26250 (N_26250,N_24040,N_25532);
and U26251 (N_26251,N_25712,N_25029);
and U26252 (N_26252,N_24024,N_24551);
and U26253 (N_26253,N_25031,N_25738);
and U26254 (N_26254,N_24294,N_25603);
xnor U26255 (N_26255,N_25536,N_25422);
or U26256 (N_26256,N_25447,N_25106);
or U26257 (N_26257,N_24665,N_24133);
xnor U26258 (N_26258,N_24545,N_24497);
and U26259 (N_26259,N_24029,N_25001);
nand U26260 (N_26260,N_25226,N_24618);
or U26261 (N_26261,N_25389,N_24944);
nand U26262 (N_26262,N_24215,N_24157);
xnor U26263 (N_26263,N_24097,N_25848);
or U26264 (N_26264,N_25792,N_24743);
nand U26265 (N_26265,N_24973,N_24017);
nand U26266 (N_26266,N_25757,N_25527);
or U26267 (N_26267,N_24109,N_25686);
or U26268 (N_26268,N_25665,N_24056);
nand U26269 (N_26269,N_25895,N_24519);
nand U26270 (N_26270,N_25944,N_25328);
nor U26271 (N_26271,N_25915,N_25737);
xnor U26272 (N_26272,N_25721,N_24898);
xor U26273 (N_26273,N_25007,N_24739);
nand U26274 (N_26274,N_24916,N_24680);
or U26275 (N_26275,N_25714,N_24151);
or U26276 (N_26276,N_24226,N_25716);
and U26277 (N_26277,N_25644,N_25883);
nand U26278 (N_26278,N_24562,N_25195);
nor U26279 (N_26279,N_24922,N_24275);
or U26280 (N_26280,N_25517,N_25974);
nand U26281 (N_26281,N_24049,N_24948);
xor U26282 (N_26282,N_24965,N_25776);
nand U26283 (N_26283,N_24549,N_24554);
or U26284 (N_26284,N_24643,N_24574);
xor U26285 (N_26285,N_24397,N_24896);
xnor U26286 (N_26286,N_24746,N_24464);
and U26287 (N_26287,N_25089,N_25528);
and U26288 (N_26288,N_24880,N_25854);
nand U26289 (N_26289,N_25318,N_24441);
nor U26290 (N_26290,N_25925,N_25047);
nor U26291 (N_26291,N_25857,N_25989);
xor U26292 (N_26292,N_25051,N_25599);
nor U26293 (N_26293,N_25027,N_25562);
or U26294 (N_26294,N_25513,N_24127);
xor U26295 (N_26295,N_24804,N_25884);
nand U26296 (N_26296,N_25663,N_25948);
nor U26297 (N_26297,N_24585,N_25952);
xnor U26298 (N_26298,N_25041,N_24947);
and U26299 (N_26299,N_24828,N_25300);
xor U26300 (N_26300,N_25127,N_24112);
nor U26301 (N_26301,N_24366,N_24742);
and U26302 (N_26302,N_25748,N_24679);
xor U26303 (N_26303,N_25042,N_25789);
nor U26304 (N_26304,N_25060,N_24309);
or U26305 (N_26305,N_25015,N_25586);
or U26306 (N_26306,N_25840,N_25846);
nand U26307 (N_26307,N_25997,N_24520);
nor U26308 (N_26308,N_24402,N_25133);
nor U26309 (N_26309,N_24971,N_25208);
xor U26310 (N_26310,N_24489,N_24262);
nor U26311 (N_26311,N_25967,N_24284);
nand U26312 (N_26312,N_24420,N_24125);
nand U26313 (N_26313,N_24048,N_24897);
xnor U26314 (N_26314,N_24940,N_25174);
or U26315 (N_26315,N_25275,N_25550);
or U26316 (N_26316,N_24527,N_25524);
nor U26317 (N_26317,N_25248,N_25203);
and U26318 (N_26318,N_24426,N_24223);
nor U26319 (N_26319,N_24392,N_25486);
nand U26320 (N_26320,N_25151,N_24851);
nor U26321 (N_26321,N_24513,N_25864);
nor U26322 (N_26322,N_25755,N_24755);
xnor U26323 (N_26323,N_25858,N_24409);
or U26324 (N_26324,N_25544,N_24320);
or U26325 (N_26325,N_24338,N_24599);
nand U26326 (N_26326,N_25606,N_24507);
and U26327 (N_26327,N_24787,N_25279);
xnor U26328 (N_26328,N_25028,N_25192);
nor U26329 (N_26329,N_24774,N_24924);
or U26330 (N_26330,N_24243,N_25498);
or U26331 (N_26331,N_24544,N_25233);
nor U26332 (N_26332,N_25917,N_24737);
nor U26333 (N_26333,N_25623,N_24490);
xnor U26334 (N_26334,N_25657,N_25410);
xnor U26335 (N_26335,N_24480,N_25908);
and U26336 (N_26336,N_24772,N_25972);
or U26337 (N_26337,N_25088,N_25288);
and U26338 (N_26338,N_25315,N_25520);
xor U26339 (N_26339,N_25143,N_24396);
xnor U26340 (N_26340,N_24870,N_25829);
nor U26341 (N_26341,N_25432,N_24183);
nor U26342 (N_26342,N_24376,N_24857);
nor U26343 (N_26343,N_25276,N_24076);
xnor U26344 (N_26344,N_24894,N_24416);
nand U26345 (N_26345,N_25308,N_25119);
or U26346 (N_26346,N_25676,N_24266);
and U26347 (N_26347,N_24345,N_24867);
and U26348 (N_26348,N_24521,N_25220);
and U26349 (N_26349,N_25342,N_25307);
nand U26350 (N_26350,N_24368,N_25678);
or U26351 (N_26351,N_24522,N_25000);
nor U26352 (N_26352,N_25056,N_25138);
and U26353 (N_26353,N_25092,N_24970);
and U26354 (N_26354,N_24845,N_24234);
xnor U26355 (N_26355,N_24928,N_25648);
and U26356 (N_26356,N_24107,N_24196);
xnor U26357 (N_26357,N_24820,N_25333);
nor U26358 (N_26358,N_24869,N_25684);
xnor U26359 (N_26359,N_25885,N_24359);
and U26360 (N_26360,N_24756,N_24635);
xnor U26361 (N_26361,N_25380,N_25052);
xor U26362 (N_26362,N_25379,N_25638);
nor U26363 (N_26363,N_24765,N_24252);
nand U26364 (N_26364,N_24572,N_25785);
nand U26365 (N_26365,N_24199,N_24375);
and U26366 (N_26366,N_25832,N_25823);
nor U26367 (N_26367,N_25863,N_24483);
nor U26368 (N_26368,N_24891,N_24773);
nand U26369 (N_26369,N_24206,N_24931);
xor U26370 (N_26370,N_25078,N_24289);
and U26371 (N_26371,N_24115,N_24137);
nor U26372 (N_26372,N_24978,N_25655);
nand U26373 (N_26373,N_25242,N_24512);
and U26374 (N_26374,N_25515,N_25104);
nor U26375 (N_26375,N_24594,N_25805);
or U26376 (N_26376,N_25055,N_24265);
xnor U26377 (N_26377,N_24710,N_25193);
nor U26378 (N_26378,N_24187,N_24579);
and U26379 (N_26379,N_25334,N_25535);
or U26380 (N_26380,N_24877,N_24646);
or U26381 (N_26381,N_24317,N_25167);
nor U26382 (N_26382,N_25639,N_24169);
and U26383 (N_26383,N_25583,N_25085);
nor U26384 (N_26384,N_25329,N_24003);
nor U26385 (N_26385,N_24731,N_24475);
and U26386 (N_26386,N_24563,N_25627);
nor U26387 (N_26387,N_24404,N_24913);
xnor U26388 (N_26388,N_25257,N_24391);
nor U26389 (N_26389,N_24631,N_25409);
or U26390 (N_26390,N_24647,N_25450);
xnor U26391 (N_26391,N_24567,N_24603);
nand U26392 (N_26392,N_25355,N_25869);
or U26393 (N_26393,N_24316,N_24209);
xor U26394 (N_26394,N_24690,N_24511);
nand U26395 (N_26395,N_24678,N_24529);
nor U26396 (N_26396,N_25809,N_25926);
xor U26397 (N_26397,N_24691,N_24800);
nor U26398 (N_26398,N_25280,N_25299);
xnor U26399 (N_26399,N_25630,N_24837);
and U26400 (N_26400,N_24451,N_24403);
nand U26401 (N_26401,N_25752,N_25555);
and U26402 (N_26402,N_24984,N_25980);
or U26403 (N_26403,N_24909,N_25212);
xor U26404 (N_26404,N_24010,N_25622);
nand U26405 (N_26405,N_25020,N_25122);
and U26406 (N_26406,N_25093,N_24822);
nor U26407 (N_26407,N_24925,N_24805);
and U26408 (N_26408,N_24689,N_25510);
xor U26409 (N_26409,N_25667,N_25330);
nand U26410 (N_26410,N_24580,N_24190);
nand U26411 (N_26411,N_24168,N_24827);
xor U26412 (N_26412,N_24531,N_25474);
nor U26413 (N_26413,N_24933,N_24829);
xor U26414 (N_26414,N_24791,N_24129);
or U26415 (N_26415,N_24292,N_25990);
nand U26416 (N_26416,N_24575,N_25601);
nor U26417 (N_26417,N_25247,N_25018);
xor U26418 (N_26418,N_24474,N_25596);
and U26419 (N_26419,N_24304,N_24538);
nor U26420 (N_26420,N_25102,N_24188);
and U26421 (N_26421,N_24461,N_25747);
or U26422 (N_26422,N_24227,N_24117);
xor U26423 (N_26423,N_24939,N_24267);
xor U26424 (N_26424,N_24446,N_24950);
nand U26425 (N_26425,N_24516,N_24514);
and U26426 (N_26426,N_25250,N_24171);
xnor U26427 (N_26427,N_24072,N_24695);
and U26428 (N_26428,N_24164,N_25292);
and U26429 (N_26429,N_25136,N_24182);
nor U26430 (N_26430,N_24429,N_24417);
or U26431 (N_26431,N_24026,N_25888);
nand U26432 (N_26432,N_24659,N_24071);
nor U26433 (N_26433,N_24581,N_24279);
xor U26434 (N_26434,N_25256,N_24034);
or U26435 (N_26435,N_24090,N_25481);
and U26436 (N_26436,N_25425,N_25530);
nand U26437 (N_26437,N_24788,N_24886);
nor U26438 (N_26438,N_25694,N_25701);
nor U26439 (N_26439,N_25921,N_24493);
nor U26440 (N_26440,N_24378,N_24178);
or U26441 (N_26441,N_25381,N_24134);
xnor U26442 (N_26442,N_25278,N_25664);
nor U26443 (N_26443,N_24834,N_24840);
nand U26444 (N_26444,N_24036,N_24943);
nor U26445 (N_26445,N_25229,N_24005);
nor U26446 (N_26446,N_24702,N_24839);
nand U26447 (N_26447,N_24260,N_24110);
nand U26448 (N_26448,N_24208,N_25604);
or U26449 (N_26449,N_25343,N_24786);
nor U26450 (N_26450,N_25795,N_24901);
nand U26451 (N_26451,N_24254,N_25831);
and U26452 (N_26452,N_24655,N_25698);
or U26453 (N_26453,N_24566,N_25107);
and U26454 (N_26454,N_24729,N_24525);
and U26455 (N_26455,N_24430,N_24242);
xnor U26456 (N_26456,N_24161,N_24253);
nand U26457 (N_26457,N_24675,N_25224);
nor U26458 (N_26458,N_24321,N_24748);
xor U26459 (N_26459,N_24921,N_24256);
nand U26460 (N_26460,N_24020,N_25268);
xor U26461 (N_26461,N_25431,N_25181);
and U26462 (N_26462,N_25505,N_25945);
nand U26463 (N_26463,N_25575,N_24160);
and U26464 (N_26464,N_24273,N_24467);
nand U26465 (N_26465,N_24670,N_24263);
xnor U26466 (N_26466,N_24433,N_25977);
and U26467 (N_26467,N_24067,N_25853);
nand U26468 (N_26468,N_24699,N_25983);
xnor U26469 (N_26469,N_24101,N_25637);
or U26470 (N_26470,N_24098,N_25019);
nor U26471 (N_26471,N_24398,N_24821);
nand U26472 (N_26472,N_24006,N_25674);
and U26473 (N_26473,N_25651,N_24795);
nand U26474 (N_26474,N_25468,N_24749);
xor U26475 (N_26475,N_24613,N_24228);
xor U26476 (N_26476,N_25734,N_25580);
and U26477 (N_26477,N_24672,N_24701);
and U26478 (N_26478,N_24308,N_25696);
nor U26479 (N_26479,N_25086,N_25539);
and U26480 (N_26480,N_24590,N_25084);
and U26481 (N_26481,N_24607,N_24175);
nor U26482 (N_26482,N_24314,N_24332);
nand U26483 (N_26483,N_25838,N_24912);
xnor U26484 (N_26484,N_25514,N_24698);
and U26485 (N_26485,N_24660,N_24197);
or U26486 (N_26486,N_24584,N_25495);
nor U26487 (N_26487,N_24453,N_24593);
or U26488 (N_26488,N_25534,N_25780);
or U26489 (N_26489,N_24344,N_24186);
nor U26490 (N_26490,N_24623,N_24759);
or U26491 (N_26491,N_25825,N_25341);
and U26492 (N_26492,N_25321,N_25609);
nand U26493 (N_26493,N_24445,N_25588);
nand U26494 (N_26494,N_25083,N_25146);
and U26495 (N_26495,N_25383,N_25236);
nor U26496 (N_26496,N_24022,N_25661);
or U26497 (N_26497,N_24324,N_24866);
or U26498 (N_26498,N_24553,N_25843);
xnor U26499 (N_26499,N_24414,N_25435);
nand U26500 (N_26500,N_25511,N_24074);
and U26501 (N_26501,N_24638,N_24360);
nor U26502 (N_26502,N_25641,N_25076);
nor U26503 (N_26503,N_24974,N_24606);
nor U26504 (N_26504,N_25004,N_24751);
or U26505 (N_26505,N_25336,N_25640);
xor U26506 (N_26506,N_24918,N_25096);
nand U26507 (N_26507,N_24524,N_24899);
xor U26508 (N_26508,N_25178,N_24220);
nor U26509 (N_26509,N_24019,N_25062);
nand U26510 (N_26510,N_24092,N_24124);
xnor U26511 (N_26511,N_25719,N_24761);
and U26512 (N_26512,N_25867,N_25852);
xor U26513 (N_26513,N_24248,N_25260);
nor U26514 (N_26514,N_24103,N_24423);
and U26515 (N_26515,N_24733,N_25169);
nor U26516 (N_26516,N_25540,N_25109);
nor U26517 (N_26517,N_24419,N_25660);
and U26518 (N_26518,N_25024,N_24300);
xor U26519 (N_26519,N_25898,N_24315);
nand U26520 (N_26520,N_25475,N_24784);
nor U26521 (N_26521,N_24487,N_24615);
nor U26522 (N_26522,N_25746,N_24712);
nand U26523 (N_26523,N_24148,N_24803);
nor U26524 (N_26524,N_24179,N_24807);
and U26525 (N_26525,N_24238,N_25199);
or U26526 (N_26526,N_25469,N_25509);
nand U26527 (N_26527,N_24121,N_25756);
nor U26528 (N_26528,N_24952,N_25628);
xor U26529 (N_26529,N_24961,N_24624);
xor U26530 (N_26530,N_24473,N_25956);
nor U26531 (N_26531,N_24873,N_24619);
nand U26532 (N_26532,N_25680,N_25467);
nor U26533 (N_26533,N_24013,N_24858);
nor U26534 (N_26534,N_24766,N_24704);
and U26535 (N_26535,N_24601,N_24232);
or U26536 (N_26536,N_25584,N_25058);
and U26537 (N_26537,N_24162,N_24650);
nor U26538 (N_26538,N_25814,N_24166);
and U26539 (N_26539,N_25688,N_24058);
xnor U26540 (N_26540,N_24149,N_24862);
xnor U26541 (N_26541,N_25162,N_24611);
nand U26542 (N_26542,N_24485,N_25163);
nand U26543 (N_26543,N_25548,N_25799);
nand U26544 (N_26544,N_25636,N_24768);
nor U26545 (N_26545,N_25907,N_25168);
and U26546 (N_26546,N_25304,N_24608);
xor U26547 (N_26547,N_25670,N_24686);
nor U26548 (N_26548,N_24953,N_24167);
nand U26549 (N_26549,N_24833,N_25081);
nor U26550 (N_26550,N_24210,N_25354);
nor U26551 (N_26551,N_24364,N_24705);
xor U26552 (N_26552,N_24333,N_25371);
and U26553 (N_26553,N_25444,N_25793);
nand U26554 (N_26554,N_25070,N_24337);
nor U26555 (N_26555,N_24841,N_24671);
nor U26556 (N_26556,N_25834,N_25362);
nand U26557 (N_26557,N_25504,N_25097);
xor U26558 (N_26558,N_25352,N_25177);
or U26559 (N_26559,N_24823,N_24449);
nand U26560 (N_26560,N_24658,N_24985);
and U26561 (N_26561,N_24977,N_24636);
xnor U26562 (N_26562,N_24271,N_24986);
and U26563 (N_26563,N_25781,N_24331);
nor U26564 (N_26564,N_25611,N_25459);
xor U26565 (N_26565,N_25733,N_25059);
and U26566 (N_26566,N_25496,N_25132);
and U26567 (N_26567,N_24105,N_25272);
xor U26568 (N_26568,N_24249,N_24233);
and U26569 (N_26569,N_25115,N_25428);
nor U26570 (N_26570,N_25191,N_25541);
or U26571 (N_26571,N_24393,N_25693);
nor U26572 (N_26572,N_25740,N_25166);
or U26573 (N_26573,N_24990,N_24630);
xnor U26574 (N_26574,N_24431,N_24547);
and U26575 (N_26575,N_25301,N_24384);
xor U26576 (N_26576,N_24797,N_25978);
nor U26577 (N_26577,N_24214,N_24666);
nor U26578 (N_26578,N_25629,N_25437);
nand U26579 (N_26579,N_24302,N_25073);
and U26580 (N_26580,N_25125,N_24676);
and U26581 (N_26581,N_25079,N_24099);
nand U26582 (N_26582,N_24889,N_25635);
nor U26583 (N_26583,N_24230,N_24815);
nand U26584 (N_26584,N_25659,N_25791);
xor U26585 (N_26585,N_25827,N_25142);
xnor U26586 (N_26586,N_25263,N_24439);
or U26587 (N_26587,N_24673,N_24086);
and U26588 (N_26588,N_24358,N_24711);
nor U26589 (N_26589,N_25361,N_25900);
nor U26590 (N_26590,N_24734,N_25008);
and U26591 (N_26591,N_24730,N_24652);
or U26592 (N_26592,N_25267,N_25187);
xnor U26593 (N_26593,N_24741,N_24421);
xor U26594 (N_26594,N_25506,N_25427);
or U26595 (N_26595,N_25842,N_25871);
xor U26596 (N_26596,N_24083,N_25982);
or U26597 (N_26597,N_25996,N_25223);
nand U26598 (N_26598,N_25128,N_25186);
xor U26599 (N_26599,N_24041,N_25441);
or U26600 (N_26600,N_24476,N_24900);
nand U26601 (N_26601,N_24425,N_25443);
nand U26602 (N_26602,N_25554,N_25295);
nor U26603 (N_26603,N_25429,N_24735);
nand U26604 (N_26604,N_24883,N_25006);
and U26605 (N_26605,N_25820,N_25744);
xnor U26606 (N_26606,N_25730,N_25464);
nand U26607 (N_26607,N_25397,N_24077);
and U26608 (N_26608,N_25101,N_25283);
or U26609 (N_26609,N_25095,N_25421);
or U26610 (N_26610,N_24369,N_24216);
xor U26611 (N_26611,N_24814,N_25416);
nor U26612 (N_26612,N_24592,N_24073);
or U26613 (N_26613,N_25349,N_25438);
and U26614 (N_26614,N_24108,N_24991);
nor U26615 (N_26615,N_24876,N_25164);
or U26616 (N_26616,N_25892,N_25501);
nor U26617 (N_26617,N_25836,N_25576);
and U26618 (N_26618,N_25523,N_24539);
and U26619 (N_26619,N_25277,N_24696);
and U26620 (N_26620,N_24736,N_25597);
nor U26621 (N_26621,N_25889,N_25011);
nand U26622 (N_26622,N_25204,N_25987);
nor U26623 (N_26623,N_25209,N_25452);
or U26624 (N_26624,N_24945,N_24796);
and U26625 (N_26625,N_25771,N_25802);
nand U26626 (N_26626,N_25891,N_24568);
or U26627 (N_26627,N_25434,N_24502);
or U26628 (N_26628,N_25175,N_25672);
and U26629 (N_26629,N_25893,N_24027);
and U26630 (N_26630,N_25614,N_25353);
xnor U26631 (N_26631,N_24357,N_25742);
xor U26632 (N_26632,N_24764,N_24622);
nor U26633 (N_26633,N_25904,N_24640);
or U26634 (N_26634,N_25766,N_24793);
xnor U26635 (N_26635,N_24958,N_24914);
nand U26636 (N_26636,N_25881,N_25139);
nand U26637 (N_26637,N_24296,N_24158);
and U26638 (N_26638,N_25565,N_25332);
or U26639 (N_26639,N_24715,N_24856);
and U26640 (N_26640,N_24340,N_24504);
nand U26641 (N_26641,N_24963,N_24625);
nor U26642 (N_26642,N_25417,N_24247);
nor U26643 (N_26643,N_24923,N_25217);
nor U26644 (N_26644,N_24463,N_25679);
nor U26645 (N_26645,N_25916,N_24202);
and U26646 (N_26646,N_25847,N_24588);
or U26647 (N_26647,N_25913,N_24153);
nor U26648 (N_26648,N_25965,N_24185);
nand U26649 (N_26649,N_24861,N_24930);
or U26650 (N_26650,N_25188,N_25141);
or U26651 (N_26651,N_24503,N_25582);
nor U26652 (N_26652,N_25608,N_25105);
nor U26653 (N_26653,N_24257,N_25666);
or U26654 (N_26654,N_24937,N_25992);
nand U26655 (N_26655,N_24838,N_24053);
nor U26656 (N_26656,N_24849,N_24683);
xnor U26657 (N_26657,N_25477,N_24802);
xnor U26658 (N_26658,N_25706,N_25243);
nand U26659 (N_26659,N_25763,N_25130);
or U26660 (N_26660,N_25285,N_24246);
xnor U26661 (N_26661,N_25099,N_24462);
xor U26662 (N_26662,N_25940,N_25057);
and U26663 (N_26663,N_25726,N_25561);
xnor U26664 (N_26664,N_24334,N_24468);
nand U26665 (N_26665,N_24159,N_24025);
nand U26666 (N_26666,N_24221,N_25699);
xor U26667 (N_26667,N_25581,N_25729);
or U26668 (N_26668,N_24050,N_24583);
xnor U26669 (N_26669,N_24035,N_24510);
nand U26670 (N_26670,N_25590,N_24395);
or U26671 (N_26671,N_24106,N_25430);
and U26672 (N_26672,N_24059,N_25794);
nand U26673 (N_26673,N_24471,N_24959);
xnor U26674 (N_26674,N_25984,N_25228);
nor U26675 (N_26675,N_24750,N_24968);
and U26676 (N_26676,N_24455,N_25845);
nand U26677 (N_26677,N_25874,N_24605);
and U26678 (N_26678,N_24123,N_25296);
xnor U26679 (N_26679,N_24365,N_24667);
or U26680 (N_26680,N_24720,N_24460);
xnor U26681 (N_26681,N_25305,N_25516);
nand U26682 (N_26682,N_24448,N_25074);
nand U26683 (N_26683,N_24173,N_24355);
nor U26684 (N_26684,N_24887,N_25491);
and U26685 (N_26685,N_24614,N_25811);
nand U26686 (N_26686,N_25014,N_25390);
and U26687 (N_26687,N_25179,N_25859);
and U26688 (N_26688,N_25796,N_24775);
and U26689 (N_26689,N_24217,N_25947);
or U26690 (N_26690,N_25201,N_24039);
xnor U26691 (N_26691,N_25198,N_25578);
xor U26692 (N_26692,N_24782,N_25546);
nor U26693 (N_26693,N_25399,N_24801);
or U26694 (N_26694,N_25113,N_25316);
and U26695 (N_26695,N_24138,N_25800);
xor U26696 (N_26696,N_24962,N_25317);
or U26697 (N_26697,N_25215,N_24654);
nor U26698 (N_26698,N_25289,N_24917);
nor U26699 (N_26699,N_25975,N_25615);
nor U26700 (N_26700,N_24385,N_24960);
nor U26701 (N_26701,N_25384,N_25281);
and U26702 (N_26702,N_24767,N_25244);
xor U26703 (N_26703,N_25731,N_24498);
nand U26704 (N_26704,N_24383,N_24656);
nand U26705 (N_26705,N_24850,N_25662);
or U26706 (N_26706,N_24612,N_25957);
xor U26707 (N_26707,N_24546,N_25160);
nor U26708 (N_26708,N_25877,N_25968);
nand U26709 (N_26709,N_24728,N_25314);
nand U26710 (N_26710,N_25394,N_25981);
xor U26711 (N_26711,N_24119,N_25108);
nor U26712 (N_26712,N_24726,N_24055);
xor U26713 (N_26713,N_24282,N_25720);
xor U26714 (N_26714,N_25922,N_25879);
nor U26715 (N_26715,N_25502,N_25753);
xor U26716 (N_26716,N_24287,N_24009);
nor U26717 (N_26717,N_24484,N_24609);
nor U26718 (N_26718,N_25261,N_24628);
and U26719 (N_26719,N_25988,N_24412);
nor U26720 (N_26720,N_25995,N_24543);
nor U26721 (N_26721,N_24653,N_24060);
xnor U26722 (N_26722,N_25351,N_24093);
nor U26723 (N_26723,N_25216,N_24180);
xor U26724 (N_26724,N_25993,N_25700);
nor U26725 (N_26725,N_24637,N_25643);
xor U26726 (N_26726,N_24335,N_25054);
or U26727 (N_26727,N_25758,N_24043);
nor U26728 (N_26728,N_24578,N_25741);
and U26729 (N_26729,N_24934,N_25165);
and U26730 (N_26730,N_25451,N_24285);
nand U26731 (N_26731,N_24816,N_24322);
nand U26732 (N_26732,N_25479,N_24763);
nor U26733 (N_26733,N_24054,N_24374);
nand U26734 (N_26734,N_24176,N_25327);
or U26735 (N_26735,N_25594,N_24576);
nor U26736 (N_26736,N_24277,N_24377);
and U26737 (N_26737,N_25692,N_24852);
and U26738 (N_26738,N_24339,N_24231);
nor U26739 (N_26739,N_24235,N_25110);
xor U26740 (N_26740,N_25497,N_24269);
xnor U26741 (N_26741,N_25754,N_25503);
and U26742 (N_26742,N_25009,N_24570);
xor U26743 (N_26743,N_24205,N_25071);
and U26744 (N_26744,N_25844,N_25413);
and U26745 (N_26745,N_24842,N_24481);
or U26746 (N_26746,N_25035,N_24405);
nand U26747 (N_26747,N_25787,N_25759);
nand U26748 (N_26748,N_24437,N_24152);
and U26749 (N_26749,N_25238,N_24600);
and U26750 (N_26750,N_25114,N_24014);
nor U26751 (N_26751,N_25920,N_24740);
and U26752 (N_26752,N_25456,N_25424);
and U26753 (N_26753,N_24018,N_25454);
nand U26754 (N_26754,N_25218,N_25703);
xor U26755 (N_26755,N_25872,N_24596);
xnor U26756 (N_26756,N_25222,N_24347);
xnor U26757 (N_26757,N_24203,N_24548);
xnor U26758 (N_26758,N_25485,N_24598);
and U26759 (N_26759,N_24102,N_24255);
and U26760 (N_26760,N_24486,N_25566);
nand U26761 (N_26761,N_25023,N_24972);
nand U26762 (N_26762,N_24354,N_24361);
xor U26763 (N_26763,N_24932,N_25436);
nor U26764 (N_26764,N_25617,N_24983);
or U26765 (N_26765,N_25722,N_24505);
or U26766 (N_26766,N_25839,N_25725);
or U26767 (N_26767,N_25231,N_25841);
and U26768 (N_26768,N_24492,N_25556);
or U26769 (N_26769,N_25090,N_24532);
nor U26770 (N_26770,N_25476,N_24988);
xnor U26771 (N_26771,N_24888,N_25072);
nand U26772 (N_26772,N_25010,N_24855);
nor U26773 (N_26773,N_25025,N_25013);
nor U26774 (N_26774,N_24371,N_25324);
or U26775 (N_26775,N_24132,N_24996);
nand U26776 (N_26776,N_25259,N_25938);
nor U26777 (N_26777,N_25140,N_24798);
and U26778 (N_26778,N_24979,N_25249);
or U26779 (N_26779,N_24341,N_25487);
and U26780 (N_26780,N_24552,N_25559);
nor U26781 (N_26781,N_24065,N_25442);
nor U26782 (N_26782,N_25439,N_24506);
or U26783 (N_26783,N_24094,N_25649);
nor U26784 (N_26784,N_25695,N_24557);
nor U26785 (N_26785,N_24571,N_25214);
and U26786 (N_26786,N_25388,N_24949);
nand U26787 (N_26787,N_25673,N_25866);
or U26788 (N_26788,N_25717,N_25046);
xnor U26789 (N_26789,N_24685,N_25710);
xnor U26790 (N_26790,N_24663,N_25650);
nor U26791 (N_26791,N_25145,N_25563);
nand U26792 (N_26792,N_24031,N_24194);
or U26793 (N_26793,N_24410,N_25264);
and U26794 (N_26794,N_24719,N_24200);
and U26795 (N_26795,N_25038,N_25387);
and U26796 (N_26796,N_24762,N_25147);
and U26797 (N_26797,N_24770,N_25906);
xor U26798 (N_26798,N_24589,N_24682);
xnor U26799 (N_26799,N_24708,N_25373);
xor U26800 (N_26800,N_25325,N_24415);
nand U26801 (N_26801,N_25392,N_24935);
nand U26802 (N_26802,N_25310,N_24470);
and U26803 (N_26803,N_24477,N_24047);
and U26804 (N_26804,N_24536,N_25471);
nand U26805 (N_26805,N_25878,N_24718);
or U26806 (N_26806,N_25739,N_25998);
xnor U26807 (N_26807,N_25157,N_25488);
or U26808 (N_26808,N_24586,N_24951);
nor U26809 (N_26809,N_24472,N_24879);
nor U26810 (N_26810,N_24987,N_25850);
and U26811 (N_26811,N_24198,N_25103);
nor U26812 (N_26812,N_24781,N_24438);
nor U26813 (N_26813,N_24070,N_25518);
and U26814 (N_26814,N_24998,N_25813);
xor U26815 (N_26815,N_24693,N_25798);
xor U26816 (N_26816,N_24620,N_24488);
and U26817 (N_26817,N_25807,N_25455);
nor U26818 (N_26818,N_24478,N_24662);
or U26819 (N_26819,N_25564,N_25685);
or U26820 (N_26820,N_24399,N_25762);
or U26821 (N_26821,N_24015,N_24111);
xnor U26822 (N_26822,N_25533,N_25570);
nand U26823 (N_26823,N_25985,N_24813);
nand U26824 (N_26824,N_25408,N_25819);
or U26825 (N_26825,N_25919,N_24966);
or U26826 (N_26826,N_25942,N_25691);
and U26827 (N_26827,N_25708,N_24794);
or U26828 (N_26828,N_25923,N_24558);
or U26829 (N_26829,N_25449,N_24926);
nor U26830 (N_26830,N_25875,N_25210);
nor U26831 (N_26831,N_24435,N_24745);
nand U26832 (N_26832,N_25400,N_24387);
and U26833 (N_26833,N_24844,N_25531);
and U26834 (N_26834,N_25902,N_24422);
nand U26835 (N_26835,N_25493,N_24677);
nand U26836 (N_26836,N_25466,N_24350);
nand U26837 (N_26837,N_25345,N_25821);
nor U26838 (N_26838,N_24920,N_25851);
or U26839 (N_26839,N_25930,N_24902);
or U26840 (N_26840,N_24051,N_25625);
and U26841 (N_26841,N_24351,N_25723);
nand U26842 (N_26842,N_25339,N_24418);
nand U26843 (N_26843,N_25291,N_24836);
nor U26844 (N_26844,N_25797,N_24632);
nand U26845 (N_26845,N_25568,N_24370);
and U26846 (N_26846,N_25669,N_24057);
nor U26847 (N_26847,N_24669,N_24868);
nor U26848 (N_26848,N_25525,N_25287);
and U26849 (N_26849,N_25129,N_25856);
xnor U26850 (N_26850,N_24104,N_24542);
nor U26851 (N_26851,N_25765,N_24244);
and U26852 (N_26852,N_24118,N_25607);
and U26853 (N_26853,N_24236,N_24401);
nand U26854 (N_26854,N_25033,N_24725);
nor U26855 (N_26855,N_25121,N_25911);
xor U26856 (N_26856,N_24982,N_24095);
xnor U26857 (N_26857,N_25068,N_25393);
and U26858 (N_26858,N_24343,N_24241);
xnor U26859 (N_26859,N_25849,N_25172);
nor U26860 (N_26860,N_24245,N_24174);
nor U26861 (N_26861,N_25241,N_25012);
nor U26862 (N_26862,N_24135,N_24792);
nand U26863 (N_26863,N_24496,N_25273);
xor U26864 (N_26864,N_25743,N_25833);
xor U26865 (N_26865,N_25350,N_24626);
nor U26866 (N_26866,N_25161,N_25284);
nand U26867 (N_26867,N_24604,N_24724);
nand U26868 (N_26868,N_25415,N_24980);
and U26869 (N_26869,N_25551,N_24799);
xor U26870 (N_26870,N_24250,N_25293);
nor U26871 (N_26871,N_25207,N_25773);
nand U26872 (N_26872,N_24874,N_24535);
xor U26873 (N_26873,N_24442,N_25775);
and U26874 (N_26874,N_24261,N_25235);
nand U26875 (N_26875,N_25595,N_25298);
nor U26876 (N_26876,N_25358,N_25647);
or U26877 (N_26877,N_24700,N_24212);
or U26878 (N_26878,N_24780,N_25890);
nor U26879 (N_26879,N_25111,N_24778);
nor U26880 (N_26880,N_24444,N_24616);
xnor U26881 (N_26881,N_24184,N_24144);
nor U26882 (N_26882,N_25616,N_24388);
xor U26883 (N_26883,N_25171,N_24278);
xor U26884 (N_26884,N_25445,N_25927);
xnor U26885 (N_26885,N_25405,N_24597);
or U26886 (N_26886,N_25905,N_24064);
or U26887 (N_26887,N_24499,N_25153);
or U26888 (N_26888,N_24318,N_25270);
or U26889 (N_26889,N_24927,N_24033);
nor U26890 (N_26890,N_24713,N_24518);
or U26891 (N_26891,N_24413,N_25116);
and U26892 (N_26892,N_25134,N_25282);
and U26893 (N_26893,N_24434,N_24028);
or U26894 (N_26894,N_25297,N_24509);
nand U26895 (N_26895,N_24229,N_25837);
or U26896 (N_26896,N_25709,N_24846);
and U26897 (N_26897,N_24872,N_25937);
nor U26898 (N_26898,N_24494,N_25702);
or U26899 (N_26899,N_24021,N_25715);
xnor U26900 (N_26900,N_25184,N_25973);
nor U26901 (N_26901,N_24703,N_25567);
nand U26902 (N_26902,N_24561,N_24177);
nor U26903 (N_26903,N_25326,N_25039);
nor U26904 (N_26904,N_25017,N_25240);
nor U26905 (N_26905,N_24684,N_24154);
xnor U26906 (N_26906,N_24452,N_24714);
and U26907 (N_26907,N_25100,N_24085);
nand U26908 (N_26908,N_24835,N_25152);
or U26909 (N_26909,N_24440,N_24938);
and U26910 (N_26910,N_25170,N_25899);
and U26911 (N_26911,N_24610,N_24113);
and U26912 (N_26912,N_24465,N_25598);
or U26913 (N_26913,N_25828,N_25537);
nor U26914 (N_26914,N_25126,N_24957);
and U26915 (N_26915,N_25366,N_25322);
or U26916 (N_26916,N_24994,N_24150);
xnor U26917 (N_26917,N_25407,N_25044);
or U26918 (N_26918,N_25420,N_25955);
or U26919 (N_26919,N_24976,N_24629);
xnor U26920 (N_26920,N_25569,N_25148);
xor U26921 (N_26921,N_24313,N_24352);
and U26922 (N_26922,N_25571,N_24323);
and U26923 (N_26923,N_25697,N_24141);
xnor U26924 (N_26924,N_25303,N_24268);
xor U26925 (N_26925,N_25266,N_24280);
nor U26926 (N_26926,N_25232,N_24919);
nor U26927 (N_26927,N_24681,N_25080);
nand U26928 (N_26928,N_25067,N_25592);
or U26929 (N_26929,N_24291,N_24760);
or U26930 (N_26930,N_25994,N_24295);
and U26931 (N_26931,N_25117,N_24582);
nor U26932 (N_26932,N_25376,N_25589);
or U26933 (N_26933,N_24326,N_25262);
nand U26934 (N_26934,N_24089,N_25718);
or U26935 (N_26935,N_25529,N_25457);
and U26936 (N_26936,N_24533,N_24559);
or U26937 (N_26937,N_25778,N_24379);
or U26938 (N_26938,N_25767,N_25182);
nand U26939 (N_26939,N_25395,N_24427);
nor U26940 (N_26940,N_25690,N_25876);
and U26941 (N_26941,N_25124,N_24560);
xor U26942 (N_26942,N_24752,N_24810);
xnor U26943 (N_26943,N_25040,N_25870);
nand U26944 (N_26944,N_25219,N_25573);
and U26945 (N_26945,N_24079,N_24372);
nand U26946 (N_26946,N_25557,N_24649);
nand U26947 (N_26947,N_25835,N_25602);
xor U26948 (N_26948,N_25591,N_25382);
xnor U26949 (N_26949,N_24457,N_25135);
nor U26950 (N_26950,N_25176,N_25286);
and U26951 (N_26951,N_24311,N_25830);
xor U26952 (N_26952,N_25462,N_25861);
nor U26953 (N_26953,N_25745,N_25453);
nand U26954 (N_26954,N_25489,N_25239);
nand U26955 (N_26955,N_24272,N_25806);
and U26956 (N_26956,N_25862,N_25727);
nand U26957 (N_26957,N_24727,N_24312);
nand U26958 (N_26958,N_25547,N_24895);
nand U26959 (N_26959,N_24651,N_24785);
xor U26960 (N_26960,N_25246,N_25552);
nor U26961 (N_26961,N_25412,N_25631);
nand U26962 (N_26962,N_24325,N_25587);
nand U26963 (N_26963,N_24929,N_25613);
or U26964 (N_26964,N_25221,N_25656);
nand U26965 (N_26965,N_24225,N_25970);
nand U26966 (N_26966,N_25360,N_24373);
or U26967 (N_26967,N_24330,N_25816);
nand U26968 (N_26968,N_24864,N_24694);
or U26969 (N_26969,N_24163,N_25946);
nor U26970 (N_26970,N_25912,N_24875);
and U26971 (N_26971,N_24170,N_25269);
nand U26972 (N_26972,N_24709,N_24738);
nor U26973 (N_26973,N_25309,N_25377);
nand U26974 (N_26974,N_25205,N_24910);
xor U26975 (N_26975,N_24757,N_24139);
nor U26976 (N_26976,N_25860,N_24290);
or U26977 (N_26977,N_25155,N_25784);
and U26978 (N_26978,N_25370,N_25234);
nand U26979 (N_26979,N_24657,N_24052);
or U26980 (N_26980,N_24789,N_24819);
nand U26981 (N_26981,N_24032,N_24063);
xnor U26982 (N_26982,N_25897,N_25050);
nand U26983 (N_26983,N_24156,N_24878);
nor U26984 (N_26984,N_24456,N_25931);
nand U26985 (N_26985,N_25961,N_25094);
and U26986 (N_26986,N_25519,N_24744);
and U26987 (N_26987,N_25402,N_25750);
nor U26988 (N_26988,N_24147,N_24342);
nor U26989 (N_26989,N_24046,N_25954);
xnor U26990 (N_26990,N_24540,N_25824);
nor U26991 (N_26991,N_24030,N_24407);
xnor U26992 (N_26992,N_24128,N_24011);
and U26993 (N_26993,N_24955,N_25482);
and U26994 (N_26994,N_25865,N_24826);
xnor U26995 (N_26995,N_25180,N_25098);
or U26996 (N_26996,N_24012,N_25396);
nor U26997 (N_26997,N_25632,N_24120);
nor U26998 (N_26998,N_24999,N_24264);
nand U26999 (N_26999,N_24565,N_25986);
xor U27000 (N_27000,N_25351,N_25055);
nor U27001 (N_27001,N_24862,N_25508);
and U27002 (N_27002,N_25878,N_25815);
nor U27003 (N_27003,N_25157,N_24365);
nand U27004 (N_27004,N_24253,N_25948);
nor U27005 (N_27005,N_25841,N_24648);
nand U27006 (N_27006,N_24442,N_25845);
nor U27007 (N_27007,N_25909,N_24437);
nand U27008 (N_27008,N_25932,N_25807);
nor U27009 (N_27009,N_24521,N_25805);
nand U27010 (N_27010,N_25778,N_24969);
nand U27011 (N_27011,N_24263,N_25456);
xor U27012 (N_27012,N_24822,N_25559);
nor U27013 (N_27013,N_25973,N_25546);
or U27014 (N_27014,N_25185,N_24293);
nor U27015 (N_27015,N_24139,N_25798);
or U27016 (N_27016,N_25204,N_24194);
nor U27017 (N_27017,N_24119,N_24922);
nand U27018 (N_27018,N_25053,N_25425);
nor U27019 (N_27019,N_25113,N_25878);
xnor U27020 (N_27020,N_24021,N_25126);
or U27021 (N_27021,N_24781,N_25704);
xor U27022 (N_27022,N_24225,N_25792);
xnor U27023 (N_27023,N_25888,N_24545);
xor U27024 (N_27024,N_25284,N_24785);
nand U27025 (N_27025,N_25206,N_24572);
xor U27026 (N_27026,N_24230,N_25938);
or U27027 (N_27027,N_25467,N_24618);
xnor U27028 (N_27028,N_25813,N_25295);
and U27029 (N_27029,N_24888,N_24845);
and U27030 (N_27030,N_25505,N_25925);
and U27031 (N_27031,N_24918,N_24963);
xnor U27032 (N_27032,N_24808,N_25173);
or U27033 (N_27033,N_25843,N_25953);
nand U27034 (N_27034,N_24649,N_24077);
nor U27035 (N_27035,N_24871,N_25047);
or U27036 (N_27036,N_25731,N_25796);
and U27037 (N_27037,N_24021,N_24539);
nor U27038 (N_27038,N_24801,N_25403);
and U27039 (N_27039,N_24368,N_24806);
xor U27040 (N_27040,N_25882,N_25952);
nand U27041 (N_27041,N_25810,N_24857);
nor U27042 (N_27042,N_24495,N_24811);
nor U27043 (N_27043,N_25342,N_24302);
xor U27044 (N_27044,N_24186,N_25669);
or U27045 (N_27045,N_24576,N_24758);
nand U27046 (N_27046,N_24220,N_24660);
and U27047 (N_27047,N_25145,N_25935);
and U27048 (N_27048,N_25958,N_24558);
nand U27049 (N_27049,N_24980,N_25489);
nand U27050 (N_27050,N_24909,N_25369);
and U27051 (N_27051,N_24193,N_24049);
nand U27052 (N_27052,N_24156,N_24649);
xnor U27053 (N_27053,N_24363,N_24427);
nand U27054 (N_27054,N_24994,N_25286);
xnor U27055 (N_27055,N_24740,N_24872);
nor U27056 (N_27056,N_25509,N_25658);
nand U27057 (N_27057,N_25735,N_24852);
nor U27058 (N_27058,N_24073,N_24237);
nand U27059 (N_27059,N_24830,N_25708);
or U27060 (N_27060,N_25881,N_25495);
nor U27061 (N_27061,N_25496,N_25033);
xnor U27062 (N_27062,N_24701,N_24814);
or U27063 (N_27063,N_24390,N_25854);
nor U27064 (N_27064,N_24878,N_24828);
and U27065 (N_27065,N_24096,N_25827);
and U27066 (N_27066,N_24806,N_24683);
and U27067 (N_27067,N_25079,N_25481);
and U27068 (N_27068,N_24621,N_24423);
and U27069 (N_27069,N_25216,N_25468);
and U27070 (N_27070,N_25418,N_25767);
nor U27071 (N_27071,N_24694,N_25967);
or U27072 (N_27072,N_25479,N_24242);
and U27073 (N_27073,N_24620,N_24565);
and U27074 (N_27074,N_25929,N_24929);
xor U27075 (N_27075,N_24378,N_25957);
nor U27076 (N_27076,N_25621,N_25557);
nand U27077 (N_27077,N_24502,N_24349);
nor U27078 (N_27078,N_24246,N_24823);
nor U27079 (N_27079,N_25294,N_24525);
xnor U27080 (N_27080,N_24907,N_25233);
and U27081 (N_27081,N_25037,N_25247);
and U27082 (N_27082,N_24924,N_25448);
nor U27083 (N_27083,N_24772,N_24485);
xnor U27084 (N_27084,N_24504,N_24490);
nand U27085 (N_27085,N_24203,N_25763);
nand U27086 (N_27086,N_25067,N_24352);
nor U27087 (N_27087,N_25827,N_25458);
or U27088 (N_27088,N_24460,N_24685);
or U27089 (N_27089,N_24339,N_25040);
nor U27090 (N_27090,N_24642,N_25548);
xnor U27091 (N_27091,N_25491,N_25427);
xor U27092 (N_27092,N_25493,N_24204);
nand U27093 (N_27093,N_25801,N_24647);
nor U27094 (N_27094,N_24026,N_25902);
xor U27095 (N_27095,N_24543,N_25804);
and U27096 (N_27096,N_24650,N_24903);
nor U27097 (N_27097,N_25824,N_24682);
and U27098 (N_27098,N_25046,N_24130);
xor U27099 (N_27099,N_24701,N_24342);
nand U27100 (N_27100,N_24276,N_24831);
and U27101 (N_27101,N_25334,N_25389);
xnor U27102 (N_27102,N_25046,N_24853);
nor U27103 (N_27103,N_24395,N_24656);
or U27104 (N_27104,N_24566,N_25181);
nand U27105 (N_27105,N_24310,N_24114);
xnor U27106 (N_27106,N_24355,N_24507);
and U27107 (N_27107,N_24169,N_24624);
nor U27108 (N_27108,N_25479,N_25819);
and U27109 (N_27109,N_24301,N_25252);
and U27110 (N_27110,N_24796,N_25889);
nor U27111 (N_27111,N_25794,N_25282);
and U27112 (N_27112,N_25439,N_25393);
and U27113 (N_27113,N_25998,N_24776);
or U27114 (N_27114,N_25285,N_25929);
or U27115 (N_27115,N_24127,N_25812);
and U27116 (N_27116,N_25300,N_25977);
and U27117 (N_27117,N_25572,N_24967);
or U27118 (N_27118,N_25707,N_25120);
or U27119 (N_27119,N_24472,N_24415);
and U27120 (N_27120,N_24382,N_24545);
xor U27121 (N_27121,N_25901,N_24790);
nand U27122 (N_27122,N_25267,N_24968);
nor U27123 (N_27123,N_25863,N_24915);
nand U27124 (N_27124,N_24719,N_25864);
nor U27125 (N_27125,N_25969,N_25627);
or U27126 (N_27126,N_25345,N_25151);
nand U27127 (N_27127,N_25119,N_24000);
and U27128 (N_27128,N_25820,N_25405);
nor U27129 (N_27129,N_25162,N_24740);
and U27130 (N_27130,N_25935,N_25789);
nand U27131 (N_27131,N_25768,N_24431);
or U27132 (N_27132,N_24875,N_24124);
or U27133 (N_27133,N_24300,N_25987);
xnor U27134 (N_27134,N_24005,N_24936);
nand U27135 (N_27135,N_25914,N_24753);
or U27136 (N_27136,N_25193,N_24051);
nand U27137 (N_27137,N_25370,N_24181);
xnor U27138 (N_27138,N_24593,N_25248);
and U27139 (N_27139,N_25451,N_25814);
nor U27140 (N_27140,N_24260,N_24271);
and U27141 (N_27141,N_25460,N_25116);
nor U27142 (N_27142,N_24977,N_25244);
nor U27143 (N_27143,N_25638,N_24558);
or U27144 (N_27144,N_25593,N_24574);
and U27145 (N_27145,N_24535,N_25336);
or U27146 (N_27146,N_24328,N_24002);
nand U27147 (N_27147,N_25944,N_24129);
nor U27148 (N_27148,N_25736,N_24557);
nand U27149 (N_27149,N_25026,N_24801);
and U27150 (N_27150,N_24795,N_25819);
nand U27151 (N_27151,N_24230,N_24127);
or U27152 (N_27152,N_24690,N_25109);
xor U27153 (N_27153,N_24353,N_25141);
nor U27154 (N_27154,N_25655,N_25798);
nor U27155 (N_27155,N_24722,N_25697);
xnor U27156 (N_27156,N_24011,N_25767);
or U27157 (N_27157,N_24303,N_24975);
nand U27158 (N_27158,N_25664,N_25355);
xnor U27159 (N_27159,N_24445,N_25766);
and U27160 (N_27160,N_25407,N_25916);
or U27161 (N_27161,N_25623,N_25630);
or U27162 (N_27162,N_25020,N_25281);
or U27163 (N_27163,N_24066,N_24542);
nand U27164 (N_27164,N_24956,N_24978);
nor U27165 (N_27165,N_24629,N_24008);
xor U27166 (N_27166,N_25963,N_24535);
or U27167 (N_27167,N_25362,N_24490);
and U27168 (N_27168,N_24480,N_25947);
or U27169 (N_27169,N_25379,N_25594);
nand U27170 (N_27170,N_24355,N_25363);
nand U27171 (N_27171,N_24685,N_25055);
or U27172 (N_27172,N_25888,N_25104);
or U27173 (N_27173,N_25484,N_24214);
xnor U27174 (N_27174,N_25951,N_25131);
nand U27175 (N_27175,N_24797,N_25673);
nor U27176 (N_27176,N_25666,N_25195);
nand U27177 (N_27177,N_24457,N_24978);
nand U27178 (N_27178,N_24219,N_24700);
or U27179 (N_27179,N_24830,N_24547);
xor U27180 (N_27180,N_24507,N_24541);
nor U27181 (N_27181,N_25660,N_24557);
or U27182 (N_27182,N_25114,N_25418);
nor U27183 (N_27183,N_25623,N_24204);
or U27184 (N_27184,N_25481,N_25341);
or U27185 (N_27185,N_25749,N_25686);
and U27186 (N_27186,N_24934,N_24693);
xor U27187 (N_27187,N_25816,N_24841);
nand U27188 (N_27188,N_25056,N_25414);
xnor U27189 (N_27189,N_24841,N_24011);
or U27190 (N_27190,N_24239,N_24223);
nor U27191 (N_27191,N_24407,N_25852);
or U27192 (N_27192,N_24234,N_25654);
or U27193 (N_27193,N_24123,N_24878);
nor U27194 (N_27194,N_24128,N_24023);
nand U27195 (N_27195,N_24522,N_24695);
nor U27196 (N_27196,N_24642,N_24567);
and U27197 (N_27197,N_24092,N_24720);
nand U27198 (N_27198,N_24605,N_24846);
nor U27199 (N_27199,N_25713,N_25303);
nand U27200 (N_27200,N_25492,N_25242);
nor U27201 (N_27201,N_24618,N_25515);
and U27202 (N_27202,N_24867,N_24465);
or U27203 (N_27203,N_25099,N_25163);
xnor U27204 (N_27204,N_25411,N_25121);
nand U27205 (N_27205,N_25835,N_25359);
nor U27206 (N_27206,N_24746,N_24080);
and U27207 (N_27207,N_24025,N_24402);
or U27208 (N_27208,N_24435,N_25060);
xnor U27209 (N_27209,N_24052,N_25736);
xor U27210 (N_27210,N_25124,N_24802);
or U27211 (N_27211,N_24193,N_24427);
and U27212 (N_27212,N_25597,N_24039);
xor U27213 (N_27213,N_24808,N_24113);
xnor U27214 (N_27214,N_25404,N_25813);
nand U27215 (N_27215,N_24045,N_24605);
or U27216 (N_27216,N_24413,N_24942);
and U27217 (N_27217,N_25797,N_24979);
or U27218 (N_27218,N_25477,N_25216);
nor U27219 (N_27219,N_24469,N_25637);
nand U27220 (N_27220,N_25008,N_25396);
nand U27221 (N_27221,N_24838,N_24302);
and U27222 (N_27222,N_24208,N_24380);
or U27223 (N_27223,N_24249,N_25784);
and U27224 (N_27224,N_25108,N_24244);
nor U27225 (N_27225,N_25843,N_25332);
or U27226 (N_27226,N_25229,N_25308);
and U27227 (N_27227,N_25452,N_25577);
nor U27228 (N_27228,N_24926,N_25981);
nor U27229 (N_27229,N_25239,N_25135);
xor U27230 (N_27230,N_24503,N_25607);
xor U27231 (N_27231,N_24082,N_25282);
and U27232 (N_27232,N_25773,N_25915);
xnor U27233 (N_27233,N_25123,N_24729);
nor U27234 (N_27234,N_25790,N_25130);
or U27235 (N_27235,N_25302,N_25535);
nand U27236 (N_27236,N_25419,N_25110);
nand U27237 (N_27237,N_25945,N_25105);
and U27238 (N_27238,N_25660,N_24172);
or U27239 (N_27239,N_24529,N_24397);
or U27240 (N_27240,N_25197,N_24867);
or U27241 (N_27241,N_24565,N_24068);
or U27242 (N_27242,N_25476,N_24749);
xor U27243 (N_27243,N_24451,N_24134);
xnor U27244 (N_27244,N_25196,N_25351);
nor U27245 (N_27245,N_25122,N_24626);
nand U27246 (N_27246,N_24982,N_24758);
and U27247 (N_27247,N_24508,N_25911);
nor U27248 (N_27248,N_25194,N_25652);
or U27249 (N_27249,N_24976,N_24511);
nand U27250 (N_27250,N_24428,N_25776);
or U27251 (N_27251,N_25653,N_25000);
nand U27252 (N_27252,N_25659,N_25358);
nand U27253 (N_27253,N_24960,N_24267);
xnor U27254 (N_27254,N_24145,N_25547);
or U27255 (N_27255,N_24690,N_25987);
nand U27256 (N_27256,N_24488,N_25334);
and U27257 (N_27257,N_24119,N_25261);
or U27258 (N_27258,N_25769,N_25822);
xor U27259 (N_27259,N_24031,N_24420);
xor U27260 (N_27260,N_25882,N_24468);
or U27261 (N_27261,N_24754,N_25301);
xor U27262 (N_27262,N_25355,N_25580);
xnor U27263 (N_27263,N_25096,N_24039);
nand U27264 (N_27264,N_25426,N_25660);
nor U27265 (N_27265,N_25607,N_24605);
nor U27266 (N_27266,N_24334,N_24281);
or U27267 (N_27267,N_25593,N_24770);
nor U27268 (N_27268,N_25048,N_24862);
or U27269 (N_27269,N_24679,N_25406);
or U27270 (N_27270,N_25991,N_24180);
nor U27271 (N_27271,N_25826,N_24299);
or U27272 (N_27272,N_24872,N_24838);
xor U27273 (N_27273,N_24496,N_25723);
and U27274 (N_27274,N_25631,N_25198);
and U27275 (N_27275,N_25435,N_25429);
or U27276 (N_27276,N_24685,N_24731);
or U27277 (N_27277,N_25568,N_25411);
nand U27278 (N_27278,N_25332,N_24344);
nand U27279 (N_27279,N_25314,N_25824);
and U27280 (N_27280,N_24552,N_24857);
or U27281 (N_27281,N_25928,N_25701);
nor U27282 (N_27282,N_24848,N_25712);
xnor U27283 (N_27283,N_24978,N_25536);
or U27284 (N_27284,N_24543,N_24742);
or U27285 (N_27285,N_25654,N_25709);
xor U27286 (N_27286,N_24309,N_24052);
xnor U27287 (N_27287,N_25678,N_25099);
and U27288 (N_27288,N_24104,N_24911);
and U27289 (N_27289,N_25176,N_25962);
or U27290 (N_27290,N_25546,N_24775);
xor U27291 (N_27291,N_25604,N_25340);
and U27292 (N_27292,N_24405,N_24700);
nand U27293 (N_27293,N_24580,N_25239);
xnor U27294 (N_27294,N_24331,N_25658);
and U27295 (N_27295,N_24033,N_25806);
xor U27296 (N_27296,N_25165,N_25776);
or U27297 (N_27297,N_24581,N_25412);
nand U27298 (N_27298,N_25097,N_25932);
nand U27299 (N_27299,N_25384,N_24271);
or U27300 (N_27300,N_25123,N_25883);
nor U27301 (N_27301,N_25042,N_24536);
nor U27302 (N_27302,N_25484,N_25097);
or U27303 (N_27303,N_25210,N_24121);
nand U27304 (N_27304,N_25963,N_25246);
xnor U27305 (N_27305,N_25202,N_25737);
or U27306 (N_27306,N_25123,N_25410);
and U27307 (N_27307,N_25867,N_24860);
xnor U27308 (N_27308,N_25625,N_24579);
and U27309 (N_27309,N_25282,N_24662);
nor U27310 (N_27310,N_24763,N_25764);
nand U27311 (N_27311,N_24377,N_24500);
nand U27312 (N_27312,N_25022,N_25672);
and U27313 (N_27313,N_25292,N_25549);
xnor U27314 (N_27314,N_25008,N_25945);
and U27315 (N_27315,N_25181,N_24457);
and U27316 (N_27316,N_25855,N_25568);
nand U27317 (N_27317,N_24163,N_24097);
nor U27318 (N_27318,N_25893,N_25200);
xnor U27319 (N_27319,N_24838,N_24842);
xor U27320 (N_27320,N_25212,N_24288);
xor U27321 (N_27321,N_24794,N_25794);
nand U27322 (N_27322,N_25013,N_25800);
or U27323 (N_27323,N_25707,N_25855);
and U27324 (N_27324,N_25097,N_25510);
xnor U27325 (N_27325,N_25482,N_25832);
or U27326 (N_27326,N_25763,N_25531);
xnor U27327 (N_27327,N_24523,N_24795);
nand U27328 (N_27328,N_24950,N_24772);
and U27329 (N_27329,N_25241,N_24901);
nor U27330 (N_27330,N_25093,N_25476);
xnor U27331 (N_27331,N_24040,N_24853);
nand U27332 (N_27332,N_25262,N_25960);
xnor U27333 (N_27333,N_25046,N_24672);
nand U27334 (N_27334,N_24797,N_25501);
or U27335 (N_27335,N_25039,N_24087);
nand U27336 (N_27336,N_25830,N_25214);
or U27337 (N_27337,N_24272,N_25956);
nand U27338 (N_27338,N_24790,N_25565);
xnor U27339 (N_27339,N_25611,N_24566);
and U27340 (N_27340,N_25267,N_25176);
or U27341 (N_27341,N_25621,N_24324);
nor U27342 (N_27342,N_25499,N_25506);
or U27343 (N_27343,N_25901,N_24127);
nor U27344 (N_27344,N_24462,N_25039);
or U27345 (N_27345,N_24922,N_24810);
xor U27346 (N_27346,N_25913,N_25964);
nand U27347 (N_27347,N_24850,N_25576);
or U27348 (N_27348,N_25796,N_25542);
nor U27349 (N_27349,N_24521,N_24576);
xnor U27350 (N_27350,N_24593,N_25690);
nand U27351 (N_27351,N_25486,N_24065);
or U27352 (N_27352,N_24212,N_24397);
nand U27353 (N_27353,N_25478,N_25087);
nor U27354 (N_27354,N_25792,N_25576);
nor U27355 (N_27355,N_24031,N_24813);
nor U27356 (N_27356,N_25551,N_24801);
nor U27357 (N_27357,N_25220,N_24540);
and U27358 (N_27358,N_25141,N_24876);
or U27359 (N_27359,N_25332,N_25433);
nand U27360 (N_27360,N_25268,N_25896);
and U27361 (N_27361,N_24264,N_24696);
nor U27362 (N_27362,N_24881,N_25403);
nand U27363 (N_27363,N_24073,N_24315);
or U27364 (N_27364,N_25173,N_25748);
xnor U27365 (N_27365,N_24217,N_24303);
xor U27366 (N_27366,N_24208,N_24849);
nand U27367 (N_27367,N_24804,N_25667);
and U27368 (N_27368,N_24521,N_24471);
or U27369 (N_27369,N_25359,N_25875);
nor U27370 (N_27370,N_24882,N_24763);
xor U27371 (N_27371,N_25091,N_25396);
xor U27372 (N_27372,N_25307,N_25287);
or U27373 (N_27373,N_24994,N_25415);
nand U27374 (N_27374,N_25925,N_25492);
xor U27375 (N_27375,N_25392,N_24787);
xor U27376 (N_27376,N_24230,N_25469);
xnor U27377 (N_27377,N_24679,N_25557);
nor U27378 (N_27378,N_24568,N_24913);
and U27379 (N_27379,N_24438,N_25801);
nand U27380 (N_27380,N_24558,N_25060);
nor U27381 (N_27381,N_24917,N_24905);
and U27382 (N_27382,N_25576,N_24769);
nor U27383 (N_27383,N_24393,N_25350);
or U27384 (N_27384,N_24859,N_24134);
and U27385 (N_27385,N_25164,N_25848);
and U27386 (N_27386,N_24919,N_24340);
nand U27387 (N_27387,N_24420,N_25539);
xnor U27388 (N_27388,N_24172,N_24292);
or U27389 (N_27389,N_25885,N_25240);
xnor U27390 (N_27390,N_24255,N_24282);
nand U27391 (N_27391,N_25193,N_24235);
nand U27392 (N_27392,N_24864,N_25263);
and U27393 (N_27393,N_25190,N_24112);
or U27394 (N_27394,N_25450,N_24300);
and U27395 (N_27395,N_25877,N_24603);
or U27396 (N_27396,N_25136,N_24099);
nand U27397 (N_27397,N_25968,N_25293);
nand U27398 (N_27398,N_24893,N_24016);
or U27399 (N_27399,N_24884,N_25287);
nor U27400 (N_27400,N_24610,N_24500);
or U27401 (N_27401,N_24900,N_24548);
or U27402 (N_27402,N_24507,N_25733);
nor U27403 (N_27403,N_24524,N_25083);
nor U27404 (N_27404,N_24603,N_25163);
or U27405 (N_27405,N_25359,N_25482);
nor U27406 (N_27406,N_24069,N_25170);
or U27407 (N_27407,N_25182,N_25927);
nor U27408 (N_27408,N_25537,N_24905);
xor U27409 (N_27409,N_25888,N_24613);
xor U27410 (N_27410,N_25011,N_24884);
and U27411 (N_27411,N_25354,N_25432);
or U27412 (N_27412,N_24620,N_24896);
or U27413 (N_27413,N_25998,N_24204);
and U27414 (N_27414,N_24819,N_24665);
nor U27415 (N_27415,N_25202,N_24891);
nor U27416 (N_27416,N_25918,N_25114);
nand U27417 (N_27417,N_24980,N_24618);
or U27418 (N_27418,N_25722,N_25031);
nor U27419 (N_27419,N_24908,N_25690);
and U27420 (N_27420,N_24148,N_24312);
nand U27421 (N_27421,N_24217,N_25656);
nor U27422 (N_27422,N_24213,N_24374);
and U27423 (N_27423,N_25835,N_24600);
xnor U27424 (N_27424,N_24259,N_24401);
and U27425 (N_27425,N_25800,N_24429);
or U27426 (N_27426,N_24195,N_25153);
and U27427 (N_27427,N_25057,N_24245);
or U27428 (N_27428,N_25506,N_24190);
nand U27429 (N_27429,N_25082,N_25959);
nand U27430 (N_27430,N_24884,N_25006);
and U27431 (N_27431,N_25495,N_24256);
nor U27432 (N_27432,N_24216,N_25237);
nand U27433 (N_27433,N_24604,N_25336);
or U27434 (N_27434,N_24618,N_24379);
or U27435 (N_27435,N_25008,N_24885);
or U27436 (N_27436,N_24984,N_24214);
nand U27437 (N_27437,N_24108,N_25911);
xnor U27438 (N_27438,N_24564,N_24028);
nor U27439 (N_27439,N_24254,N_24293);
or U27440 (N_27440,N_25378,N_25501);
xnor U27441 (N_27441,N_24826,N_24966);
xnor U27442 (N_27442,N_25079,N_24000);
nor U27443 (N_27443,N_24127,N_24248);
and U27444 (N_27444,N_24869,N_25216);
xor U27445 (N_27445,N_25267,N_24859);
and U27446 (N_27446,N_24409,N_25965);
and U27447 (N_27447,N_25626,N_24790);
and U27448 (N_27448,N_24420,N_25615);
nand U27449 (N_27449,N_25261,N_24729);
or U27450 (N_27450,N_25097,N_25685);
xor U27451 (N_27451,N_24091,N_24666);
xnor U27452 (N_27452,N_24845,N_25627);
xor U27453 (N_27453,N_25773,N_24737);
nor U27454 (N_27454,N_25929,N_25825);
or U27455 (N_27455,N_25536,N_25317);
or U27456 (N_27456,N_24397,N_25375);
and U27457 (N_27457,N_25047,N_25752);
xnor U27458 (N_27458,N_24174,N_24013);
or U27459 (N_27459,N_24741,N_24206);
or U27460 (N_27460,N_24748,N_24214);
xor U27461 (N_27461,N_24670,N_24828);
or U27462 (N_27462,N_25204,N_25228);
nor U27463 (N_27463,N_25914,N_25503);
nand U27464 (N_27464,N_25494,N_25956);
nand U27465 (N_27465,N_24115,N_24018);
nand U27466 (N_27466,N_24197,N_24971);
or U27467 (N_27467,N_25370,N_24814);
nand U27468 (N_27468,N_25824,N_24738);
nand U27469 (N_27469,N_25477,N_24725);
nor U27470 (N_27470,N_25719,N_25986);
nand U27471 (N_27471,N_24574,N_24562);
and U27472 (N_27472,N_25878,N_24992);
xor U27473 (N_27473,N_24467,N_25264);
nand U27474 (N_27474,N_25363,N_24625);
xor U27475 (N_27475,N_25431,N_25242);
xnor U27476 (N_27476,N_25810,N_25464);
nand U27477 (N_27477,N_24551,N_24035);
nand U27478 (N_27478,N_25345,N_24531);
nor U27479 (N_27479,N_24835,N_25533);
or U27480 (N_27480,N_25660,N_24696);
xnor U27481 (N_27481,N_24342,N_24359);
or U27482 (N_27482,N_24840,N_25168);
and U27483 (N_27483,N_25113,N_25594);
nand U27484 (N_27484,N_25428,N_25970);
xor U27485 (N_27485,N_24006,N_24557);
and U27486 (N_27486,N_24397,N_25262);
nand U27487 (N_27487,N_24462,N_25686);
nor U27488 (N_27488,N_25198,N_25589);
or U27489 (N_27489,N_24079,N_24395);
nand U27490 (N_27490,N_24575,N_25997);
xnor U27491 (N_27491,N_25962,N_24098);
or U27492 (N_27492,N_24585,N_25732);
xnor U27493 (N_27493,N_25136,N_25749);
nor U27494 (N_27494,N_24425,N_24090);
xnor U27495 (N_27495,N_24646,N_24063);
or U27496 (N_27496,N_24630,N_25899);
or U27497 (N_27497,N_24573,N_24830);
xor U27498 (N_27498,N_24920,N_24950);
or U27499 (N_27499,N_25660,N_24946);
nand U27500 (N_27500,N_25222,N_25849);
nor U27501 (N_27501,N_25271,N_24890);
nor U27502 (N_27502,N_25070,N_24029);
nand U27503 (N_27503,N_25295,N_25822);
xor U27504 (N_27504,N_24543,N_24005);
xnor U27505 (N_27505,N_24524,N_24734);
nand U27506 (N_27506,N_25786,N_24603);
nor U27507 (N_27507,N_25664,N_24244);
and U27508 (N_27508,N_24923,N_24538);
or U27509 (N_27509,N_24869,N_25192);
nor U27510 (N_27510,N_25992,N_25900);
or U27511 (N_27511,N_25618,N_25441);
nor U27512 (N_27512,N_25731,N_24793);
nor U27513 (N_27513,N_24042,N_25497);
xor U27514 (N_27514,N_25901,N_24427);
nor U27515 (N_27515,N_25624,N_24880);
and U27516 (N_27516,N_24388,N_24389);
xor U27517 (N_27517,N_24791,N_25135);
or U27518 (N_27518,N_24226,N_24336);
nand U27519 (N_27519,N_25144,N_24595);
or U27520 (N_27520,N_25104,N_24509);
xnor U27521 (N_27521,N_25191,N_25740);
and U27522 (N_27522,N_24884,N_24717);
xor U27523 (N_27523,N_25673,N_25612);
and U27524 (N_27524,N_24805,N_24963);
and U27525 (N_27525,N_24363,N_25321);
or U27526 (N_27526,N_25771,N_25147);
xnor U27527 (N_27527,N_24434,N_25993);
nand U27528 (N_27528,N_25154,N_24096);
nand U27529 (N_27529,N_25645,N_24668);
or U27530 (N_27530,N_25827,N_25910);
and U27531 (N_27531,N_24673,N_24981);
nand U27532 (N_27532,N_25685,N_25585);
xnor U27533 (N_27533,N_25266,N_25654);
nor U27534 (N_27534,N_24993,N_25901);
nor U27535 (N_27535,N_25739,N_25163);
or U27536 (N_27536,N_25798,N_24865);
xor U27537 (N_27537,N_25075,N_24447);
and U27538 (N_27538,N_24144,N_25534);
or U27539 (N_27539,N_25344,N_25867);
nand U27540 (N_27540,N_24107,N_24396);
xnor U27541 (N_27541,N_25821,N_25884);
or U27542 (N_27542,N_24860,N_25093);
nor U27543 (N_27543,N_24394,N_24300);
or U27544 (N_27544,N_24175,N_24934);
xnor U27545 (N_27545,N_25903,N_24719);
or U27546 (N_27546,N_25684,N_25840);
xnor U27547 (N_27547,N_24916,N_24671);
nor U27548 (N_27548,N_24412,N_24118);
nand U27549 (N_27549,N_24801,N_25919);
nor U27550 (N_27550,N_25262,N_25591);
nor U27551 (N_27551,N_24612,N_24447);
nor U27552 (N_27552,N_24751,N_24357);
xor U27553 (N_27553,N_24611,N_24643);
and U27554 (N_27554,N_25918,N_24303);
nor U27555 (N_27555,N_24947,N_25474);
nand U27556 (N_27556,N_25288,N_25684);
nor U27557 (N_27557,N_24264,N_25076);
nor U27558 (N_27558,N_24941,N_24585);
nor U27559 (N_27559,N_25716,N_24025);
nand U27560 (N_27560,N_24317,N_24086);
nor U27561 (N_27561,N_24398,N_24519);
nor U27562 (N_27562,N_24764,N_24858);
xnor U27563 (N_27563,N_25945,N_24225);
nand U27564 (N_27564,N_24841,N_25443);
or U27565 (N_27565,N_24653,N_24305);
xor U27566 (N_27566,N_25932,N_24317);
nor U27567 (N_27567,N_25978,N_24809);
nand U27568 (N_27568,N_25482,N_24933);
nand U27569 (N_27569,N_24352,N_25141);
xor U27570 (N_27570,N_25199,N_24263);
nor U27571 (N_27571,N_25082,N_25784);
or U27572 (N_27572,N_25774,N_24301);
or U27573 (N_27573,N_24093,N_24510);
nand U27574 (N_27574,N_24198,N_24518);
or U27575 (N_27575,N_25324,N_24585);
and U27576 (N_27576,N_24953,N_25624);
or U27577 (N_27577,N_25766,N_24389);
and U27578 (N_27578,N_24129,N_24534);
xor U27579 (N_27579,N_25620,N_25195);
xor U27580 (N_27580,N_25496,N_24437);
nor U27581 (N_27581,N_24794,N_24121);
and U27582 (N_27582,N_24440,N_25152);
and U27583 (N_27583,N_25234,N_25597);
or U27584 (N_27584,N_25204,N_24760);
nand U27585 (N_27585,N_24871,N_24547);
or U27586 (N_27586,N_25179,N_25392);
or U27587 (N_27587,N_25568,N_24877);
or U27588 (N_27588,N_24636,N_24787);
or U27589 (N_27589,N_25927,N_25251);
nand U27590 (N_27590,N_25994,N_25392);
nor U27591 (N_27591,N_24029,N_24360);
xnor U27592 (N_27592,N_25372,N_24194);
xor U27593 (N_27593,N_24576,N_25659);
nand U27594 (N_27594,N_25240,N_25841);
and U27595 (N_27595,N_24421,N_24368);
xor U27596 (N_27596,N_25635,N_24690);
or U27597 (N_27597,N_24063,N_25012);
and U27598 (N_27598,N_24114,N_24434);
and U27599 (N_27599,N_25940,N_24567);
and U27600 (N_27600,N_25055,N_25791);
xor U27601 (N_27601,N_25662,N_25018);
nor U27602 (N_27602,N_24546,N_25933);
and U27603 (N_27603,N_24618,N_25155);
nand U27604 (N_27604,N_25834,N_25040);
and U27605 (N_27605,N_25198,N_24395);
or U27606 (N_27606,N_25817,N_25621);
xor U27607 (N_27607,N_24818,N_24873);
nor U27608 (N_27608,N_24012,N_24801);
xor U27609 (N_27609,N_24033,N_25884);
nand U27610 (N_27610,N_25736,N_25210);
or U27611 (N_27611,N_25089,N_25736);
or U27612 (N_27612,N_25520,N_25230);
or U27613 (N_27613,N_24116,N_25269);
nor U27614 (N_27614,N_24791,N_24071);
nand U27615 (N_27615,N_24987,N_24386);
and U27616 (N_27616,N_25812,N_25698);
nor U27617 (N_27617,N_24980,N_24882);
and U27618 (N_27618,N_25968,N_25860);
nor U27619 (N_27619,N_25948,N_24823);
nor U27620 (N_27620,N_24540,N_25660);
nand U27621 (N_27621,N_25321,N_25093);
or U27622 (N_27622,N_24382,N_24483);
nor U27623 (N_27623,N_25595,N_25927);
and U27624 (N_27624,N_25717,N_24958);
nand U27625 (N_27625,N_24032,N_25334);
xor U27626 (N_27626,N_25140,N_24390);
xor U27627 (N_27627,N_24240,N_25814);
nor U27628 (N_27628,N_24793,N_25845);
and U27629 (N_27629,N_25843,N_25819);
nand U27630 (N_27630,N_25165,N_24476);
or U27631 (N_27631,N_24516,N_25276);
nand U27632 (N_27632,N_24613,N_25084);
or U27633 (N_27633,N_24548,N_25931);
xor U27634 (N_27634,N_24264,N_25441);
or U27635 (N_27635,N_24077,N_24039);
and U27636 (N_27636,N_24383,N_25686);
nor U27637 (N_27637,N_24949,N_24720);
xnor U27638 (N_27638,N_25269,N_25280);
nand U27639 (N_27639,N_24987,N_25458);
xnor U27640 (N_27640,N_24986,N_24806);
and U27641 (N_27641,N_24844,N_24757);
nor U27642 (N_27642,N_24532,N_24937);
nor U27643 (N_27643,N_24205,N_25399);
nand U27644 (N_27644,N_25017,N_24422);
or U27645 (N_27645,N_25093,N_24220);
xor U27646 (N_27646,N_24454,N_25902);
nor U27647 (N_27647,N_24761,N_24808);
or U27648 (N_27648,N_25235,N_24426);
xor U27649 (N_27649,N_25044,N_25472);
xor U27650 (N_27650,N_25094,N_25357);
and U27651 (N_27651,N_24122,N_24729);
nor U27652 (N_27652,N_24619,N_25166);
or U27653 (N_27653,N_25816,N_25095);
nor U27654 (N_27654,N_24395,N_24432);
nand U27655 (N_27655,N_24490,N_25328);
nand U27656 (N_27656,N_25024,N_25455);
or U27657 (N_27657,N_24137,N_24000);
and U27658 (N_27658,N_25207,N_24502);
nand U27659 (N_27659,N_25233,N_25160);
and U27660 (N_27660,N_24253,N_24430);
nor U27661 (N_27661,N_25215,N_24407);
xor U27662 (N_27662,N_24465,N_24594);
or U27663 (N_27663,N_25811,N_24341);
nor U27664 (N_27664,N_24255,N_24552);
nor U27665 (N_27665,N_25937,N_25323);
nand U27666 (N_27666,N_25766,N_24334);
nor U27667 (N_27667,N_24454,N_24304);
xor U27668 (N_27668,N_24412,N_25398);
and U27669 (N_27669,N_25688,N_25934);
and U27670 (N_27670,N_24239,N_25888);
xor U27671 (N_27671,N_24765,N_24976);
nor U27672 (N_27672,N_24474,N_25789);
nor U27673 (N_27673,N_24042,N_25215);
and U27674 (N_27674,N_24102,N_25935);
xnor U27675 (N_27675,N_25718,N_25341);
or U27676 (N_27676,N_24063,N_24566);
and U27677 (N_27677,N_25617,N_25209);
or U27678 (N_27678,N_25532,N_25020);
nand U27679 (N_27679,N_25879,N_24571);
xnor U27680 (N_27680,N_25256,N_25223);
or U27681 (N_27681,N_24139,N_25657);
nand U27682 (N_27682,N_25313,N_25718);
nor U27683 (N_27683,N_24503,N_25099);
xor U27684 (N_27684,N_25312,N_25805);
nand U27685 (N_27685,N_24288,N_24072);
nor U27686 (N_27686,N_25523,N_25559);
nand U27687 (N_27687,N_25061,N_24456);
xor U27688 (N_27688,N_25112,N_25631);
nor U27689 (N_27689,N_25848,N_25551);
and U27690 (N_27690,N_24849,N_24914);
xnor U27691 (N_27691,N_25736,N_25235);
nand U27692 (N_27692,N_24467,N_25995);
nand U27693 (N_27693,N_25754,N_24129);
nand U27694 (N_27694,N_25326,N_25340);
or U27695 (N_27695,N_24247,N_24610);
nand U27696 (N_27696,N_24123,N_24792);
nand U27697 (N_27697,N_24845,N_25400);
and U27698 (N_27698,N_24120,N_24023);
xor U27699 (N_27699,N_24174,N_25817);
and U27700 (N_27700,N_25978,N_24023);
or U27701 (N_27701,N_24156,N_24923);
nor U27702 (N_27702,N_24296,N_24698);
nor U27703 (N_27703,N_25944,N_25521);
and U27704 (N_27704,N_25563,N_24102);
and U27705 (N_27705,N_25433,N_25659);
nor U27706 (N_27706,N_25675,N_24811);
xor U27707 (N_27707,N_24598,N_24588);
nand U27708 (N_27708,N_25499,N_24328);
and U27709 (N_27709,N_24816,N_24966);
or U27710 (N_27710,N_25960,N_24071);
nor U27711 (N_27711,N_25341,N_25589);
xor U27712 (N_27712,N_24386,N_25346);
or U27713 (N_27713,N_25953,N_24026);
or U27714 (N_27714,N_24313,N_24520);
xnor U27715 (N_27715,N_24340,N_24729);
or U27716 (N_27716,N_24036,N_25115);
and U27717 (N_27717,N_25713,N_25530);
or U27718 (N_27718,N_24396,N_24865);
nand U27719 (N_27719,N_24020,N_24507);
or U27720 (N_27720,N_25352,N_24583);
or U27721 (N_27721,N_25679,N_25952);
xor U27722 (N_27722,N_24109,N_25630);
xor U27723 (N_27723,N_24139,N_24023);
or U27724 (N_27724,N_24790,N_25687);
or U27725 (N_27725,N_25391,N_25093);
nand U27726 (N_27726,N_24524,N_24010);
xor U27727 (N_27727,N_24848,N_25337);
or U27728 (N_27728,N_24936,N_25135);
xnor U27729 (N_27729,N_25737,N_25361);
or U27730 (N_27730,N_25014,N_25990);
or U27731 (N_27731,N_24374,N_24732);
nor U27732 (N_27732,N_25849,N_24866);
xor U27733 (N_27733,N_24192,N_25249);
xnor U27734 (N_27734,N_24763,N_24620);
or U27735 (N_27735,N_24301,N_24319);
xnor U27736 (N_27736,N_24221,N_25650);
nor U27737 (N_27737,N_24151,N_24427);
xor U27738 (N_27738,N_25770,N_25135);
nand U27739 (N_27739,N_24002,N_25221);
or U27740 (N_27740,N_25540,N_24235);
nor U27741 (N_27741,N_24623,N_25993);
nor U27742 (N_27742,N_25255,N_25318);
nor U27743 (N_27743,N_25744,N_24695);
nand U27744 (N_27744,N_24301,N_24450);
nor U27745 (N_27745,N_24129,N_24464);
nor U27746 (N_27746,N_25241,N_24482);
and U27747 (N_27747,N_24644,N_25260);
and U27748 (N_27748,N_25018,N_24854);
xnor U27749 (N_27749,N_24438,N_24710);
or U27750 (N_27750,N_25328,N_25776);
or U27751 (N_27751,N_24969,N_25979);
xnor U27752 (N_27752,N_25451,N_24558);
or U27753 (N_27753,N_24892,N_25368);
nand U27754 (N_27754,N_25219,N_24777);
or U27755 (N_27755,N_24472,N_25273);
nor U27756 (N_27756,N_24690,N_24958);
or U27757 (N_27757,N_25304,N_25171);
nor U27758 (N_27758,N_25714,N_24849);
nand U27759 (N_27759,N_24018,N_25834);
xnor U27760 (N_27760,N_25569,N_25844);
nor U27761 (N_27761,N_25074,N_24616);
or U27762 (N_27762,N_25207,N_25992);
xor U27763 (N_27763,N_25395,N_24413);
and U27764 (N_27764,N_24248,N_25866);
and U27765 (N_27765,N_25739,N_25945);
and U27766 (N_27766,N_24646,N_24205);
and U27767 (N_27767,N_25892,N_25614);
nor U27768 (N_27768,N_25242,N_25410);
nand U27769 (N_27769,N_25588,N_25090);
nand U27770 (N_27770,N_24226,N_25634);
or U27771 (N_27771,N_25353,N_25065);
or U27772 (N_27772,N_25179,N_25295);
nor U27773 (N_27773,N_24300,N_24571);
or U27774 (N_27774,N_25562,N_25190);
nand U27775 (N_27775,N_24180,N_25605);
and U27776 (N_27776,N_24571,N_25361);
nor U27777 (N_27777,N_25753,N_25265);
nor U27778 (N_27778,N_25454,N_24597);
or U27779 (N_27779,N_25787,N_24792);
xor U27780 (N_27780,N_25150,N_24509);
and U27781 (N_27781,N_24298,N_24923);
xnor U27782 (N_27782,N_25489,N_25773);
nor U27783 (N_27783,N_24298,N_24170);
and U27784 (N_27784,N_25998,N_25561);
nor U27785 (N_27785,N_24873,N_24773);
nand U27786 (N_27786,N_24517,N_24525);
and U27787 (N_27787,N_25807,N_25464);
nand U27788 (N_27788,N_25230,N_25174);
or U27789 (N_27789,N_24564,N_25962);
nand U27790 (N_27790,N_25806,N_24289);
nand U27791 (N_27791,N_25234,N_25358);
xnor U27792 (N_27792,N_25310,N_24937);
nor U27793 (N_27793,N_24698,N_25880);
or U27794 (N_27794,N_25932,N_24684);
nand U27795 (N_27795,N_25121,N_24317);
and U27796 (N_27796,N_24462,N_24353);
or U27797 (N_27797,N_25902,N_24150);
nor U27798 (N_27798,N_25876,N_25211);
nor U27799 (N_27799,N_25319,N_24947);
nor U27800 (N_27800,N_24725,N_25087);
xnor U27801 (N_27801,N_25891,N_25253);
nand U27802 (N_27802,N_25134,N_25474);
or U27803 (N_27803,N_25894,N_24947);
nor U27804 (N_27804,N_25203,N_25164);
xnor U27805 (N_27805,N_25992,N_25212);
nand U27806 (N_27806,N_25918,N_24060);
or U27807 (N_27807,N_25599,N_25422);
nand U27808 (N_27808,N_25160,N_24659);
xnor U27809 (N_27809,N_24602,N_24632);
nand U27810 (N_27810,N_25194,N_24352);
and U27811 (N_27811,N_24014,N_25614);
and U27812 (N_27812,N_25365,N_24960);
or U27813 (N_27813,N_25086,N_25816);
xnor U27814 (N_27814,N_24464,N_25658);
xnor U27815 (N_27815,N_25649,N_25836);
and U27816 (N_27816,N_24612,N_25944);
nand U27817 (N_27817,N_25748,N_25095);
xnor U27818 (N_27818,N_25439,N_25900);
or U27819 (N_27819,N_25365,N_24998);
or U27820 (N_27820,N_25587,N_25139);
xnor U27821 (N_27821,N_24364,N_25710);
nand U27822 (N_27822,N_24290,N_24649);
xor U27823 (N_27823,N_24101,N_24478);
xor U27824 (N_27824,N_24854,N_25597);
or U27825 (N_27825,N_24804,N_25608);
or U27826 (N_27826,N_24261,N_24716);
and U27827 (N_27827,N_24379,N_25573);
or U27828 (N_27828,N_24552,N_24314);
or U27829 (N_27829,N_25005,N_24638);
nor U27830 (N_27830,N_24701,N_24305);
nand U27831 (N_27831,N_25731,N_25419);
xor U27832 (N_27832,N_24931,N_24492);
nor U27833 (N_27833,N_24313,N_25928);
and U27834 (N_27834,N_24546,N_25366);
and U27835 (N_27835,N_25211,N_25238);
and U27836 (N_27836,N_24693,N_24118);
xnor U27837 (N_27837,N_25466,N_25392);
nand U27838 (N_27838,N_24214,N_24150);
xor U27839 (N_27839,N_25461,N_25099);
nor U27840 (N_27840,N_24730,N_25687);
and U27841 (N_27841,N_25264,N_25663);
or U27842 (N_27842,N_24486,N_24186);
or U27843 (N_27843,N_24229,N_25422);
nand U27844 (N_27844,N_24085,N_25842);
nor U27845 (N_27845,N_25059,N_25184);
nor U27846 (N_27846,N_24482,N_24001);
or U27847 (N_27847,N_25467,N_25115);
xor U27848 (N_27848,N_24739,N_24735);
and U27849 (N_27849,N_25301,N_24111);
xor U27850 (N_27850,N_24956,N_24215);
and U27851 (N_27851,N_24750,N_24705);
and U27852 (N_27852,N_25592,N_25036);
and U27853 (N_27853,N_25083,N_24532);
nor U27854 (N_27854,N_25050,N_25674);
and U27855 (N_27855,N_24480,N_25495);
and U27856 (N_27856,N_24753,N_25539);
nand U27857 (N_27857,N_25692,N_24254);
nor U27858 (N_27858,N_25152,N_24411);
and U27859 (N_27859,N_24197,N_24718);
xor U27860 (N_27860,N_25605,N_25892);
nand U27861 (N_27861,N_24497,N_24914);
and U27862 (N_27862,N_25742,N_25540);
nand U27863 (N_27863,N_25174,N_24363);
and U27864 (N_27864,N_24602,N_25086);
nor U27865 (N_27865,N_25947,N_24490);
nor U27866 (N_27866,N_24938,N_24600);
nand U27867 (N_27867,N_25740,N_25502);
xnor U27868 (N_27868,N_24275,N_24072);
xnor U27869 (N_27869,N_25862,N_24041);
nand U27870 (N_27870,N_25279,N_24175);
nor U27871 (N_27871,N_24010,N_24992);
and U27872 (N_27872,N_24276,N_25307);
or U27873 (N_27873,N_24420,N_24239);
xnor U27874 (N_27874,N_24904,N_25404);
nand U27875 (N_27875,N_25390,N_24256);
nand U27876 (N_27876,N_25027,N_25549);
nand U27877 (N_27877,N_24503,N_25037);
xnor U27878 (N_27878,N_24269,N_25727);
and U27879 (N_27879,N_25828,N_25137);
xnor U27880 (N_27880,N_25237,N_24829);
or U27881 (N_27881,N_25074,N_25024);
nor U27882 (N_27882,N_25837,N_25414);
or U27883 (N_27883,N_25741,N_25753);
nand U27884 (N_27884,N_25646,N_25471);
or U27885 (N_27885,N_24658,N_24836);
or U27886 (N_27886,N_25688,N_25917);
nor U27887 (N_27887,N_24112,N_25303);
nand U27888 (N_27888,N_24892,N_25143);
nor U27889 (N_27889,N_25020,N_24923);
nor U27890 (N_27890,N_25341,N_25566);
xnor U27891 (N_27891,N_25765,N_24761);
xnor U27892 (N_27892,N_24035,N_24829);
or U27893 (N_27893,N_24499,N_25515);
xnor U27894 (N_27894,N_25045,N_25721);
and U27895 (N_27895,N_24118,N_24734);
xor U27896 (N_27896,N_25131,N_25463);
and U27897 (N_27897,N_25285,N_24682);
xor U27898 (N_27898,N_24004,N_24898);
nand U27899 (N_27899,N_24238,N_24615);
xnor U27900 (N_27900,N_25483,N_24600);
xnor U27901 (N_27901,N_24357,N_25700);
xor U27902 (N_27902,N_24181,N_24604);
nor U27903 (N_27903,N_25963,N_24294);
nand U27904 (N_27904,N_25719,N_24212);
or U27905 (N_27905,N_24303,N_24706);
or U27906 (N_27906,N_24319,N_25372);
and U27907 (N_27907,N_24443,N_25308);
nor U27908 (N_27908,N_25447,N_24061);
nor U27909 (N_27909,N_24079,N_24741);
and U27910 (N_27910,N_25229,N_24132);
nand U27911 (N_27911,N_24140,N_24936);
xnor U27912 (N_27912,N_24647,N_25292);
nor U27913 (N_27913,N_24435,N_24939);
nor U27914 (N_27914,N_25221,N_24658);
nand U27915 (N_27915,N_24334,N_25970);
or U27916 (N_27916,N_24853,N_24253);
and U27917 (N_27917,N_25255,N_24506);
xnor U27918 (N_27918,N_24047,N_25068);
nand U27919 (N_27919,N_24460,N_24383);
xnor U27920 (N_27920,N_24806,N_24892);
and U27921 (N_27921,N_25565,N_24891);
and U27922 (N_27922,N_24195,N_25559);
nand U27923 (N_27923,N_24165,N_24646);
xnor U27924 (N_27924,N_24593,N_24021);
nand U27925 (N_27925,N_24979,N_25717);
nand U27926 (N_27926,N_25326,N_25632);
nand U27927 (N_27927,N_24900,N_25941);
nand U27928 (N_27928,N_25128,N_25395);
nand U27929 (N_27929,N_24822,N_24488);
nor U27930 (N_27930,N_24577,N_25184);
nand U27931 (N_27931,N_24548,N_24065);
nand U27932 (N_27932,N_25639,N_24686);
and U27933 (N_27933,N_25732,N_24364);
nor U27934 (N_27934,N_25142,N_24641);
and U27935 (N_27935,N_25610,N_24732);
or U27936 (N_27936,N_24399,N_25030);
and U27937 (N_27937,N_24999,N_24620);
and U27938 (N_27938,N_24481,N_24744);
xor U27939 (N_27939,N_25727,N_25328);
and U27940 (N_27940,N_24075,N_25392);
nor U27941 (N_27941,N_24998,N_25005);
or U27942 (N_27942,N_25936,N_25678);
and U27943 (N_27943,N_25320,N_24909);
and U27944 (N_27944,N_25027,N_24256);
or U27945 (N_27945,N_24417,N_25114);
xor U27946 (N_27946,N_24324,N_24838);
nor U27947 (N_27947,N_24118,N_25393);
nor U27948 (N_27948,N_25715,N_24090);
or U27949 (N_27949,N_25489,N_24836);
xor U27950 (N_27950,N_24128,N_24470);
or U27951 (N_27951,N_25324,N_25061);
xnor U27952 (N_27952,N_24814,N_25991);
or U27953 (N_27953,N_25067,N_25740);
nand U27954 (N_27954,N_24022,N_24838);
or U27955 (N_27955,N_25787,N_25313);
and U27956 (N_27956,N_25516,N_24072);
nor U27957 (N_27957,N_24358,N_24222);
nor U27958 (N_27958,N_24674,N_25083);
or U27959 (N_27959,N_25113,N_24617);
or U27960 (N_27960,N_25298,N_25046);
and U27961 (N_27961,N_25373,N_24897);
nor U27962 (N_27962,N_24960,N_24998);
nor U27963 (N_27963,N_24797,N_24393);
and U27964 (N_27964,N_24168,N_25928);
xor U27965 (N_27965,N_25393,N_24237);
xor U27966 (N_27966,N_25068,N_25468);
nor U27967 (N_27967,N_25766,N_24394);
xnor U27968 (N_27968,N_24271,N_25421);
nor U27969 (N_27969,N_25325,N_25629);
or U27970 (N_27970,N_25787,N_24280);
nand U27971 (N_27971,N_24776,N_24635);
and U27972 (N_27972,N_25139,N_24389);
nand U27973 (N_27973,N_24458,N_24744);
nand U27974 (N_27974,N_24459,N_24659);
and U27975 (N_27975,N_25501,N_24618);
and U27976 (N_27976,N_25467,N_25148);
nor U27977 (N_27977,N_24088,N_25210);
and U27978 (N_27978,N_25507,N_24830);
nand U27979 (N_27979,N_25348,N_24603);
or U27980 (N_27980,N_25922,N_25566);
and U27981 (N_27981,N_25397,N_25444);
nand U27982 (N_27982,N_25862,N_25954);
nor U27983 (N_27983,N_24473,N_24450);
nor U27984 (N_27984,N_24947,N_25182);
nand U27985 (N_27985,N_25319,N_25871);
and U27986 (N_27986,N_24397,N_24961);
nand U27987 (N_27987,N_25468,N_24856);
and U27988 (N_27988,N_25814,N_25892);
or U27989 (N_27989,N_25725,N_25602);
or U27990 (N_27990,N_24031,N_25317);
nand U27991 (N_27991,N_25180,N_24933);
xor U27992 (N_27992,N_25100,N_25922);
nand U27993 (N_27993,N_25804,N_25802);
xnor U27994 (N_27994,N_24797,N_25093);
xnor U27995 (N_27995,N_25640,N_25523);
and U27996 (N_27996,N_24959,N_25609);
and U27997 (N_27997,N_24652,N_24741);
and U27998 (N_27998,N_25467,N_24084);
and U27999 (N_27999,N_25602,N_25054);
nand U28000 (N_28000,N_26424,N_27073);
xor U28001 (N_28001,N_26731,N_27784);
xnor U28002 (N_28002,N_26537,N_26127);
xor U28003 (N_28003,N_26565,N_27843);
nand U28004 (N_28004,N_27469,N_27295);
or U28005 (N_28005,N_26704,N_26784);
nand U28006 (N_28006,N_27506,N_27879);
or U28007 (N_28007,N_27373,N_27017);
nand U28008 (N_28008,N_26927,N_26665);
and U28009 (N_28009,N_27076,N_27361);
and U28010 (N_28010,N_26336,N_26305);
nand U28011 (N_28011,N_26155,N_26102);
nor U28012 (N_28012,N_27712,N_26641);
and U28013 (N_28013,N_27253,N_26572);
nor U28014 (N_28014,N_27386,N_27819);
or U28015 (N_28015,N_27226,N_27065);
nand U28016 (N_28016,N_27875,N_27481);
nor U28017 (N_28017,N_26004,N_26380);
nand U28018 (N_28018,N_26893,N_26835);
xor U28019 (N_28019,N_26575,N_27929);
nand U28020 (N_28020,N_26212,N_27865);
and U28021 (N_28021,N_26753,N_26171);
nor U28022 (N_28022,N_27938,N_27293);
nor U28023 (N_28023,N_27093,N_27086);
or U28024 (N_28024,N_26685,N_26216);
nor U28025 (N_28025,N_26861,N_27381);
nor U28026 (N_28026,N_27070,N_26110);
nor U28027 (N_28027,N_27135,N_27264);
nor U28028 (N_28028,N_27905,N_26323);
nor U28029 (N_28029,N_26454,N_27384);
nor U28030 (N_28030,N_26053,N_26787);
or U28031 (N_28031,N_26369,N_27155);
xor U28032 (N_28032,N_26334,N_27857);
xor U28033 (N_28033,N_26453,N_26374);
or U28034 (N_28034,N_26942,N_26697);
or U28035 (N_28035,N_27051,N_26031);
nor U28036 (N_28036,N_27870,N_26436);
and U28037 (N_28037,N_26002,N_26370);
or U28038 (N_28038,N_26802,N_27651);
nor U28039 (N_28039,N_27650,N_27802);
xor U28040 (N_28040,N_26388,N_26748);
xor U28041 (N_28041,N_27926,N_26187);
nor U28042 (N_28042,N_26863,N_27636);
and U28043 (N_28043,N_26017,N_27113);
and U28044 (N_28044,N_26325,N_26023);
nor U28045 (N_28045,N_27511,N_26656);
nand U28046 (N_28046,N_26426,N_26885);
xnor U28047 (N_28047,N_27727,N_27431);
or U28048 (N_28048,N_26905,N_26610);
nor U28049 (N_28049,N_27700,N_27593);
or U28050 (N_28050,N_26159,N_26399);
nor U28051 (N_28051,N_26383,N_27831);
and U28052 (N_28052,N_27250,N_27907);
nor U28053 (N_28053,N_26793,N_27062);
or U28054 (N_28054,N_27358,N_27847);
nand U28055 (N_28055,N_27932,N_27614);
nand U28056 (N_28056,N_27467,N_27595);
xnor U28057 (N_28057,N_27818,N_27861);
xor U28058 (N_28058,N_26214,N_26098);
and U28059 (N_28059,N_27188,N_27441);
or U28060 (N_28060,N_27437,N_27222);
nor U28061 (N_28061,N_26706,N_27478);
xnor U28062 (N_28062,N_27805,N_27309);
or U28063 (N_28063,N_27344,N_26006);
nand U28064 (N_28064,N_27207,N_27339);
nand U28065 (N_28065,N_27710,N_27670);
nor U28066 (N_28066,N_26547,N_27356);
nor U28067 (N_28067,N_26373,N_26649);
xnor U28068 (N_28068,N_27814,N_26149);
and U28069 (N_28069,N_27349,N_27759);
and U28070 (N_28070,N_27797,N_26157);
nand U28071 (N_28071,N_27883,N_27448);
xor U28072 (N_28072,N_27761,N_27044);
nor U28073 (N_28073,N_26496,N_26766);
and U28074 (N_28074,N_26672,N_27045);
or U28075 (N_28075,N_27007,N_27308);
nand U28076 (N_28076,N_27732,N_26939);
nor U28077 (N_28077,N_26526,N_27137);
xnor U28078 (N_28078,N_27800,N_26679);
and U28079 (N_28079,N_27443,N_26810);
nor U28080 (N_28080,N_27164,N_27669);
nand U28081 (N_28081,N_27778,N_26936);
or U28082 (N_28082,N_26930,N_27081);
xnor U28083 (N_28083,N_27083,N_26594);
and U28084 (N_28084,N_26949,N_27615);
and U28085 (N_28085,N_27860,N_27816);
and U28086 (N_28086,N_26191,N_27176);
and U28087 (N_28087,N_26099,N_27647);
nor U28088 (N_28088,N_26966,N_27106);
and U28089 (N_28089,N_27713,N_26488);
nor U28090 (N_28090,N_27584,N_27195);
xor U28091 (N_28091,N_26777,N_26176);
or U28092 (N_28092,N_26612,N_27234);
and U28093 (N_28093,N_26137,N_26283);
or U28094 (N_28094,N_27413,N_27403);
and U28095 (N_28095,N_26328,N_26164);
or U28096 (N_28096,N_27163,N_27180);
xnor U28097 (N_28097,N_27142,N_26479);
nor U28098 (N_28098,N_26993,N_26534);
xor U28099 (N_28099,N_27125,N_27366);
xor U28100 (N_28100,N_27069,N_27617);
and U28101 (N_28101,N_27578,N_26446);
or U28102 (N_28102,N_26846,N_26552);
or U28103 (N_28103,N_27987,N_26347);
xor U28104 (N_28104,N_26838,N_27791);
and U28105 (N_28105,N_27054,N_26103);
xnor U28106 (N_28106,N_27733,N_27368);
xnor U28107 (N_28107,N_27406,N_27360);
nand U28108 (N_28108,N_27644,N_26541);
xor U28109 (N_28109,N_26986,N_26184);
xor U28110 (N_28110,N_26756,N_26686);
and U28111 (N_28111,N_26544,N_26282);
nor U28112 (N_28112,N_26958,N_26460);
nand U28113 (N_28113,N_26108,N_26307);
or U28114 (N_28114,N_26177,N_26293);
nor U28115 (N_28115,N_27322,N_26145);
or U28116 (N_28116,N_26985,N_26548);
nor U28117 (N_28117,N_27558,N_27502);
or U28118 (N_28118,N_27191,N_27346);
and U28119 (N_28119,N_27154,N_27648);
or U28120 (N_28120,N_27130,N_26324);
and U28121 (N_28121,N_26186,N_26485);
nand U28122 (N_28122,N_27653,N_27983);
nand U28123 (N_28123,N_27256,N_26476);
and U28124 (N_28124,N_26068,N_27399);
or U28125 (N_28125,N_27451,N_26249);
nand U28126 (N_28126,N_26082,N_26915);
nand U28127 (N_28127,N_27876,N_26759);
and U28128 (N_28128,N_26409,N_27618);
or U28129 (N_28129,N_26979,N_26058);
nand U28130 (N_28130,N_27335,N_27535);
nand U28131 (N_28131,N_26983,N_26524);
and U28132 (N_28132,N_27553,N_26218);
nor U28133 (N_28133,N_27904,N_26111);
or U28134 (N_28134,N_27931,N_26921);
nand U28135 (N_28135,N_27056,N_26188);
nand U28136 (N_28136,N_26754,N_27462);
nor U28137 (N_28137,N_27807,N_26900);
or U28138 (N_28138,N_27991,N_27075);
nor U28139 (N_28139,N_26288,N_27012);
and U28140 (N_28140,N_27064,N_26878);
xor U28141 (N_28141,N_26363,N_26126);
and U28142 (N_28142,N_26616,N_26167);
xor U28143 (N_28143,N_27949,N_26521);
nand U28144 (N_28144,N_26340,N_26296);
or U28145 (N_28145,N_26350,N_26318);
and U28146 (N_28146,N_27930,N_27059);
and U28147 (N_28147,N_27786,N_26179);
nor U28148 (N_28148,N_27171,N_27245);
nor U28149 (N_28149,N_26493,N_26841);
or U28150 (N_28150,N_27216,N_27785);
or U28151 (N_28151,N_26830,N_27579);
xnor U28152 (N_28152,N_26243,N_26258);
and U28153 (N_28153,N_26107,N_27992);
or U28154 (N_28154,N_26267,N_27205);
nand U28155 (N_28155,N_26505,N_27503);
nor U28156 (N_28156,N_27019,N_26408);
or U28157 (N_28157,N_27436,N_27912);
or U28158 (N_28158,N_27375,N_27129);
and U28159 (N_28159,N_26783,N_26634);
or U28160 (N_28160,N_26069,N_26281);
xnor U28161 (N_28161,N_27960,N_27353);
xor U28162 (N_28162,N_27474,N_26509);
or U28163 (N_28163,N_27189,N_26302);
nor U28164 (N_28164,N_27783,N_26019);
and U28165 (N_28165,N_27835,N_27951);
nand U28166 (N_28166,N_26445,N_26448);
or U28167 (N_28167,N_27588,N_26236);
nand U28168 (N_28168,N_26892,N_27116);
or U28169 (N_28169,N_27661,N_27925);
or U28170 (N_28170,N_26684,N_26129);
and U28171 (N_28171,N_27167,N_27817);
and U28172 (N_28172,N_26312,N_27998);
xor U28173 (N_28173,N_26471,N_27838);
or U28174 (N_28174,N_26175,N_27911);
xor U28175 (N_28175,N_26590,N_26842);
and U28176 (N_28176,N_27539,N_27336);
and U28177 (N_28177,N_26554,N_27048);
xnor U28178 (N_28178,N_27978,N_27852);
xnor U28179 (N_28179,N_26928,N_26173);
xnor U28180 (N_28180,N_26911,N_26086);
nand U28181 (N_28181,N_27283,N_27480);
xnor U28182 (N_28182,N_26276,N_27745);
nand U28183 (N_28183,N_27881,N_27694);
nand U28184 (N_28184,N_26192,N_27412);
nor U28185 (N_28185,N_26403,N_26333);
and U28186 (N_28186,N_26196,N_27679);
nor U28187 (N_28187,N_27763,N_27340);
nor U28188 (N_28188,N_27173,N_27776);
nand U28189 (N_28189,N_27418,N_26361);
or U28190 (N_28190,N_26235,N_27590);
or U28191 (N_28191,N_27976,N_26286);
nand U28192 (N_28192,N_26709,N_26331);
nand U28193 (N_28193,N_27587,N_27799);
xnor U28194 (N_28194,N_27550,N_26113);
nor U28195 (N_28195,N_27668,N_26978);
xnor U28196 (N_28196,N_27488,N_26732);
and U28197 (N_28197,N_26583,N_26193);
nor U28198 (N_28198,N_27545,N_27787);
nor U28199 (N_28199,N_27994,N_27476);
xor U28200 (N_28200,N_26353,N_27767);
nand U28201 (N_28201,N_26502,N_27301);
and U28202 (N_28202,N_26495,N_27552);
and U28203 (N_28203,N_26848,N_26545);
nand U28204 (N_28204,N_26938,N_26750);
xor U28205 (N_28205,N_27215,N_27836);
xor U28206 (N_28206,N_27306,N_26944);
nand U28207 (N_28207,N_26886,N_27842);
nor U28208 (N_28208,N_26007,N_26996);
nand U28209 (N_28209,N_27898,N_27049);
nor U28210 (N_28210,N_27908,N_27722);
nor U28211 (N_28211,N_27919,N_27655);
or U28212 (N_28212,N_26934,N_26794);
and U28213 (N_28213,N_26392,N_27546);
nor U28214 (N_28214,N_26628,N_27863);
nand U28215 (N_28215,N_26675,N_26116);
nand U28216 (N_28216,N_27260,N_27554);
nor U28217 (N_28217,N_26571,N_27294);
nand U28218 (N_28218,N_26504,N_27633);
nand U28219 (N_28219,N_26217,N_26459);
and U28220 (N_28220,N_26974,N_27702);
nand U28221 (N_28221,N_26132,N_27193);
xor U28222 (N_28222,N_27989,N_26077);
nand U28223 (N_28223,N_26028,N_27209);
nand U28224 (N_28224,N_27878,N_26051);
xor U28225 (N_28225,N_26608,N_27082);
xor U28226 (N_28226,N_27496,N_27198);
nand U28227 (N_28227,N_27956,N_27594);
nor U28228 (N_28228,N_27933,N_26751);
xnor U28229 (N_28229,N_27072,N_27122);
nand U28230 (N_28230,N_26024,N_27407);
nand U28231 (N_28231,N_27498,N_27156);
and U28232 (N_28232,N_26566,N_27683);
xor U28233 (N_28233,N_26382,N_26160);
and U28234 (N_28234,N_26876,N_27867);
xnor U28235 (N_28235,N_26523,N_26564);
or U28236 (N_28236,N_27228,N_27832);
or U28237 (N_28237,N_26584,N_27147);
nand U28238 (N_28238,N_27471,N_26860);
xor U28239 (N_28239,N_27034,N_26385);
nor U28240 (N_28240,N_27757,N_27280);
nand U28241 (N_28241,N_26278,N_26642);
or U28242 (N_28242,N_26128,N_27258);
xor U28243 (N_28243,N_27459,N_26531);
nor U28244 (N_28244,N_27078,N_26755);
or U28245 (N_28245,N_27362,N_26600);
nor U28246 (N_28246,N_26412,N_26183);
and U28247 (N_28247,N_26669,N_27909);
xnor U28248 (N_28248,N_27846,N_27004);
and U28249 (N_28249,N_27442,N_27940);
nand U28250 (N_28250,N_26744,N_27887);
nand U28251 (N_28251,N_27747,N_27916);
nand U28252 (N_28252,N_26648,N_27149);
xnor U28253 (N_28253,N_27782,N_26952);
nor U28254 (N_28254,N_27127,N_27533);
xnor U28255 (N_28255,N_26659,N_26617);
nand U28256 (N_28256,N_26849,N_27828);
nand U28257 (N_28257,N_26094,N_27305);
and U28258 (N_28258,N_27411,N_26620);
nand U28259 (N_28259,N_27845,N_27482);
nand U28260 (N_28260,N_26390,N_26394);
nor U28261 (N_28261,N_26255,N_27825);
and U28262 (N_28262,N_27131,N_26873);
and U28263 (N_28263,N_26297,N_27024);
nand U28264 (N_28264,N_27603,N_27434);
xor U28265 (N_28265,N_27500,N_26015);
nand U28266 (N_28266,N_26239,N_26883);
or U28267 (N_28267,N_27058,N_27141);
and U28268 (N_28268,N_27212,N_26664);
and U28269 (N_28269,N_27257,N_26712);
xor U28270 (N_28270,N_27374,N_27133);
and U28271 (N_28271,N_27756,N_27641);
or U28272 (N_28272,N_26260,N_26419);
and U28273 (N_28273,N_27066,N_26304);
xor U28274 (N_28274,N_27897,N_26317);
or U28275 (N_28275,N_27580,N_26428);
or U28276 (N_28276,N_26761,N_27858);
nor U28277 (N_28277,N_27543,N_27401);
xor U28278 (N_28278,N_27068,N_26055);
or U28279 (N_28279,N_26976,N_27225);
or U28280 (N_28280,N_26854,N_26377);
nor U28281 (N_28281,N_26977,N_27914);
xor U28282 (N_28282,N_26633,N_27321);
nor U28283 (N_28283,N_26042,N_26152);
and U28284 (N_28284,N_27332,N_26487);
and U28285 (N_28285,N_26461,N_26513);
or U28286 (N_28286,N_26158,N_26062);
nand U28287 (N_28287,N_26968,N_26231);
nor U28288 (N_28288,N_26889,N_26725);
or U28289 (N_28289,N_26533,N_27900);
nand U28290 (N_28290,N_26769,N_27917);
nor U28291 (N_28291,N_27510,N_27853);
and U28292 (N_28292,N_27598,N_27150);
or U28293 (N_28293,N_27248,N_26225);
and U28294 (N_28294,N_27018,N_27415);
or U28295 (N_28295,N_27682,N_27709);
xnor U28296 (N_28296,N_26210,N_26821);
nor U28297 (N_28297,N_27145,N_27087);
and U28298 (N_28298,N_26730,N_27052);
nand U28299 (N_28299,N_27118,N_27888);
and U28300 (N_28300,N_26064,N_26840);
nor U28301 (N_28301,N_27667,N_27788);
or U28302 (N_28302,N_26970,N_27972);
xnor U28303 (N_28303,N_27096,N_26011);
or U28304 (N_28304,N_27270,N_27906);
and U28305 (N_28305,N_27774,N_26497);
xor U28306 (N_28306,N_26964,N_26945);
or U28307 (N_28307,N_27859,N_27798);
nor U28308 (N_28308,N_27158,N_27996);
nor U28309 (N_28309,N_27479,N_26563);
and U28310 (N_28310,N_27752,N_26457);
and U28311 (N_28311,N_27963,N_27313);
xor U28312 (N_28312,N_26018,N_26035);
nand U28313 (N_28313,N_27117,N_26715);
nor U28314 (N_28314,N_27760,N_26988);
nand U28315 (N_28315,N_27796,N_27564);
or U28316 (N_28316,N_27291,N_27589);
and U28317 (N_28317,N_27182,N_27530);
nand U28318 (N_28318,N_26527,N_27014);
xnor U28319 (N_28319,N_26395,N_27273);
nor U28320 (N_28320,N_26814,N_26462);
nand U28321 (N_28321,N_27955,N_26681);
or U28322 (N_28322,N_27296,N_26598);
xnor U28323 (N_28323,N_26919,N_26559);
or U28324 (N_28324,N_26711,N_27604);
xor U28325 (N_28325,N_26588,N_26441);
and U28326 (N_28326,N_27329,N_27562);
or U28327 (N_28327,N_27187,N_27674);
and U28328 (N_28328,N_26615,N_26582);
or U28329 (N_28329,N_26314,N_26950);
xor U28330 (N_28330,N_26067,N_27977);
and U28331 (N_28331,N_26096,N_27043);
or U28332 (N_28332,N_27720,N_27608);
nor U28333 (N_28333,N_26875,N_27357);
nand U28334 (N_28334,N_27626,N_26010);
nand U28335 (N_28335,N_26285,N_27822);
or U28336 (N_28336,N_27707,N_26494);
or U28337 (N_28337,N_26718,N_26105);
nand U28338 (N_28338,N_26658,N_27902);
xor U28339 (N_28339,N_27862,N_27197);
and U28340 (N_28340,N_26003,N_27526);
or U28341 (N_28341,N_26894,N_27941);
or U28342 (N_28342,N_27023,N_27008);
and U28343 (N_28343,N_27490,N_26991);
or U28344 (N_28344,N_26182,N_26827);
nand U28345 (N_28345,N_26951,N_27020);
or U28346 (N_28346,N_26095,N_27923);
and U28347 (N_28347,N_26279,N_27586);
and U28348 (N_28348,N_26813,N_26029);
and U28349 (N_28349,N_27027,N_26039);
nor U28350 (N_28350,N_27492,N_26234);
nor U28351 (N_28351,N_26728,N_26902);
xor U28352 (N_28352,N_26817,N_26351);
and U28353 (N_28353,N_26301,N_26417);
or U28354 (N_28354,N_27962,N_27241);
nand U28355 (N_28355,N_27277,N_27591);
xor U28356 (N_28356,N_26063,N_26389);
nand U28357 (N_28357,N_26578,N_27328);
and U28358 (N_28358,N_27247,N_27943);
nand U28359 (N_28359,N_26933,N_26240);
and U28360 (N_28360,N_27246,N_26677);
nor U28361 (N_28361,N_27334,N_27851);
xnor U28362 (N_28362,N_26667,N_26908);
xnor U28363 (N_28363,N_26367,N_26808);
xnor U28364 (N_28364,N_26178,N_26972);
nand U28365 (N_28365,N_26984,N_27728);
and U28366 (N_28366,N_27190,N_26008);
xnor U28367 (N_28367,N_26960,N_27893);
nand U28368 (N_28368,N_26078,N_26506);
nand U28369 (N_28369,N_27186,N_27534);
nand U28370 (N_28370,N_27192,N_26346);
xnor U28371 (N_28371,N_27810,N_26912);
and U28372 (N_28372,N_27809,N_26273);
and U28373 (N_28373,N_27676,N_26238);
nand U28374 (N_28374,N_27903,N_26573);
and U28375 (N_28375,N_26291,N_27988);
nor U28376 (N_28376,N_26427,N_27687);
nand U28377 (N_28377,N_26200,N_26083);
nor U28378 (N_28378,N_27744,N_27445);
and U28379 (N_28379,N_27077,N_27120);
xnor U28380 (N_28380,N_26514,N_26593);
nor U28381 (N_28381,N_27529,N_27457);
xor U28382 (N_28382,N_27491,N_27566);
or U28383 (N_28383,N_27542,N_26717);
nor U28384 (N_28384,N_27446,N_27153);
or U28385 (N_28385,N_26166,N_27772);
and U28386 (N_28386,N_27243,N_26473);
xor U28387 (N_28387,N_27741,N_26115);
nand U28388 (N_28388,N_26655,N_26515);
xor U28389 (N_28389,N_27416,N_26219);
nand U28390 (N_28390,N_27821,N_27622);
or U28391 (N_28391,N_26118,N_27544);
nor U28392 (N_28392,N_27298,N_26376);
nor U28393 (N_28393,N_27515,N_26671);
nor U28394 (N_28394,N_26364,N_26070);
and U28395 (N_28395,N_26190,N_26980);
xor U28396 (N_28396,N_27168,N_26737);
and U28397 (N_28397,N_27850,N_27547);
nand U28398 (N_28398,N_26226,N_26466);
xnor U28399 (N_28399,N_27612,N_26532);
and U28400 (N_28400,N_27629,N_27029);
and U28401 (N_28401,N_26757,N_26562);
xnor U28402 (N_28402,N_26580,N_27556);
xor U28403 (N_28403,N_27691,N_27265);
or U28404 (N_28404,N_27826,N_26603);
and U28405 (N_28405,N_27954,N_26909);
xnor U28406 (N_28406,N_26269,N_27990);
nor U28407 (N_28407,N_27487,N_27119);
nand U28408 (N_28408,N_27704,N_27675);
nor U28409 (N_28409,N_27706,N_27729);
or U28410 (N_28410,N_27725,N_26136);
and U28411 (N_28411,N_27123,N_26591);
or U28412 (N_28412,N_26185,N_27948);
xnor U28413 (N_28413,N_27218,N_27229);
and U28414 (N_28414,N_27035,N_27477);
nand U28415 (N_28415,N_26792,N_26901);
nor U28416 (N_28416,N_27395,N_26740);
nand U28417 (N_28417,N_26081,N_26499);
nand U28418 (N_28418,N_27016,N_26680);
and U28419 (N_28419,N_26844,N_26089);
and U28420 (N_28420,N_27743,N_26696);
xor U28421 (N_28421,N_27946,N_26539);
or U28422 (N_28422,N_26907,N_26780);
nand U28423 (N_28423,N_26402,N_27061);
nand U28424 (N_28424,N_27607,N_27179);
or U28425 (N_28425,N_27521,N_26644);
xnor U28426 (N_28426,N_27178,N_27494);
and U28427 (N_28427,N_26246,N_27465);
or U28428 (N_28428,N_26943,N_26043);
xor U28429 (N_28429,N_27868,N_26887);
or U28430 (N_28430,N_27032,N_26021);
xor U28431 (N_28431,N_27272,N_26148);
nor U28432 (N_28432,N_26271,N_27238);
nand U28433 (N_28433,N_26799,N_26335);
and U28434 (N_28434,N_27697,N_26119);
or U28435 (N_28435,N_27400,N_26474);
xor U28436 (N_28436,N_27677,N_27646);
nand U28437 (N_28437,N_26440,N_26091);
nor U28438 (N_28438,N_27690,N_26154);
nor U28439 (N_28439,N_26000,N_27512);
and U28440 (N_28440,N_27200,N_27936);
nor U28441 (N_28441,N_27950,N_26880);
or U28442 (N_28442,N_26903,N_27316);
nor U28443 (N_28443,N_27582,N_26037);
and U28444 (N_28444,N_26843,N_26768);
nand U28445 (N_28445,N_27486,N_26061);
or U28446 (N_28446,N_27762,N_27924);
or U28447 (N_28447,N_27765,N_26822);
nor U28448 (N_28448,N_27516,N_27185);
nor U28449 (N_28449,N_26619,N_27703);
and U28450 (N_28450,N_26311,N_27249);
xnor U28451 (N_28451,N_26956,N_26222);
nand U28452 (N_28452,N_27428,N_26057);
nand U28453 (N_28453,N_27753,N_26967);
and U28454 (N_28454,N_27255,N_26451);
nor U28455 (N_28455,N_27665,N_27686);
or U28456 (N_28456,N_27639,N_26646);
nor U28457 (N_28457,N_26881,N_26241);
or U28458 (N_28458,N_27281,N_26606);
xnor U28459 (N_28459,N_27723,N_26447);
or U28460 (N_28460,N_27880,N_27021);
and U28461 (N_28461,N_27874,N_27995);
or U28462 (N_28462,N_26857,N_26244);
nor U28463 (N_28463,N_27746,N_26773);
or U28464 (N_28464,N_27750,N_27354);
xnor U28465 (N_28465,N_27177,N_26651);
nor U28466 (N_28466,N_26801,N_27110);
nand U28467 (N_28467,N_27731,N_26073);
nand U28468 (N_28468,N_27263,N_26101);
or U28469 (N_28469,N_27997,N_27770);
and U28470 (N_28470,N_27557,N_26948);
nand U28471 (N_28471,N_27261,N_27751);
nor U28472 (N_28472,N_27953,N_26125);
nor U28473 (N_28473,N_26404,N_26072);
xnor U28474 (N_28474,N_26992,N_27806);
or U28475 (N_28475,N_26144,N_26341);
or U28476 (N_28476,N_27681,N_26345);
nand U28477 (N_28477,N_27433,N_27551);
nor U28478 (N_28478,N_27312,N_26501);
xor U28479 (N_28479,N_26708,N_26250);
nor U28480 (N_28480,N_26692,N_27678);
or U28481 (N_28481,N_26026,N_27203);
or U28482 (N_28482,N_26925,N_26270);
or U28483 (N_28483,N_27327,N_27775);
xor U28484 (N_28484,N_26629,N_27097);
nor U28485 (N_28485,N_27872,N_26577);
nor U28486 (N_28486,N_27037,N_26492);
xnor U28487 (N_28487,N_27705,N_26862);
and U28488 (N_28488,N_26726,N_27755);
nand U28489 (N_28489,N_26483,N_26391);
and U28490 (N_28490,N_27895,N_27808);
xnor U28491 (N_28491,N_26468,N_26981);
nor U28492 (N_28492,N_26609,N_26439);
nand U28493 (N_28493,N_26469,N_26422);
or U28494 (N_28494,N_27297,N_27532);
or U28495 (N_28495,N_27517,N_26356);
xnor U28496 (N_28496,N_27599,N_26371);
xor U28497 (N_28497,N_26438,N_26087);
xnor U28498 (N_28498,N_27157,N_26811);
nor U28499 (N_28499,N_26044,N_26997);
xnor U28500 (N_28500,N_26172,N_27952);
nor U28501 (N_28501,N_27271,N_27314);
nor U28502 (N_28502,N_26033,N_27559);
nor U28503 (N_28503,N_27033,N_27408);
and U28504 (N_28504,N_26001,N_27438);
nor U28505 (N_28505,N_27624,N_27625);
xnor U28506 (N_28506,N_27126,N_26147);
or U28507 (N_28507,N_27719,N_27970);
or U28508 (N_28508,N_26449,N_27343);
nand U28509 (N_28509,N_26498,N_27605);
or U28510 (N_28510,N_27139,N_26174);
and U28511 (N_28511,N_26785,N_26994);
or U28512 (N_28512,N_27585,N_26618);
or U28513 (N_28513,N_26772,N_27734);
or U28514 (N_28514,N_26530,N_26798);
nand U28515 (N_28515,N_26831,N_27779);
nor U28516 (N_28516,N_27456,N_26198);
nand U28517 (N_28517,N_27473,N_27922);
nand U28518 (N_28518,N_27947,N_26396);
nand U28519 (N_28519,N_26112,N_27758);
and U28520 (N_28520,N_27421,N_26229);
nor U28521 (N_28521,N_26071,N_26989);
or U28522 (N_28522,N_26670,N_26433);
nor U28523 (N_28523,N_27716,N_27230);
or U28524 (N_28524,N_26660,N_27320);
xnor U28525 (N_28525,N_27227,N_27310);
nor U28526 (N_28526,N_27285,N_26969);
and U28527 (N_28527,N_27523,N_27402);
nand U28528 (N_28528,N_27387,N_26215);
or U28529 (N_28529,N_27439,N_27030);
nor U28530 (N_28530,N_27561,N_26349);
xor U28531 (N_28531,N_27921,N_27080);
and U28532 (N_28532,N_26771,N_27302);
nor U28533 (N_28533,N_27513,N_26330);
nand U28534 (N_28534,N_26678,N_27392);
or U28535 (N_28535,N_26005,N_26975);
and U28536 (N_28536,N_26607,N_26877);
and U28537 (N_28537,N_26481,N_26247);
nor U28538 (N_28538,N_27409,N_27262);
nand U28539 (N_28539,N_26957,N_27627);
nand U28540 (N_28540,N_26856,N_26140);
nand U28541 (N_28541,N_26213,N_27036);
nand U28542 (N_28542,N_26904,N_26084);
nor U28543 (N_28543,N_26625,N_26899);
nor U28544 (N_28544,N_27689,N_27444);
or U28545 (N_28545,N_27333,N_27107);
and U28546 (N_28546,N_26700,N_27568);
and U28547 (N_28547,N_27204,N_26315);
nand U28548 (N_28548,N_27531,N_26721);
nor U28549 (N_28549,N_27645,N_27284);
and U28550 (N_28550,N_26774,N_26729);
and U28551 (N_28551,N_27183,N_27251);
nor U28552 (N_28552,N_27606,N_26195);
xor U28553 (N_28553,N_26066,N_26429);
and U28554 (N_28554,N_26227,N_26106);
or U28555 (N_28555,N_27672,N_27520);
and U28556 (N_28556,N_26657,N_26248);
and U28557 (N_28557,N_26516,N_27640);
nand U28558 (N_28558,N_26253,N_27768);
nor U28559 (N_28559,N_27074,N_26682);
or U28560 (N_28560,N_27538,N_27159);
xnor U28561 (N_28561,N_26163,N_26987);
and U28562 (N_28562,N_27514,N_27601);
and U28563 (N_28563,N_27792,N_27342);
nor U28564 (N_28564,N_27664,N_26569);
nor U28565 (N_28565,N_26022,N_26941);
and U28566 (N_28566,N_27528,N_26027);
xor U28567 (N_28567,N_27737,N_26917);
or U28568 (N_28568,N_27967,N_26202);
xnor U28569 (N_28569,N_27570,N_27958);
xnor U28570 (N_28570,N_26816,N_26931);
nand U28571 (N_28571,N_26828,N_27449);
nor U28572 (N_28572,N_27696,N_27470);
and U28573 (N_28573,N_27405,N_26458);
or U28574 (N_28574,N_26245,N_27315);
and U28575 (N_28575,N_26170,N_27985);
xor U28576 (N_28576,N_26401,N_27969);
xor U28577 (N_28577,N_26543,N_27508);
and U28578 (N_28578,N_27913,N_27658);
and U28579 (N_28579,N_27896,N_26074);
nand U28580 (N_28580,N_27435,N_26384);
xnor U28581 (N_28581,N_26169,N_26257);
xor U28582 (N_28582,N_27920,N_27174);
xor U28583 (N_28583,N_26359,N_26268);
xor U28584 (N_28584,N_26701,N_26254);
xnor U28585 (N_28585,N_27856,N_27337);
xnor U28586 (N_28586,N_26542,N_27091);
nand U28587 (N_28587,N_27011,N_26032);
nand U28588 (N_28588,N_26261,N_27304);
or U28589 (N_28589,N_27583,N_26054);
and U28590 (N_28590,N_26668,N_27965);
nand U28591 (N_28591,N_26770,N_27370);
and U28592 (N_28592,N_26865,N_26638);
nand U28593 (N_28593,N_26971,N_26805);
and U28594 (N_28594,N_26558,N_26561);
xor U28595 (N_28595,N_26437,N_26251);
or U28596 (N_28596,N_26040,N_27244);
nor U28597 (N_28597,N_27038,N_26557);
nand U28598 (N_28598,N_27472,N_27440);
xnor U28599 (N_28599,N_27892,N_26151);
or U28600 (N_28600,N_26742,N_27221);
xor U28601 (N_28601,N_26643,N_27864);
nor U28602 (N_28602,N_26060,N_27871);
xnor U28603 (N_28603,N_27202,N_26475);
and U28604 (N_28604,N_26674,N_26386);
xnor U28605 (N_28605,N_27282,N_26209);
xor U28606 (N_28606,N_26745,N_27928);
nor U28607 (N_28607,N_26430,N_27430);
nand U28608 (N_28608,N_27391,N_26233);
and U28609 (N_28609,N_26699,N_26150);
xnor U28610 (N_28610,N_26012,N_26631);
nand U28611 (N_28611,N_26122,N_26546);
nor U28612 (N_28612,N_27420,N_27942);
or U28613 (N_28613,N_27351,N_27764);
nor U28614 (N_28614,N_27427,N_26199);
nor U28615 (N_28615,N_27964,N_26688);
or U28616 (N_28616,N_27397,N_26423);
and U28617 (N_28617,N_27780,N_27827);
xor U28618 (N_28618,N_26747,N_26207);
xnor U28619 (N_28619,N_27447,N_26228);
and U28620 (N_28620,N_27602,N_26898);
nand U28621 (N_28621,N_27934,N_27609);
or U28622 (N_28622,N_27208,N_26372);
and U28623 (N_28623,N_27596,N_27882);
or U28624 (N_28624,N_26973,N_27338);
and U28625 (N_28625,N_26895,N_27522);
nor U28626 (N_28626,N_26597,N_27383);
nor U28627 (N_28627,N_27957,N_26852);
and U28628 (N_28628,N_27112,N_26906);
nor U28629 (N_28629,N_27986,N_27592);
nor U28630 (N_28630,N_26525,N_27649);
nand U28631 (N_28631,N_27781,N_27695);
nor U28632 (N_28632,N_26553,N_27981);
nor U28633 (N_28633,N_26418,N_26640);
or U28634 (N_28634,N_27039,N_26321);
nand U28635 (N_28635,N_26507,N_27266);
or U28636 (N_28636,N_27220,N_26491);
xor U28637 (N_28637,N_26352,N_26826);
xnor U28638 (N_28638,N_27289,N_27466);
nand U28639 (N_28639,N_26818,N_26549);
xor U28640 (N_28640,N_27026,N_26824);
nor U28641 (N_28641,N_27028,N_26647);
nor U28642 (N_28642,N_26421,N_26259);
and U28643 (N_28643,N_27146,N_26280);
nand U28644 (N_28644,N_27688,N_26693);
or U28645 (N_28645,N_26274,N_26326);
or U28646 (N_28646,N_26104,N_27453);
nor U28647 (N_28647,N_27365,N_26605);
nand U28648 (N_28648,N_27324,N_26139);
nand U28649 (N_28649,N_26632,N_26411);
nor U28650 (N_28650,N_26832,N_27715);
nor U28651 (N_28651,N_27548,N_26540);
and U28652 (N_28652,N_27915,N_26809);
nand U28653 (N_28653,N_26850,N_27572);
nor U28654 (N_28654,N_27485,N_26845);
nand U28655 (N_28655,N_27345,N_27540);
nand U28656 (N_28656,N_26752,N_26834);
nand U28657 (N_28657,N_26009,N_27194);
nand U28658 (N_28658,N_27162,N_26707);
nand U28659 (N_28659,N_27359,N_26237);
and U28660 (N_28660,N_26079,N_26300);
and U28661 (N_28661,N_26758,N_26738);
xor U28662 (N_28662,N_27721,N_26360);
or U28663 (N_28663,N_26637,N_26653);
xor U28664 (N_28664,N_26041,N_26538);
nand U28665 (N_28665,N_27458,N_27777);
or U28666 (N_28666,N_27372,N_26627);
xnor U28667 (N_28667,N_27053,N_26080);
and U28668 (N_28668,N_27060,N_26796);
nand U28669 (N_28669,N_26478,N_26398);
and U28670 (N_28670,N_26716,N_27840);
nor U28671 (N_28671,N_27815,N_27259);
nand U28672 (N_28672,N_26626,N_27005);
and U28673 (N_28673,N_27652,N_26414);
nor U28674 (N_28674,N_26884,N_27055);
and U28675 (N_28675,N_27015,N_26162);
nor U28676 (N_28676,N_26733,N_27143);
nor U28677 (N_28677,N_26292,N_27378);
and U28678 (N_28678,N_26791,N_26735);
and U28679 (N_28679,N_26630,N_27993);
nand U28680 (N_28680,N_27611,N_27736);
or U28681 (N_28681,N_26666,N_27555);
xnor U28682 (N_28682,N_26923,N_26076);
and U28683 (N_28683,N_26443,N_26432);
nand U28684 (N_28684,N_26407,N_26635);
or U28685 (N_28685,N_27352,N_26954);
nand U28686 (N_28686,N_26922,N_26604);
nand U28687 (N_28687,N_26581,N_26963);
nand U28688 (N_28688,N_27140,N_27394);
and U28689 (N_28689,N_26518,N_26463);
and U28690 (N_28690,N_27869,N_27311);
nand U28691 (N_28691,N_27549,N_26959);
nor U28692 (N_28692,N_27206,N_27396);
nor U28693 (N_28693,N_26940,N_27041);
nand U28694 (N_28694,N_26511,N_26998);
and U28695 (N_28695,N_26536,N_26464);
nand U28696 (N_28696,N_27376,N_27974);
nor U28697 (N_28697,N_27377,N_27422);
nor U28698 (N_28698,N_26025,N_27899);
nand U28699 (N_28699,N_26661,N_26743);
nand U28700 (N_28700,N_27886,N_26639);
and U28701 (N_28701,N_26142,N_27254);
xnor U28702 (N_28702,N_26090,N_27837);
nor U28703 (N_28703,N_26654,N_26425);
nand U28704 (N_28704,N_26265,N_26294);
nor U28705 (N_28705,N_27812,N_26789);
nor U28706 (N_28706,N_27463,N_27569);
and U28707 (N_28707,N_26723,N_27701);
nor U28708 (N_28708,N_27223,N_27656);
nand U28709 (N_28709,N_26224,N_26556);
and U28710 (N_28710,N_26413,N_27484);
nor U28711 (N_28711,N_26263,N_27673);
and U28712 (N_28712,N_27279,N_26316);
and U28713 (N_28713,N_26309,N_27468);
nand U28714 (N_28714,N_27499,N_26870);
nor U28715 (N_28715,N_27268,N_26358);
nor U28716 (N_28716,N_26313,N_27303);
nand U28717 (N_28717,N_26990,N_26036);
or U28718 (N_28718,N_26092,N_27654);
and U28719 (N_28719,N_27717,N_27201);
xnor U28720 (N_28720,N_27820,N_26576);
nor U28721 (N_28721,N_26803,N_26691);
and U28722 (N_28722,N_27410,N_26047);
and U28723 (N_28723,N_26882,N_26866);
and U28724 (N_28724,N_27979,N_26763);
nand U28725 (N_28725,N_26277,N_27001);
nand U28726 (N_28726,N_27666,N_26613);
nand U28727 (N_28727,N_26477,N_27169);
nor U28728 (N_28728,N_26916,N_26853);
xor U28729 (N_28729,N_27749,N_27698);
nand U28730 (N_28730,N_26056,N_26713);
xor U28731 (N_28731,N_26775,N_27105);
and U28732 (N_28732,N_26965,N_27455);
nor U28733 (N_28733,N_26705,N_27144);
or U28734 (N_28734,N_27748,N_26470);
xor U28735 (N_28735,N_26702,N_27331);
nor U28736 (N_28736,N_26306,N_27849);
nand U28737 (N_28737,N_26223,N_27114);
nor U28738 (N_28738,N_26045,N_27684);
and U28739 (N_28739,N_27050,N_27927);
nand U28740 (N_28740,N_26365,N_27497);
and U28741 (N_28741,N_27236,N_26764);
and U28742 (N_28742,N_27450,N_27663);
nand U28743 (N_28743,N_26181,N_26962);
xnor U28744 (N_28744,N_27935,N_26663);
xnor U28745 (N_28745,N_27839,N_26332);
nand U28746 (N_28746,N_26587,N_26052);
and U28747 (N_28747,N_27240,N_27945);
or U28748 (N_28748,N_26806,N_27769);
or U28749 (N_28749,N_26455,N_26100);
or U28750 (N_28750,N_26130,N_27610);
nor U28751 (N_28751,N_27090,N_26602);
xnor U28752 (N_28752,N_26528,N_27382);
or U28753 (N_28753,N_26308,N_26555);
nor U28754 (N_28754,N_26013,N_26189);
nor U28755 (N_28755,N_27108,N_27278);
nand U28756 (N_28756,N_26415,N_26320);
or U28757 (N_28757,N_27619,N_27371);
nor U28758 (N_28758,N_27326,N_27771);
xnor U28759 (N_28759,N_26232,N_26503);
nand U28760 (N_28760,N_26579,N_27095);
or U28761 (N_28761,N_26982,N_27982);
or U28762 (N_28762,N_27010,N_26075);
or U28763 (N_28763,N_27094,N_26121);
and U28764 (N_28764,N_27855,N_27623);
or U28765 (N_28765,N_27597,N_26741);
nor U28766 (N_28766,N_26790,N_26357);
nor U28767 (N_28767,N_27891,N_27866);
or U28768 (N_28768,N_26109,N_27973);
or U28769 (N_28769,N_27693,N_26393);
or U28770 (N_28770,N_27565,N_26093);
nor U28771 (N_28771,N_27388,N_27460);
or U28772 (N_28772,N_26955,N_26165);
nor U28773 (N_28773,N_27848,N_26135);
nor U28774 (N_28774,N_26937,N_26614);
and U28775 (N_28775,N_26120,N_27638);
xnor U28776 (N_28776,N_27642,N_27489);
xor U28777 (N_28777,N_26703,N_26867);
and U28778 (N_28778,N_26319,N_26890);
or U28779 (N_28779,N_27031,N_27844);
nor U28780 (N_28780,N_26508,N_26918);
nand U28781 (N_28781,N_26355,N_27057);
nor U28782 (N_28782,N_26180,N_26676);
nor U28783 (N_28783,N_26570,N_26624);
or U28784 (N_28784,N_26467,N_27219);
and U28785 (N_28785,N_26059,N_27109);
nor U28786 (N_28786,N_26623,N_26872);
and U28787 (N_28787,N_27999,N_26085);
xor U28788 (N_28788,N_27801,N_27877);
nor U28789 (N_28789,N_26327,N_26746);
xor U28790 (N_28790,N_26387,N_27009);
or U28791 (N_28791,N_26611,N_27237);
nand U28792 (N_28792,N_27184,N_27730);
and U28793 (N_28793,N_26289,N_27711);
and U28794 (N_28794,N_26858,N_27873);
nor U28795 (N_28795,N_26897,N_27111);
xnor U28796 (N_28796,N_26522,N_27134);
or U28797 (N_28797,N_27299,N_26156);
and U28798 (N_28798,N_26924,N_26201);
nor U28799 (N_28799,N_27239,N_27475);
nand U28800 (N_28800,N_27461,N_26490);
or U28801 (N_28801,N_27323,N_26134);
nand U28802 (N_28802,N_26420,N_26208);
or U28803 (N_28803,N_27084,N_27138);
xor U28804 (N_28804,N_26204,N_26456);
xnor U28805 (N_28805,N_26368,N_27577);
nor U28806 (N_28806,N_26779,N_27417);
xnor U28807 (N_28807,N_26695,N_26714);
nand U28808 (N_28808,N_27918,N_26284);
or U28809 (N_28809,N_27347,N_26143);
and U28810 (N_28810,N_26815,N_27170);
and U28811 (N_28811,N_27419,N_26535);
nor U28812 (N_28812,N_26762,N_26337);
nand U28813 (N_28813,N_27726,N_26168);
or U28814 (N_28814,N_26153,N_27735);
or U28815 (N_28815,N_26953,N_27181);
nor U28816 (N_28816,N_27196,N_27754);
xnor U28817 (N_28817,N_27136,N_27939);
nor U28818 (N_28818,N_26275,N_27276);
and U28819 (N_28819,N_27794,N_27884);
nor U28820 (N_28820,N_27635,N_27414);
or U28821 (N_28821,N_27286,N_26290);
and U28822 (N_28822,N_27854,N_26298);
nand U28823 (N_28823,N_26690,N_26864);
xnor U28824 (N_28824,N_26482,N_27724);
nor U28825 (N_28825,N_26820,N_27275);
or U28826 (N_28826,N_26694,N_27104);
nand U28827 (N_28827,N_27232,N_27317);
or U28828 (N_28828,N_26434,N_27789);
or U28829 (N_28829,N_27067,N_27124);
and U28830 (N_28830,N_26416,N_27235);
nor U28831 (N_28831,N_27288,N_26804);
nand U28832 (N_28832,N_27092,N_26891);
xor U28833 (N_28833,N_26961,N_27132);
nand U28834 (N_28834,N_26836,N_26935);
or U28835 (N_28835,N_26203,N_27390);
and U28836 (N_28836,N_27890,N_26833);
nand U28837 (N_28837,N_26344,N_27637);
nand U28838 (N_28838,N_27426,N_26592);
nand U28839 (N_28839,N_27959,N_27657);
nor U28840 (N_28840,N_27089,N_26765);
nor U28841 (N_28841,N_27398,N_27040);
nor U28842 (N_28842,N_27269,N_27984);
nand U28843 (N_28843,N_27507,N_27563);
xor U28844 (N_28844,N_27574,N_26450);
or U28845 (N_28845,N_26859,N_27660);
nor U28846 (N_28846,N_26839,N_27575);
xnor U28847 (N_28847,N_26366,N_26117);
or U28848 (N_28848,N_27600,N_27424);
xnor U28849 (N_28849,N_27003,N_26689);
xor U28850 (N_28850,N_27432,N_26776);
nor U28851 (N_28851,N_26295,N_26484);
xnor U28852 (N_28852,N_27103,N_26339);
nor U28853 (N_28853,N_26375,N_27423);
or U28854 (N_28854,N_27330,N_26807);
xnor U28855 (N_28855,N_27389,N_26879);
nor U28856 (N_28856,N_26266,N_27527);
or U28857 (N_28857,N_27699,N_26397);
nand U28858 (N_28858,N_27319,N_26512);
nand U28859 (N_28859,N_27576,N_27350);
and U28860 (N_28860,N_27631,N_27252);
and U28861 (N_28861,N_27738,N_26131);
nand U28862 (N_28862,N_27233,N_27231);
nor U28863 (N_28863,N_27047,N_27620);
nand U28864 (N_28864,N_26161,N_27128);
nand U28865 (N_28865,N_26673,N_27161);
xor U28866 (N_28866,N_27099,N_27525);
nor U28867 (N_28867,N_27505,N_26338);
nand U28868 (N_28868,N_26724,N_26560);
nor U28869 (N_28869,N_27613,N_27537);
nand U28870 (N_28870,N_26896,N_27823);
nand U28871 (N_28871,N_26823,N_26486);
or U28872 (N_28872,N_26829,N_27079);
or U28873 (N_28873,N_27560,N_27740);
xnor U28874 (N_28874,N_26914,N_27901);
or U28875 (N_28875,N_27483,N_27790);
or U28876 (N_28876,N_27536,N_27364);
nand U28877 (N_28877,N_26211,N_26727);
and U28878 (N_28878,N_27148,N_27966);
or U28879 (N_28879,N_27630,N_27274);
xnor U28880 (N_28880,N_27214,N_27355);
nor U28881 (N_28881,N_27100,N_26855);
xor U28882 (N_28882,N_27509,N_27224);
or U28883 (N_28883,N_27971,N_26303);
and U28884 (N_28884,N_26264,N_26310);
and U28885 (N_28885,N_26205,N_26946);
nor U28886 (N_28886,N_26206,N_27363);
nand U28887 (N_28887,N_26065,N_27910);
and U28888 (N_28888,N_26868,N_27085);
or U28889 (N_28889,N_27454,N_27101);
nand U28890 (N_28890,N_27292,N_26652);
xnor U28891 (N_28891,N_26381,N_26342);
or U28892 (N_28892,N_26739,N_26343);
nand U28893 (N_28893,N_26252,N_26030);
nor U28894 (N_28894,N_26230,N_27404);
nand U28895 (N_28895,N_26194,N_27002);
and U28896 (N_28896,N_27115,N_27714);
or U28897 (N_28897,N_27841,N_26683);
and U28898 (N_28898,N_27307,N_26322);
or U28899 (N_28899,N_26256,N_27616);
nand U28900 (N_28900,N_27718,N_27829);
nand U28901 (N_28901,N_26550,N_27571);
nor U28902 (N_28902,N_27242,N_26088);
nand U28903 (N_28903,N_27937,N_27739);
or U28904 (N_28904,N_27166,N_27518);
or U28905 (N_28905,N_27121,N_26348);
xnor U28906 (N_28906,N_26014,N_27318);
nand U28907 (N_28907,N_26114,N_27567);
or U28908 (N_28908,N_26995,N_27573);
nor U28909 (N_28909,N_26287,N_26472);
or U28910 (N_28910,N_27813,N_26141);
and U28911 (N_28911,N_27063,N_26520);
nor U28912 (N_28912,N_26767,N_26586);
xor U28913 (N_28913,N_27172,N_26123);
or U28914 (N_28914,N_27367,N_26020);
nor U28915 (N_28915,N_26034,N_26049);
nand U28916 (N_28916,N_26444,N_26800);
and U28917 (N_28917,N_27501,N_27175);
xnor U28918 (N_28918,N_27385,N_27210);
nand U28919 (N_28919,N_26662,N_26272);
nor U28920 (N_28920,N_26910,N_26480);
xnor U28921 (N_28921,N_27803,N_27025);
or U28922 (N_28922,N_26622,N_27504);
or U28923 (N_28923,N_26888,N_27643);
xnor U28924 (N_28924,N_27325,N_27944);
xor U28925 (N_28925,N_26920,N_26146);
nor U28926 (N_28926,N_27300,N_27006);
xor U28927 (N_28927,N_26050,N_26406);
nand U28928 (N_28928,N_27000,N_27961);
or U28929 (N_28929,N_27013,N_26947);
or U28930 (N_28930,N_26435,N_26929);
xnor U28931 (N_28931,N_26795,N_26197);
or U28932 (N_28932,N_27042,N_27524);
nor U28933 (N_28933,N_26687,N_27519);
xor U28934 (N_28934,N_26760,N_26329);
nor U28935 (N_28935,N_27464,N_26452);
or U28936 (N_28936,N_27102,N_26221);
nor U28937 (N_28937,N_26405,N_26574);
xnor U28938 (N_28938,N_27685,N_27393);
or U28939 (N_28939,N_27495,N_27541);
and U28940 (N_28940,N_26529,N_27217);
nand U28941 (N_28941,N_27834,N_26048);
or U28942 (N_28942,N_27267,N_27581);
or U28943 (N_28943,N_26599,N_27199);
xnor U28944 (N_28944,N_27811,N_26837);
nand U28945 (N_28945,N_26362,N_26354);
and U28946 (N_28946,N_26567,N_26016);
xor U28947 (N_28947,N_26138,N_27379);
or U28948 (N_28948,N_26489,N_27833);
or U28949 (N_28949,N_27621,N_27425);
xor U28950 (N_28950,N_26847,N_27071);
nand U28951 (N_28951,N_26719,N_26851);
or U28952 (N_28952,N_26038,N_27151);
and U28953 (N_28953,N_27830,N_27968);
or U28954 (N_28954,N_27885,N_27894);
and U28955 (N_28955,N_26400,N_27671);
or U28956 (N_28956,N_26786,N_27766);
or U28957 (N_28957,N_26596,N_26734);
nand U28958 (N_28958,N_26913,N_26782);
nand U28959 (N_28959,N_26410,N_26551);
or U28960 (N_28960,N_27793,N_26825);
nor U28961 (N_28961,N_27213,N_26500);
and U28962 (N_28962,N_26926,N_26442);
nor U28963 (N_28963,N_27795,N_27287);
or U28964 (N_28964,N_26517,N_27152);
nor U28965 (N_28965,N_27680,N_27211);
or U28966 (N_28966,N_27046,N_26589);
xnor U28967 (N_28967,N_27348,N_26220);
and U28968 (N_28968,N_27341,N_26097);
and U28969 (N_28969,N_27708,N_26046);
nand U28970 (N_28970,N_27369,N_26133);
and U28971 (N_28971,N_26262,N_26650);
nand U28972 (N_28972,N_27165,N_26698);
nor U28973 (N_28973,N_27290,N_27659);
nor U28974 (N_28974,N_27493,N_26645);
or U28975 (N_28975,N_26736,N_26431);
and U28976 (N_28976,N_27975,N_27662);
and U28977 (N_28977,N_26621,N_26720);
and U28978 (N_28978,N_26636,N_27380);
or U28979 (N_28979,N_26510,N_27632);
nand U28980 (N_28980,N_26585,N_26932);
nand U28981 (N_28981,N_26781,N_26778);
xor U28982 (N_28982,N_27889,N_27692);
and U28983 (N_28983,N_26710,N_26722);
nor U28984 (N_28984,N_26797,N_26999);
nand U28985 (N_28985,N_27098,N_26819);
or U28986 (N_28986,N_27452,N_27824);
or U28987 (N_28987,N_26299,N_27429);
xnor U28988 (N_28988,N_26595,N_26568);
and U28989 (N_28989,N_27980,N_26379);
nor U28990 (N_28990,N_27628,N_26601);
and U28991 (N_28991,N_26812,N_26465);
or U28992 (N_28992,N_27022,N_27742);
or U28993 (N_28993,N_26869,N_26871);
or U28994 (N_28994,N_26788,N_27804);
xnor U28995 (N_28995,N_26124,N_27773);
or U28996 (N_28996,N_26749,N_26242);
nand U28997 (N_28997,N_27160,N_26874);
and U28998 (N_28998,N_27634,N_26519);
xnor U28999 (N_28999,N_27088,N_26378);
or U29000 (N_29000,N_26808,N_26302);
and U29001 (N_29001,N_26966,N_27589);
nand U29002 (N_29002,N_27571,N_27956);
or U29003 (N_29003,N_26651,N_27251);
and U29004 (N_29004,N_26293,N_26635);
xor U29005 (N_29005,N_26334,N_26552);
xor U29006 (N_29006,N_27252,N_27596);
nand U29007 (N_29007,N_26463,N_26466);
nand U29008 (N_29008,N_27410,N_27740);
xor U29009 (N_29009,N_26687,N_26427);
or U29010 (N_29010,N_26728,N_26291);
nand U29011 (N_29011,N_26345,N_27016);
and U29012 (N_29012,N_27336,N_27363);
and U29013 (N_29013,N_27445,N_26699);
and U29014 (N_29014,N_27813,N_26567);
nor U29015 (N_29015,N_27642,N_27447);
nor U29016 (N_29016,N_26979,N_27212);
nand U29017 (N_29017,N_27323,N_27362);
or U29018 (N_29018,N_26380,N_27392);
or U29019 (N_29019,N_26330,N_26548);
nor U29020 (N_29020,N_26805,N_27572);
nor U29021 (N_29021,N_26256,N_27442);
or U29022 (N_29022,N_27280,N_26893);
xnor U29023 (N_29023,N_27976,N_26092);
or U29024 (N_29024,N_26558,N_26245);
and U29025 (N_29025,N_26708,N_27396);
and U29026 (N_29026,N_26899,N_26787);
or U29027 (N_29027,N_27436,N_27357);
nor U29028 (N_29028,N_26963,N_26950);
or U29029 (N_29029,N_27780,N_26088);
or U29030 (N_29030,N_26029,N_27273);
and U29031 (N_29031,N_27806,N_26963);
nor U29032 (N_29032,N_27526,N_26276);
xnor U29033 (N_29033,N_26587,N_26083);
xnor U29034 (N_29034,N_26710,N_27838);
nand U29035 (N_29035,N_26359,N_27024);
xor U29036 (N_29036,N_26615,N_26629);
or U29037 (N_29037,N_26382,N_26171);
nand U29038 (N_29038,N_27968,N_27005);
or U29039 (N_29039,N_26671,N_27162);
xnor U29040 (N_29040,N_27924,N_26988);
xor U29041 (N_29041,N_27622,N_26368);
nor U29042 (N_29042,N_26701,N_27550);
xnor U29043 (N_29043,N_26792,N_26432);
and U29044 (N_29044,N_26171,N_26811);
nor U29045 (N_29045,N_27987,N_26360);
xor U29046 (N_29046,N_27400,N_27890);
or U29047 (N_29047,N_27636,N_26236);
or U29048 (N_29048,N_26753,N_26135);
xor U29049 (N_29049,N_27631,N_26738);
nor U29050 (N_29050,N_27323,N_27087);
nor U29051 (N_29051,N_27001,N_27162);
nand U29052 (N_29052,N_26697,N_27499);
or U29053 (N_29053,N_27301,N_26232);
nand U29054 (N_29054,N_27030,N_27128);
and U29055 (N_29055,N_26012,N_27503);
xnor U29056 (N_29056,N_27875,N_27498);
or U29057 (N_29057,N_26714,N_27933);
xor U29058 (N_29058,N_26088,N_27633);
xor U29059 (N_29059,N_26246,N_26974);
xnor U29060 (N_29060,N_26783,N_27258);
nor U29061 (N_29061,N_26963,N_26180);
and U29062 (N_29062,N_27822,N_27800);
or U29063 (N_29063,N_27237,N_27192);
or U29064 (N_29064,N_26238,N_26599);
nor U29065 (N_29065,N_27335,N_26901);
nand U29066 (N_29066,N_27206,N_26065);
and U29067 (N_29067,N_27162,N_26234);
xor U29068 (N_29068,N_26809,N_26870);
nor U29069 (N_29069,N_26974,N_26827);
nor U29070 (N_29070,N_27668,N_27493);
xor U29071 (N_29071,N_27536,N_27133);
or U29072 (N_29072,N_27638,N_27004);
and U29073 (N_29073,N_26876,N_27131);
xor U29074 (N_29074,N_26606,N_26534);
xor U29075 (N_29075,N_27992,N_26719);
nand U29076 (N_29076,N_26819,N_26785);
nand U29077 (N_29077,N_27439,N_26933);
nand U29078 (N_29078,N_27447,N_26776);
nor U29079 (N_29079,N_26173,N_26941);
xor U29080 (N_29080,N_27822,N_26875);
nor U29081 (N_29081,N_26957,N_27657);
xnor U29082 (N_29082,N_27848,N_26759);
nand U29083 (N_29083,N_26408,N_27088);
xnor U29084 (N_29084,N_27029,N_26913);
and U29085 (N_29085,N_26934,N_27552);
nor U29086 (N_29086,N_27739,N_26377);
nor U29087 (N_29087,N_26729,N_26557);
and U29088 (N_29088,N_27903,N_27398);
and U29089 (N_29089,N_27395,N_27479);
or U29090 (N_29090,N_26187,N_27043);
nor U29091 (N_29091,N_26118,N_26965);
nor U29092 (N_29092,N_27823,N_27014);
nand U29093 (N_29093,N_26804,N_27959);
xnor U29094 (N_29094,N_26236,N_27721);
and U29095 (N_29095,N_26865,N_27708);
xnor U29096 (N_29096,N_26789,N_27677);
nand U29097 (N_29097,N_27298,N_27175);
or U29098 (N_29098,N_27651,N_26399);
xnor U29099 (N_29099,N_26829,N_27166);
nand U29100 (N_29100,N_26076,N_26532);
or U29101 (N_29101,N_26245,N_26866);
and U29102 (N_29102,N_27004,N_27205);
and U29103 (N_29103,N_26625,N_26013);
xor U29104 (N_29104,N_26592,N_26245);
xnor U29105 (N_29105,N_27001,N_26854);
nor U29106 (N_29106,N_27147,N_26615);
nor U29107 (N_29107,N_26292,N_26852);
nor U29108 (N_29108,N_26085,N_26003);
or U29109 (N_29109,N_27942,N_27896);
xnor U29110 (N_29110,N_26207,N_26354);
nand U29111 (N_29111,N_26251,N_26585);
and U29112 (N_29112,N_26678,N_27266);
or U29113 (N_29113,N_27487,N_26492);
nand U29114 (N_29114,N_26949,N_26468);
and U29115 (N_29115,N_26379,N_26667);
nor U29116 (N_29116,N_26648,N_27968);
nor U29117 (N_29117,N_26838,N_26087);
nor U29118 (N_29118,N_26765,N_27971);
nand U29119 (N_29119,N_27063,N_27171);
and U29120 (N_29120,N_27426,N_26983);
nand U29121 (N_29121,N_27656,N_27058);
or U29122 (N_29122,N_27333,N_27020);
and U29123 (N_29123,N_27562,N_27049);
and U29124 (N_29124,N_27291,N_27778);
nor U29125 (N_29125,N_26273,N_27873);
and U29126 (N_29126,N_26822,N_27588);
and U29127 (N_29127,N_27240,N_26853);
and U29128 (N_29128,N_27553,N_26398);
and U29129 (N_29129,N_26983,N_26130);
or U29130 (N_29130,N_26045,N_26066);
and U29131 (N_29131,N_26764,N_26471);
nor U29132 (N_29132,N_26181,N_27270);
and U29133 (N_29133,N_27245,N_26230);
xor U29134 (N_29134,N_26302,N_27906);
nand U29135 (N_29135,N_27346,N_26167);
or U29136 (N_29136,N_27825,N_26489);
or U29137 (N_29137,N_27837,N_26966);
and U29138 (N_29138,N_26903,N_26225);
and U29139 (N_29139,N_27764,N_27524);
xor U29140 (N_29140,N_26937,N_26461);
nand U29141 (N_29141,N_26772,N_27814);
and U29142 (N_29142,N_26529,N_26440);
and U29143 (N_29143,N_27019,N_27710);
nor U29144 (N_29144,N_27699,N_27475);
nor U29145 (N_29145,N_26407,N_27078);
xor U29146 (N_29146,N_27676,N_26842);
nor U29147 (N_29147,N_26491,N_26661);
xor U29148 (N_29148,N_26604,N_27078);
nand U29149 (N_29149,N_27122,N_27149);
nand U29150 (N_29150,N_26954,N_27202);
nand U29151 (N_29151,N_27709,N_27956);
xor U29152 (N_29152,N_27842,N_26374);
nand U29153 (N_29153,N_27203,N_27670);
and U29154 (N_29154,N_27436,N_27973);
and U29155 (N_29155,N_26530,N_27084);
nor U29156 (N_29156,N_26113,N_27762);
or U29157 (N_29157,N_27366,N_26897);
or U29158 (N_29158,N_27036,N_26612);
or U29159 (N_29159,N_27620,N_27750);
and U29160 (N_29160,N_26067,N_26271);
nor U29161 (N_29161,N_27830,N_27308);
nor U29162 (N_29162,N_26298,N_27993);
or U29163 (N_29163,N_26949,N_27553);
xor U29164 (N_29164,N_26801,N_26469);
and U29165 (N_29165,N_26198,N_27313);
xnor U29166 (N_29166,N_26698,N_26902);
or U29167 (N_29167,N_26679,N_27827);
or U29168 (N_29168,N_27467,N_26740);
or U29169 (N_29169,N_26249,N_27796);
and U29170 (N_29170,N_26933,N_27102);
and U29171 (N_29171,N_27327,N_26937);
xnor U29172 (N_29172,N_26875,N_27329);
xor U29173 (N_29173,N_26005,N_26903);
nand U29174 (N_29174,N_27805,N_26284);
nand U29175 (N_29175,N_27500,N_26713);
xnor U29176 (N_29176,N_26101,N_26912);
xor U29177 (N_29177,N_26841,N_27826);
nand U29178 (N_29178,N_26940,N_27789);
and U29179 (N_29179,N_27976,N_27158);
or U29180 (N_29180,N_26160,N_27870);
xnor U29181 (N_29181,N_27281,N_27426);
nor U29182 (N_29182,N_26378,N_26179);
nor U29183 (N_29183,N_26894,N_26915);
nor U29184 (N_29184,N_27646,N_27364);
nand U29185 (N_29185,N_27081,N_26969);
or U29186 (N_29186,N_27731,N_26180);
nand U29187 (N_29187,N_26623,N_26660);
and U29188 (N_29188,N_26174,N_27658);
nor U29189 (N_29189,N_27908,N_26749);
xnor U29190 (N_29190,N_27570,N_26613);
xnor U29191 (N_29191,N_26620,N_27208);
xor U29192 (N_29192,N_26770,N_27234);
nor U29193 (N_29193,N_27756,N_26473);
nor U29194 (N_29194,N_26209,N_26864);
nor U29195 (N_29195,N_27595,N_26787);
nand U29196 (N_29196,N_26000,N_27921);
or U29197 (N_29197,N_26530,N_27200);
nand U29198 (N_29198,N_27659,N_26117);
and U29199 (N_29199,N_26442,N_26299);
xnor U29200 (N_29200,N_26004,N_26258);
and U29201 (N_29201,N_27504,N_27104);
nand U29202 (N_29202,N_26984,N_26779);
or U29203 (N_29203,N_27415,N_27476);
and U29204 (N_29204,N_26722,N_26078);
and U29205 (N_29205,N_27326,N_27028);
nand U29206 (N_29206,N_27944,N_26005);
nand U29207 (N_29207,N_26890,N_26113);
or U29208 (N_29208,N_26351,N_26433);
nand U29209 (N_29209,N_26651,N_27296);
nor U29210 (N_29210,N_27761,N_26522);
and U29211 (N_29211,N_27954,N_27714);
xor U29212 (N_29212,N_26606,N_27721);
or U29213 (N_29213,N_26560,N_27010);
nand U29214 (N_29214,N_27280,N_26578);
nand U29215 (N_29215,N_26378,N_26307);
xor U29216 (N_29216,N_27547,N_26993);
xor U29217 (N_29217,N_26982,N_26950);
nor U29218 (N_29218,N_26682,N_26808);
and U29219 (N_29219,N_27813,N_26895);
nand U29220 (N_29220,N_26349,N_27643);
nor U29221 (N_29221,N_26410,N_26458);
xnor U29222 (N_29222,N_27444,N_26867);
nand U29223 (N_29223,N_27595,N_26577);
and U29224 (N_29224,N_26932,N_26851);
nor U29225 (N_29225,N_27692,N_26215);
xor U29226 (N_29226,N_27986,N_26015);
xor U29227 (N_29227,N_27703,N_27069);
and U29228 (N_29228,N_27872,N_26727);
nand U29229 (N_29229,N_26897,N_27238);
xor U29230 (N_29230,N_26509,N_26635);
or U29231 (N_29231,N_27986,N_27636);
xor U29232 (N_29232,N_26971,N_26795);
nor U29233 (N_29233,N_27111,N_27483);
and U29234 (N_29234,N_26396,N_26107);
xnor U29235 (N_29235,N_26330,N_27597);
nor U29236 (N_29236,N_27672,N_27616);
xor U29237 (N_29237,N_27004,N_27316);
nor U29238 (N_29238,N_26416,N_27739);
and U29239 (N_29239,N_26872,N_26452);
and U29240 (N_29240,N_26412,N_27237);
and U29241 (N_29241,N_26086,N_26405);
nand U29242 (N_29242,N_27739,N_26744);
nor U29243 (N_29243,N_26336,N_26871);
nor U29244 (N_29244,N_26836,N_26812);
or U29245 (N_29245,N_26212,N_26764);
nand U29246 (N_29246,N_26474,N_27898);
nor U29247 (N_29247,N_27382,N_27146);
or U29248 (N_29248,N_27992,N_26516);
nor U29249 (N_29249,N_27376,N_27508);
or U29250 (N_29250,N_27437,N_27036);
and U29251 (N_29251,N_27650,N_26632);
nand U29252 (N_29252,N_26565,N_26308);
and U29253 (N_29253,N_27736,N_26302);
and U29254 (N_29254,N_27609,N_26717);
nand U29255 (N_29255,N_27464,N_27475);
xor U29256 (N_29256,N_26727,N_26084);
xor U29257 (N_29257,N_27493,N_26216);
and U29258 (N_29258,N_27560,N_26156);
xor U29259 (N_29259,N_26542,N_26324);
xnor U29260 (N_29260,N_26682,N_26746);
or U29261 (N_29261,N_26992,N_26585);
nor U29262 (N_29262,N_27608,N_27075);
and U29263 (N_29263,N_27335,N_26545);
xor U29264 (N_29264,N_27918,N_26187);
nand U29265 (N_29265,N_26020,N_27175);
xnor U29266 (N_29266,N_27577,N_26395);
xor U29267 (N_29267,N_27058,N_26446);
or U29268 (N_29268,N_27348,N_26812);
xnor U29269 (N_29269,N_27984,N_27632);
or U29270 (N_29270,N_26201,N_26031);
xnor U29271 (N_29271,N_27826,N_26545);
or U29272 (N_29272,N_26943,N_26567);
nand U29273 (N_29273,N_27653,N_27094);
nand U29274 (N_29274,N_27795,N_26265);
and U29275 (N_29275,N_27408,N_27536);
nand U29276 (N_29276,N_26048,N_26532);
nor U29277 (N_29277,N_27677,N_26249);
and U29278 (N_29278,N_27802,N_26537);
xor U29279 (N_29279,N_26334,N_26492);
or U29280 (N_29280,N_26614,N_26003);
and U29281 (N_29281,N_27798,N_27578);
nand U29282 (N_29282,N_26220,N_27694);
and U29283 (N_29283,N_27778,N_26951);
nor U29284 (N_29284,N_26027,N_26014);
and U29285 (N_29285,N_27448,N_27558);
nor U29286 (N_29286,N_27784,N_26236);
nor U29287 (N_29287,N_27630,N_26910);
and U29288 (N_29288,N_26257,N_27348);
and U29289 (N_29289,N_27842,N_27989);
nor U29290 (N_29290,N_26776,N_27299);
or U29291 (N_29291,N_26017,N_26610);
nor U29292 (N_29292,N_26508,N_27024);
or U29293 (N_29293,N_26010,N_26892);
xor U29294 (N_29294,N_27321,N_26673);
nor U29295 (N_29295,N_26235,N_27927);
nor U29296 (N_29296,N_27540,N_27716);
and U29297 (N_29297,N_27598,N_26090);
and U29298 (N_29298,N_26906,N_26644);
and U29299 (N_29299,N_27129,N_26840);
and U29300 (N_29300,N_27304,N_26658);
nand U29301 (N_29301,N_26569,N_27324);
xor U29302 (N_29302,N_26645,N_27441);
nand U29303 (N_29303,N_27977,N_26718);
nor U29304 (N_29304,N_26672,N_27426);
or U29305 (N_29305,N_27682,N_27774);
xor U29306 (N_29306,N_27525,N_27086);
or U29307 (N_29307,N_27485,N_27351);
or U29308 (N_29308,N_27575,N_27279);
or U29309 (N_29309,N_26962,N_27356);
nor U29310 (N_29310,N_27035,N_27564);
nor U29311 (N_29311,N_27092,N_27655);
or U29312 (N_29312,N_26227,N_26907);
xnor U29313 (N_29313,N_26446,N_27306);
nand U29314 (N_29314,N_26049,N_27371);
and U29315 (N_29315,N_26813,N_27963);
or U29316 (N_29316,N_26237,N_26798);
nand U29317 (N_29317,N_26078,N_27403);
nand U29318 (N_29318,N_26991,N_27257);
nor U29319 (N_29319,N_26186,N_26374);
or U29320 (N_29320,N_27279,N_27876);
nand U29321 (N_29321,N_26610,N_26656);
and U29322 (N_29322,N_26632,N_27658);
xnor U29323 (N_29323,N_27193,N_26542);
xnor U29324 (N_29324,N_27641,N_26321);
and U29325 (N_29325,N_26791,N_26337);
xnor U29326 (N_29326,N_26615,N_26256);
or U29327 (N_29327,N_26951,N_27378);
nand U29328 (N_29328,N_26631,N_26991);
and U29329 (N_29329,N_27959,N_27209);
or U29330 (N_29330,N_26069,N_27433);
or U29331 (N_29331,N_27069,N_27496);
nand U29332 (N_29332,N_26691,N_27050);
xor U29333 (N_29333,N_27873,N_27560);
xor U29334 (N_29334,N_27185,N_26874);
nand U29335 (N_29335,N_27621,N_27183);
or U29336 (N_29336,N_27499,N_26292);
and U29337 (N_29337,N_26734,N_27013);
and U29338 (N_29338,N_27031,N_27215);
xor U29339 (N_29339,N_26091,N_26347);
xor U29340 (N_29340,N_26301,N_26364);
or U29341 (N_29341,N_26844,N_26093);
and U29342 (N_29342,N_27350,N_26051);
xnor U29343 (N_29343,N_27768,N_26424);
nor U29344 (N_29344,N_26604,N_27414);
or U29345 (N_29345,N_26113,N_27295);
or U29346 (N_29346,N_26375,N_26268);
xnor U29347 (N_29347,N_26100,N_26031);
or U29348 (N_29348,N_27189,N_26516);
and U29349 (N_29349,N_26939,N_26632);
nor U29350 (N_29350,N_27633,N_27193);
or U29351 (N_29351,N_26526,N_27481);
xor U29352 (N_29352,N_26439,N_26118);
xnor U29353 (N_29353,N_27246,N_27720);
and U29354 (N_29354,N_26099,N_27474);
nand U29355 (N_29355,N_27983,N_27908);
and U29356 (N_29356,N_26523,N_26761);
nand U29357 (N_29357,N_26280,N_27796);
nand U29358 (N_29358,N_27567,N_27243);
nor U29359 (N_29359,N_26954,N_26996);
and U29360 (N_29360,N_26172,N_27224);
or U29361 (N_29361,N_26863,N_26728);
or U29362 (N_29362,N_27729,N_26816);
nand U29363 (N_29363,N_26678,N_26851);
nand U29364 (N_29364,N_27036,N_26296);
nor U29365 (N_29365,N_27374,N_26659);
nand U29366 (N_29366,N_27307,N_27650);
or U29367 (N_29367,N_26785,N_27422);
nor U29368 (N_29368,N_27526,N_26311);
xor U29369 (N_29369,N_26602,N_27191);
nand U29370 (N_29370,N_26732,N_26309);
xor U29371 (N_29371,N_27714,N_27350);
nor U29372 (N_29372,N_26343,N_27172);
xor U29373 (N_29373,N_26534,N_27701);
nor U29374 (N_29374,N_26579,N_27505);
and U29375 (N_29375,N_27707,N_26965);
nand U29376 (N_29376,N_26334,N_27221);
nand U29377 (N_29377,N_26660,N_27344);
nand U29378 (N_29378,N_26562,N_27000);
or U29379 (N_29379,N_26805,N_26849);
nor U29380 (N_29380,N_27132,N_26396);
xor U29381 (N_29381,N_26187,N_26527);
and U29382 (N_29382,N_27783,N_27427);
or U29383 (N_29383,N_26619,N_27533);
nand U29384 (N_29384,N_27490,N_27600);
nand U29385 (N_29385,N_26192,N_26919);
or U29386 (N_29386,N_26346,N_27321);
or U29387 (N_29387,N_27546,N_26025);
nand U29388 (N_29388,N_26457,N_26600);
or U29389 (N_29389,N_27854,N_27301);
nand U29390 (N_29390,N_26010,N_26695);
or U29391 (N_29391,N_27143,N_27222);
nor U29392 (N_29392,N_27717,N_27443);
and U29393 (N_29393,N_27388,N_27271);
and U29394 (N_29394,N_26914,N_27543);
xor U29395 (N_29395,N_27582,N_26834);
nor U29396 (N_29396,N_27351,N_26886);
nor U29397 (N_29397,N_27245,N_27410);
or U29398 (N_29398,N_26519,N_27990);
and U29399 (N_29399,N_27227,N_27811);
nand U29400 (N_29400,N_27187,N_26274);
nor U29401 (N_29401,N_27686,N_26538);
nand U29402 (N_29402,N_27006,N_26684);
and U29403 (N_29403,N_27855,N_27283);
nor U29404 (N_29404,N_26642,N_26690);
xnor U29405 (N_29405,N_26520,N_27022);
nand U29406 (N_29406,N_27019,N_27435);
nand U29407 (N_29407,N_26139,N_26325);
xnor U29408 (N_29408,N_26461,N_27641);
nand U29409 (N_29409,N_26635,N_27502);
or U29410 (N_29410,N_26559,N_26788);
nor U29411 (N_29411,N_26068,N_26024);
nand U29412 (N_29412,N_27413,N_26657);
and U29413 (N_29413,N_27353,N_26037);
and U29414 (N_29414,N_27131,N_27063);
nor U29415 (N_29415,N_26690,N_26203);
or U29416 (N_29416,N_27554,N_26491);
or U29417 (N_29417,N_26537,N_27181);
xor U29418 (N_29418,N_27947,N_26095);
nand U29419 (N_29419,N_27896,N_26856);
and U29420 (N_29420,N_26007,N_26525);
and U29421 (N_29421,N_26781,N_26032);
nor U29422 (N_29422,N_26660,N_26211);
and U29423 (N_29423,N_26378,N_26578);
and U29424 (N_29424,N_26955,N_27986);
or U29425 (N_29425,N_27514,N_27360);
or U29426 (N_29426,N_26736,N_26336);
and U29427 (N_29427,N_27612,N_26125);
nor U29428 (N_29428,N_26808,N_27404);
nand U29429 (N_29429,N_26187,N_26661);
and U29430 (N_29430,N_26962,N_26801);
nand U29431 (N_29431,N_27979,N_27902);
xnor U29432 (N_29432,N_26948,N_26305);
and U29433 (N_29433,N_26904,N_26465);
nand U29434 (N_29434,N_27176,N_27348);
nand U29435 (N_29435,N_26886,N_26456);
nor U29436 (N_29436,N_27148,N_26535);
xnor U29437 (N_29437,N_26871,N_26785);
nor U29438 (N_29438,N_27525,N_27773);
nor U29439 (N_29439,N_27127,N_27472);
nand U29440 (N_29440,N_26069,N_26711);
xnor U29441 (N_29441,N_27559,N_27475);
nand U29442 (N_29442,N_26578,N_27139);
nor U29443 (N_29443,N_26486,N_27419);
xnor U29444 (N_29444,N_26227,N_27302);
and U29445 (N_29445,N_27692,N_26742);
nand U29446 (N_29446,N_27070,N_26884);
nor U29447 (N_29447,N_26420,N_26937);
nor U29448 (N_29448,N_27114,N_27365);
nor U29449 (N_29449,N_27405,N_26086);
or U29450 (N_29450,N_27144,N_26385);
and U29451 (N_29451,N_27495,N_27687);
nor U29452 (N_29452,N_26253,N_26252);
nand U29453 (N_29453,N_26334,N_27200);
or U29454 (N_29454,N_26248,N_27676);
nand U29455 (N_29455,N_27482,N_27749);
xnor U29456 (N_29456,N_27609,N_27517);
and U29457 (N_29457,N_26823,N_27906);
xor U29458 (N_29458,N_26926,N_26736);
nand U29459 (N_29459,N_26450,N_26233);
xor U29460 (N_29460,N_27833,N_27038);
nand U29461 (N_29461,N_26848,N_26728);
xor U29462 (N_29462,N_27701,N_26181);
nand U29463 (N_29463,N_26015,N_26048);
or U29464 (N_29464,N_27426,N_26506);
nand U29465 (N_29465,N_27809,N_26412);
nor U29466 (N_29466,N_26171,N_26010);
nand U29467 (N_29467,N_26049,N_27235);
and U29468 (N_29468,N_27280,N_26966);
nor U29469 (N_29469,N_26289,N_27091);
and U29470 (N_29470,N_27714,N_26745);
and U29471 (N_29471,N_27042,N_27924);
nor U29472 (N_29472,N_26380,N_26746);
nand U29473 (N_29473,N_26578,N_26630);
or U29474 (N_29474,N_27932,N_26753);
xnor U29475 (N_29475,N_27735,N_27154);
xor U29476 (N_29476,N_27583,N_26769);
and U29477 (N_29477,N_27111,N_27043);
xnor U29478 (N_29478,N_26626,N_27139);
or U29479 (N_29479,N_26766,N_27947);
and U29480 (N_29480,N_27572,N_26722);
nand U29481 (N_29481,N_27726,N_26471);
nor U29482 (N_29482,N_26084,N_26896);
and U29483 (N_29483,N_27069,N_27980);
xnor U29484 (N_29484,N_27799,N_27035);
nand U29485 (N_29485,N_27150,N_27072);
nor U29486 (N_29486,N_27071,N_27544);
or U29487 (N_29487,N_26706,N_26484);
nand U29488 (N_29488,N_27817,N_27221);
nor U29489 (N_29489,N_26790,N_26737);
or U29490 (N_29490,N_26914,N_27612);
xnor U29491 (N_29491,N_27913,N_26569);
xnor U29492 (N_29492,N_27391,N_26797);
xnor U29493 (N_29493,N_27549,N_26632);
nand U29494 (N_29494,N_26096,N_27291);
and U29495 (N_29495,N_27309,N_26418);
nand U29496 (N_29496,N_27308,N_26636);
or U29497 (N_29497,N_27819,N_27448);
and U29498 (N_29498,N_26932,N_27814);
and U29499 (N_29499,N_27476,N_27286);
nor U29500 (N_29500,N_27451,N_26817);
nor U29501 (N_29501,N_27974,N_27692);
and U29502 (N_29502,N_27934,N_26050);
and U29503 (N_29503,N_27184,N_26235);
and U29504 (N_29504,N_27190,N_27904);
xor U29505 (N_29505,N_26370,N_27786);
nor U29506 (N_29506,N_27716,N_26286);
and U29507 (N_29507,N_27298,N_26271);
and U29508 (N_29508,N_27375,N_26462);
xor U29509 (N_29509,N_26460,N_26632);
or U29510 (N_29510,N_27611,N_26815);
nor U29511 (N_29511,N_27329,N_26742);
nand U29512 (N_29512,N_26284,N_26925);
nand U29513 (N_29513,N_26547,N_26711);
xnor U29514 (N_29514,N_26944,N_27525);
nand U29515 (N_29515,N_27658,N_26425);
xnor U29516 (N_29516,N_26546,N_27059);
nand U29517 (N_29517,N_27844,N_27194);
nand U29518 (N_29518,N_26611,N_27049);
nor U29519 (N_29519,N_26548,N_27564);
xor U29520 (N_29520,N_26323,N_26003);
nand U29521 (N_29521,N_27224,N_26909);
and U29522 (N_29522,N_26895,N_26471);
and U29523 (N_29523,N_27566,N_26009);
xor U29524 (N_29524,N_27120,N_26564);
nor U29525 (N_29525,N_26289,N_27462);
or U29526 (N_29526,N_27457,N_26422);
xnor U29527 (N_29527,N_27611,N_27251);
or U29528 (N_29528,N_26946,N_26321);
or U29529 (N_29529,N_26263,N_26930);
and U29530 (N_29530,N_27573,N_27307);
nand U29531 (N_29531,N_26473,N_27558);
nor U29532 (N_29532,N_27117,N_26260);
nand U29533 (N_29533,N_26977,N_26897);
or U29534 (N_29534,N_26998,N_26220);
nor U29535 (N_29535,N_26692,N_26754);
xnor U29536 (N_29536,N_27038,N_27899);
and U29537 (N_29537,N_27799,N_26523);
and U29538 (N_29538,N_26317,N_27072);
and U29539 (N_29539,N_26225,N_26412);
nor U29540 (N_29540,N_27784,N_26052);
xor U29541 (N_29541,N_27412,N_27839);
nand U29542 (N_29542,N_26721,N_27865);
xor U29543 (N_29543,N_26871,N_27963);
xor U29544 (N_29544,N_26825,N_27561);
nor U29545 (N_29545,N_27323,N_26800);
and U29546 (N_29546,N_27919,N_26469);
or U29547 (N_29547,N_27900,N_26415);
or U29548 (N_29548,N_26865,N_26858);
xor U29549 (N_29549,N_27539,N_27885);
and U29550 (N_29550,N_27800,N_26388);
xnor U29551 (N_29551,N_27217,N_26742);
xor U29552 (N_29552,N_26833,N_27727);
xor U29553 (N_29553,N_27415,N_26765);
xnor U29554 (N_29554,N_27023,N_26884);
nand U29555 (N_29555,N_26052,N_27974);
and U29556 (N_29556,N_27988,N_27372);
nor U29557 (N_29557,N_26981,N_26743);
nor U29558 (N_29558,N_27746,N_26362);
xor U29559 (N_29559,N_27008,N_26326);
nor U29560 (N_29560,N_26118,N_26960);
xor U29561 (N_29561,N_27894,N_27130);
nor U29562 (N_29562,N_26380,N_26083);
xnor U29563 (N_29563,N_27589,N_26964);
or U29564 (N_29564,N_27408,N_26207);
nand U29565 (N_29565,N_27885,N_26029);
or U29566 (N_29566,N_27933,N_26044);
and U29567 (N_29567,N_26773,N_27377);
nor U29568 (N_29568,N_26666,N_26406);
nand U29569 (N_29569,N_27208,N_27528);
nor U29570 (N_29570,N_27377,N_27916);
nand U29571 (N_29571,N_27346,N_26999);
nor U29572 (N_29572,N_27828,N_27530);
xor U29573 (N_29573,N_26573,N_26332);
or U29574 (N_29574,N_26229,N_27994);
or U29575 (N_29575,N_27888,N_26455);
nand U29576 (N_29576,N_27330,N_27695);
and U29577 (N_29577,N_27268,N_26630);
xor U29578 (N_29578,N_27234,N_26577);
nand U29579 (N_29579,N_26003,N_27682);
and U29580 (N_29580,N_26429,N_27902);
and U29581 (N_29581,N_27338,N_26372);
nand U29582 (N_29582,N_27061,N_26302);
and U29583 (N_29583,N_27269,N_27016);
and U29584 (N_29584,N_26172,N_26555);
nand U29585 (N_29585,N_26290,N_26694);
and U29586 (N_29586,N_26819,N_27122);
and U29587 (N_29587,N_27773,N_27036);
nor U29588 (N_29588,N_27151,N_26736);
nor U29589 (N_29589,N_27309,N_27002);
xnor U29590 (N_29590,N_26971,N_27787);
and U29591 (N_29591,N_26573,N_27277);
nand U29592 (N_29592,N_26289,N_27241);
xnor U29593 (N_29593,N_26092,N_26299);
or U29594 (N_29594,N_27076,N_26753);
nor U29595 (N_29595,N_26596,N_27057);
and U29596 (N_29596,N_26080,N_27220);
or U29597 (N_29597,N_27448,N_27035);
nor U29598 (N_29598,N_26850,N_26582);
and U29599 (N_29599,N_27490,N_26458);
nor U29600 (N_29600,N_27657,N_26116);
and U29601 (N_29601,N_26149,N_27788);
and U29602 (N_29602,N_27799,N_27237);
nor U29603 (N_29603,N_26503,N_26676);
nand U29604 (N_29604,N_26625,N_27205);
xnor U29605 (N_29605,N_26556,N_27694);
nor U29606 (N_29606,N_26754,N_27186);
and U29607 (N_29607,N_26989,N_27086);
xnor U29608 (N_29608,N_26214,N_27748);
and U29609 (N_29609,N_26119,N_26487);
and U29610 (N_29610,N_27852,N_26459);
and U29611 (N_29611,N_26470,N_27866);
and U29612 (N_29612,N_27197,N_26279);
nor U29613 (N_29613,N_27898,N_27697);
and U29614 (N_29614,N_26553,N_27521);
nand U29615 (N_29615,N_26830,N_26380);
and U29616 (N_29616,N_26950,N_26898);
and U29617 (N_29617,N_27802,N_27315);
nor U29618 (N_29618,N_26578,N_27682);
nor U29619 (N_29619,N_27476,N_26984);
and U29620 (N_29620,N_27187,N_27410);
xnor U29621 (N_29621,N_26498,N_26904);
nand U29622 (N_29622,N_27636,N_27134);
nand U29623 (N_29623,N_27517,N_27146);
nor U29624 (N_29624,N_26902,N_27174);
nor U29625 (N_29625,N_26334,N_27540);
nand U29626 (N_29626,N_27251,N_26723);
nor U29627 (N_29627,N_27834,N_27886);
or U29628 (N_29628,N_26454,N_26748);
or U29629 (N_29629,N_26130,N_27887);
nand U29630 (N_29630,N_27660,N_27108);
and U29631 (N_29631,N_26083,N_26779);
and U29632 (N_29632,N_26199,N_26108);
nor U29633 (N_29633,N_26654,N_26730);
and U29634 (N_29634,N_27190,N_26719);
nor U29635 (N_29635,N_26907,N_26905);
or U29636 (N_29636,N_26883,N_27149);
or U29637 (N_29637,N_27014,N_26039);
nand U29638 (N_29638,N_26111,N_26852);
and U29639 (N_29639,N_26983,N_26299);
and U29640 (N_29640,N_26536,N_26959);
and U29641 (N_29641,N_26806,N_26206);
and U29642 (N_29642,N_26261,N_26773);
and U29643 (N_29643,N_26820,N_27588);
nand U29644 (N_29644,N_26342,N_26877);
xor U29645 (N_29645,N_27060,N_26340);
nand U29646 (N_29646,N_27039,N_26364);
nand U29647 (N_29647,N_26464,N_26783);
nor U29648 (N_29648,N_26241,N_27299);
and U29649 (N_29649,N_26643,N_26276);
nor U29650 (N_29650,N_26103,N_26948);
xor U29651 (N_29651,N_27779,N_27163);
and U29652 (N_29652,N_26827,N_26950);
or U29653 (N_29653,N_26631,N_26026);
or U29654 (N_29654,N_27588,N_27655);
nand U29655 (N_29655,N_26402,N_27499);
and U29656 (N_29656,N_27698,N_27004);
and U29657 (N_29657,N_27774,N_27978);
nor U29658 (N_29658,N_26917,N_27628);
or U29659 (N_29659,N_26184,N_27439);
or U29660 (N_29660,N_26204,N_26352);
or U29661 (N_29661,N_26945,N_27319);
nand U29662 (N_29662,N_26733,N_26392);
nand U29663 (N_29663,N_26144,N_26744);
nand U29664 (N_29664,N_26352,N_27769);
nor U29665 (N_29665,N_27964,N_26329);
or U29666 (N_29666,N_27685,N_27244);
xor U29667 (N_29667,N_26657,N_26157);
nor U29668 (N_29668,N_27390,N_26517);
nand U29669 (N_29669,N_27623,N_27956);
and U29670 (N_29670,N_27399,N_26869);
nand U29671 (N_29671,N_26857,N_26963);
and U29672 (N_29672,N_27571,N_27910);
or U29673 (N_29673,N_27943,N_26138);
xor U29674 (N_29674,N_26978,N_26993);
or U29675 (N_29675,N_26992,N_27856);
and U29676 (N_29676,N_26257,N_26058);
nor U29677 (N_29677,N_27673,N_26713);
nor U29678 (N_29678,N_27855,N_27415);
or U29679 (N_29679,N_26463,N_27378);
xnor U29680 (N_29680,N_26378,N_26997);
or U29681 (N_29681,N_26701,N_26480);
xnor U29682 (N_29682,N_27329,N_27477);
nand U29683 (N_29683,N_26226,N_27480);
or U29684 (N_29684,N_26514,N_26723);
nor U29685 (N_29685,N_26547,N_26707);
and U29686 (N_29686,N_27679,N_26974);
xnor U29687 (N_29687,N_27152,N_26616);
nand U29688 (N_29688,N_27097,N_27370);
nor U29689 (N_29689,N_26504,N_27679);
and U29690 (N_29690,N_26485,N_26879);
nand U29691 (N_29691,N_27494,N_26652);
nor U29692 (N_29692,N_26975,N_27839);
nor U29693 (N_29693,N_26317,N_26084);
nor U29694 (N_29694,N_27033,N_26916);
xor U29695 (N_29695,N_26156,N_27832);
or U29696 (N_29696,N_26744,N_27660);
nand U29697 (N_29697,N_27522,N_26397);
or U29698 (N_29698,N_27608,N_27033);
or U29699 (N_29699,N_26171,N_26644);
nor U29700 (N_29700,N_26787,N_27307);
or U29701 (N_29701,N_26816,N_26219);
or U29702 (N_29702,N_26933,N_26489);
or U29703 (N_29703,N_27417,N_26008);
or U29704 (N_29704,N_27386,N_27239);
or U29705 (N_29705,N_27137,N_26705);
nand U29706 (N_29706,N_26936,N_26922);
or U29707 (N_29707,N_26664,N_26851);
nor U29708 (N_29708,N_27828,N_27248);
and U29709 (N_29709,N_27612,N_26729);
or U29710 (N_29710,N_26612,N_26462);
nor U29711 (N_29711,N_27474,N_27084);
xor U29712 (N_29712,N_26666,N_27882);
nand U29713 (N_29713,N_27915,N_26326);
xnor U29714 (N_29714,N_27524,N_27791);
nand U29715 (N_29715,N_27196,N_26591);
nand U29716 (N_29716,N_27003,N_26402);
or U29717 (N_29717,N_26796,N_26616);
xnor U29718 (N_29718,N_27853,N_26767);
xnor U29719 (N_29719,N_26431,N_26815);
xor U29720 (N_29720,N_26945,N_26305);
or U29721 (N_29721,N_26443,N_27790);
xor U29722 (N_29722,N_26751,N_27030);
xnor U29723 (N_29723,N_26406,N_27098);
xor U29724 (N_29724,N_27073,N_27927);
xnor U29725 (N_29725,N_26888,N_26796);
nand U29726 (N_29726,N_27311,N_27554);
or U29727 (N_29727,N_26453,N_26059);
or U29728 (N_29728,N_27747,N_27340);
and U29729 (N_29729,N_26884,N_27063);
nor U29730 (N_29730,N_27049,N_27906);
xnor U29731 (N_29731,N_26182,N_27471);
nor U29732 (N_29732,N_26578,N_27389);
and U29733 (N_29733,N_26487,N_26144);
and U29734 (N_29734,N_26958,N_27861);
and U29735 (N_29735,N_26680,N_27720);
nor U29736 (N_29736,N_26629,N_27747);
nand U29737 (N_29737,N_26838,N_26289);
xor U29738 (N_29738,N_26182,N_27352);
and U29739 (N_29739,N_27473,N_27167);
xnor U29740 (N_29740,N_26324,N_27937);
or U29741 (N_29741,N_27563,N_26058);
and U29742 (N_29742,N_27928,N_27358);
nand U29743 (N_29743,N_27830,N_27426);
or U29744 (N_29744,N_27721,N_27379);
nor U29745 (N_29745,N_27417,N_26666);
and U29746 (N_29746,N_27560,N_27966);
nand U29747 (N_29747,N_26555,N_26457);
nand U29748 (N_29748,N_27616,N_27957);
nor U29749 (N_29749,N_27653,N_26745);
nand U29750 (N_29750,N_26860,N_26814);
nand U29751 (N_29751,N_26802,N_27069);
nand U29752 (N_29752,N_27886,N_27079);
and U29753 (N_29753,N_26941,N_27716);
nand U29754 (N_29754,N_26187,N_27263);
nand U29755 (N_29755,N_26811,N_26031);
nor U29756 (N_29756,N_27408,N_26374);
or U29757 (N_29757,N_27293,N_26998);
xnor U29758 (N_29758,N_26132,N_26771);
xor U29759 (N_29759,N_27782,N_26938);
xor U29760 (N_29760,N_27061,N_26056);
or U29761 (N_29761,N_27196,N_26081);
or U29762 (N_29762,N_27980,N_27872);
nor U29763 (N_29763,N_27283,N_26627);
xnor U29764 (N_29764,N_27403,N_26982);
or U29765 (N_29765,N_26409,N_27644);
or U29766 (N_29766,N_26362,N_26585);
nor U29767 (N_29767,N_27220,N_27388);
xnor U29768 (N_29768,N_26135,N_27371);
nor U29769 (N_29769,N_26603,N_26678);
nor U29770 (N_29770,N_26249,N_26763);
or U29771 (N_29771,N_27703,N_27762);
xnor U29772 (N_29772,N_27736,N_27076);
xnor U29773 (N_29773,N_27686,N_27974);
xnor U29774 (N_29774,N_26441,N_27183);
xor U29775 (N_29775,N_26865,N_27282);
nand U29776 (N_29776,N_27739,N_26179);
or U29777 (N_29777,N_26660,N_26100);
nand U29778 (N_29778,N_27430,N_27496);
and U29779 (N_29779,N_27134,N_26204);
xor U29780 (N_29780,N_26810,N_27105);
and U29781 (N_29781,N_27977,N_26107);
xor U29782 (N_29782,N_26101,N_27583);
xnor U29783 (N_29783,N_27099,N_27730);
nand U29784 (N_29784,N_26043,N_26308);
or U29785 (N_29785,N_27903,N_26595);
nand U29786 (N_29786,N_26804,N_26721);
nand U29787 (N_29787,N_26992,N_26924);
or U29788 (N_29788,N_27610,N_27490);
xnor U29789 (N_29789,N_27067,N_26245);
nand U29790 (N_29790,N_26127,N_26563);
nand U29791 (N_29791,N_26628,N_27697);
nand U29792 (N_29792,N_27996,N_26229);
or U29793 (N_29793,N_26603,N_27537);
xor U29794 (N_29794,N_26474,N_26051);
xor U29795 (N_29795,N_27025,N_27523);
nand U29796 (N_29796,N_26380,N_27054);
nor U29797 (N_29797,N_26467,N_27581);
nand U29798 (N_29798,N_27909,N_27534);
xor U29799 (N_29799,N_26272,N_27709);
or U29800 (N_29800,N_26326,N_27350);
or U29801 (N_29801,N_27018,N_26174);
or U29802 (N_29802,N_26282,N_27495);
nand U29803 (N_29803,N_26587,N_26120);
or U29804 (N_29804,N_26502,N_27639);
and U29805 (N_29805,N_27058,N_27352);
or U29806 (N_29806,N_26641,N_26488);
xor U29807 (N_29807,N_27661,N_27147);
nand U29808 (N_29808,N_27406,N_26785);
or U29809 (N_29809,N_26732,N_27033);
and U29810 (N_29810,N_27941,N_26527);
xnor U29811 (N_29811,N_27888,N_26625);
xor U29812 (N_29812,N_26531,N_27483);
nand U29813 (N_29813,N_27985,N_26879);
and U29814 (N_29814,N_27728,N_26130);
xnor U29815 (N_29815,N_27021,N_26440);
and U29816 (N_29816,N_26155,N_27085);
xnor U29817 (N_29817,N_26893,N_27353);
or U29818 (N_29818,N_27865,N_27997);
and U29819 (N_29819,N_27537,N_26112);
or U29820 (N_29820,N_27620,N_26183);
nand U29821 (N_29821,N_27904,N_27208);
nand U29822 (N_29822,N_27421,N_26553);
or U29823 (N_29823,N_26812,N_26949);
nor U29824 (N_29824,N_27117,N_26476);
xor U29825 (N_29825,N_26173,N_26348);
nor U29826 (N_29826,N_26207,N_27624);
or U29827 (N_29827,N_26602,N_26605);
and U29828 (N_29828,N_26752,N_26038);
and U29829 (N_29829,N_26633,N_26584);
xor U29830 (N_29830,N_27599,N_27659);
nand U29831 (N_29831,N_27210,N_26749);
xor U29832 (N_29832,N_26236,N_27026);
nand U29833 (N_29833,N_26764,N_27316);
nand U29834 (N_29834,N_27241,N_26367);
xor U29835 (N_29835,N_26246,N_27966);
nor U29836 (N_29836,N_26040,N_26164);
or U29837 (N_29837,N_27294,N_26720);
and U29838 (N_29838,N_27069,N_27488);
and U29839 (N_29839,N_27148,N_26443);
nor U29840 (N_29840,N_26416,N_27385);
xor U29841 (N_29841,N_26505,N_26572);
or U29842 (N_29842,N_26989,N_26301);
xor U29843 (N_29843,N_27295,N_26854);
or U29844 (N_29844,N_26484,N_26904);
nand U29845 (N_29845,N_26907,N_27549);
and U29846 (N_29846,N_26449,N_26346);
and U29847 (N_29847,N_26637,N_27621);
or U29848 (N_29848,N_26165,N_27573);
or U29849 (N_29849,N_26615,N_26653);
nand U29850 (N_29850,N_26628,N_27112);
and U29851 (N_29851,N_27268,N_27146);
xnor U29852 (N_29852,N_27615,N_26460);
xor U29853 (N_29853,N_27944,N_26930);
nand U29854 (N_29854,N_27924,N_26127);
and U29855 (N_29855,N_27007,N_27167);
or U29856 (N_29856,N_26753,N_27565);
xnor U29857 (N_29857,N_26236,N_26671);
or U29858 (N_29858,N_26438,N_27565);
nand U29859 (N_29859,N_26869,N_26489);
xor U29860 (N_29860,N_26021,N_27799);
xor U29861 (N_29861,N_26286,N_27028);
and U29862 (N_29862,N_27970,N_26533);
nand U29863 (N_29863,N_27191,N_27450);
or U29864 (N_29864,N_27409,N_27517);
nand U29865 (N_29865,N_26492,N_26566);
xor U29866 (N_29866,N_26409,N_26759);
or U29867 (N_29867,N_27928,N_26362);
nor U29868 (N_29868,N_27664,N_27052);
or U29869 (N_29869,N_27381,N_26819);
nor U29870 (N_29870,N_26381,N_27964);
nand U29871 (N_29871,N_27777,N_27435);
or U29872 (N_29872,N_26281,N_26589);
and U29873 (N_29873,N_26338,N_26481);
and U29874 (N_29874,N_26966,N_26458);
nand U29875 (N_29875,N_27306,N_27222);
xor U29876 (N_29876,N_27383,N_27877);
nor U29877 (N_29877,N_26395,N_27470);
nor U29878 (N_29878,N_27916,N_26973);
and U29879 (N_29879,N_26476,N_26824);
nand U29880 (N_29880,N_27172,N_26336);
or U29881 (N_29881,N_26343,N_26249);
nor U29882 (N_29882,N_26960,N_26046);
or U29883 (N_29883,N_27618,N_27785);
nand U29884 (N_29884,N_26596,N_27118);
nor U29885 (N_29885,N_27848,N_27056);
xnor U29886 (N_29886,N_27342,N_26222);
nor U29887 (N_29887,N_26728,N_26276);
and U29888 (N_29888,N_27164,N_27814);
nand U29889 (N_29889,N_26019,N_27722);
xnor U29890 (N_29890,N_26785,N_26901);
and U29891 (N_29891,N_27017,N_26773);
nor U29892 (N_29892,N_27086,N_27777);
and U29893 (N_29893,N_26084,N_27932);
xor U29894 (N_29894,N_27132,N_26415);
xnor U29895 (N_29895,N_26163,N_27266);
and U29896 (N_29896,N_27042,N_27295);
nand U29897 (N_29897,N_27425,N_27710);
or U29898 (N_29898,N_27094,N_26889);
xor U29899 (N_29899,N_26885,N_27825);
xnor U29900 (N_29900,N_26813,N_26820);
and U29901 (N_29901,N_26548,N_27168);
or U29902 (N_29902,N_27265,N_27108);
nor U29903 (N_29903,N_26007,N_27037);
nand U29904 (N_29904,N_26272,N_26003);
or U29905 (N_29905,N_26547,N_26689);
or U29906 (N_29906,N_26323,N_26031);
and U29907 (N_29907,N_26517,N_26913);
and U29908 (N_29908,N_27634,N_27467);
and U29909 (N_29909,N_26462,N_26395);
nand U29910 (N_29910,N_27467,N_27350);
nor U29911 (N_29911,N_27685,N_27425);
nor U29912 (N_29912,N_26765,N_26325);
and U29913 (N_29913,N_26264,N_27967);
nand U29914 (N_29914,N_26975,N_26314);
or U29915 (N_29915,N_26222,N_26885);
nor U29916 (N_29916,N_27437,N_26860);
xor U29917 (N_29917,N_26650,N_27537);
nand U29918 (N_29918,N_27985,N_26955);
or U29919 (N_29919,N_27316,N_27172);
and U29920 (N_29920,N_26394,N_26306);
nor U29921 (N_29921,N_27104,N_26325);
or U29922 (N_29922,N_27168,N_26461);
or U29923 (N_29923,N_26741,N_26204);
nand U29924 (N_29924,N_26283,N_26656);
xnor U29925 (N_29925,N_27919,N_26193);
or U29926 (N_29926,N_26448,N_26941);
or U29927 (N_29927,N_26969,N_26356);
nand U29928 (N_29928,N_27893,N_27838);
nand U29929 (N_29929,N_27653,N_27116);
or U29930 (N_29930,N_27878,N_26043);
or U29931 (N_29931,N_26937,N_26713);
nor U29932 (N_29932,N_26043,N_26885);
and U29933 (N_29933,N_26730,N_27455);
or U29934 (N_29934,N_26049,N_26862);
nand U29935 (N_29935,N_26976,N_26973);
nand U29936 (N_29936,N_27564,N_26367);
and U29937 (N_29937,N_26988,N_27451);
or U29938 (N_29938,N_26299,N_27459);
nor U29939 (N_29939,N_26505,N_26445);
and U29940 (N_29940,N_27258,N_27198);
or U29941 (N_29941,N_27588,N_27995);
nor U29942 (N_29942,N_27164,N_27664);
nand U29943 (N_29943,N_27024,N_27208);
or U29944 (N_29944,N_26505,N_27440);
nor U29945 (N_29945,N_26709,N_27047);
xnor U29946 (N_29946,N_27665,N_27374);
nand U29947 (N_29947,N_27739,N_27896);
xnor U29948 (N_29948,N_26445,N_27245);
and U29949 (N_29949,N_26959,N_26932);
nor U29950 (N_29950,N_26682,N_27447);
or U29951 (N_29951,N_27827,N_26850);
nand U29952 (N_29952,N_27906,N_27758);
nand U29953 (N_29953,N_27893,N_26216);
or U29954 (N_29954,N_27789,N_26522);
nor U29955 (N_29955,N_27740,N_26147);
and U29956 (N_29956,N_26903,N_26115);
or U29957 (N_29957,N_26488,N_27198);
and U29958 (N_29958,N_26213,N_26652);
and U29959 (N_29959,N_27808,N_26643);
nand U29960 (N_29960,N_27573,N_27039);
xnor U29961 (N_29961,N_26533,N_27597);
and U29962 (N_29962,N_27041,N_27091);
or U29963 (N_29963,N_27230,N_26395);
xor U29964 (N_29964,N_26331,N_26772);
and U29965 (N_29965,N_27055,N_26835);
nand U29966 (N_29966,N_26648,N_27736);
nand U29967 (N_29967,N_26991,N_27643);
xnor U29968 (N_29968,N_26096,N_26595);
and U29969 (N_29969,N_27872,N_27088);
or U29970 (N_29970,N_26303,N_27734);
nand U29971 (N_29971,N_27864,N_26582);
and U29972 (N_29972,N_27640,N_27184);
xor U29973 (N_29973,N_26614,N_27348);
and U29974 (N_29974,N_27429,N_26690);
and U29975 (N_29975,N_26842,N_27889);
nor U29976 (N_29976,N_27606,N_26649);
or U29977 (N_29977,N_27438,N_27792);
nor U29978 (N_29978,N_26379,N_27901);
nor U29979 (N_29979,N_26307,N_26687);
or U29980 (N_29980,N_27151,N_27442);
xnor U29981 (N_29981,N_26812,N_26341);
xnor U29982 (N_29982,N_26454,N_26199);
or U29983 (N_29983,N_27854,N_26573);
xnor U29984 (N_29984,N_27063,N_26010);
nor U29985 (N_29985,N_26620,N_26250);
or U29986 (N_29986,N_26694,N_26988);
nor U29987 (N_29987,N_26614,N_27555);
xnor U29988 (N_29988,N_27285,N_27617);
and U29989 (N_29989,N_26716,N_27124);
nor U29990 (N_29990,N_27166,N_27414);
xnor U29991 (N_29991,N_26802,N_26213);
nand U29992 (N_29992,N_27375,N_26311);
or U29993 (N_29993,N_26921,N_26901);
nor U29994 (N_29994,N_27685,N_27833);
and U29995 (N_29995,N_26884,N_27643);
or U29996 (N_29996,N_26733,N_26917);
nor U29997 (N_29997,N_27084,N_27705);
nand U29998 (N_29998,N_27688,N_26471);
xor U29999 (N_29999,N_27185,N_27949);
or U30000 (N_30000,N_28066,N_29098);
and U30001 (N_30001,N_28409,N_29773);
xnor U30002 (N_30002,N_29457,N_28114);
nand U30003 (N_30003,N_28273,N_28426);
xor U30004 (N_30004,N_29170,N_29000);
nand U30005 (N_30005,N_29958,N_29908);
or U30006 (N_30006,N_29453,N_29533);
or U30007 (N_30007,N_29735,N_29705);
or U30008 (N_30008,N_28124,N_29720);
and U30009 (N_30009,N_28744,N_29850);
and U30010 (N_30010,N_28282,N_29291);
or U30011 (N_30011,N_29848,N_29650);
or U30012 (N_30012,N_29346,N_28210);
nor U30013 (N_30013,N_28693,N_29407);
nor U30014 (N_30014,N_28177,N_28142);
xor U30015 (N_30015,N_28859,N_28002);
xnor U30016 (N_30016,N_29334,N_29825);
xor U30017 (N_30017,N_29587,N_29575);
nor U30018 (N_30018,N_28986,N_28216);
or U30019 (N_30019,N_29066,N_29903);
nor U30020 (N_30020,N_29838,N_28025);
xnor U30021 (N_30021,N_29294,N_28224);
xor U30022 (N_30022,N_28331,N_28886);
or U30023 (N_30023,N_29040,N_28536);
or U30024 (N_30024,N_29865,N_29785);
and U30025 (N_30025,N_29237,N_29555);
xnor U30026 (N_30026,N_28607,N_29123);
and U30027 (N_30027,N_28497,N_29916);
or U30028 (N_30028,N_29975,N_28975);
and U30029 (N_30029,N_29623,N_28213);
and U30030 (N_30030,N_29015,N_28288);
nand U30031 (N_30031,N_28326,N_28082);
nor U30032 (N_30032,N_29100,N_28593);
xor U30033 (N_30033,N_28814,N_28220);
nand U30034 (N_30034,N_28932,N_29350);
nand U30035 (N_30035,N_29444,N_29665);
nand U30036 (N_30036,N_28931,N_29791);
and U30037 (N_30037,N_28184,N_28881);
and U30038 (N_30038,N_29948,N_28329);
and U30039 (N_30039,N_29298,N_29034);
nor U30040 (N_30040,N_28261,N_29551);
xor U30041 (N_30041,N_29487,N_28334);
or U30042 (N_30042,N_28139,N_28543);
xor U30043 (N_30043,N_28992,N_28767);
nor U30044 (N_30044,N_28472,N_28550);
nor U30045 (N_30045,N_29120,N_28257);
nor U30046 (N_30046,N_29099,N_29065);
nand U30047 (N_30047,N_29780,N_29790);
xnor U30048 (N_30048,N_28447,N_29414);
and U30049 (N_30049,N_28519,N_28157);
xnor U30050 (N_30050,N_28839,N_28529);
nand U30051 (N_30051,N_29235,N_28999);
nand U30052 (N_30052,N_28285,N_28454);
or U30053 (N_30053,N_28908,N_28777);
or U30054 (N_30054,N_29523,N_29259);
nand U30055 (N_30055,N_28278,N_28978);
nor U30056 (N_30056,N_29658,N_29894);
or U30057 (N_30057,N_28422,N_29244);
xnor U30058 (N_30058,N_29549,N_29163);
xnor U30059 (N_30059,N_28858,N_29987);
xnor U30060 (N_30060,N_29499,N_28164);
or U30061 (N_30061,N_28949,N_29655);
nor U30062 (N_30062,N_28874,N_28463);
nor U30063 (N_30063,N_29546,N_29153);
nand U30064 (N_30064,N_28009,N_29342);
xnor U30065 (N_30065,N_29925,N_29620);
nand U30066 (N_30066,N_29101,N_29857);
nand U30067 (N_30067,N_29193,N_29363);
or U30068 (N_30068,N_29602,N_29915);
and U30069 (N_30069,N_29880,N_29969);
nand U30070 (N_30070,N_28465,N_28227);
nor U30071 (N_30071,N_29743,N_29030);
nor U30072 (N_30072,N_29608,N_29766);
nand U30073 (N_30073,N_29741,N_29370);
nand U30074 (N_30074,N_29074,N_28580);
xor U30075 (N_30075,N_29971,N_28651);
nor U30076 (N_30076,N_29822,N_29859);
xor U30077 (N_30077,N_28035,N_29717);
or U30078 (N_30078,N_28205,N_29049);
nand U30079 (N_30079,N_29393,N_28170);
nand U30080 (N_30080,N_28926,N_28330);
xnor U30081 (N_30081,N_29621,N_29902);
nor U30082 (N_30082,N_29212,N_29185);
or U30083 (N_30083,N_28517,N_29321);
and U30084 (N_30084,N_28522,N_29891);
xor U30085 (N_30085,N_29315,N_29796);
and U30086 (N_30086,N_29669,N_28145);
nand U30087 (N_30087,N_28609,N_28392);
nand U30088 (N_30088,N_28880,N_29973);
and U30089 (N_30089,N_29371,N_28462);
xor U30090 (N_30090,N_29028,N_29698);
or U30091 (N_30091,N_29784,N_29612);
or U30092 (N_30092,N_29113,N_28789);
nor U30093 (N_30093,N_28716,N_29464);
nand U30094 (N_30094,N_29919,N_29323);
and U30095 (N_30095,N_29861,N_29386);
nor U30096 (N_30096,N_29823,N_28831);
or U30097 (N_30097,N_28531,N_28923);
and U30098 (N_30098,N_28364,N_29484);
or U30099 (N_30099,N_28322,N_29277);
and U30100 (N_30100,N_29438,N_28102);
or U30101 (N_30101,N_29316,N_28953);
nand U30102 (N_30102,N_28402,N_29164);
xnor U30103 (N_30103,N_29428,N_28351);
nor U30104 (N_30104,N_29813,N_29461);
or U30105 (N_30105,N_29318,N_28407);
xor U30106 (N_30106,N_28732,N_28306);
xnor U30107 (N_30107,N_28456,N_28692);
nor U30108 (N_30108,N_28361,N_29086);
or U30109 (N_30109,N_28386,N_28628);
nand U30110 (N_30110,N_29189,N_29899);
nand U30111 (N_30111,N_28059,N_28741);
and U30112 (N_30112,N_29467,N_29826);
xor U30113 (N_30113,N_29656,N_28235);
or U30114 (N_30114,N_29430,N_28501);
xnor U30115 (N_30115,N_28676,N_29754);
nand U30116 (N_30116,N_29327,N_29645);
and U30117 (N_30117,N_29095,N_29128);
or U30118 (N_30118,N_28044,N_28650);
nor U30119 (N_30119,N_29554,N_28682);
and U30120 (N_30120,N_28806,N_28724);
or U30121 (N_30121,N_28662,N_29686);
xnor U30122 (N_30122,N_28622,N_28547);
nand U30123 (N_30123,N_28250,N_28939);
nor U30124 (N_30124,N_28918,N_28199);
and U30125 (N_30125,N_28352,N_28730);
or U30126 (N_30126,N_28981,N_28803);
and U30127 (N_30127,N_29243,N_28299);
and U30128 (N_30128,N_29172,N_29075);
nand U30129 (N_30129,N_29409,N_29357);
xor U30130 (N_30130,N_28538,N_29425);
and U30131 (N_30131,N_28238,N_29141);
or U30132 (N_30132,N_29572,N_28838);
nor U30133 (N_30133,N_29520,N_29437);
nand U30134 (N_30134,N_29330,N_28921);
nor U30135 (N_30135,N_29732,N_29625);
nor U30136 (N_30136,N_28566,N_28188);
or U30137 (N_30137,N_29675,N_28968);
nor U30138 (N_30138,N_28093,N_29692);
xor U30139 (N_30139,N_28075,N_29198);
nand U30140 (N_30140,N_28892,N_28208);
or U30141 (N_30141,N_28153,N_28324);
and U30142 (N_30142,N_29498,N_28756);
nor U30143 (N_30143,N_29423,N_28868);
nor U30144 (N_30144,N_29362,N_28759);
xnor U30145 (N_30145,N_29068,N_28267);
nand U30146 (N_30146,N_29694,N_29797);
or U30147 (N_30147,N_29283,N_29521);
nand U30148 (N_30148,N_29904,N_28961);
nand U30149 (N_30149,N_28414,N_29261);
nor U30150 (N_30150,N_28408,N_28841);
and U30151 (N_30151,N_29562,N_28180);
or U30152 (N_30152,N_28011,N_28496);
nor U30153 (N_30153,N_29154,N_29308);
nand U30154 (N_30154,N_28980,N_28239);
and U30155 (N_30155,N_28680,N_28191);
nor U30156 (N_30156,N_28976,N_28029);
or U30157 (N_30157,N_28530,N_29905);
and U30158 (N_30158,N_28576,N_29677);
nand U30159 (N_30159,N_28490,N_28010);
nand U30160 (N_30160,N_28200,N_29538);
xor U30161 (N_30161,N_29045,N_28370);
nor U30162 (N_30162,N_28190,N_29455);
xnor U30163 (N_30163,N_29800,N_29365);
nor U30164 (N_30164,N_28254,N_28509);
and U30165 (N_30165,N_28620,N_28482);
and U30166 (N_30166,N_28726,N_28865);
nand U30167 (N_30167,N_29389,N_28721);
nor U30168 (N_30168,N_29273,N_28668);
or U30169 (N_30169,N_29684,N_29936);
nor U30170 (N_30170,N_29553,N_28192);
or U30171 (N_30171,N_28440,N_28819);
nor U30172 (N_30172,N_29026,N_28901);
and U30173 (N_30173,N_29087,N_29661);
or U30174 (N_30174,N_28610,N_29395);
nor U30175 (N_30175,N_29238,N_29188);
nand U30176 (N_30176,N_29872,N_29006);
or U30177 (N_30177,N_29269,N_29347);
and U30178 (N_30178,N_29060,N_28132);
or U30179 (N_30179,N_29264,N_28665);
nand U30180 (N_30180,N_28018,N_29944);
nor U30181 (N_30181,N_29685,N_29771);
or U30182 (N_30182,N_29814,N_29080);
and U30183 (N_30183,N_29585,N_28753);
nor U30184 (N_30184,N_29664,N_29618);
and U30185 (N_30185,N_28479,N_28373);
or U30186 (N_30186,N_28061,N_28301);
or U30187 (N_30187,N_29509,N_28141);
xor U30188 (N_30188,N_28222,N_28935);
and U30189 (N_30189,N_28270,N_28760);
and U30190 (N_30190,N_28277,N_28037);
xor U30191 (N_30191,N_28768,N_29319);
and U30192 (N_30192,N_29847,N_28106);
and U30193 (N_30193,N_29740,N_29485);
and U30194 (N_30194,N_28051,N_29260);
nand U30195 (N_30195,N_29292,N_28050);
and U30196 (N_30196,N_28451,N_29274);
nand U30197 (N_30197,N_29184,N_28335);
or U30198 (N_30198,N_28209,N_29898);
nor U30199 (N_30199,N_29793,N_28657);
xor U30200 (N_30200,N_28098,N_29950);
nand U30201 (N_30201,N_29358,N_29832);
and U30202 (N_30202,N_29419,N_28390);
nor U30203 (N_30203,N_29882,N_28644);
nor U30204 (N_30204,N_28601,N_29781);
xnor U30205 (N_30205,N_29079,N_29886);
nor U30206 (N_30206,N_29312,N_29426);
or U30207 (N_30207,N_29256,N_28954);
xnor U30208 (N_30208,N_29054,N_28274);
and U30209 (N_30209,N_29081,N_29938);
nor U30210 (N_30210,N_28175,N_28007);
and U30211 (N_30211,N_28342,N_28090);
xnor U30212 (N_30212,N_29439,N_28832);
nor U30213 (N_30213,N_29951,N_29631);
nand U30214 (N_30214,N_29736,N_28070);
nor U30215 (N_30215,N_29515,N_28129);
nand U30216 (N_30216,N_29531,N_29728);
nand U30217 (N_30217,N_29765,N_29206);
or U30218 (N_30218,N_29820,N_29276);
xor U30219 (N_30219,N_28927,N_28749);
nand U30220 (N_30220,N_28537,N_29992);
or U30221 (N_30221,N_29476,N_28424);
xor U30222 (N_30222,N_29854,N_29402);
xnor U30223 (N_30223,N_29897,N_29452);
or U30224 (N_30224,N_29042,N_28535);
and U30225 (N_30225,N_29932,N_28187);
nand U30226 (N_30226,N_28378,N_28582);
xnor U30227 (N_30227,N_28323,N_29460);
or U30228 (N_30228,N_28169,N_28336);
nand U30229 (N_30229,N_29116,N_29048);
xor U30230 (N_30230,N_29768,N_29615);
and U30231 (N_30231,N_28242,N_28000);
nand U30232 (N_30232,N_28138,N_28340);
and U30233 (N_30233,N_29345,N_28718);
nor U30234 (N_30234,N_28183,N_29328);
nand U30235 (N_30235,N_29988,N_29607);
nor U30236 (N_30236,N_29084,N_28856);
xor U30237 (N_30237,N_28572,N_29536);
nand U30238 (N_30238,N_28486,N_29415);
xor U30239 (N_30239,N_29734,N_29199);
or U30240 (N_30240,N_28967,N_28052);
nand U30241 (N_30241,N_29778,N_29159);
or U30242 (N_30242,N_28673,N_29842);
and U30243 (N_30243,N_29144,N_28325);
nand U30244 (N_30244,N_29456,N_28775);
nand U30245 (N_30245,N_28885,N_29436);
nor U30246 (N_30246,N_29610,N_29494);
or U30247 (N_30247,N_29433,N_28597);
xnor U30248 (N_30248,N_29954,N_29912);
nor U30249 (N_30249,N_28743,N_28211);
nand U30250 (N_30250,N_28108,N_29716);
nand U30251 (N_30251,N_28605,N_29879);
nand U30252 (N_30252,N_28684,N_29566);
and U30253 (N_30253,N_29939,N_29809);
xor U30254 (N_30254,N_29666,N_28508);
or U30255 (N_30255,N_29731,N_28964);
nand U30256 (N_30256,N_29941,N_28160);
nand U30257 (N_30257,N_29480,N_29351);
and U30258 (N_30258,N_28688,N_29094);
nand U30259 (N_30259,N_28232,N_28487);
nor U30260 (N_30260,N_28715,N_29552);
and U30261 (N_30261,N_29031,N_29638);
nor U30262 (N_30262,N_28608,N_29795);
nor U30263 (N_30263,N_29794,N_29300);
nand U30264 (N_30264,N_28128,N_28930);
and U30265 (N_30265,N_29176,N_29588);
nor U30266 (N_30266,N_28779,N_28307);
nor U30267 (N_30267,N_29182,N_28989);
nand U30268 (N_30268,N_28339,N_28649);
and U30269 (N_30269,N_28548,N_28646);
nand U30270 (N_30270,N_29935,N_29712);
or U30271 (N_30271,N_29600,N_28006);
xnor U30272 (N_30272,N_29746,N_28687);
xnor U30273 (N_30273,N_29753,N_28023);
nor U30274 (N_30274,N_29601,N_29282);
or U30275 (N_30275,N_29751,N_28393);
and U30276 (N_30276,N_28925,N_29076);
and U30277 (N_30277,N_28505,N_28864);
or U30278 (N_30278,N_29018,N_28558);
or U30279 (N_30279,N_29671,N_28249);
or U30280 (N_30280,N_29895,N_29338);
nand U30281 (N_30281,N_28846,N_29937);
xor U30282 (N_30282,N_28912,N_28068);
xnor U30283 (N_30283,N_29632,N_28984);
or U30284 (N_30284,N_28540,N_28404);
nand U30285 (N_30285,N_28381,N_28906);
nor U30286 (N_30286,N_28406,N_29413);
and U30287 (N_30287,N_29417,N_28659);
and U30288 (N_30288,N_28573,N_28642);
xor U30289 (N_30289,N_28998,N_28416);
nor U30290 (N_30290,N_29896,N_28761);
xor U30291 (N_30291,N_28481,N_29096);
xnor U30292 (N_30292,N_29225,N_29285);
nor U30293 (N_30293,N_28127,N_29210);
and U30294 (N_30294,N_28845,N_28368);
xnor U30295 (N_30295,N_29077,N_29577);
and U30296 (N_30296,N_29392,N_28467);
nor U30297 (N_30297,N_28638,N_28251);
nor U30298 (N_30298,N_28816,N_29770);
nand U30299 (N_30299,N_28577,N_29254);
nor U30300 (N_30300,N_29642,N_28510);
or U30301 (N_30301,N_29910,N_29876);
nor U30302 (N_30302,N_29482,N_28419);
and U30303 (N_30303,N_28281,N_28396);
nand U30304 (N_30304,N_28765,N_28742);
nand U30305 (N_30305,N_28258,N_29802);
xor U30306 (N_30306,N_29483,N_28950);
nor U30307 (N_30307,N_28498,N_29541);
and U30308 (N_30308,N_28204,N_28438);
nor U30309 (N_30309,N_29940,N_29724);
nor U30310 (N_30310,N_29332,N_29372);
nor U30311 (N_30311,N_28105,N_28941);
xnor U30312 (N_30312,N_29401,N_28488);
and U30313 (N_30313,N_29512,N_28896);
or U30314 (N_30314,N_29616,N_29550);
nor U30315 (N_30315,N_29364,N_28604);
and U30316 (N_30316,N_29636,N_28174);
nand U30317 (N_30317,N_28613,N_29477);
or U30318 (N_30318,N_29090,N_28116);
or U30319 (N_30319,N_29445,N_29829);
and U30320 (N_30320,N_29667,N_28700);
nand U30321 (N_30321,N_28300,N_28740);
or U30322 (N_30322,N_29474,N_29107);
nand U30323 (N_30323,N_29548,N_29534);
and U30324 (N_30324,N_28219,N_28195);
nor U30325 (N_30325,N_28713,N_28872);
or U30326 (N_30326,N_29858,N_28444);
or U30327 (N_30327,N_29257,N_29394);
nand U30328 (N_30328,N_29267,N_29178);
xor U30329 (N_30329,N_28221,N_29376);
nand U30330 (N_30330,N_28624,N_29725);
or U30331 (N_30331,N_29173,N_28725);
nor U30332 (N_30332,N_29381,N_28372);
xnor U30333 (N_30333,N_29703,N_28264);
and U30334 (N_30334,N_28985,N_28122);
and U30335 (N_30335,N_28842,N_29752);
and U30336 (N_30336,N_29134,N_28499);
or U30337 (N_30337,N_28395,N_28942);
nor U30338 (N_30338,N_28988,N_29320);
or U30339 (N_30339,N_29002,N_28049);
or U30340 (N_30340,N_28148,N_28778);
or U30341 (N_30341,N_29673,N_29043);
or U30342 (N_30342,N_28997,N_29124);
and U30343 (N_30343,N_29982,N_29535);
nor U30344 (N_30344,N_28965,N_29668);
nand U30345 (N_30345,N_29085,N_28963);
nor U30346 (N_30346,N_29258,N_29967);
xnor U30347 (N_30347,N_28786,N_29819);
or U30348 (N_30348,N_29216,N_29873);
nor U30349 (N_30349,N_28674,N_29447);
or U30350 (N_30350,N_29730,N_29408);
xnor U30351 (N_30351,N_28347,N_28476);
and U30352 (N_30352,N_29605,N_28707);
xor U30353 (N_30353,N_29375,N_28924);
and U30354 (N_30354,N_29434,N_28561);
and U30355 (N_30355,N_29041,N_28389);
nand U30356 (N_30356,N_29037,N_29091);
nand U30357 (N_30357,N_29831,N_29652);
or U30358 (N_30358,N_28581,N_29296);
xnor U30359 (N_30359,N_28256,N_29690);
nand U30360 (N_30360,N_28748,N_29962);
nand U30361 (N_30361,N_29776,N_29166);
nand U30362 (N_30362,N_29877,N_29889);
nor U30363 (N_30363,N_28592,N_28111);
nor U30364 (N_30364,N_29335,N_28015);
nand U30365 (N_30365,N_29231,N_28943);
and U30366 (N_30366,N_29744,N_28354);
xnor U30367 (N_30367,N_28751,N_29676);
nand U30368 (N_30368,N_29197,N_28729);
nand U30369 (N_30369,N_29595,N_29012);
and U30370 (N_30370,N_29949,N_29108);
and U30371 (N_30371,N_29493,N_29022);
and U30372 (N_30372,N_29567,N_29025);
xnor U30373 (N_30373,N_28060,N_28194);
nand U30374 (N_30374,N_28647,N_29885);
nor U30375 (N_30375,N_28246,N_28722);
and U30376 (N_30376,N_28783,N_28584);
nand U30377 (N_30377,N_28553,N_29475);
nand U30378 (N_30378,N_29278,N_29624);
nor U30379 (N_30379,N_29815,N_28552);
nor U30380 (N_30380,N_28425,N_28969);
xnor U30381 (N_30381,N_29110,N_29405);
or U30382 (N_30382,N_29830,N_28828);
nor U30383 (N_30383,N_28539,N_28720);
or U30384 (N_30384,N_28631,N_28310);
nor U30385 (N_30385,N_28947,N_29069);
nand U30386 (N_30386,N_29369,N_29262);
xnor U30387 (N_30387,N_29637,N_28046);
and U30388 (N_30388,N_28888,N_29827);
or U30389 (N_30389,N_29367,N_28327);
and U30390 (N_30390,N_29646,N_28709);
and U30391 (N_30391,N_29868,N_28279);
or U30392 (N_30392,N_28080,N_29119);
nor U30393 (N_30393,N_29317,N_29726);
and U30394 (N_30394,N_29853,N_28664);
or U30395 (N_30395,N_28661,N_28712);
nor U30396 (N_30396,N_28627,N_29855);
and U30397 (N_30397,N_28683,N_28792);
and U30398 (N_30398,N_29497,N_29053);
or U30399 (N_30399,N_28915,N_29050);
nor U30400 (N_30400,N_28436,N_29036);
or U30401 (N_30401,N_28109,N_28866);
xnor U30402 (N_30402,N_28030,N_29047);
or U30403 (N_30403,N_29146,N_29789);
and U30404 (N_30404,N_28589,N_28136);
nor U30405 (N_30405,N_28995,N_29556);
xnor U30406 (N_30406,N_28889,N_29016);
and U30407 (N_30407,N_28830,N_29996);
nor U30408 (N_30408,N_29748,N_29126);
nand U30409 (N_30409,N_29103,N_29488);
nor U30410 (N_30410,N_29930,N_29183);
nor U30411 (N_30411,N_28168,N_29921);
and U30412 (N_30412,N_29662,N_29451);
xor U30413 (N_30413,N_29757,N_28648);
nor U30414 (N_30414,N_29023,N_29174);
nor U30415 (N_30415,N_29568,N_28694);
nor U30416 (N_30416,N_28144,N_28067);
xor U30417 (N_30417,N_28384,N_28265);
or U30418 (N_30418,N_28036,N_29510);
or U30419 (N_30419,N_29617,N_28849);
or U30420 (N_30420,N_29303,N_29241);
nand U30421 (N_30421,N_29884,N_29530);
nand U30422 (N_30422,N_28317,N_28933);
nor U30423 (N_30423,N_29200,N_29311);
and U30424 (N_30424,N_28379,N_28269);
and U30425 (N_30425,N_28096,N_28152);
nor U30426 (N_30426,N_29305,N_28296);
nor U30427 (N_30427,N_29496,N_29598);
nor U30428 (N_30428,N_28672,N_29729);
nand U30429 (N_30429,N_29804,N_29704);
nor U30430 (N_30430,N_29309,N_28911);
and U30431 (N_30431,N_28365,N_28367);
nand U30432 (N_30432,N_29398,N_28196);
and U30433 (N_30433,N_28863,N_28994);
or U30434 (N_30434,N_28787,N_29805);
xor U30435 (N_30435,N_29129,N_28240);
and U30436 (N_30436,N_28745,N_28433);
and U30437 (N_30437,N_29514,N_28355);
nand U30438 (N_30438,N_29251,N_28520);
or U30439 (N_30439,N_29192,N_29380);
xnor U30440 (N_30440,N_29301,N_28869);
and U30441 (N_30441,N_28003,N_29738);
xor U30442 (N_30442,N_28181,N_28477);
nand U30443 (N_30443,N_28179,N_28328);
nor U30444 (N_30444,N_28614,N_28103);
nand U30445 (N_30445,N_28883,N_29325);
and U30446 (N_30446,N_29112,N_28401);
and U30447 (N_30447,N_29500,N_28588);
xnor U30448 (N_30448,N_28574,N_28356);
nand U30449 (N_30449,N_29024,N_28972);
nor U30450 (N_30450,N_29786,N_29481);
xnor U30451 (N_30451,N_28226,N_28893);
xnor U30452 (N_30452,N_29239,N_28701);
nor U30453 (N_30453,N_29466,N_29088);
xnor U30454 (N_30454,N_29670,N_28033);
and U30455 (N_30455,N_29966,N_29293);
and U30456 (N_30456,N_28147,N_28788);
nand U30457 (N_30457,N_29106,N_29522);
xor U30458 (N_30458,N_28795,N_29203);
or U30459 (N_30459,N_28137,N_28822);
nand U30460 (N_30460,N_28791,N_29155);
nor U30461 (N_30461,N_28554,N_28360);
xnor U30462 (N_30462,N_29343,N_29078);
or U30463 (N_30463,N_28185,N_28057);
nand U30464 (N_30464,N_29974,N_28442);
nand U30465 (N_30465,N_28675,N_29570);
nand U30466 (N_30466,N_29593,N_29927);
and U30467 (N_30467,N_29529,N_28844);
nor U30468 (N_30468,N_28708,N_29719);
nor U30469 (N_30469,N_29339,N_29366);
or U30470 (N_30470,N_29102,N_28758);
nor U30471 (N_30471,N_29573,N_28432);
nand U30472 (N_30472,N_28303,N_28769);
nand U30473 (N_30473,N_28810,N_28115);
and U30474 (N_30474,N_29945,N_28807);
or U30475 (N_30475,N_28271,N_28189);
nand U30476 (N_30476,N_29862,N_29242);
and U30477 (N_30477,N_28366,N_29150);
and U30478 (N_30478,N_29574,N_28375);
and U30479 (N_30479,N_28056,N_29639);
nor U30480 (N_30480,N_28542,N_28236);
or U30481 (N_30481,N_29377,N_29972);
and U30482 (N_30482,N_29918,N_28417);
or U30483 (N_30483,N_28836,N_29250);
xnor U30484 (N_30484,N_29416,N_28289);
and U30485 (N_30485,N_28053,N_28871);
and U30486 (N_30486,N_29418,N_28678);
xnor U30487 (N_30487,N_29633,N_29863);
xnor U30488 (N_30488,N_29777,N_28891);
nand U30489 (N_30489,N_28039,N_29067);
nand U30490 (N_30490,N_28909,N_29833);
xor U30491 (N_30491,N_28086,N_29582);
or U30492 (N_30492,N_29630,N_28853);
and U30493 (N_30493,N_28076,N_28171);
nor U30494 (N_30494,N_28085,N_28956);
xnor U30495 (N_30495,N_28824,N_29539);
xor U30496 (N_30496,N_28385,N_29266);
or U30497 (N_30497,N_28974,N_28799);
nand U30498 (N_30498,N_29845,N_28217);
nor U30499 (N_30499,N_29115,N_29818);
and U30500 (N_30500,N_28736,N_28818);
xnor U30501 (N_30501,N_29013,N_28387);
nand U30502 (N_30502,N_28996,N_28471);
and U30503 (N_30503,N_28895,N_28523);
xnor U30504 (N_30504,N_29479,N_28699);
nor U30505 (N_30505,N_29852,N_29222);
xnor U30506 (N_30506,N_28727,N_29219);
nand U30507 (N_30507,N_29526,N_28772);
xor U30508 (N_30508,N_29644,N_28645);
or U30509 (N_30509,N_29986,N_29458);
nor U30510 (N_30510,N_28570,N_28321);
nand U30511 (N_30511,N_29157,N_28095);
xnor U30512 (N_30512,N_29787,N_29286);
and U30513 (N_30513,N_28653,N_29687);
xor U30514 (N_30514,N_29991,N_28506);
nor U30515 (N_30515,N_29265,N_28557);
and U30516 (N_30516,N_28443,N_28371);
or U30517 (N_30517,N_29397,N_29767);
nand U30518 (N_30518,N_28504,N_28919);
or U30519 (N_30519,N_28248,N_28877);
nor U30520 (N_30520,N_28212,N_29289);
or U30521 (N_30521,N_28193,N_29368);
xor U30522 (N_30522,N_29341,N_28163);
xor U30523 (N_30523,N_29224,N_28502);
nor U30524 (N_30524,N_28630,N_28565);
nand U30525 (N_30525,N_28591,N_28514);
or U30526 (N_30526,N_28418,N_28920);
nand U30527 (N_30527,N_28429,N_28245);
and U30528 (N_30528,N_28415,N_28469);
nand U30529 (N_30529,N_29135,N_28134);
nor U30530 (N_30530,N_29387,N_29981);
xnor U30531 (N_30531,N_28750,N_29190);
nor U30532 (N_30532,N_29122,N_28166);
nor U30533 (N_30533,N_28619,N_28879);
and U30534 (N_30534,N_28024,N_28012);
and U30535 (N_30535,N_28294,N_28237);
nor U30536 (N_30536,N_28827,N_29839);
nor U30537 (N_30537,N_29214,N_28623);
nor U30538 (N_30538,N_28855,N_29281);
xor U30539 (N_30539,N_29353,N_29892);
xor U30540 (N_30540,N_29609,N_29378);
or U30541 (N_30541,N_29275,N_29486);
xnor U30542 (N_30542,N_29217,N_28617);
or U30543 (N_30543,N_28446,N_29761);
or U30544 (N_30544,N_28097,N_28119);
and U30545 (N_30545,N_29240,N_28640);
nand U30546 (N_30546,N_29942,N_29161);
and U30547 (N_30547,N_29431,N_29721);
nor U30548 (N_30548,N_28977,N_28423);
nor U30549 (N_30549,N_29340,N_28733);
or U30550 (N_30550,N_29020,N_28437);
nor U30551 (N_30551,N_28862,N_29329);
nor U30552 (N_30552,N_28887,N_29816);
nand U30553 (N_30553,N_28399,N_29643);
nor U30554 (N_30554,N_29976,N_29411);
xnor U30555 (N_30555,N_28705,N_29931);
or U30556 (N_30556,N_28731,N_28639);
or U30557 (N_30557,N_28062,N_29691);
and U30558 (N_30558,N_29959,N_29569);
or U30559 (N_30559,N_29651,N_28154);
nand U30560 (N_30560,N_29009,N_28629);
nand U30561 (N_30561,N_28120,N_29384);
nand U30562 (N_30562,N_28234,N_28677);
nand U30563 (N_30563,N_29900,N_29968);
xor U30564 (N_30564,N_29232,N_28940);
and U30565 (N_30565,N_28110,N_29856);
xnor U30566 (N_30566,N_28867,N_29177);
nand U30567 (N_30567,N_28280,N_28316);
and U30568 (N_30568,N_29326,N_29614);
xnor U30569 (N_30569,N_29145,N_29764);
or U30570 (N_30570,N_28228,N_28875);
or U30571 (N_30571,N_28290,N_28696);
or U30572 (N_30572,N_28840,N_29131);
nand U30573 (N_30573,N_29578,N_29348);
nand U30574 (N_30574,N_29055,N_29680);
nor U30575 (N_30575,N_28723,N_29956);
nand U30576 (N_30576,N_28706,N_29980);
and U30577 (N_30577,N_28586,N_28669);
xnor U30578 (N_30578,N_29540,N_28562);
nand U30579 (N_30579,N_28491,N_28241);
or U30580 (N_30580,N_29169,N_29727);
xnor U30581 (N_30581,N_29089,N_28805);
xnor U30582 (N_30582,N_28847,N_29205);
xor U30583 (N_30583,N_28074,N_28873);
nand U30584 (N_30584,N_28971,N_28133);
xnor U30585 (N_30585,N_29011,N_29230);
nor U30586 (N_30586,N_28671,N_29870);
or U30587 (N_30587,N_28843,N_29801);
nand U30588 (N_30588,N_28774,N_28599);
and U30589 (N_30589,N_28910,N_28808);
and U30590 (N_30590,N_29151,N_29571);
xnor U30591 (N_30591,N_29194,N_28594);
nand U30592 (N_30592,N_28560,N_29118);
or U30593 (N_30593,N_29213,N_28876);
and U30594 (N_30594,N_29689,N_28014);
or U30595 (N_30595,N_28081,N_29779);
nor U30596 (N_30596,N_28013,N_29688);
nand U30597 (N_30597,N_28521,N_28031);
xor U30598 (N_30598,N_28430,N_29933);
xnor U30599 (N_30599,N_29207,N_29064);
xor U30600 (N_30600,N_28612,N_29501);
nor U30601 (N_30601,N_29459,N_29634);
or U30602 (N_30602,N_29626,N_29970);
or U30603 (N_30603,N_28341,N_28991);
xor U30604 (N_30604,N_28559,N_29180);
xor U30605 (N_30605,N_29017,N_28230);
and U30606 (N_30606,N_29558,N_28634);
nor U30607 (N_30607,N_28155,N_28315);
nor U30608 (N_30608,N_29071,N_29304);
or U30609 (N_30609,N_28473,N_28266);
or U30610 (N_30610,N_29700,N_29288);
nand U30611 (N_30611,N_28259,N_29137);
nand U30612 (N_30612,N_28679,N_29629);
xor U30613 (N_30613,N_29824,N_28345);
xnor U30614 (N_30614,N_29111,N_29513);
xnor U30615 (N_30615,N_29590,N_29997);
xor U30616 (N_30616,N_28578,N_28092);
and U30617 (N_30617,N_29249,N_28796);
nor U30618 (N_30618,N_28541,N_29465);
or U30619 (N_30619,N_29679,N_28434);
nor U30620 (N_30620,N_28349,N_28817);
nor U30621 (N_30621,N_29152,N_28641);
or U30622 (N_30622,N_28455,N_28973);
and U30623 (N_30623,N_29563,N_28460);
nand U30624 (N_30624,N_29769,N_29061);
nor U30625 (N_30625,N_28040,N_28099);
nor U30626 (N_30626,N_29875,N_29527);
or U30627 (N_30627,N_29943,N_28917);
or U30628 (N_30628,N_29313,N_28689);
and U30629 (N_30629,N_29599,N_28602);
xor U30630 (N_30630,N_29817,N_28861);
xor U30631 (N_30631,N_29410,N_28149);
xor U30632 (N_30632,N_29783,N_29774);
nor U30633 (N_30633,N_28207,N_28957);
nor U30634 (N_30634,N_28088,N_29307);
and U30635 (N_30635,N_28159,N_29297);
xnor U30636 (N_30636,N_28203,N_28427);
or U30637 (N_30637,N_29469,N_29663);
nand U30638 (N_30638,N_29762,N_29149);
nor U30639 (N_30639,N_29263,N_29462);
or U30640 (N_30640,N_29995,N_28632);
nand U30641 (N_30641,N_28717,N_28766);
nor U30642 (N_30642,N_28870,N_29010);
nand U30643 (N_30643,N_29739,N_29641);
xor U30644 (N_30644,N_29385,N_28439);
and U30645 (N_30645,N_29105,N_28058);
or U30646 (N_30646,N_29955,N_29127);
xnor U30647 (N_30647,N_28546,N_28172);
xor U30648 (N_30648,N_29707,N_29635);
nand U30649 (N_30649,N_29349,N_29056);
xor U30650 (N_30650,N_28857,N_28685);
nand U30651 (N_30651,N_28763,N_29674);
or U30652 (N_30652,N_29537,N_28276);
nor U30653 (N_30653,N_29532,N_28936);
or U30654 (N_30654,N_28231,N_29442);
and U30655 (N_30655,N_29139,N_29195);
nor U30656 (N_30656,N_29589,N_28958);
or U30657 (N_30657,N_28215,N_29807);
and U30658 (N_30658,N_28494,N_28480);
nor U30659 (N_30659,N_29506,N_29391);
nand U30660 (N_30660,N_29792,N_28292);
nor U30661 (N_30661,N_29653,N_29104);
and U30662 (N_30662,N_29373,N_29489);
or U30663 (N_30663,N_28516,N_28982);
or U30664 (N_30664,N_29983,N_28348);
nor U30665 (N_30665,N_29763,N_28125);
or U30666 (N_30666,N_29140,N_29603);
nor U30667 (N_30667,N_29424,N_28403);
or U30668 (N_30668,N_28951,N_28391);
nor U30669 (N_30669,N_29035,N_29782);
and U30670 (N_30670,N_29701,N_28987);
nand U30671 (N_30671,N_28860,N_28660);
or U30672 (N_30672,N_29355,N_29001);
nand U30673 (N_30673,N_29117,N_29502);
nor U30674 (N_30674,N_29913,N_28776);
or U30675 (N_30675,N_29519,N_29382);
or U30676 (N_30676,N_28534,N_28293);
nor U30677 (N_30677,N_29271,N_28513);
xor U30678 (N_30678,N_29014,N_29396);
nand U30679 (N_30679,N_29960,N_28955);
nand U30680 (N_30680,N_28063,N_28268);
and U30681 (N_30681,N_28636,N_29306);
or U30682 (N_30682,N_29874,N_28287);
and U30683 (N_30683,N_28474,N_29547);
nor U30684 (N_30684,N_28555,N_28017);
or U30685 (N_30685,N_29907,N_29171);
nand U30686 (N_30686,N_29491,N_29597);
nand U30687 (N_30687,N_28771,N_28616);
nor U30688 (N_30688,N_29749,N_29659);
nor U30689 (N_30689,N_29742,N_29864);
xnor U30690 (N_30690,N_28412,N_28794);
and U30691 (N_30691,N_29208,N_28489);
or U30692 (N_30692,N_28595,N_28945);
xnor U30693 (N_30693,N_29503,N_28711);
or U30694 (N_30694,N_28851,N_28475);
nand U30695 (N_30695,N_29928,N_28398);
nand U30696 (N_30696,N_28042,N_28358);
xnor U30697 (N_30697,N_28143,N_28357);
and U30698 (N_30698,N_29733,N_28146);
and U30699 (N_30699,N_28284,N_28286);
nand U30700 (N_30700,N_29559,N_29881);
or U30701 (N_30701,N_28654,N_29204);
nand U30702 (N_30702,N_28551,N_28902);
nor U30703 (N_30703,N_28135,N_28083);
or U30704 (N_30704,N_29835,N_29888);
xnor U30705 (N_30705,N_29083,N_28703);
nand U30706 (N_30706,N_29611,N_28702);
or U30707 (N_30707,N_29072,N_29070);
nor U30708 (N_30708,N_28728,N_29706);
nand U30709 (N_30709,N_29799,N_28983);
nor U30710 (N_30710,N_28113,N_29846);
nand U30711 (N_30711,N_29400,N_29561);
nand U30712 (N_30712,N_29887,N_28739);
xor U30713 (N_30713,N_29229,N_29114);
and U30714 (N_30714,N_28457,N_29403);
nand U30715 (N_30715,N_28311,N_28054);
nor U30716 (N_30716,N_29248,N_28637);
or U30717 (N_30717,N_28821,N_29429);
nand U30718 (N_30718,N_28045,N_29454);
or U30719 (N_30719,N_29211,N_29156);
and U30720 (N_30720,N_29989,N_29678);
or U30721 (N_30721,N_29287,N_29201);
or U30722 (N_30722,N_28162,N_29682);
nor U30723 (N_30723,N_29906,N_28691);
or U30724 (N_30724,N_29406,N_29542);
or U30725 (N_30725,N_28104,N_29755);
xnor U30726 (N_30726,N_28123,N_29019);
xnor U30727 (N_30727,N_28089,N_28319);
nand U30728 (N_30728,N_28253,N_29468);
nand U30729 (N_30729,N_29021,N_29628);
nand U30730 (N_30730,N_29255,N_28218);
and U30731 (N_30731,N_29843,N_29580);
and U30732 (N_30732,N_28394,N_29422);
nand U30733 (N_30733,N_28666,N_28829);
nand U30734 (N_30734,N_28690,N_28338);
or U30735 (N_30735,N_29798,N_28878);
nor U30736 (N_30736,N_29133,N_29811);
xor U30737 (N_30737,N_28283,N_29007);
xor U30738 (N_30738,N_28966,N_29947);
or U30739 (N_30739,N_29361,N_28308);
nand U30740 (N_30740,N_28421,N_29683);
xnor U30741 (N_30741,N_29545,N_28946);
xor U30742 (N_30742,N_28483,N_28959);
xor U30743 (N_30743,N_29702,N_28882);
and U30744 (N_30744,N_28507,N_29961);
nand U30745 (N_30745,N_29565,N_29756);
nand U30746 (N_30746,N_28618,N_29978);
and U30747 (N_30747,N_29883,N_29412);
xor U30748 (N_30748,N_28852,N_28603);
nand U30749 (N_30749,N_29672,N_28781);
and U30750 (N_30750,N_29310,N_28518);
and U30751 (N_30751,N_28515,N_28449);
nand U30752 (N_30752,N_29165,N_29508);
and U30753 (N_30753,N_28633,N_28485);
nand U30754 (N_30754,N_28382,N_28894);
nor U30755 (N_30755,N_28359,N_29640);
xnor U30756 (N_30756,N_29227,N_29860);
and U30757 (N_30757,N_29337,N_28201);
nor U30758 (N_30758,N_28747,N_28611);
nand U30759 (N_30759,N_29964,N_28079);
or U30760 (N_30760,N_28837,N_29867);
or U30761 (N_30761,N_28118,N_29849);
and U30762 (N_30762,N_28038,N_28197);
xor U30763 (N_30763,N_29158,N_29223);
nor U30764 (N_30764,N_29866,N_29354);
nor U30765 (N_30765,N_28670,N_28346);
nand U30766 (N_30766,N_29226,N_29093);
nand U30767 (N_30767,N_28126,N_28907);
xor U30768 (N_30768,N_28527,N_29027);
nand U30769 (N_30769,N_29379,N_29709);
nand U30770 (N_30770,N_28008,N_28350);
or U30771 (N_30771,N_28314,N_29994);
nand U30772 (N_30772,N_29837,N_29302);
xnor U30773 (N_30773,N_28428,N_29125);
and U30774 (N_30774,N_29051,N_29657);
nand U30775 (N_30775,N_29985,N_29052);
xnor U30776 (N_30776,N_28320,N_29926);
nand U30777 (N_30777,N_29490,N_28503);
xnor U30778 (N_30778,N_28313,N_28388);
nor U30779 (N_30779,N_28150,N_28156);
and U30780 (N_30780,N_29871,N_28780);
and U30781 (N_30781,N_28929,N_28698);
and U30782 (N_30782,N_28484,N_29953);
and U30783 (N_30783,N_29252,N_28028);
nor U30784 (N_30784,N_29008,N_28596);
and U30785 (N_30785,N_29160,N_29383);
xor U30786 (N_30786,N_28071,N_29427);
xor U30787 (N_30787,N_28165,N_28064);
and U30788 (N_30788,N_29473,N_29890);
xnor U30789 (N_30789,N_28470,N_28970);
or U30790 (N_30790,N_29594,N_28101);
nor U30791 (N_30791,N_28545,N_29033);
and U30792 (N_30792,N_29758,N_29524);
nand U30793 (N_30793,N_28448,N_28714);
and U30794 (N_30794,N_28225,N_29697);
or U30795 (N_30795,N_28511,N_28734);
xnor U30796 (N_30796,N_29699,N_29922);
nor U30797 (N_30797,N_28938,N_28032);
nand U30798 (N_30798,N_28084,N_28445);
and U30799 (N_30799,N_29649,N_29044);
nor U30800 (N_30800,N_28021,N_29627);
xnor U30801 (N_30801,N_29923,N_29138);
and U30802 (N_30802,N_29516,N_29187);
nor U30803 (N_30803,N_28600,N_29073);
or U30804 (N_30804,N_28532,N_28948);
xor U30805 (N_30805,N_28850,N_29723);
xnor U30806 (N_30806,N_28797,N_29869);
nor U30807 (N_30807,N_29057,N_29440);
nand U30808 (N_30808,N_29901,N_28087);
or U30809 (N_30809,N_28979,N_29450);
nor U30810 (N_30810,N_29543,N_29747);
or U30811 (N_30811,N_28652,N_29421);
and U30812 (N_30812,N_29284,N_28461);
or U30813 (N_30813,N_28223,N_28626);
nand U30814 (N_30814,N_28934,N_28065);
xor U30815 (N_30815,N_29920,N_28615);
or U30816 (N_30816,N_29648,N_28112);
or U30817 (N_30817,N_29234,N_29039);
and U30818 (N_30818,N_28297,N_29390);
or U30819 (N_30819,N_29696,N_28383);
nand U30820 (N_30820,N_28585,N_29245);
nand U30821 (N_30821,N_28825,N_29909);
nor U30822 (N_30822,N_29576,N_29147);
nor U30823 (N_30823,N_28078,N_29708);
or U30824 (N_30824,N_28782,N_28272);
xor U30825 (N_30825,N_28130,N_29324);
nand U30826 (N_30826,N_29993,N_28140);
nor U30827 (N_30827,N_29314,N_29082);
or U30828 (N_30828,N_29760,N_28900);
nor U30829 (N_30829,N_29715,N_29718);
nor U30830 (N_30830,N_29990,N_28377);
xor U30831 (N_30831,N_28410,N_29695);
xnor U30832 (N_30832,N_28468,N_29495);
nand U30833 (N_30833,N_28019,N_29878);
nand U30834 (N_30834,N_28380,N_28043);
xor U30835 (N_30835,N_29713,N_29604);
and U30836 (N_30836,N_28944,N_29714);
and U30837 (N_30837,N_28304,N_28563);
or U30838 (N_30838,N_28754,N_29803);
and U30839 (N_30839,N_29253,N_28990);
nor U30840 (N_30840,N_29142,N_28214);
or U30841 (N_30841,N_29821,N_28450);
nor U30842 (N_30842,N_29097,N_29722);
nor U30843 (N_30843,N_28312,N_29191);
xor U30844 (N_30844,N_28773,N_29336);
nor U30845 (N_30845,N_28400,N_28478);
nor U30846 (N_30846,N_28022,N_29359);
xnor U30847 (N_30847,N_29812,N_28100);
xnor U30848 (N_30848,N_28151,N_29745);
xor U30849 (N_30849,N_29270,N_29038);
and U30850 (N_30850,N_29472,N_29591);
nand U30851 (N_30851,N_28621,N_28291);
and U30852 (N_30852,N_29834,N_29005);
xnor U30853 (N_30853,N_29840,N_28571);
xor U30854 (N_30854,N_29505,N_29130);
nor U30855 (N_30855,N_28809,N_29934);
and U30856 (N_30856,N_29544,N_28229);
or U30857 (N_30857,N_29470,N_28041);
nor U30858 (N_30858,N_29525,N_28452);
and U30859 (N_30859,N_28757,N_28922);
and U30860 (N_30860,N_28663,N_28525);
nand U30861 (N_30861,N_29202,N_28161);
or U30862 (N_30862,N_28027,N_29841);
and U30863 (N_30863,N_28913,N_29750);
and U30864 (N_30864,N_28158,N_28247);
nor U30865 (N_30865,N_28544,N_29167);
nor U30866 (N_30866,N_28492,N_29851);
nor U30867 (N_30867,N_29109,N_29528);
nor U30868 (N_30868,N_28524,N_29492);
and U30869 (N_30869,N_28500,N_29143);
and U30870 (N_30870,N_29352,N_29246);
nand U30871 (N_30871,N_29233,N_28533);
nor U30872 (N_30872,N_28738,N_29435);
nand U30873 (N_30873,N_28459,N_29399);
nand U30874 (N_30874,N_28804,N_28526);
xor U30875 (N_30875,N_29693,N_28579);
nand U30876 (N_30876,N_28420,N_28295);
nand U30877 (N_30877,N_29660,N_28173);
nor U30878 (N_30878,N_29004,N_28411);
and U30879 (N_30879,N_29914,N_29517);
nor U30880 (N_30880,N_28686,N_28362);
nand U30881 (N_30881,N_29478,N_28764);
or U30882 (N_30882,N_28575,N_29441);
or U30883 (N_30883,N_28337,N_29581);
and U30884 (N_30884,N_29221,N_29917);
and U30885 (N_30885,N_28719,N_29092);
nand U30886 (N_30886,N_28755,N_28363);
xor U30887 (N_30887,N_29148,N_28904);
xnor U30888 (N_30888,N_28275,N_28658);
xor U30889 (N_30889,N_28244,N_28512);
xor U30890 (N_30890,N_28263,N_29181);
or U30891 (N_30891,N_29929,N_29979);
or U30892 (N_30892,N_28826,N_28233);
nor U30893 (N_30893,N_29810,N_29218);
xor U30894 (N_30894,N_29136,N_28752);
nor U30895 (N_30895,N_28903,N_29586);
xnor U30896 (N_30896,N_29984,N_28587);
nor U30897 (N_30897,N_29063,N_29175);
nand U30898 (N_30898,N_28854,N_28020);
and U30899 (N_30899,N_29374,N_28801);
xor U30900 (N_30900,N_28564,N_28962);
nor U30901 (N_30901,N_28567,N_29443);
xor U30902 (N_30902,N_29121,N_29471);
or U30903 (N_30903,N_29333,N_28811);
xor U30904 (N_30904,N_28528,N_29356);
xnor U30905 (N_30905,N_28704,N_29596);
or U30906 (N_30906,N_28790,N_28305);
xnor U30907 (N_30907,N_29432,N_28916);
or U30908 (N_30908,N_28784,N_28458);
xor U30909 (N_30909,N_29518,N_28899);
and U30910 (N_30910,N_28262,N_28464);
and U30911 (N_30911,N_29236,N_29507);
and U30912 (N_30912,N_28833,N_29759);
xnor U30913 (N_30913,N_28435,N_28569);
nand U30914 (N_30914,N_29977,N_29946);
xnor U30915 (N_30915,N_28815,N_29179);
xor U30916 (N_30916,N_28405,N_29280);
xnor U30917 (N_30917,N_28182,N_28431);
xnor U30918 (N_30918,N_29322,N_28047);
xnor U30919 (N_30919,N_28167,N_28077);
nor U30920 (N_30920,N_28897,N_29446);
nand U30921 (N_30921,N_28413,N_29247);
nor U30922 (N_30922,N_28005,N_28374);
and U30923 (N_30923,N_28823,N_29998);
and U30924 (N_30924,N_28697,N_29168);
and U30925 (N_30925,N_28583,N_28094);
nor U30926 (N_30926,N_28800,N_29420);
or U30927 (N_30927,N_28813,N_28309);
and U30928 (N_30928,N_28016,N_28121);
nor U30929 (N_30929,N_28710,N_29999);
xnor U30930 (N_30930,N_28441,N_28004);
and U30931 (N_30931,N_28905,N_29965);
nor U30932 (N_30932,N_29808,N_29162);
nand U30933 (N_30933,N_29613,N_28667);
nor U30934 (N_30934,N_29775,N_28073);
xnor U30935 (N_30935,N_29463,N_28048);
or U30936 (N_30936,N_29186,N_28376);
and U30937 (N_30937,N_28802,N_29622);
nand U30938 (N_30938,N_29360,N_29062);
nand U30939 (N_30939,N_28343,N_28055);
nand U30940 (N_30940,N_28001,N_28834);
and U30941 (N_30941,N_28466,N_28091);
and U30942 (N_30942,N_29963,N_28890);
xnor U30943 (N_30943,N_29772,N_29046);
nand U30944 (N_30944,N_29619,N_29647);
nand U30945 (N_30945,N_29893,N_28069);
nand U30946 (N_30946,N_28914,N_29003);
and U30947 (N_30947,N_28117,N_29404);
xnor U30948 (N_30948,N_28453,N_28952);
nand U30949 (N_30949,N_28397,N_29272);
nand U30950 (N_30950,N_29583,N_29344);
or U30951 (N_30951,N_29504,N_28206);
nor U30952 (N_30952,N_28333,N_29788);
nor U30953 (N_30953,N_28176,N_29952);
nor U30954 (N_30954,N_28960,N_28318);
and U30955 (N_30955,N_29584,N_28298);
xnor U30956 (N_30956,N_28735,N_29924);
and U30957 (N_30957,N_28131,N_29911);
xor U30958 (N_30958,N_29957,N_28243);
xnor U30959 (N_30959,N_28798,N_28635);
and U30960 (N_30960,N_29029,N_28034);
xnor U30961 (N_30961,N_28625,N_28202);
or U30962 (N_30962,N_29331,N_29059);
xor U30963 (N_30963,N_28770,N_28186);
and U30964 (N_30964,N_29295,N_28353);
nand U30965 (N_30965,N_28344,N_28178);
and U30966 (N_30966,N_29448,N_29032);
or U30967 (N_30967,N_28737,N_28762);
and U30968 (N_30968,N_29579,N_29711);
nor U30969 (N_30969,N_29828,N_29737);
xnor U30970 (N_30970,N_29710,N_29511);
and U30971 (N_30971,N_28848,N_29279);
and U30972 (N_30972,N_29268,N_29215);
nand U30973 (N_30973,N_28302,N_29564);
nor U30974 (N_30974,N_29836,N_29844);
or U30975 (N_30975,N_29228,N_28072);
nor U30976 (N_30976,N_29654,N_28785);
nand U30977 (N_30977,N_28937,N_28332);
xor U30978 (N_30978,N_29806,N_28255);
nor U30979 (N_30979,N_29388,N_28369);
nand U30980 (N_30980,N_29449,N_28026);
nand U30981 (N_30981,N_28252,N_29209);
or U30982 (N_30982,N_28656,N_28695);
or U30983 (N_30983,N_28549,N_28495);
nor U30984 (N_30984,N_28598,N_28812);
xor U30985 (N_30985,N_29132,N_29606);
xor U30986 (N_30986,N_28568,N_28681);
xnor U30987 (N_30987,N_28993,N_28793);
xnor U30988 (N_30988,N_28898,N_29681);
nand U30989 (N_30989,N_28820,N_28493);
nor U30990 (N_30990,N_28928,N_28107);
and U30991 (N_30991,N_29557,N_29196);
and U30992 (N_30992,N_29299,N_28590);
nor U30993 (N_30993,N_28643,N_28556);
or U30994 (N_30994,N_29220,N_28884);
nand U30995 (N_30995,N_28655,N_28198);
nor U30996 (N_30996,N_29560,N_29058);
or U30997 (N_30997,N_28606,N_28746);
xnor U30998 (N_30998,N_28835,N_29592);
or U30999 (N_30999,N_28260,N_29290);
or U31000 (N_31000,N_28923,N_29071);
nand U31001 (N_31001,N_29906,N_29336);
xnor U31002 (N_31002,N_28389,N_28164);
and U31003 (N_31003,N_28040,N_29957);
or U31004 (N_31004,N_29611,N_28117);
nor U31005 (N_31005,N_29804,N_28372);
or U31006 (N_31006,N_29839,N_28554);
nor U31007 (N_31007,N_29820,N_28030);
xor U31008 (N_31008,N_29275,N_29978);
nor U31009 (N_31009,N_29370,N_28946);
and U31010 (N_31010,N_28217,N_28741);
and U31011 (N_31011,N_29024,N_29815);
xor U31012 (N_31012,N_28329,N_28581);
xor U31013 (N_31013,N_29588,N_29845);
nand U31014 (N_31014,N_29709,N_28245);
nand U31015 (N_31015,N_28342,N_28820);
and U31016 (N_31016,N_29605,N_29376);
nand U31017 (N_31017,N_29727,N_29964);
nand U31018 (N_31018,N_29611,N_29889);
xnor U31019 (N_31019,N_28111,N_29604);
nand U31020 (N_31020,N_28140,N_29974);
or U31021 (N_31021,N_28259,N_28957);
or U31022 (N_31022,N_28436,N_28141);
nand U31023 (N_31023,N_28299,N_29463);
xor U31024 (N_31024,N_29696,N_29163);
and U31025 (N_31025,N_28382,N_28388);
or U31026 (N_31026,N_28353,N_29256);
xnor U31027 (N_31027,N_28826,N_29397);
nor U31028 (N_31028,N_28445,N_29122);
nor U31029 (N_31029,N_29676,N_29390);
or U31030 (N_31030,N_28595,N_28344);
nand U31031 (N_31031,N_28897,N_29048);
or U31032 (N_31032,N_29578,N_29907);
xnor U31033 (N_31033,N_28759,N_29959);
and U31034 (N_31034,N_28156,N_28129);
xor U31035 (N_31035,N_28038,N_28125);
nor U31036 (N_31036,N_28924,N_29311);
and U31037 (N_31037,N_29967,N_29718);
xor U31038 (N_31038,N_28294,N_28492);
and U31039 (N_31039,N_29620,N_29795);
nor U31040 (N_31040,N_28169,N_28792);
or U31041 (N_31041,N_28877,N_28939);
or U31042 (N_31042,N_28981,N_28423);
or U31043 (N_31043,N_29612,N_28090);
xnor U31044 (N_31044,N_29654,N_28401);
nor U31045 (N_31045,N_29196,N_28985);
nor U31046 (N_31046,N_28483,N_29721);
or U31047 (N_31047,N_28450,N_29070);
nand U31048 (N_31048,N_28359,N_28086);
nand U31049 (N_31049,N_28238,N_29198);
and U31050 (N_31050,N_29583,N_29613);
or U31051 (N_31051,N_29515,N_29179);
or U31052 (N_31052,N_29462,N_28649);
xnor U31053 (N_31053,N_28444,N_28792);
and U31054 (N_31054,N_28595,N_29657);
or U31055 (N_31055,N_29575,N_29827);
and U31056 (N_31056,N_29105,N_28688);
nand U31057 (N_31057,N_28478,N_29056);
and U31058 (N_31058,N_28532,N_29962);
nand U31059 (N_31059,N_28607,N_28526);
xnor U31060 (N_31060,N_28042,N_29769);
or U31061 (N_31061,N_28152,N_29578);
nand U31062 (N_31062,N_29031,N_28983);
nand U31063 (N_31063,N_28676,N_29653);
nor U31064 (N_31064,N_29327,N_28089);
nor U31065 (N_31065,N_28170,N_29329);
xnor U31066 (N_31066,N_28611,N_28952);
and U31067 (N_31067,N_28328,N_29149);
xor U31068 (N_31068,N_29910,N_29216);
or U31069 (N_31069,N_29936,N_29339);
and U31070 (N_31070,N_29916,N_29652);
or U31071 (N_31071,N_29914,N_29691);
and U31072 (N_31072,N_28545,N_29224);
xor U31073 (N_31073,N_28679,N_28912);
and U31074 (N_31074,N_29585,N_29137);
xor U31075 (N_31075,N_28825,N_29294);
nor U31076 (N_31076,N_28180,N_29357);
nor U31077 (N_31077,N_29012,N_29813);
nor U31078 (N_31078,N_29102,N_28496);
nor U31079 (N_31079,N_29322,N_28759);
nand U31080 (N_31080,N_29126,N_28652);
or U31081 (N_31081,N_29250,N_29537);
nor U31082 (N_31082,N_29620,N_28355);
nor U31083 (N_31083,N_28151,N_28202);
nand U31084 (N_31084,N_28861,N_29390);
and U31085 (N_31085,N_29608,N_28198);
and U31086 (N_31086,N_28734,N_29333);
nand U31087 (N_31087,N_29064,N_29108);
nor U31088 (N_31088,N_28559,N_28986);
nor U31089 (N_31089,N_29222,N_29282);
xnor U31090 (N_31090,N_29501,N_29869);
and U31091 (N_31091,N_28469,N_29341);
xor U31092 (N_31092,N_29376,N_28770);
xor U31093 (N_31093,N_29252,N_29467);
or U31094 (N_31094,N_28304,N_29667);
nand U31095 (N_31095,N_29937,N_28838);
nor U31096 (N_31096,N_28360,N_29242);
nand U31097 (N_31097,N_29949,N_29098);
and U31098 (N_31098,N_29805,N_28754);
xnor U31099 (N_31099,N_28116,N_29886);
nor U31100 (N_31100,N_29026,N_29979);
xor U31101 (N_31101,N_29265,N_29058);
and U31102 (N_31102,N_29843,N_29592);
and U31103 (N_31103,N_28962,N_29275);
or U31104 (N_31104,N_28277,N_28004);
and U31105 (N_31105,N_29346,N_29972);
nand U31106 (N_31106,N_29843,N_28574);
nand U31107 (N_31107,N_29215,N_28587);
xor U31108 (N_31108,N_28814,N_29087);
nand U31109 (N_31109,N_28254,N_29102);
and U31110 (N_31110,N_29602,N_29757);
nand U31111 (N_31111,N_28892,N_29406);
nor U31112 (N_31112,N_29610,N_28983);
nor U31113 (N_31113,N_29082,N_28506);
or U31114 (N_31114,N_29784,N_28142);
xor U31115 (N_31115,N_29949,N_28533);
nand U31116 (N_31116,N_29305,N_29760);
nand U31117 (N_31117,N_28168,N_29958);
xnor U31118 (N_31118,N_28855,N_28311);
and U31119 (N_31119,N_28065,N_28366);
nor U31120 (N_31120,N_29920,N_28930);
xnor U31121 (N_31121,N_28475,N_29778);
nor U31122 (N_31122,N_29547,N_29427);
nand U31123 (N_31123,N_28873,N_28048);
xnor U31124 (N_31124,N_29721,N_29934);
or U31125 (N_31125,N_29027,N_28554);
xnor U31126 (N_31126,N_28849,N_28022);
xnor U31127 (N_31127,N_29788,N_29616);
nand U31128 (N_31128,N_28207,N_29395);
xnor U31129 (N_31129,N_28149,N_29374);
nor U31130 (N_31130,N_28314,N_28230);
nand U31131 (N_31131,N_29703,N_28074);
or U31132 (N_31132,N_29762,N_28530);
xor U31133 (N_31133,N_28084,N_28783);
nand U31134 (N_31134,N_29683,N_29988);
nand U31135 (N_31135,N_28284,N_28481);
nand U31136 (N_31136,N_29531,N_29024);
nor U31137 (N_31137,N_29977,N_29173);
or U31138 (N_31138,N_28671,N_28193);
nand U31139 (N_31139,N_28801,N_29525);
xor U31140 (N_31140,N_28468,N_28392);
or U31141 (N_31141,N_28771,N_28033);
nor U31142 (N_31142,N_29727,N_29104);
nor U31143 (N_31143,N_29922,N_29805);
nand U31144 (N_31144,N_29463,N_28102);
or U31145 (N_31145,N_29369,N_29746);
and U31146 (N_31146,N_29089,N_28215);
nor U31147 (N_31147,N_28831,N_28089);
xor U31148 (N_31148,N_29579,N_29450);
nor U31149 (N_31149,N_29286,N_28345);
nor U31150 (N_31150,N_29955,N_28094);
nand U31151 (N_31151,N_29047,N_28772);
nor U31152 (N_31152,N_29855,N_29192);
xor U31153 (N_31153,N_29734,N_29828);
and U31154 (N_31154,N_29660,N_29387);
or U31155 (N_31155,N_29089,N_29731);
nand U31156 (N_31156,N_28458,N_28923);
xnor U31157 (N_31157,N_29230,N_29019);
nor U31158 (N_31158,N_29642,N_29462);
and U31159 (N_31159,N_28812,N_29223);
or U31160 (N_31160,N_29952,N_29320);
or U31161 (N_31161,N_28135,N_29122);
or U31162 (N_31162,N_29527,N_28792);
or U31163 (N_31163,N_28660,N_29161);
and U31164 (N_31164,N_28612,N_28064);
nand U31165 (N_31165,N_28029,N_28156);
xor U31166 (N_31166,N_29606,N_28847);
and U31167 (N_31167,N_28533,N_29520);
or U31168 (N_31168,N_28209,N_29628);
nand U31169 (N_31169,N_29278,N_28498);
nor U31170 (N_31170,N_28091,N_28065);
nand U31171 (N_31171,N_28880,N_29248);
nand U31172 (N_31172,N_28265,N_28589);
nor U31173 (N_31173,N_28037,N_28093);
and U31174 (N_31174,N_28622,N_29172);
xor U31175 (N_31175,N_28999,N_29865);
xnor U31176 (N_31176,N_28933,N_29195);
nor U31177 (N_31177,N_29331,N_28096);
nor U31178 (N_31178,N_28203,N_29719);
and U31179 (N_31179,N_29631,N_28105);
nand U31180 (N_31180,N_29882,N_28301);
and U31181 (N_31181,N_29334,N_29591);
nor U31182 (N_31182,N_28547,N_28562);
nand U31183 (N_31183,N_29704,N_29648);
nand U31184 (N_31184,N_28267,N_28323);
and U31185 (N_31185,N_28736,N_29672);
nand U31186 (N_31186,N_29444,N_28824);
nor U31187 (N_31187,N_29297,N_28477);
or U31188 (N_31188,N_29713,N_29075);
nand U31189 (N_31189,N_28062,N_29895);
nand U31190 (N_31190,N_29528,N_29792);
nor U31191 (N_31191,N_28082,N_28630);
nand U31192 (N_31192,N_28966,N_28436);
nand U31193 (N_31193,N_28740,N_28920);
or U31194 (N_31194,N_28620,N_29593);
nor U31195 (N_31195,N_29993,N_28249);
and U31196 (N_31196,N_28168,N_29968);
nor U31197 (N_31197,N_28202,N_28248);
nor U31198 (N_31198,N_28802,N_28136);
nor U31199 (N_31199,N_28841,N_29172);
or U31200 (N_31200,N_29409,N_29539);
and U31201 (N_31201,N_28255,N_29397);
nand U31202 (N_31202,N_28908,N_28655);
xor U31203 (N_31203,N_29064,N_29448);
or U31204 (N_31204,N_29530,N_28328);
and U31205 (N_31205,N_29067,N_29502);
or U31206 (N_31206,N_28637,N_29788);
nor U31207 (N_31207,N_28376,N_29271);
nand U31208 (N_31208,N_28145,N_28373);
xnor U31209 (N_31209,N_29961,N_29061);
xnor U31210 (N_31210,N_28904,N_28784);
xor U31211 (N_31211,N_28807,N_29633);
and U31212 (N_31212,N_29500,N_28267);
nor U31213 (N_31213,N_29642,N_29867);
or U31214 (N_31214,N_29400,N_28987);
or U31215 (N_31215,N_28153,N_28704);
nor U31216 (N_31216,N_28401,N_28259);
and U31217 (N_31217,N_29106,N_28550);
and U31218 (N_31218,N_29818,N_29850);
nand U31219 (N_31219,N_28624,N_29597);
nand U31220 (N_31220,N_28617,N_28511);
and U31221 (N_31221,N_29752,N_29841);
nor U31222 (N_31222,N_29202,N_29097);
and U31223 (N_31223,N_28019,N_29380);
and U31224 (N_31224,N_29525,N_28666);
nand U31225 (N_31225,N_28299,N_29200);
xnor U31226 (N_31226,N_29198,N_29095);
and U31227 (N_31227,N_28411,N_29596);
and U31228 (N_31228,N_28577,N_29079);
and U31229 (N_31229,N_29366,N_28710);
nor U31230 (N_31230,N_29900,N_28293);
and U31231 (N_31231,N_28162,N_28725);
xor U31232 (N_31232,N_28016,N_28308);
nor U31233 (N_31233,N_29390,N_28872);
nand U31234 (N_31234,N_28763,N_28364);
nor U31235 (N_31235,N_28013,N_29800);
xnor U31236 (N_31236,N_29027,N_28031);
nand U31237 (N_31237,N_28805,N_29479);
nand U31238 (N_31238,N_28801,N_28864);
and U31239 (N_31239,N_29142,N_28940);
xnor U31240 (N_31240,N_29639,N_28761);
xor U31241 (N_31241,N_28147,N_29317);
nor U31242 (N_31242,N_28845,N_28302);
xnor U31243 (N_31243,N_29706,N_28118);
nor U31244 (N_31244,N_29446,N_28284);
nand U31245 (N_31245,N_29179,N_28296);
xnor U31246 (N_31246,N_29138,N_28122);
nand U31247 (N_31247,N_29245,N_28208);
nand U31248 (N_31248,N_28866,N_29643);
nand U31249 (N_31249,N_28393,N_28728);
or U31250 (N_31250,N_28204,N_29167);
nor U31251 (N_31251,N_28964,N_29503);
xnor U31252 (N_31252,N_28791,N_28959);
nand U31253 (N_31253,N_28976,N_29231);
or U31254 (N_31254,N_29299,N_28158);
and U31255 (N_31255,N_29845,N_28978);
and U31256 (N_31256,N_28389,N_28187);
xor U31257 (N_31257,N_28254,N_28661);
and U31258 (N_31258,N_28200,N_28763);
nand U31259 (N_31259,N_29623,N_29421);
nor U31260 (N_31260,N_29472,N_28895);
and U31261 (N_31261,N_29838,N_29733);
and U31262 (N_31262,N_29321,N_28360);
nand U31263 (N_31263,N_28535,N_29008);
xnor U31264 (N_31264,N_28257,N_28757);
nand U31265 (N_31265,N_29348,N_29878);
or U31266 (N_31266,N_28395,N_28249);
and U31267 (N_31267,N_28889,N_28322);
or U31268 (N_31268,N_29623,N_29152);
and U31269 (N_31269,N_28797,N_28043);
or U31270 (N_31270,N_28253,N_28851);
xor U31271 (N_31271,N_29349,N_28565);
nor U31272 (N_31272,N_29652,N_29098);
or U31273 (N_31273,N_28771,N_28927);
nand U31274 (N_31274,N_29144,N_29559);
nor U31275 (N_31275,N_28305,N_28777);
or U31276 (N_31276,N_28545,N_28202);
nor U31277 (N_31277,N_29177,N_28544);
and U31278 (N_31278,N_29689,N_28602);
xnor U31279 (N_31279,N_29755,N_28971);
and U31280 (N_31280,N_29185,N_29350);
nand U31281 (N_31281,N_28315,N_29716);
nor U31282 (N_31282,N_28955,N_29633);
nor U31283 (N_31283,N_28443,N_28630);
xnor U31284 (N_31284,N_28205,N_29486);
nor U31285 (N_31285,N_28133,N_29399);
or U31286 (N_31286,N_29620,N_29176);
nor U31287 (N_31287,N_28122,N_29396);
or U31288 (N_31288,N_28831,N_28686);
and U31289 (N_31289,N_28472,N_29503);
xnor U31290 (N_31290,N_29221,N_29968);
nor U31291 (N_31291,N_29338,N_28299);
nor U31292 (N_31292,N_29439,N_29313);
nand U31293 (N_31293,N_28761,N_28294);
xnor U31294 (N_31294,N_29400,N_29892);
nor U31295 (N_31295,N_29053,N_28460);
nor U31296 (N_31296,N_28547,N_29524);
and U31297 (N_31297,N_28017,N_28002);
nor U31298 (N_31298,N_29480,N_28579);
nor U31299 (N_31299,N_28213,N_29462);
or U31300 (N_31300,N_28892,N_29574);
xnor U31301 (N_31301,N_28896,N_29591);
nand U31302 (N_31302,N_29115,N_29108);
nand U31303 (N_31303,N_28028,N_29508);
and U31304 (N_31304,N_29580,N_29501);
or U31305 (N_31305,N_29816,N_28944);
nor U31306 (N_31306,N_29440,N_29941);
xor U31307 (N_31307,N_28562,N_29866);
and U31308 (N_31308,N_29103,N_28069);
and U31309 (N_31309,N_28319,N_28868);
or U31310 (N_31310,N_29409,N_28373);
xnor U31311 (N_31311,N_29274,N_29099);
and U31312 (N_31312,N_28390,N_28137);
and U31313 (N_31313,N_29788,N_29246);
nor U31314 (N_31314,N_28878,N_28512);
or U31315 (N_31315,N_29469,N_28416);
or U31316 (N_31316,N_29897,N_29990);
nor U31317 (N_31317,N_29458,N_29768);
or U31318 (N_31318,N_29773,N_28748);
nor U31319 (N_31319,N_29656,N_28423);
or U31320 (N_31320,N_29758,N_29350);
and U31321 (N_31321,N_28335,N_28256);
and U31322 (N_31322,N_28954,N_29272);
nor U31323 (N_31323,N_28257,N_28661);
or U31324 (N_31324,N_29828,N_29493);
and U31325 (N_31325,N_28400,N_29490);
and U31326 (N_31326,N_29031,N_28267);
nor U31327 (N_31327,N_29601,N_28977);
nand U31328 (N_31328,N_28212,N_29492);
nor U31329 (N_31329,N_29324,N_28334);
nand U31330 (N_31330,N_29126,N_28996);
nand U31331 (N_31331,N_28063,N_29093);
and U31332 (N_31332,N_28849,N_28402);
and U31333 (N_31333,N_29528,N_28028);
xor U31334 (N_31334,N_29279,N_29238);
and U31335 (N_31335,N_28298,N_28621);
nor U31336 (N_31336,N_29210,N_29481);
nand U31337 (N_31337,N_29030,N_28056);
xnor U31338 (N_31338,N_29563,N_28692);
or U31339 (N_31339,N_29144,N_28735);
nand U31340 (N_31340,N_28999,N_28636);
nor U31341 (N_31341,N_28432,N_29904);
and U31342 (N_31342,N_29687,N_28343);
and U31343 (N_31343,N_28184,N_29185);
xor U31344 (N_31344,N_29246,N_28766);
or U31345 (N_31345,N_28761,N_29367);
xor U31346 (N_31346,N_29053,N_29086);
nand U31347 (N_31347,N_28033,N_28169);
and U31348 (N_31348,N_29102,N_29699);
and U31349 (N_31349,N_28363,N_28533);
nand U31350 (N_31350,N_28014,N_28370);
or U31351 (N_31351,N_28211,N_29402);
xnor U31352 (N_31352,N_28201,N_29890);
or U31353 (N_31353,N_29924,N_29915);
or U31354 (N_31354,N_28680,N_28206);
nand U31355 (N_31355,N_28781,N_29905);
and U31356 (N_31356,N_29255,N_28016);
nor U31357 (N_31357,N_29157,N_28404);
or U31358 (N_31358,N_28827,N_29101);
and U31359 (N_31359,N_28730,N_28593);
and U31360 (N_31360,N_28945,N_29861);
nor U31361 (N_31361,N_29289,N_28752);
and U31362 (N_31362,N_29017,N_29763);
or U31363 (N_31363,N_29198,N_28237);
nor U31364 (N_31364,N_28550,N_28952);
or U31365 (N_31365,N_29050,N_28564);
or U31366 (N_31366,N_29028,N_29390);
or U31367 (N_31367,N_29863,N_29551);
xnor U31368 (N_31368,N_28488,N_29351);
nand U31369 (N_31369,N_28032,N_28470);
nor U31370 (N_31370,N_28517,N_28850);
and U31371 (N_31371,N_28968,N_29986);
nand U31372 (N_31372,N_29697,N_29041);
and U31373 (N_31373,N_28433,N_29204);
and U31374 (N_31374,N_29509,N_29337);
or U31375 (N_31375,N_28381,N_29332);
and U31376 (N_31376,N_29889,N_29516);
or U31377 (N_31377,N_28589,N_29354);
and U31378 (N_31378,N_29942,N_29714);
nand U31379 (N_31379,N_29732,N_28675);
and U31380 (N_31380,N_29806,N_28366);
nor U31381 (N_31381,N_28274,N_28352);
nand U31382 (N_31382,N_28989,N_29958);
nor U31383 (N_31383,N_29205,N_28683);
and U31384 (N_31384,N_29483,N_28302);
nand U31385 (N_31385,N_29543,N_29944);
or U31386 (N_31386,N_28342,N_29665);
or U31387 (N_31387,N_28527,N_29934);
nor U31388 (N_31388,N_28287,N_29290);
xnor U31389 (N_31389,N_28452,N_28407);
nor U31390 (N_31390,N_29317,N_29581);
xor U31391 (N_31391,N_28822,N_29757);
nand U31392 (N_31392,N_28180,N_29602);
nor U31393 (N_31393,N_29419,N_29800);
nand U31394 (N_31394,N_28196,N_29839);
nand U31395 (N_31395,N_29878,N_29068);
or U31396 (N_31396,N_29629,N_28870);
nand U31397 (N_31397,N_29864,N_29921);
nor U31398 (N_31398,N_29785,N_29974);
xor U31399 (N_31399,N_28234,N_29000);
nand U31400 (N_31400,N_28300,N_29022);
nand U31401 (N_31401,N_28410,N_28980);
nor U31402 (N_31402,N_29469,N_29343);
nand U31403 (N_31403,N_28538,N_29827);
and U31404 (N_31404,N_28875,N_28849);
xor U31405 (N_31405,N_28115,N_28149);
nor U31406 (N_31406,N_29848,N_28418);
and U31407 (N_31407,N_28903,N_28464);
xnor U31408 (N_31408,N_29766,N_29236);
nand U31409 (N_31409,N_29500,N_28356);
nor U31410 (N_31410,N_28309,N_28120);
and U31411 (N_31411,N_28089,N_28823);
nand U31412 (N_31412,N_28295,N_29498);
or U31413 (N_31413,N_29504,N_29163);
or U31414 (N_31414,N_29046,N_29007);
or U31415 (N_31415,N_29760,N_28586);
xnor U31416 (N_31416,N_28686,N_29095);
and U31417 (N_31417,N_29939,N_28577);
or U31418 (N_31418,N_29056,N_29763);
nor U31419 (N_31419,N_28461,N_29117);
or U31420 (N_31420,N_29453,N_29135);
and U31421 (N_31421,N_29437,N_29868);
or U31422 (N_31422,N_29231,N_28228);
or U31423 (N_31423,N_29609,N_28028);
or U31424 (N_31424,N_28025,N_29887);
nand U31425 (N_31425,N_29169,N_28800);
nor U31426 (N_31426,N_29846,N_29405);
nor U31427 (N_31427,N_29353,N_29276);
nand U31428 (N_31428,N_29795,N_29057);
nand U31429 (N_31429,N_29499,N_29291);
nor U31430 (N_31430,N_28548,N_29626);
nand U31431 (N_31431,N_29172,N_28467);
and U31432 (N_31432,N_29478,N_28079);
or U31433 (N_31433,N_28517,N_28263);
nand U31434 (N_31434,N_29589,N_28123);
and U31435 (N_31435,N_28024,N_29928);
nand U31436 (N_31436,N_29858,N_29536);
nor U31437 (N_31437,N_28572,N_28054);
or U31438 (N_31438,N_29092,N_28065);
nand U31439 (N_31439,N_29188,N_29560);
or U31440 (N_31440,N_29319,N_29121);
and U31441 (N_31441,N_28498,N_28279);
xnor U31442 (N_31442,N_29113,N_28139);
or U31443 (N_31443,N_29063,N_29872);
and U31444 (N_31444,N_28042,N_29981);
or U31445 (N_31445,N_28293,N_28736);
nor U31446 (N_31446,N_29596,N_28563);
nor U31447 (N_31447,N_29202,N_28608);
nor U31448 (N_31448,N_29936,N_28382);
nand U31449 (N_31449,N_28460,N_28232);
nand U31450 (N_31450,N_29447,N_29936);
and U31451 (N_31451,N_29136,N_28223);
nand U31452 (N_31452,N_29750,N_29677);
nor U31453 (N_31453,N_28610,N_29053);
nand U31454 (N_31454,N_28292,N_28029);
or U31455 (N_31455,N_28621,N_29451);
xnor U31456 (N_31456,N_28702,N_29626);
and U31457 (N_31457,N_28113,N_28093);
and U31458 (N_31458,N_28655,N_29495);
nand U31459 (N_31459,N_29629,N_29161);
nand U31460 (N_31460,N_29318,N_28910);
xor U31461 (N_31461,N_29615,N_29904);
nor U31462 (N_31462,N_29545,N_29850);
and U31463 (N_31463,N_28784,N_28482);
nor U31464 (N_31464,N_28607,N_29802);
nand U31465 (N_31465,N_28501,N_29914);
nand U31466 (N_31466,N_29307,N_29394);
and U31467 (N_31467,N_28464,N_29512);
or U31468 (N_31468,N_28776,N_29683);
and U31469 (N_31469,N_28953,N_28408);
xnor U31470 (N_31470,N_28991,N_28191);
xnor U31471 (N_31471,N_28418,N_28003);
or U31472 (N_31472,N_28350,N_28395);
xor U31473 (N_31473,N_29979,N_28157);
or U31474 (N_31474,N_28913,N_29027);
or U31475 (N_31475,N_28455,N_29230);
and U31476 (N_31476,N_28740,N_29957);
xnor U31477 (N_31477,N_29314,N_28713);
nor U31478 (N_31478,N_29251,N_29167);
nor U31479 (N_31479,N_28912,N_29184);
xor U31480 (N_31480,N_29429,N_29949);
xnor U31481 (N_31481,N_28024,N_29270);
nand U31482 (N_31482,N_28206,N_29235);
or U31483 (N_31483,N_28687,N_28444);
nor U31484 (N_31484,N_29591,N_28136);
or U31485 (N_31485,N_29161,N_29211);
or U31486 (N_31486,N_29970,N_29203);
xnor U31487 (N_31487,N_29582,N_29301);
and U31488 (N_31488,N_28184,N_29207);
xor U31489 (N_31489,N_28884,N_28278);
xor U31490 (N_31490,N_28966,N_28710);
nor U31491 (N_31491,N_29924,N_28011);
xnor U31492 (N_31492,N_29808,N_29101);
nor U31493 (N_31493,N_29030,N_28320);
nand U31494 (N_31494,N_29619,N_28464);
nand U31495 (N_31495,N_29608,N_29306);
and U31496 (N_31496,N_29313,N_28181);
xnor U31497 (N_31497,N_28848,N_29211);
and U31498 (N_31498,N_28091,N_29965);
nor U31499 (N_31499,N_29989,N_29436);
nor U31500 (N_31500,N_28149,N_29904);
nor U31501 (N_31501,N_28814,N_28194);
nor U31502 (N_31502,N_29875,N_28391);
nand U31503 (N_31503,N_28539,N_29597);
nand U31504 (N_31504,N_28363,N_29594);
and U31505 (N_31505,N_29595,N_28785);
xor U31506 (N_31506,N_29662,N_28238);
and U31507 (N_31507,N_28568,N_29543);
nand U31508 (N_31508,N_29046,N_28717);
nand U31509 (N_31509,N_29610,N_28381);
xnor U31510 (N_31510,N_28118,N_28427);
nor U31511 (N_31511,N_28853,N_29093);
nor U31512 (N_31512,N_29165,N_29780);
xor U31513 (N_31513,N_28465,N_28275);
and U31514 (N_31514,N_29089,N_29889);
or U31515 (N_31515,N_28032,N_29609);
and U31516 (N_31516,N_28531,N_28249);
nor U31517 (N_31517,N_28957,N_28817);
or U31518 (N_31518,N_29162,N_29027);
or U31519 (N_31519,N_28290,N_28218);
or U31520 (N_31520,N_28347,N_28348);
nand U31521 (N_31521,N_28825,N_28141);
nand U31522 (N_31522,N_29197,N_29088);
nor U31523 (N_31523,N_29771,N_28757);
nor U31524 (N_31524,N_28906,N_28097);
nand U31525 (N_31525,N_29431,N_28506);
xor U31526 (N_31526,N_28863,N_28142);
and U31527 (N_31527,N_28202,N_29380);
or U31528 (N_31528,N_29880,N_29538);
nand U31529 (N_31529,N_29332,N_29044);
and U31530 (N_31530,N_28552,N_29491);
or U31531 (N_31531,N_28596,N_29484);
or U31532 (N_31532,N_28810,N_29119);
nand U31533 (N_31533,N_28611,N_28517);
nor U31534 (N_31534,N_28870,N_29232);
xor U31535 (N_31535,N_29661,N_28220);
nand U31536 (N_31536,N_29006,N_29673);
nor U31537 (N_31537,N_28625,N_29654);
and U31538 (N_31538,N_28261,N_29601);
and U31539 (N_31539,N_28725,N_28172);
nand U31540 (N_31540,N_29647,N_29465);
nand U31541 (N_31541,N_29060,N_29327);
xnor U31542 (N_31542,N_28576,N_29515);
nand U31543 (N_31543,N_28435,N_29018);
nand U31544 (N_31544,N_29795,N_28917);
xnor U31545 (N_31545,N_29274,N_28620);
xor U31546 (N_31546,N_29960,N_28309);
nor U31547 (N_31547,N_28523,N_29447);
nand U31548 (N_31548,N_29317,N_28851);
or U31549 (N_31549,N_28636,N_29128);
nor U31550 (N_31550,N_29568,N_28657);
or U31551 (N_31551,N_28521,N_29853);
nand U31552 (N_31552,N_28470,N_29381);
and U31553 (N_31553,N_28665,N_28077);
xor U31554 (N_31554,N_29734,N_28338);
and U31555 (N_31555,N_28023,N_28461);
xor U31556 (N_31556,N_29610,N_29116);
and U31557 (N_31557,N_28097,N_29606);
nor U31558 (N_31558,N_29651,N_29381);
nor U31559 (N_31559,N_28107,N_28102);
or U31560 (N_31560,N_28692,N_28896);
or U31561 (N_31561,N_28656,N_29332);
and U31562 (N_31562,N_28333,N_28036);
and U31563 (N_31563,N_28331,N_28204);
or U31564 (N_31564,N_28355,N_28887);
or U31565 (N_31565,N_28891,N_29630);
nor U31566 (N_31566,N_29070,N_29947);
and U31567 (N_31567,N_29412,N_29726);
or U31568 (N_31568,N_28497,N_28558);
nor U31569 (N_31569,N_29244,N_28228);
nor U31570 (N_31570,N_29225,N_29728);
and U31571 (N_31571,N_28956,N_28701);
and U31572 (N_31572,N_28711,N_28885);
and U31573 (N_31573,N_29062,N_28286);
or U31574 (N_31574,N_29584,N_29528);
xor U31575 (N_31575,N_29066,N_28131);
nand U31576 (N_31576,N_29762,N_29616);
or U31577 (N_31577,N_29439,N_29003);
nor U31578 (N_31578,N_29528,N_29348);
nor U31579 (N_31579,N_29366,N_29003);
or U31580 (N_31580,N_29214,N_28355);
and U31581 (N_31581,N_28039,N_28120);
xor U31582 (N_31582,N_28446,N_28966);
nor U31583 (N_31583,N_28133,N_29602);
xnor U31584 (N_31584,N_28530,N_28233);
nand U31585 (N_31585,N_29218,N_28486);
nand U31586 (N_31586,N_29252,N_29329);
nor U31587 (N_31587,N_28810,N_28065);
xnor U31588 (N_31588,N_28729,N_28301);
nand U31589 (N_31589,N_29889,N_29878);
xor U31590 (N_31590,N_29297,N_28454);
xnor U31591 (N_31591,N_29592,N_29269);
or U31592 (N_31592,N_29778,N_29510);
and U31593 (N_31593,N_29314,N_28560);
nand U31594 (N_31594,N_29546,N_28702);
nand U31595 (N_31595,N_28766,N_28475);
xor U31596 (N_31596,N_28231,N_28427);
or U31597 (N_31597,N_29770,N_29866);
or U31598 (N_31598,N_28390,N_28859);
xor U31599 (N_31599,N_28914,N_28122);
or U31600 (N_31600,N_29561,N_28000);
or U31601 (N_31601,N_28904,N_29517);
or U31602 (N_31602,N_28316,N_28775);
nor U31603 (N_31603,N_29497,N_28857);
or U31604 (N_31604,N_28964,N_28816);
nor U31605 (N_31605,N_28617,N_28837);
xnor U31606 (N_31606,N_29813,N_29606);
or U31607 (N_31607,N_29041,N_28775);
nor U31608 (N_31608,N_28785,N_29785);
and U31609 (N_31609,N_28733,N_28803);
nor U31610 (N_31610,N_29762,N_28823);
nor U31611 (N_31611,N_28137,N_29693);
xnor U31612 (N_31612,N_28349,N_28515);
nand U31613 (N_31613,N_29233,N_28239);
nor U31614 (N_31614,N_29112,N_29990);
nand U31615 (N_31615,N_28247,N_29421);
xnor U31616 (N_31616,N_28133,N_29959);
xnor U31617 (N_31617,N_28618,N_29408);
and U31618 (N_31618,N_28929,N_28591);
or U31619 (N_31619,N_28666,N_28815);
nor U31620 (N_31620,N_29902,N_28659);
and U31621 (N_31621,N_28194,N_28503);
nor U31622 (N_31622,N_28203,N_28341);
xor U31623 (N_31623,N_28820,N_29423);
xor U31624 (N_31624,N_28348,N_28211);
xor U31625 (N_31625,N_29953,N_29151);
or U31626 (N_31626,N_29230,N_29391);
or U31627 (N_31627,N_29272,N_28271);
nand U31628 (N_31628,N_28838,N_29812);
nor U31629 (N_31629,N_29117,N_29879);
xor U31630 (N_31630,N_29104,N_28795);
nor U31631 (N_31631,N_29947,N_29051);
xor U31632 (N_31632,N_29111,N_29676);
nor U31633 (N_31633,N_28625,N_28299);
and U31634 (N_31634,N_29819,N_29162);
nand U31635 (N_31635,N_29504,N_29999);
xor U31636 (N_31636,N_28255,N_28158);
nand U31637 (N_31637,N_29757,N_29971);
or U31638 (N_31638,N_28708,N_29848);
nor U31639 (N_31639,N_28081,N_28463);
nand U31640 (N_31640,N_28282,N_28126);
and U31641 (N_31641,N_29182,N_28730);
and U31642 (N_31642,N_28447,N_28613);
nor U31643 (N_31643,N_29549,N_29964);
nor U31644 (N_31644,N_29475,N_28322);
nor U31645 (N_31645,N_29811,N_28549);
and U31646 (N_31646,N_29287,N_28024);
xnor U31647 (N_31647,N_29716,N_28086);
nand U31648 (N_31648,N_29244,N_28310);
nand U31649 (N_31649,N_29379,N_29791);
or U31650 (N_31650,N_29633,N_28682);
and U31651 (N_31651,N_28649,N_29775);
nor U31652 (N_31652,N_29240,N_28512);
nand U31653 (N_31653,N_28539,N_28392);
nor U31654 (N_31654,N_29758,N_28986);
xnor U31655 (N_31655,N_29825,N_29880);
and U31656 (N_31656,N_29746,N_29039);
xor U31657 (N_31657,N_29546,N_28550);
nand U31658 (N_31658,N_28622,N_28305);
xnor U31659 (N_31659,N_28508,N_28564);
nand U31660 (N_31660,N_28782,N_28700);
and U31661 (N_31661,N_28288,N_28747);
nand U31662 (N_31662,N_29873,N_28977);
and U31663 (N_31663,N_29217,N_29823);
or U31664 (N_31664,N_29290,N_29436);
nor U31665 (N_31665,N_29764,N_29630);
and U31666 (N_31666,N_29429,N_28952);
xor U31667 (N_31667,N_28843,N_28278);
xor U31668 (N_31668,N_28245,N_29309);
xnor U31669 (N_31669,N_29777,N_29144);
and U31670 (N_31670,N_28380,N_29962);
or U31671 (N_31671,N_28414,N_29250);
xnor U31672 (N_31672,N_29254,N_29838);
xor U31673 (N_31673,N_29358,N_28271);
or U31674 (N_31674,N_28175,N_28201);
xor U31675 (N_31675,N_28821,N_29485);
xnor U31676 (N_31676,N_29391,N_29601);
or U31677 (N_31677,N_28812,N_28415);
nand U31678 (N_31678,N_29531,N_28336);
nor U31679 (N_31679,N_29411,N_29332);
and U31680 (N_31680,N_28661,N_28958);
nand U31681 (N_31681,N_29249,N_29101);
nor U31682 (N_31682,N_29874,N_29659);
nor U31683 (N_31683,N_28176,N_29825);
or U31684 (N_31684,N_29471,N_28275);
or U31685 (N_31685,N_29227,N_28451);
nor U31686 (N_31686,N_28593,N_29225);
xnor U31687 (N_31687,N_29965,N_29497);
nand U31688 (N_31688,N_29197,N_29676);
and U31689 (N_31689,N_29607,N_28958);
and U31690 (N_31690,N_29167,N_29133);
or U31691 (N_31691,N_28922,N_28750);
and U31692 (N_31692,N_29565,N_28524);
nor U31693 (N_31693,N_29112,N_29870);
and U31694 (N_31694,N_29804,N_29512);
nor U31695 (N_31695,N_28121,N_29625);
xor U31696 (N_31696,N_28148,N_28861);
or U31697 (N_31697,N_28625,N_29583);
nand U31698 (N_31698,N_29283,N_28018);
xor U31699 (N_31699,N_28479,N_29846);
nor U31700 (N_31700,N_29185,N_28213);
xnor U31701 (N_31701,N_28549,N_28401);
nand U31702 (N_31702,N_28749,N_28699);
nand U31703 (N_31703,N_29391,N_29287);
xnor U31704 (N_31704,N_28781,N_28151);
and U31705 (N_31705,N_29399,N_29113);
xnor U31706 (N_31706,N_29392,N_28733);
and U31707 (N_31707,N_28564,N_28850);
or U31708 (N_31708,N_28102,N_29958);
xor U31709 (N_31709,N_28688,N_28730);
nand U31710 (N_31710,N_29243,N_29967);
and U31711 (N_31711,N_29947,N_28686);
xor U31712 (N_31712,N_29921,N_29347);
xor U31713 (N_31713,N_29300,N_28733);
or U31714 (N_31714,N_28086,N_29292);
or U31715 (N_31715,N_28956,N_29177);
nand U31716 (N_31716,N_29553,N_28262);
xor U31717 (N_31717,N_29195,N_28860);
nand U31718 (N_31718,N_28509,N_29501);
nor U31719 (N_31719,N_29784,N_28043);
nand U31720 (N_31720,N_28694,N_29687);
nand U31721 (N_31721,N_28869,N_29826);
or U31722 (N_31722,N_28737,N_29764);
or U31723 (N_31723,N_28353,N_28288);
or U31724 (N_31724,N_29457,N_28445);
xor U31725 (N_31725,N_28829,N_28481);
or U31726 (N_31726,N_28893,N_29276);
or U31727 (N_31727,N_28200,N_29119);
or U31728 (N_31728,N_28090,N_28636);
or U31729 (N_31729,N_28920,N_29211);
xor U31730 (N_31730,N_28956,N_28066);
nand U31731 (N_31731,N_28039,N_29815);
nor U31732 (N_31732,N_28652,N_28668);
xor U31733 (N_31733,N_28370,N_28809);
xnor U31734 (N_31734,N_29766,N_29915);
nand U31735 (N_31735,N_28607,N_29653);
xor U31736 (N_31736,N_28244,N_29912);
xnor U31737 (N_31737,N_28809,N_29577);
nand U31738 (N_31738,N_29008,N_29881);
and U31739 (N_31739,N_28429,N_28712);
xor U31740 (N_31740,N_29288,N_29433);
and U31741 (N_31741,N_28799,N_28115);
xor U31742 (N_31742,N_29601,N_28774);
xor U31743 (N_31743,N_28147,N_28539);
xnor U31744 (N_31744,N_29523,N_28427);
nand U31745 (N_31745,N_29976,N_28286);
xnor U31746 (N_31746,N_29411,N_29009);
xor U31747 (N_31747,N_28470,N_29358);
and U31748 (N_31748,N_28507,N_28671);
or U31749 (N_31749,N_28709,N_29849);
nand U31750 (N_31750,N_28067,N_28651);
or U31751 (N_31751,N_29586,N_29748);
nand U31752 (N_31752,N_28055,N_28144);
and U31753 (N_31753,N_28151,N_29828);
nand U31754 (N_31754,N_28799,N_29943);
nand U31755 (N_31755,N_29425,N_29297);
or U31756 (N_31756,N_28957,N_29290);
or U31757 (N_31757,N_29122,N_28088);
nand U31758 (N_31758,N_28980,N_28804);
and U31759 (N_31759,N_29820,N_29603);
nand U31760 (N_31760,N_29674,N_28498);
nor U31761 (N_31761,N_28608,N_28139);
xnor U31762 (N_31762,N_29492,N_29357);
nor U31763 (N_31763,N_29498,N_28438);
or U31764 (N_31764,N_28651,N_28392);
xnor U31765 (N_31765,N_28638,N_28221);
nor U31766 (N_31766,N_29406,N_28943);
and U31767 (N_31767,N_29283,N_28919);
and U31768 (N_31768,N_28696,N_28128);
nand U31769 (N_31769,N_29507,N_29972);
nand U31770 (N_31770,N_28067,N_28430);
nand U31771 (N_31771,N_29549,N_28772);
and U31772 (N_31772,N_29918,N_29635);
xor U31773 (N_31773,N_29989,N_28728);
and U31774 (N_31774,N_29469,N_28510);
xnor U31775 (N_31775,N_29212,N_29385);
or U31776 (N_31776,N_28675,N_28807);
xnor U31777 (N_31777,N_28687,N_28565);
or U31778 (N_31778,N_28798,N_29875);
or U31779 (N_31779,N_28343,N_28318);
nand U31780 (N_31780,N_28151,N_29358);
and U31781 (N_31781,N_29609,N_29223);
nand U31782 (N_31782,N_29207,N_28084);
xor U31783 (N_31783,N_29835,N_29531);
xor U31784 (N_31784,N_28286,N_29508);
and U31785 (N_31785,N_28331,N_29067);
or U31786 (N_31786,N_29917,N_28452);
xnor U31787 (N_31787,N_29327,N_28181);
and U31788 (N_31788,N_28425,N_29896);
nand U31789 (N_31789,N_29605,N_28503);
nand U31790 (N_31790,N_28436,N_28819);
nand U31791 (N_31791,N_28751,N_28733);
xnor U31792 (N_31792,N_29703,N_28639);
and U31793 (N_31793,N_28050,N_29259);
nor U31794 (N_31794,N_29089,N_29466);
or U31795 (N_31795,N_28003,N_29381);
and U31796 (N_31796,N_29657,N_29431);
or U31797 (N_31797,N_29204,N_28611);
xor U31798 (N_31798,N_28360,N_28936);
nor U31799 (N_31799,N_29142,N_29855);
xnor U31800 (N_31800,N_28985,N_28398);
nor U31801 (N_31801,N_29811,N_28100);
xnor U31802 (N_31802,N_28773,N_28921);
or U31803 (N_31803,N_28152,N_29546);
xnor U31804 (N_31804,N_28175,N_28581);
nand U31805 (N_31805,N_29943,N_29355);
nor U31806 (N_31806,N_29046,N_29672);
xnor U31807 (N_31807,N_29211,N_29753);
nor U31808 (N_31808,N_29639,N_29480);
xnor U31809 (N_31809,N_28338,N_29773);
xor U31810 (N_31810,N_29994,N_29426);
xnor U31811 (N_31811,N_28990,N_28617);
and U31812 (N_31812,N_28303,N_28773);
nor U31813 (N_31813,N_29512,N_29508);
and U31814 (N_31814,N_29093,N_28827);
xor U31815 (N_31815,N_28756,N_28885);
nor U31816 (N_31816,N_28447,N_28953);
xor U31817 (N_31817,N_29957,N_29172);
and U31818 (N_31818,N_28058,N_28071);
xor U31819 (N_31819,N_28550,N_28685);
xor U31820 (N_31820,N_28417,N_29114);
or U31821 (N_31821,N_29810,N_29385);
or U31822 (N_31822,N_28501,N_29834);
xnor U31823 (N_31823,N_29504,N_29141);
xnor U31824 (N_31824,N_28638,N_28137);
nand U31825 (N_31825,N_28237,N_28776);
or U31826 (N_31826,N_28356,N_29065);
nor U31827 (N_31827,N_29953,N_28849);
nor U31828 (N_31828,N_28538,N_29555);
nor U31829 (N_31829,N_28787,N_29906);
nor U31830 (N_31830,N_29662,N_29784);
xor U31831 (N_31831,N_29762,N_28935);
nor U31832 (N_31832,N_29816,N_29771);
and U31833 (N_31833,N_29489,N_28482);
xnor U31834 (N_31834,N_28825,N_29884);
xor U31835 (N_31835,N_29491,N_28285);
and U31836 (N_31836,N_29178,N_29717);
nor U31837 (N_31837,N_28580,N_29675);
xnor U31838 (N_31838,N_28016,N_28887);
or U31839 (N_31839,N_28111,N_28112);
or U31840 (N_31840,N_29496,N_28714);
or U31841 (N_31841,N_28669,N_28652);
nand U31842 (N_31842,N_29096,N_28525);
nand U31843 (N_31843,N_29078,N_29370);
nor U31844 (N_31844,N_29280,N_28625);
xor U31845 (N_31845,N_28488,N_29750);
nand U31846 (N_31846,N_28912,N_28517);
xor U31847 (N_31847,N_29766,N_28549);
nor U31848 (N_31848,N_28643,N_29612);
xnor U31849 (N_31849,N_29433,N_29859);
xnor U31850 (N_31850,N_29891,N_28987);
nor U31851 (N_31851,N_29840,N_29039);
and U31852 (N_31852,N_29675,N_29225);
nand U31853 (N_31853,N_28732,N_29371);
and U31854 (N_31854,N_28280,N_28526);
xor U31855 (N_31855,N_28596,N_29725);
and U31856 (N_31856,N_28906,N_28623);
and U31857 (N_31857,N_28018,N_29204);
nor U31858 (N_31858,N_29071,N_29910);
and U31859 (N_31859,N_29949,N_29774);
and U31860 (N_31860,N_28750,N_29948);
nand U31861 (N_31861,N_28633,N_29955);
nand U31862 (N_31862,N_29130,N_29523);
or U31863 (N_31863,N_28816,N_28848);
nand U31864 (N_31864,N_28792,N_28648);
nor U31865 (N_31865,N_29382,N_28705);
nor U31866 (N_31866,N_29626,N_28519);
and U31867 (N_31867,N_28252,N_28535);
nor U31868 (N_31868,N_28323,N_28875);
xor U31869 (N_31869,N_29808,N_28231);
or U31870 (N_31870,N_29149,N_29049);
nor U31871 (N_31871,N_29322,N_28725);
nor U31872 (N_31872,N_29625,N_28008);
nand U31873 (N_31873,N_29646,N_28458);
xnor U31874 (N_31874,N_29669,N_28829);
or U31875 (N_31875,N_28143,N_29248);
nand U31876 (N_31876,N_28212,N_29740);
xnor U31877 (N_31877,N_28443,N_29773);
nand U31878 (N_31878,N_29250,N_28999);
nor U31879 (N_31879,N_29939,N_28966);
xor U31880 (N_31880,N_28762,N_29113);
or U31881 (N_31881,N_28391,N_29134);
xnor U31882 (N_31882,N_28015,N_29693);
nand U31883 (N_31883,N_29192,N_29345);
and U31884 (N_31884,N_29429,N_29774);
nand U31885 (N_31885,N_29217,N_29496);
xor U31886 (N_31886,N_28294,N_28507);
or U31887 (N_31887,N_28062,N_28430);
nor U31888 (N_31888,N_28203,N_28435);
xnor U31889 (N_31889,N_29759,N_29751);
or U31890 (N_31890,N_28018,N_28189);
and U31891 (N_31891,N_29352,N_28959);
xor U31892 (N_31892,N_28130,N_29357);
nor U31893 (N_31893,N_28561,N_29435);
or U31894 (N_31894,N_29515,N_28886);
or U31895 (N_31895,N_28167,N_28302);
or U31896 (N_31896,N_28148,N_28100);
nor U31897 (N_31897,N_28617,N_29127);
and U31898 (N_31898,N_28294,N_29931);
xnor U31899 (N_31899,N_28843,N_28255);
nand U31900 (N_31900,N_28527,N_28591);
nand U31901 (N_31901,N_28943,N_29450);
nand U31902 (N_31902,N_28385,N_29711);
xor U31903 (N_31903,N_29269,N_28823);
nand U31904 (N_31904,N_29680,N_28100);
and U31905 (N_31905,N_28933,N_29567);
nand U31906 (N_31906,N_29597,N_29523);
nand U31907 (N_31907,N_28423,N_29808);
nand U31908 (N_31908,N_28640,N_29414);
and U31909 (N_31909,N_28626,N_29327);
nor U31910 (N_31910,N_29805,N_29142);
xor U31911 (N_31911,N_29460,N_28994);
xor U31912 (N_31912,N_28783,N_28155);
nand U31913 (N_31913,N_28306,N_29759);
xor U31914 (N_31914,N_28307,N_29744);
xnor U31915 (N_31915,N_29571,N_28027);
xor U31916 (N_31916,N_28691,N_28751);
nand U31917 (N_31917,N_29329,N_29049);
xnor U31918 (N_31918,N_28013,N_28992);
nand U31919 (N_31919,N_29079,N_28819);
or U31920 (N_31920,N_28534,N_29646);
and U31921 (N_31921,N_28953,N_29257);
nor U31922 (N_31922,N_28544,N_29219);
or U31923 (N_31923,N_29301,N_29842);
nand U31924 (N_31924,N_29799,N_29750);
and U31925 (N_31925,N_29462,N_28499);
or U31926 (N_31926,N_29145,N_29017);
and U31927 (N_31927,N_29380,N_29207);
nor U31928 (N_31928,N_29361,N_29937);
nand U31929 (N_31929,N_29501,N_28891);
nand U31930 (N_31930,N_29784,N_28133);
nor U31931 (N_31931,N_28205,N_29578);
xnor U31932 (N_31932,N_29843,N_29062);
or U31933 (N_31933,N_29230,N_28443);
and U31934 (N_31934,N_28304,N_28949);
or U31935 (N_31935,N_28573,N_29391);
or U31936 (N_31936,N_28312,N_29611);
and U31937 (N_31937,N_28154,N_29423);
nand U31938 (N_31938,N_29866,N_28513);
or U31939 (N_31939,N_28920,N_29407);
xnor U31940 (N_31940,N_28904,N_28321);
xor U31941 (N_31941,N_29227,N_29429);
xor U31942 (N_31942,N_29025,N_28934);
and U31943 (N_31943,N_29470,N_28054);
xnor U31944 (N_31944,N_29030,N_29370);
or U31945 (N_31945,N_28957,N_28657);
or U31946 (N_31946,N_29118,N_28427);
or U31947 (N_31947,N_29266,N_29209);
or U31948 (N_31948,N_28610,N_29903);
xor U31949 (N_31949,N_29389,N_29524);
and U31950 (N_31950,N_29815,N_28161);
or U31951 (N_31951,N_29678,N_29282);
nor U31952 (N_31952,N_29232,N_28502);
nand U31953 (N_31953,N_28016,N_29834);
nor U31954 (N_31954,N_28315,N_29545);
nor U31955 (N_31955,N_28943,N_29784);
nor U31956 (N_31956,N_28745,N_29131);
nor U31957 (N_31957,N_29587,N_28232);
and U31958 (N_31958,N_29098,N_29514);
and U31959 (N_31959,N_29131,N_29204);
nor U31960 (N_31960,N_28747,N_29229);
nor U31961 (N_31961,N_28374,N_28264);
nor U31962 (N_31962,N_28382,N_28888);
nand U31963 (N_31963,N_29353,N_28836);
xnor U31964 (N_31964,N_28982,N_29236);
nor U31965 (N_31965,N_28780,N_29379);
nor U31966 (N_31966,N_28704,N_29914);
nor U31967 (N_31967,N_29738,N_28085);
and U31968 (N_31968,N_28960,N_29864);
nand U31969 (N_31969,N_29158,N_29465);
nor U31970 (N_31970,N_29805,N_29840);
nand U31971 (N_31971,N_29948,N_29199);
and U31972 (N_31972,N_28293,N_28356);
or U31973 (N_31973,N_28852,N_28025);
nand U31974 (N_31974,N_28689,N_28136);
nor U31975 (N_31975,N_28828,N_28822);
nand U31976 (N_31976,N_28206,N_29117);
nor U31977 (N_31977,N_28525,N_29841);
xnor U31978 (N_31978,N_29829,N_29388);
and U31979 (N_31979,N_29711,N_28509);
or U31980 (N_31980,N_28449,N_29599);
nor U31981 (N_31981,N_28479,N_29368);
or U31982 (N_31982,N_28356,N_29222);
or U31983 (N_31983,N_29206,N_28580);
or U31984 (N_31984,N_28781,N_29700);
nor U31985 (N_31985,N_29015,N_29424);
and U31986 (N_31986,N_28176,N_29441);
xor U31987 (N_31987,N_29923,N_29347);
nor U31988 (N_31988,N_29556,N_28204);
nand U31989 (N_31989,N_29966,N_29571);
xnor U31990 (N_31990,N_28297,N_29510);
nor U31991 (N_31991,N_28539,N_28073);
nor U31992 (N_31992,N_28681,N_29982);
xor U31993 (N_31993,N_29740,N_28531);
or U31994 (N_31994,N_29304,N_28437);
xnor U31995 (N_31995,N_29386,N_28267);
nor U31996 (N_31996,N_28289,N_29096);
or U31997 (N_31997,N_29559,N_28373);
xnor U31998 (N_31998,N_28719,N_28644);
nor U31999 (N_31999,N_29193,N_28265);
and U32000 (N_32000,N_30133,N_30485);
nand U32001 (N_32001,N_31886,N_30413);
nand U32002 (N_32002,N_30150,N_31063);
xnor U32003 (N_32003,N_31420,N_31568);
and U32004 (N_32004,N_30429,N_30299);
nand U32005 (N_32005,N_30911,N_31548);
nand U32006 (N_32006,N_30492,N_30015);
or U32007 (N_32007,N_31761,N_30262);
xnor U32008 (N_32008,N_31232,N_30422);
nand U32009 (N_32009,N_31369,N_30744);
or U32010 (N_32010,N_30444,N_31482);
nand U32011 (N_32011,N_30479,N_30063);
and U32012 (N_32012,N_30844,N_31009);
and U32013 (N_32013,N_30249,N_30938);
nand U32014 (N_32014,N_31173,N_30678);
xor U32015 (N_32015,N_31674,N_30031);
nor U32016 (N_32016,N_30724,N_30100);
xnor U32017 (N_32017,N_30443,N_31607);
nand U32018 (N_32018,N_31104,N_31090);
and U32019 (N_32019,N_31382,N_30017);
xor U32020 (N_32020,N_31948,N_30821);
nand U32021 (N_32021,N_31850,N_30189);
xnor U32022 (N_32022,N_31581,N_30318);
nor U32023 (N_32023,N_30402,N_31410);
and U32024 (N_32024,N_31363,N_31663);
and U32025 (N_32025,N_30784,N_30863);
xor U32026 (N_32026,N_31446,N_31352);
and U32027 (N_32027,N_31221,N_30054);
nand U32028 (N_32028,N_30576,N_31056);
nand U32029 (N_32029,N_30788,N_31348);
and U32030 (N_32030,N_31434,N_30549);
nor U32031 (N_32031,N_30436,N_31456);
and U32032 (N_32032,N_30459,N_30157);
and U32033 (N_32033,N_31919,N_30737);
xor U32034 (N_32034,N_31849,N_31015);
or U32035 (N_32035,N_30500,N_31159);
nand U32036 (N_32036,N_31126,N_30426);
nor U32037 (N_32037,N_31193,N_30556);
or U32038 (N_32038,N_31552,N_30193);
xor U32039 (N_32039,N_31899,N_31487);
or U32040 (N_32040,N_31987,N_31218);
and U32041 (N_32041,N_31284,N_31416);
or U32042 (N_32042,N_30277,N_31544);
nor U32043 (N_32043,N_30652,N_30503);
xnor U32044 (N_32044,N_30759,N_31388);
nor U32045 (N_32045,N_31190,N_30288);
nor U32046 (N_32046,N_30547,N_30304);
or U32047 (N_32047,N_30506,N_31319);
and U32048 (N_32048,N_30071,N_30296);
and U32049 (N_32049,N_30445,N_30581);
and U32050 (N_32050,N_31982,N_30011);
xor U32051 (N_32051,N_30648,N_30292);
xor U32052 (N_32052,N_31039,N_30397);
nor U32053 (N_32053,N_31633,N_31342);
nand U32054 (N_32054,N_31955,N_30168);
xor U32055 (N_32055,N_31317,N_30316);
xnor U32056 (N_32056,N_30416,N_31315);
and U32057 (N_32057,N_31597,N_30423);
and U32058 (N_32058,N_31207,N_31616);
xnor U32059 (N_32059,N_31244,N_31165);
nor U32060 (N_32060,N_30812,N_30018);
nor U32061 (N_32061,N_31569,N_31959);
nor U32062 (N_32062,N_30142,N_30461);
nand U32063 (N_32063,N_31102,N_30165);
nor U32064 (N_32064,N_31867,N_30213);
nor U32065 (N_32065,N_31464,N_31330);
nor U32066 (N_32066,N_30679,N_30907);
nand U32067 (N_32067,N_30879,N_31110);
or U32068 (N_32068,N_31485,N_30786);
xnor U32069 (N_32069,N_31515,N_30921);
xnor U32070 (N_32070,N_31121,N_30908);
and U32071 (N_32071,N_30517,N_31715);
nor U32072 (N_32072,N_31040,N_30792);
and U32073 (N_32073,N_31662,N_30343);
or U32074 (N_32074,N_31103,N_31801);
nor U32075 (N_32075,N_31058,N_31275);
xor U32076 (N_32076,N_31430,N_31671);
and U32077 (N_32077,N_31037,N_30686);
or U32078 (N_32078,N_30721,N_31424);
nor U32079 (N_32079,N_30362,N_31454);
or U32080 (N_32080,N_30866,N_30120);
nor U32081 (N_32081,N_31957,N_30748);
nand U32082 (N_32082,N_31089,N_30406);
nor U32083 (N_32083,N_30487,N_31326);
xor U32084 (N_32084,N_30955,N_31890);
and U32085 (N_32085,N_30962,N_30009);
xor U32086 (N_32086,N_31545,N_30127);
and U32087 (N_32087,N_31051,N_31985);
and U32088 (N_32088,N_31308,N_30123);
nor U32089 (N_32089,N_30861,N_30654);
nor U32090 (N_32090,N_31947,N_31885);
nand U32091 (N_32091,N_31175,N_31695);
and U32092 (N_32092,N_31415,N_30375);
nand U32093 (N_32093,N_31983,N_31403);
or U32094 (N_32094,N_30476,N_31478);
and U32095 (N_32095,N_31672,N_30202);
and U32096 (N_32096,N_31707,N_31293);
nand U32097 (N_32097,N_30871,N_31306);
or U32098 (N_32098,N_31543,N_31178);
and U32099 (N_32099,N_31566,N_31921);
or U32100 (N_32100,N_30135,N_30597);
and U32101 (N_32101,N_31156,N_30872);
and U32102 (N_32102,N_30950,N_30694);
nor U32103 (N_32103,N_30338,N_30876);
or U32104 (N_32104,N_30096,N_30473);
nand U32105 (N_32105,N_31018,N_30300);
xor U32106 (N_32106,N_30973,N_30892);
nor U32107 (N_32107,N_30242,N_31168);
and U32108 (N_32108,N_30245,N_31627);
and U32109 (N_32109,N_30885,N_31032);
nand U32110 (N_32110,N_31967,N_31419);
nor U32111 (N_32111,N_31523,N_31585);
xor U32112 (N_32112,N_30056,N_31473);
or U32113 (N_32113,N_31975,N_30527);
xor U32114 (N_32114,N_30488,N_30232);
or U32115 (N_32115,N_31825,N_31973);
nand U32116 (N_32116,N_30466,N_30188);
nor U32117 (N_32117,N_30779,N_30330);
or U32118 (N_32118,N_30948,N_31535);
xnor U32119 (N_32119,N_31278,N_30331);
and U32120 (N_32120,N_31337,N_31064);
nand U32121 (N_32121,N_31976,N_30642);
xor U32122 (N_32122,N_30790,N_30320);
and U32123 (N_32123,N_31316,N_30105);
nor U32124 (N_32124,N_31309,N_30037);
and U32125 (N_32125,N_31873,N_30915);
and U32126 (N_32126,N_30563,N_31996);
and U32127 (N_32127,N_30231,N_30393);
nand U32128 (N_32128,N_30477,N_30773);
or U32129 (N_32129,N_30038,N_31225);
xor U32130 (N_32130,N_30069,N_31934);
or U32131 (N_32131,N_30215,N_30968);
xor U32132 (N_32132,N_31611,N_30541);
and U32133 (N_32133,N_30042,N_30484);
nand U32134 (N_32134,N_30728,N_31276);
and U32135 (N_32135,N_31676,N_30019);
or U32136 (N_32136,N_31010,N_30496);
nand U32137 (N_32137,N_30602,N_30187);
or U32138 (N_32138,N_31577,N_31184);
nor U32139 (N_32139,N_31829,N_31839);
or U32140 (N_32140,N_30624,N_31900);
xor U32141 (N_32141,N_30794,N_31742);
nor U32142 (N_32142,N_31704,N_31786);
nand U32143 (N_32143,N_30403,N_31239);
or U32144 (N_32144,N_31368,N_31830);
and U32145 (N_32145,N_31183,N_31150);
nand U32146 (N_32146,N_30611,N_31792);
nor U32147 (N_32147,N_31272,N_31459);
and U32148 (N_32148,N_30628,N_31385);
nand U32149 (N_32149,N_30052,N_30282);
nor U32150 (N_32150,N_31865,N_30200);
nor U32151 (N_32151,N_30785,N_31914);
or U32152 (N_32152,N_31120,N_31054);
xnor U32153 (N_32153,N_30588,N_31167);
xnor U32154 (N_32154,N_30247,N_31893);
xor U32155 (N_32155,N_31367,N_30841);
or U32156 (N_32156,N_31853,N_31231);
nand U32157 (N_32157,N_31828,N_31229);
or U32158 (N_32158,N_31654,N_31359);
and U32159 (N_32159,N_30226,N_30369);
nand U32160 (N_32160,N_30224,N_31012);
or U32161 (N_32161,N_31764,N_30637);
xor U32162 (N_32162,N_30949,N_31790);
xnor U32163 (N_32163,N_31449,N_31999);
and U32164 (N_32164,N_31574,N_31860);
and U32165 (N_32165,N_31087,N_30060);
nor U32166 (N_32166,N_31818,N_31946);
nand U32167 (N_32167,N_31870,N_30162);
and U32168 (N_32168,N_31497,N_31637);
xnor U32169 (N_32169,N_30182,N_30713);
xor U32170 (N_32170,N_31595,N_30023);
nand U32171 (N_32171,N_31274,N_30591);
xnor U32172 (N_32172,N_31956,N_31992);
or U32173 (N_32173,N_31644,N_31047);
or U32174 (N_32174,N_31282,N_30222);
nand U32175 (N_32175,N_30417,N_30310);
xnor U32176 (N_32176,N_30551,N_31913);
and U32177 (N_32177,N_30380,N_30816);
nand U32178 (N_32178,N_31458,N_30904);
nor U32179 (N_32179,N_31406,N_31556);
nand U32180 (N_32180,N_31245,N_31536);
xor U32181 (N_32181,N_31608,N_30902);
nand U32182 (N_32182,N_31003,N_30837);
nor U32183 (N_32183,N_30431,N_30720);
nor U32184 (N_32184,N_31048,N_31248);
xnor U32185 (N_32185,N_30378,N_31554);
and U32186 (N_32186,N_31095,N_31409);
xnor U32187 (N_32187,N_30618,N_30146);
and U32188 (N_32188,N_30129,N_31290);
and U32189 (N_32189,N_30787,N_30176);
nor U32190 (N_32190,N_31777,N_30554);
nand U32191 (N_32191,N_31273,N_30317);
nor U32192 (N_32192,N_30057,N_31177);
xnor U32193 (N_32193,N_30817,N_30035);
or U32194 (N_32194,N_31143,N_30192);
nor U32195 (N_32195,N_30987,N_31065);
or U32196 (N_32196,N_31374,N_31270);
xnor U32197 (N_32197,N_31749,N_30522);
or U32198 (N_32198,N_31861,N_31741);
and U32199 (N_32199,N_31365,N_31318);
xnor U32200 (N_32200,N_31622,N_30099);
or U32201 (N_32201,N_30631,N_31334);
and U32202 (N_32202,N_31341,N_30004);
xnor U32203 (N_32203,N_30223,N_31132);
nand U32204 (N_32204,N_31538,N_30308);
nor U32205 (N_32205,N_30098,N_30131);
nor U32206 (N_32206,N_30287,N_30481);
nor U32207 (N_32207,N_30217,N_30428);
and U32208 (N_32208,N_31646,N_30460);
or U32209 (N_32209,N_30906,N_31289);
xor U32210 (N_32210,N_31049,N_31862);
nand U32211 (N_32211,N_30778,N_30661);
nand U32212 (N_32212,N_30960,N_31563);
nand U32213 (N_32213,N_30511,N_30513);
nand U32214 (N_32214,N_31411,N_31732);
xor U32215 (N_32215,N_30234,N_31407);
xor U32216 (N_32216,N_30977,N_31736);
and U32217 (N_32217,N_30411,N_30983);
and U32218 (N_32218,N_30881,N_31267);
or U32219 (N_32219,N_30078,N_30838);
nor U32220 (N_32220,N_30167,N_30809);
nand U32221 (N_32221,N_31857,N_31602);
nand U32222 (N_32222,N_30205,N_30064);
nor U32223 (N_32223,N_30208,N_31511);
nand U32224 (N_32224,N_30993,N_30085);
and U32225 (N_32225,N_31846,N_30598);
and U32226 (N_32226,N_30629,N_31299);
or U32227 (N_32227,N_30689,N_31811);
xnor U32228 (N_32228,N_30373,N_31522);
and U32229 (N_32229,N_31440,N_31755);
or U32230 (N_32230,N_31147,N_30260);
xnor U32231 (N_32231,N_31423,N_31029);
and U32232 (N_32232,N_31257,N_30356);
nor U32233 (N_32233,N_30890,N_30325);
xnor U32234 (N_32234,N_30566,N_30228);
nor U32235 (N_32235,N_31703,N_31149);
nor U32236 (N_32236,N_30236,N_30827);
or U32237 (N_32237,N_30824,N_31979);
xor U32238 (N_32238,N_30680,N_31370);
or U32239 (N_32239,N_31729,N_31349);
nand U32240 (N_32240,N_30329,N_31692);
nor U32241 (N_32241,N_31144,N_30593);
or U32242 (N_32242,N_30497,N_30770);
and U32243 (N_32243,N_30989,N_30735);
nand U32244 (N_32244,N_31591,N_31036);
nand U32245 (N_32245,N_30240,N_30610);
nor U32246 (N_32246,N_30692,N_31752);
xor U32247 (N_32247,N_30332,N_31224);
and U32248 (N_32248,N_31307,N_30749);
and U32249 (N_32249,N_31963,N_31437);
nor U32250 (N_32250,N_30263,N_30802);
xor U32251 (N_32251,N_31471,N_31016);
nand U32252 (N_32252,N_31803,N_30440);
and U32253 (N_32253,N_31356,N_31025);
and U32254 (N_32254,N_31137,N_31105);
xnor U32255 (N_32255,N_30280,N_31882);
and U32256 (N_32256,N_30732,N_30596);
xnor U32257 (N_32257,N_31355,N_31281);
nand U32258 (N_32258,N_30579,N_31793);
nor U32259 (N_32259,N_30276,N_30498);
and U32260 (N_32260,N_30048,N_31321);
nor U32261 (N_32261,N_30923,N_31205);
xor U32262 (N_32262,N_30243,N_30571);
nand U32263 (N_32263,N_31404,N_31966);
and U32264 (N_32264,N_30640,N_30399);
xnor U32265 (N_32265,N_30095,N_30136);
or U32266 (N_32266,N_31390,N_31808);
nand U32267 (N_32267,N_31286,N_31305);
nand U32268 (N_32268,N_31195,N_30543);
or U32269 (N_32269,N_31945,N_30857);
nor U32270 (N_32270,N_30121,N_30229);
nand U32271 (N_32271,N_31160,N_31255);
or U32272 (N_32272,N_31131,N_30183);
nor U32273 (N_32273,N_30434,N_31557);
nor U32274 (N_32274,N_30400,N_31433);
and U32275 (N_32275,N_30516,N_30185);
or U32276 (N_32276,N_30319,N_31495);
xor U32277 (N_32277,N_31773,N_30860);
nor U32278 (N_32278,N_31513,N_30722);
or U32279 (N_32279,N_30996,N_31053);
or U32280 (N_32280,N_30734,N_31797);
and U32281 (N_32281,N_30164,N_31202);
xor U32282 (N_32282,N_30177,N_31720);
or U32283 (N_32283,N_31970,N_31172);
and U32284 (N_32284,N_30261,N_30803);
or U32285 (N_32285,N_31188,N_30390);
or U32286 (N_32286,N_30580,N_31498);
and U32287 (N_32287,N_30895,N_30920);
or U32288 (N_32288,N_31520,N_30442);
nand U32289 (N_32289,N_30725,N_31649);
xnor U32290 (N_32290,N_31603,N_30561);
and U32291 (N_32291,N_30825,N_30886);
xnor U32292 (N_32292,N_30265,N_31344);
nor U32293 (N_32293,N_31869,N_30483);
or U32294 (N_32294,N_31387,N_31292);
or U32295 (N_32295,N_31550,N_30769);
xnor U32296 (N_32296,N_31558,N_30945);
nand U32297 (N_32297,N_31978,N_31117);
nor U32298 (N_32298,N_31559,N_31336);
or U32299 (N_32299,N_31429,N_30981);
xor U32300 (N_32300,N_30854,N_30791);
nand U32301 (N_32301,N_30357,N_31041);
xor U32302 (N_32302,N_31942,N_30355);
nand U32303 (N_32303,N_30621,N_30501);
or U32304 (N_32304,N_30218,N_31450);
or U32305 (N_32305,N_30917,N_31938);
or U32306 (N_32306,N_31484,N_31022);
and U32307 (N_32307,N_31954,N_30934);
xor U32308 (N_32308,N_30995,N_31743);
and U32309 (N_32309,N_30649,N_30365);
and U32310 (N_32310,N_31555,N_30457);
nand U32311 (N_32311,N_30814,N_30793);
and U32312 (N_32312,N_30194,N_31303);
xnor U32313 (N_32313,N_30106,N_31169);
or U32314 (N_32314,N_30999,N_30819);
xor U32315 (N_32315,N_30462,N_30718);
nor U32316 (N_32316,N_30062,N_30627);
or U32317 (N_32317,N_31294,N_30326);
and U32318 (N_32318,N_31926,N_30107);
xnor U32319 (N_32319,N_30586,N_31858);
or U32320 (N_32320,N_30974,N_31897);
and U32321 (N_32321,N_31066,N_31017);
nand U32322 (N_32322,N_31699,N_31468);
or U32323 (N_32323,N_30410,N_30548);
or U32324 (N_32324,N_31804,N_30540);
xor U32325 (N_32325,N_30074,N_30931);
xor U32326 (N_32326,N_30028,N_31665);
nand U32327 (N_32327,N_30697,N_31241);
xor U32328 (N_32328,N_30238,N_31546);
or U32329 (N_32329,N_30097,N_30198);
xnor U32330 (N_32330,N_30845,N_30211);
nand U32331 (N_32331,N_30274,N_31587);
and U32332 (N_32332,N_30704,N_30518);
or U32333 (N_32333,N_31194,N_31227);
and U32334 (N_32334,N_31613,N_30616);
nor U32335 (N_32335,N_31004,N_31412);
and U32336 (N_32336,N_30763,N_31991);
nand U32337 (N_32337,N_30859,N_31347);
nor U32338 (N_32338,N_30701,N_31852);
nor U32339 (N_32339,N_30926,N_31974);
xnor U32340 (N_32340,N_30374,N_30528);
xnor U32341 (N_32341,N_31961,N_30046);
nand U32342 (N_32342,N_31529,N_31211);
nor U32343 (N_32343,N_31042,N_31679);
or U32344 (N_32344,N_31969,N_31322);
nand U32345 (N_32345,N_31258,N_31619);
or U32346 (N_32346,N_31297,N_31474);
or U32347 (N_32347,N_31133,N_31837);
and U32348 (N_32348,N_31716,N_31146);
xnor U32349 (N_32349,N_31312,N_30266);
nand U32350 (N_32350,N_31684,N_30524);
and U32351 (N_32351,N_31431,N_30835);
nand U32352 (N_32352,N_30268,N_30345);
and U32353 (N_32353,N_30030,N_31686);
xor U32354 (N_32354,N_31106,N_31170);
nor U32355 (N_32355,N_31204,N_31681);
nand U32356 (N_32356,N_30252,N_31448);
nand U32357 (N_32357,N_31084,N_30740);
nand U32358 (N_32358,N_31807,N_31075);
xnor U32359 (N_32359,N_31219,N_30230);
xor U32360 (N_32360,N_31215,N_30843);
and U32361 (N_32361,N_30818,N_31453);
or U32362 (N_32362,N_31057,N_30585);
nand U32363 (N_32363,N_31779,N_31189);
xor U32364 (N_32364,N_31836,N_30149);
nor U32365 (N_32365,N_31091,N_30657);
and U32366 (N_32366,N_30978,N_30315);
nand U32367 (N_32367,N_31909,N_31614);
nor U32368 (N_32368,N_30924,N_30206);
xnor U32369 (N_32369,N_31094,N_31851);
nand U32370 (N_32370,N_30191,N_30026);
and U32371 (N_32371,N_31078,N_30255);
nand U32372 (N_32372,N_30065,N_31986);
and U32373 (N_32373,N_30010,N_30708);
xor U32374 (N_32374,N_30956,N_31514);
nand U32375 (N_32375,N_31206,N_30448);
nand U32376 (N_32376,N_31656,N_31551);
xnor U32377 (N_32377,N_31508,N_30041);
xor U32378 (N_32378,N_30337,N_30039);
nand U32379 (N_32379,N_31583,N_31894);
xnor U32380 (N_32380,N_30578,N_30542);
nor U32381 (N_32381,N_30970,N_31605);
or U32382 (N_32382,N_31020,N_31014);
nand U32383 (N_32383,N_31217,N_31351);
or U32384 (N_32384,N_31621,N_30607);
xor U32385 (N_32385,N_30612,N_31046);
nor U32386 (N_32386,N_31623,N_30303);
nor U32387 (N_32387,N_30178,N_30469);
xor U32388 (N_32388,N_30088,N_30246);
xnor U32389 (N_32389,N_31157,N_31664);
and U32390 (N_32390,N_31575,N_30148);
nand U32391 (N_32391,N_30927,N_31499);
nand U32392 (N_32392,N_31216,N_31380);
and U32393 (N_32393,N_31826,N_31254);
nor U32394 (N_32394,N_31402,N_30884);
or U32395 (N_32395,N_30644,N_30850);
nor U32396 (N_32396,N_30573,N_31725);
nand U32397 (N_32397,N_30003,N_30197);
or U32398 (N_32398,N_31570,N_30617);
nand U32399 (N_32399,N_31625,N_31972);
and U32400 (N_32400,N_30975,N_30592);
nor U32401 (N_32401,N_31197,N_30147);
and U32402 (N_32402,N_31128,N_30221);
xnor U32403 (N_32403,N_30568,N_31405);
xor U32404 (N_32404,N_31086,N_31384);
and U32405 (N_32405,N_30623,N_31162);
xnor U32406 (N_32406,N_30570,N_30874);
nand U32407 (N_32407,N_30179,N_30289);
nand U32408 (N_32408,N_30295,N_31151);
or U32409 (N_32409,N_30050,N_31845);
or U32410 (N_32410,N_31391,N_30024);
nor U32411 (N_32411,N_30614,N_30499);
nand U32412 (N_32412,N_30111,N_31951);
or U32413 (N_32413,N_31234,N_31472);
xnor U32414 (N_32414,N_30830,N_31228);
and U32415 (N_32415,N_30195,N_31669);
xor U32416 (N_32416,N_30384,N_30673);
nand U32417 (N_32417,N_30807,N_30405);
xor U32418 (N_32418,N_31636,N_30755);
and U32419 (N_32419,N_30766,N_31067);
or U32420 (N_32420,N_31791,N_31396);
and U32421 (N_32421,N_30868,N_30493);
xnor U32422 (N_32422,N_31418,N_31531);
and U32423 (N_32423,N_30630,N_30550);
or U32424 (N_32424,N_31620,N_31280);
or U32425 (N_32425,N_30601,N_30333);
or U32426 (N_32426,N_31901,N_30777);
nor U32427 (N_32427,N_31787,N_31580);
and U32428 (N_32428,N_31031,N_31876);
nor U32429 (N_32429,N_30953,N_30181);
nand U32430 (N_32430,N_31696,N_30104);
xor U32431 (N_32431,N_31589,N_31888);
nor U32432 (N_32432,N_30698,N_30716);
nor U32433 (N_32433,N_30092,N_31518);
and U32434 (N_32434,N_31953,N_31855);
xnor U32435 (N_32435,N_30335,N_31125);
and U32436 (N_32436,N_31249,N_31719);
or U32437 (N_32437,N_31806,N_30875);
nand U32438 (N_32438,N_31737,N_30723);
xnor U32439 (N_32439,N_30959,N_31230);
nand U32440 (N_32440,N_30446,N_31462);
nor U32441 (N_32441,N_31479,N_30220);
nor U32442 (N_32442,N_30767,N_30599);
nand U32443 (N_32443,N_30729,N_31813);
nor U32444 (N_32444,N_31504,N_30703);
nor U32445 (N_32445,N_31313,N_31503);
nand U32446 (N_32446,N_31944,N_31237);
and U32447 (N_32447,N_31698,N_31332);
xnor U32448 (N_32448,N_30529,N_31019);
and U32449 (N_32449,N_31422,N_30258);
nor U32450 (N_32450,N_31346,N_31373);
nor U32451 (N_32451,N_31489,N_31085);
nor U32452 (N_32452,N_31701,N_31044);
nor U32453 (N_32453,N_30301,N_30354);
nand U32454 (N_32454,N_30108,N_30151);
nand U32455 (N_32455,N_30899,N_30828);
nand U32456 (N_32456,N_30352,N_31182);
or U32457 (N_32457,N_31301,N_31599);
and U32458 (N_32458,N_30858,N_31002);
nor U32459 (N_32459,N_31812,N_30988);
nor U32460 (N_32460,N_31835,N_30622);
nor U32461 (N_32461,N_31809,N_30765);
xor U32462 (N_32462,N_31486,N_30776);
and U32463 (N_32463,N_30005,N_31768);
nand U32464 (N_32464,N_31748,N_30311);
nor U32465 (N_32465,N_30257,N_31109);
nor U32466 (N_32466,N_30203,N_30419);
or U32467 (N_32467,N_31261,N_30782);
and U32468 (N_32468,N_30947,N_31304);
and U32469 (N_32469,N_31076,N_31733);
or U32470 (N_32470,N_30801,N_30693);
nand U32471 (N_32471,N_31738,N_30437);
nand U32472 (N_32472,N_30856,N_30984);
or U32473 (N_32473,N_30075,N_30103);
or U32474 (N_32474,N_30233,N_31553);
nor U32475 (N_32475,N_31222,N_31670);
and U32476 (N_32476,N_31265,N_30327);
and U32477 (N_32477,N_31774,N_31493);
nor U32478 (N_32478,N_30738,N_30937);
nor U32479 (N_32479,N_31466,N_31148);
nor U32480 (N_32480,N_30609,N_31394);
nor U32481 (N_32481,N_30762,N_30909);
nand U32482 (N_32482,N_30992,N_30883);
nor U32483 (N_32483,N_31724,N_30253);
and U32484 (N_32484,N_31708,N_30896);
nor U32485 (N_32485,N_31868,N_30997);
nor U32486 (N_32486,N_31354,N_30334);
or U32487 (N_32487,N_31993,N_30567);
nor U32488 (N_32488,N_31874,N_31930);
and U32489 (N_32489,N_30882,N_30020);
nor U32490 (N_32490,N_30432,N_30658);
xnor U32491 (N_32491,N_30388,N_30372);
nor U32492 (N_32492,N_31176,N_30864);
and U32493 (N_32493,N_30404,N_31444);
nand U32494 (N_32494,N_30214,N_31795);
or U32495 (N_32495,N_31571,N_31122);
xnor U32496 (N_32496,N_30491,N_30368);
or U32497 (N_32497,N_30143,N_30170);
nor U32498 (N_32498,N_30867,N_30302);
nor U32499 (N_32499,N_31123,N_30196);
nand U32500 (N_32500,N_31643,N_31842);
or U32501 (N_32501,N_31141,N_30800);
nand U32502 (N_32502,N_31107,N_31628);
xnor U32503 (N_32503,N_30662,N_30672);
and U32504 (N_32504,N_30764,N_30797);
xnor U32505 (N_32505,N_30674,N_31824);
xor U32506 (N_32506,N_31537,N_31586);
xnor U32507 (N_32507,N_30025,N_30877);
nand U32508 (N_32508,N_31335,N_30395);
and U32509 (N_32509,N_31264,N_31451);
xnor U32510 (N_32510,N_30066,N_31902);
nand U32511 (N_32511,N_31939,N_30594);
nand U32512 (N_32512,N_31481,N_31099);
and U32513 (N_32513,N_31895,N_31421);
xor U32514 (N_32514,N_30606,N_30958);
and U32515 (N_32515,N_30717,N_30815);
nor U32516 (N_32516,N_31629,N_31443);
nand U32517 (N_32517,N_31590,N_31467);
and U32518 (N_32518,N_30781,N_30468);
and U32519 (N_32519,N_31924,N_30972);
nand U32520 (N_32520,N_31908,N_30954);
xor U32521 (N_32521,N_30427,N_30898);
and U32522 (N_32522,N_30430,N_30053);
nor U32523 (N_32523,N_30851,N_30952);
and U32524 (N_32524,N_30158,N_31880);
nor U32525 (N_32525,N_30472,N_30161);
or U32526 (N_32526,N_31268,N_30936);
xor U32527 (N_32527,N_30638,N_31035);
xnor U32528 (N_32528,N_30283,N_31632);
and U32529 (N_32529,N_30119,N_30577);
or U32530 (N_32530,N_31638,N_31140);
and U32531 (N_32531,N_30746,N_31889);
xor U32532 (N_32532,N_30101,N_30152);
or U32533 (N_32533,N_30639,N_30305);
or U32534 (N_32534,N_31389,N_30665);
xor U32535 (N_32535,N_30383,N_31805);
nor U32536 (N_32536,N_30387,N_31769);
xnor U32537 (N_32537,N_30747,N_30651);
or U32538 (N_32538,N_31528,N_31832);
xnor U32539 (N_32539,N_31158,N_30507);
or U32540 (N_32540,N_30965,N_31631);
nor U32541 (N_32541,N_31233,N_31989);
or U32542 (N_32542,N_30141,N_31576);
nor U32543 (N_32543,N_30306,N_31130);
nor U32544 (N_32544,N_31062,N_31612);
nand U32545 (N_32545,N_30055,N_31740);
nor U32546 (N_32546,N_30361,N_31984);
nand U32547 (N_32547,N_31350,N_30798);
nor U32548 (N_32548,N_31547,N_30163);
or U32549 (N_32549,N_31929,N_31134);
or U32550 (N_32550,N_30905,N_31030);
xor U32551 (N_32551,N_30112,N_31112);
nor U32552 (N_32552,N_30967,N_31758);
xor U32553 (N_32553,N_31936,N_31477);
xnor U32554 (N_32554,N_30710,N_31688);
or U32555 (N_32555,N_30027,N_30036);
nand U32556 (N_32556,N_30412,N_31155);
nor U32557 (N_32557,N_30682,N_30439);
nand U32558 (N_32558,N_31174,N_31376);
or U32559 (N_32559,N_31937,N_31626);
and U32560 (N_32560,N_30346,N_31775);
and U32561 (N_32561,N_31778,N_31817);
or U32562 (N_32562,N_30398,N_31541);
and U32563 (N_32563,N_30626,N_31726);
nor U32564 (N_32564,N_30942,N_31731);
xor U32565 (N_32565,N_30081,N_30450);
and U32566 (N_32566,N_31116,N_31208);
nand U32567 (N_32567,N_30001,N_31950);
nor U32568 (N_32568,N_30424,N_31310);
or U32569 (N_32569,N_31693,N_31843);
xor U32570 (N_32570,N_31788,N_31940);
or U32571 (N_32571,N_30451,N_30455);
nor U32572 (N_32572,N_31038,N_30155);
or U32573 (N_32573,N_30789,N_30901);
and U32574 (N_32574,N_30389,N_31124);
nor U32575 (N_32575,N_30966,N_30675);
nor U32576 (N_32576,N_30897,N_31080);
and U32577 (N_32577,N_31653,N_30328);
nor U32578 (N_32578,N_31023,N_30013);
nand U32579 (N_32579,N_31799,N_30562);
xnor U32580 (N_32580,N_30538,N_30731);
and U32581 (N_32581,N_30754,N_31645);
nor U32582 (N_32582,N_31300,N_31683);
or U32583 (N_32583,N_31345,N_30715);
xnor U32584 (N_32584,N_30341,N_31810);
and U32585 (N_32585,N_30826,N_31253);
or U32586 (N_32586,N_31578,N_30925);
and U32587 (N_32587,N_30862,N_30144);
xor U32588 (N_32588,N_30980,N_31366);
and U32589 (N_32589,N_31180,N_31007);
or U32590 (N_32590,N_31210,N_30553);
xor U32591 (N_32591,N_30241,N_31081);
or U32592 (N_32592,N_31651,N_31000);
nand U32593 (N_32593,N_31794,N_31838);
xnor U32594 (N_32594,N_30394,N_31465);
xor U32595 (N_32595,N_31658,N_30963);
nor U32596 (N_32596,N_31320,N_30269);
nor U32597 (N_32597,N_31127,N_31892);
xnor U32598 (N_32598,N_31166,N_31776);
nand U32599 (N_32599,N_31834,N_30209);
nand U32600 (N_32600,N_31425,N_31859);
nor U32601 (N_32601,N_30653,N_30175);
and U32602 (N_32602,N_31329,N_31302);
nor U32603 (N_32603,N_30248,N_30204);
nor U32604 (N_32604,N_31362,N_31841);
nor U32605 (N_32605,N_31516,N_31689);
xor U32606 (N_32606,N_31727,N_31910);
xor U32607 (N_32607,N_31565,N_30526);
xnor U32608 (N_32608,N_30016,N_31185);
nand U32609 (N_32609,N_30523,N_31325);
or U32610 (N_32610,N_30912,N_30558);
and U32611 (N_32611,N_30891,N_31816);
nor U32612 (N_32612,N_30285,N_31240);
nand U32613 (N_32613,N_31680,N_30741);
xor U32614 (N_32614,N_30225,N_30447);
xnor U32615 (N_32615,N_30683,N_30137);
and U32616 (N_32616,N_30464,N_30537);
or U32617 (N_32617,N_31034,N_30254);
nand U32618 (N_32618,N_30441,N_31988);
nand U32619 (N_32619,N_30180,N_30122);
nor U32620 (N_32620,N_30575,N_31718);
nor U32621 (N_32621,N_30351,N_31781);
or U32622 (N_32622,N_30349,N_31766);
xnor U32623 (N_32623,N_30264,N_31920);
or U32624 (N_32624,N_31256,N_30935);
and U32625 (N_32625,N_31428,N_31360);
nand U32626 (N_32626,N_31906,N_31070);
or U32627 (N_32627,N_30505,N_30076);
xnor U32628 (N_32628,N_30745,N_30853);
nor U32629 (N_32629,N_30298,N_31136);
xor U32630 (N_32630,N_30557,N_31161);
nor U32631 (N_32631,N_30865,N_30870);
xor U32632 (N_32632,N_30667,N_31624);
and U32633 (N_32633,N_31750,N_30083);
nand U32634 (N_32634,N_31510,N_31324);
or U32635 (N_32635,N_31502,N_30216);
nand U32636 (N_32636,N_30878,N_30750);
xor U32637 (N_32637,N_30831,N_30687);
nor U32638 (N_32638,N_30173,N_30508);
xnor U32639 (N_32639,N_31584,N_30115);
nor U32640 (N_32640,N_31734,N_30456);
or U32641 (N_32641,N_30685,N_31711);
xor U32642 (N_32642,N_30235,N_31610);
nand U32643 (N_32643,N_30820,N_30940);
or U32644 (N_32644,N_30212,N_30619);
nor U32645 (N_32645,N_31678,N_31875);
nor U32646 (N_32646,N_31925,N_30894);
or U32647 (N_32647,N_30546,N_30093);
nor U32648 (N_32648,N_30124,N_31964);
and U32649 (N_32649,N_31011,N_30363);
or U32650 (N_32650,N_30323,N_30620);
nor U32651 (N_32651,N_30145,N_30615);
nand U32652 (N_32652,N_31521,N_30842);
nand U32653 (N_32653,N_30139,N_30033);
or U32654 (N_32654,N_31746,N_30275);
and U32655 (N_32655,N_31463,N_30059);
and U32656 (N_32656,N_30590,N_31907);
and U32657 (N_32657,N_31856,N_30887);
and U32658 (N_32658,N_30153,N_31596);
nor U32659 (N_32659,N_30705,N_31960);
xor U32660 (N_32660,N_30184,N_31005);
and U32661 (N_32661,N_31118,N_31735);
xor U32662 (N_32662,N_31687,N_30916);
xor U32663 (N_32663,N_30418,N_31840);
and U32664 (N_32664,N_30067,N_30272);
xnor U32665 (N_32665,N_30166,N_30421);
and U32666 (N_32666,N_31138,N_30201);
and U32667 (N_32667,N_30660,N_31753);
or U32668 (N_32668,N_31198,N_30084);
xnor U32669 (N_32669,N_30669,N_30806);
xor U32670 (N_32670,N_30979,N_31700);
xnor U32671 (N_32671,N_30034,N_31439);
nand U32672 (N_32672,N_30077,N_30382);
or U32673 (N_32673,N_30465,N_30531);
nand U32674 (N_32674,N_31630,N_31728);
or U32675 (N_32675,N_31379,N_30359);
and U32676 (N_32676,N_30094,N_30251);
and U32677 (N_32677,N_30991,N_30544);
nand U32678 (N_32678,N_30900,N_31615);
xnor U32679 (N_32679,N_31800,N_31745);
or U32680 (N_32680,N_31582,N_31661);
nand U32681 (N_32681,N_31196,N_31968);
xnor U32682 (N_32682,N_31780,N_30140);
xor U32683 (N_32683,N_30504,N_30774);
or U32684 (N_32684,N_31785,N_30452);
and U32685 (N_32685,N_30922,N_31277);
nor U32686 (N_32686,N_30943,N_31427);
or U32687 (N_32687,N_30297,N_30379);
or U32688 (N_32688,N_31327,N_31863);
nand U32689 (N_32689,N_31668,N_30290);
xor U32690 (N_32690,N_30932,N_31714);
nor U32691 (N_32691,N_31475,N_31283);
or U32692 (N_32692,N_30756,N_30480);
nor U32693 (N_32693,N_30271,N_30348);
nor U32694 (N_32694,N_30110,N_31747);
nor U32695 (N_32695,N_31877,N_31952);
nand U32696 (N_32696,N_31026,N_30478);
nand U32697 (N_32697,N_30312,N_31098);
nand U32698 (N_32698,N_30757,N_30535);
nor U32699 (N_32699,N_30396,N_31706);
nor U32700 (N_32700,N_31483,N_31441);
nor U32701 (N_32701,N_31647,N_30939);
xnor U32702 (N_32702,N_31214,N_30314);
and U32703 (N_32703,N_31001,N_31904);
and U32704 (N_32704,N_30086,N_31833);
or U32705 (N_32705,N_30433,N_31311);
xor U32706 (N_32706,N_30367,N_30364);
or U32707 (N_32707,N_30360,N_31266);
nand U32708 (N_32708,N_31935,N_30664);
xnor U32709 (N_32709,N_31295,N_30555);
nand U32710 (N_32710,N_30587,N_30712);
and U32711 (N_32711,N_30855,N_30969);
xor U32712 (N_32712,N_30486,N_30670);
nor U32713 (N_32713,N_30377,N_31911);
nor U32714 (N_32714,N_31171,N_30267);
nor U32715 (N_32715,N_30810,N_31682);
and U32716 (N_32716,N_31922,N_31524);
or U32717 (N_32717,N_31220,N_30000);
and U32718 (N_32718,N_31872,N_31854);
and U32719 (N_32719,N_30951,N_30521);
nor U32720 (N_32720,N_31561,N_31971);
and U32721 (N_32721,N_31263,N_30643);
and U32722 (N_32722,N_31259,N_30210);
and U32723 (N_32723,N_30227,N_31532);
nand U32724 (N_32724,N_30848,N_31097);
or U32725 (N_32725,N_30339,N_31135);
or U32726 (N_32726,N_30138,N_30589);
nor U32727 (N_32727,N_31898,N_31417);
xor U32728 (N_32728,N_31639,N_30976);
xor U32729 (N_32729,N_30913,N_30040);
xor U32730 (N_32730,N_30852,N_31500);
nand U32731 (N_32731,N_31525,N_31667);
nand U32732 (N_32732,N_31476,N_30840);
nand U32733 (N_32733,N_30370,N_31338);
xnor U32734 (N_32734,N_31958,N_30391);
xor U32735 (N_32735,N_31413,N_31650);
and U32736 (N_32736,N_30780,N_30080);
and U32737 (N_32737,N_30957,N_30032);
or U32738 (N_32738,N_30449,N_31685);
or U32739 (N_32739,N_31271,N_31592);
or U32740 (N_32740,N_31756,N_30321);
and U32741 (N_32741,N_31072,N_30006);
nor U32742 (N_32742,N_31512,N_31977);
nor U32743 (N_32743,N_30510,N_31092);
xor U32744 (N_32744,N_30944,N_31896);
xor U32745 (N_32745,N_31246,N_31328);
xor U32746 (N_32746,N_31722,N_31710);
nor U32747 (N_32747,N_30650,N_31519);
nor U32748 (N_32748,N_30941,N_30495);
xnor U32749 (N_32749,N_31549,N_30742);
nand U32750 (N_32750,N_31045,N_31236);
xor U32751 (N_32751,N_31399,N_30933);
xnor U32752 (N_32752,N_31252,N_30199);
nand U32753 (N_32753,N_31386,N_30519);
and U32754 (N_32754,N_30730,N_31377);
and U32755 (N_32755,N_31050,N_31093);
or U32756 (N_32756,N_30758,N_30125);
nand U32757 (N_32757,N_31279,N_31702);
nand U32758 (N_32758,N_31343,N_31933);
or U32759 (N_32759,N_31887,N_31579);
or U32760 (N_32760,N_30259,N_31881);
or U32761 (N_32761,N_31353,N_31494);
and U32762 (N_32762,N_31760,N_30494);
nand U32763 (N_32763,N_30671,N_30930);
nand U32764 (N_32764,N_31997,N_31690);
nor U32765 (N_32765,N_30534,N_30113);
or U32766 (N_32766,N_30250,N_30336);
and U32767 (N_32767,N_31916,N_30772);
and U32768 (N_32768,N_30116,N_30425);
or U32769 (N_32769,N_31077,N_31223);
or U32770 (N_32770,N_31393,N_30279);
nand U32771 (N_32771,N_31697,N_30663);
or U32772 (N_32772,N_31187,N_30929);
nand U32773 (N_32773,N_30134,N_31823);
or U32774 (N_32774,N_31709,N_31705);
and U32775 (N_32775,N_31340,N_31226);
or U32776 (N_32776,N_30058,N_31096);
or U32777 (N_32777,N_30743,N_31530);
and U32778 (N_32778,N_31375,N_30281);
nand U32779 (N_32779,N_31212,N_31142);
or U32780 (N_32780,N_30392,N_31847);
or U32781 (N_32781,N_31397,N_30313);
and U32782 (N_32782,N_31298,N_30474);
nor U32783 (N_32783,N_30632,N_31071);
xnor U32784 (N_32784,N_30714,N_31878);
nor U32785 (N_32785,N_31657,N_30696);
or U32786 (N_32786,N_31028,N_30676);
nand U32787 (N_32787,N_30366,N_31517);
nand U32788 (N_32788,N_31339,N_30903);
and U32789 (N_32789,N_30582,N_30795);
and U32790 (N_32790,N_31073,N_31154);
nor U32791 (N_32791,N_30768,N_30572);
nand U32792 (N_32792,N_30702,N_30771);
and U32793 (N_32793,N_30174,N_30114);
xnor U32794 (N_32794,N_31822,N_30839);
nand U32795 (N_32795,N_30552,N_31981);
or U32796 (N_32796,N_31452,N_30985);
nand U32797 (N_32797,N_30045,N_30273);
and U32798 (N_32798,N_30047,N_31618);
nand U32799 (N_32799,N_31864,N_31827);
or U32800 (N_32800,N_31153,N_31436);
nand U32801 (N_32801,N_31819,N_30467);
or U32802 (N_32802,N_30634,N_31820);
and U32803 (N_32803,N_31903,N_31199);
xor U32804 (N_32804,N_30386,N_31560);
nor U32805 (N_32805,N_31371,N_31357);
nand U32806 (N_32806,N_31260,N_30172);
xor U32807 (N_32807,N_30029,N_31163);
and U32808 (N_32808,N_31712,N_31635);
or U32809 (N_32809,N_30002,N_30760);
nand U32810 (N_32810,N_31201,N_31783);
nand U32811 (N_32811,N_31013,N_30775);
and U32812 (N_32812,N_30470,N_31540);
and U32813 (N_32813,N_30799,N_30849);
and U32814 (N_32814,N_31721,N_31600);
or U32815 (N_32815,N_31186,N_30736);
xnor U32816 (N_32816,N_30869,N_30964);
and U32817 (N_32817,N_30512,N_30823);
xor U32818 (N_32818,N_30873,N_30044);
nand U32819 (N_32819,N_30415,N_30834);
nor U32820 (N_32820,N_31980,N_31079);
and U32821 (N_32821,N_31021,N_31364);
and U32822 (N_32822,N_31460,N_30482);
nor U32823 (N_32823,N_31962,N_31995);
xnor U32824 (N_32824,N_31480,N_30376);
xnor U32825 (N_32825,N_30733,N_31027);
and U32826 (N_32826,N_30914,N_31905);
or U32827 (N_32827,N_31455,N_31990);
and U32828 (N_32828,N_31496,N_30813);
or U32829 (N_32829,N_31145,N_30605);
nor U32830 (N_32830,N_31640,N_30880);
or U32831 (N_32831,N_30961,N_31111);
nor U32832 (N_32832,N_31848,N_30463);
nand U32833 (N_32833,N_31378,N_30239);
nor U32834 (N_32834,N_31572,N_31432);
xor U32835 (N_32835,N_31762,N_30128);
or U32836 (N_32836,N_30489,N_30502);
nand U32837 (N_32837,N_30109,N_30691);
nor U32838 (N_32838,N_31691,N_31043);
nor U32839 (N_32839,N_30539,N_31821);
nor U32840 (N_32840,N_31641,N_31250);
or U32841 (N_32841,N_31262,N_31100);
and U32842 (N_32842,N_31251,N_31291);
and U32843 (N_32843,N_30695,N_31943);
nand U32844 (N_32844,N_30409,N_31438);
nor U32845 (N_32845,N_30471,N_30990);
nand U32846 (N_32846,N_31372,N_31247);
or U32847 (N_32847,N_30117,N_31617);
xor U32848 (N_32848,N_31006,N_31470);
nor U32849 (N_32849,N_30986,N_30244);
nor U32850 (N_32850,N_31642,N_31789);
nand U32851 (N_32851,N_31634,N_30677);
xnor U32852 (N_32852,N_31815,N_31181);
and U32853 (N_32853,N_31772,N_30126);
and U32854 (N_32854,N_31601,N_30569);
or U32855 (N_32855,N_31717,N_30946);
xnor U32856 (N_32856,N_31108,N_31490);
and U32857 (N_32857,N_31694,N_31744);
nor U32858 (N_32858,N_31457,N_30846);
nand U32859 (N_32859,N_31119,N_30515);
nor U32860 (N_32860,N_31771,N_30829);
nand U32861 (N_32861,N_30583,N_31469);
and U32862 (N_32862,N_31358,N_30822);
nor U32863 (N_32863,N_30889,N_31593);
nor U32864 (N_32864,N_31677,N_30690);
and U32865 (N_32865,N_31088,N_31883);
nand U32866 (N_32866,N_30635,N_30256);
xnor U32867 (N_32867,N_31400,N_31492);
and U32868 (N_32868,N_30284,N_30414);
nor U32869 (N_32869,N_30603,N_31114);
nand U32870 (N_32870,N_30739,N_30560);
xnor U32871 (N_32871,N_30090,N_30207);
nand U32872 (N_32872,N_30408,N_30998);
or U32873 (N_32873,N_31203,N_30808);
and U32874 (N_32874,N_31765,N_31287);
xor U32875 (N_32875,N_31713,N_30407);
and U32876 (N_32876,N_31296,N_31866);
nand U32877 (N_32877,N_31507,N_30600);
xnor U32878 (N_32878,N_30982,N_30796);
nand U32879 (N_32879,N_30727,N_31723);
xnor U32880 (N_32880,N_31269,N_30753);
nand U32881 (N_32881,N_30190,N_30186);
nand U32882 (N_32882,N_30811,N_31501);
or U32883 (N_32883,N_30270,N_30532);
or U32884 (N_32884,N_31798,N_30309);
nand U32885 (N_32885,N_30559,N_31052);
xor U32886 (N_32886,N_31113,N_30171);
nand U32887 (N_32887,N_31831,N_30711);
nor U32888 (N_32888,N_31666,N_31802);
nand U32889 (N_32889,N_30564,N_31917);
or U32890 (N_32890,N_30699,N_31844);
or U32891 (N_32891,N_31998,N_31879);
or U32892 (N_32892,N_30910,N_30751);
nor U32893 (N_32893,N_30350,N_31243);
and U32894 (N_32894,N_31314,N_31395);
or U32895 (N_32895,N_31488,N_31200);
xor U32896 (N_32896,N_30595,N_31213);
and U32897 (N_32897,N_31759,N_31567);
and U32898 (N_32898,N_30645,N_31192);
nand U32899 (N_32899,N_30833,N_30219);
nor U32900 (N_32900,N_31573,N_30371);
or U32901 (N_32901,N_30525,N_31383);
or U32902 (N_32902,N_31152,N_30681);
xnor U32903 (N_32903,N_30918,N_31083);
nor U32904 (N_32904,N_31652,N_31739);
nand U32905 (N_32905,N_31068,N_31361);
nor U32906 (N_32906,N_30068,N_30707);
xnor U32907 (N_32907,N_30520,N_31949);
nor U32908 (N_32908,N_31101,N_30070);
xnor U32909 (N_32909,N_30545,N_31069);
xor U32910 (N_32910,N_31594,N_30533);
nor U32911 (N_32911,N_31381,N_31164);
nand U32912 (N_32912,N_30061,N_30613);
and U32913 (N_32913,N_31871,N_30647);
nor U32914 (N_32914,N_30051,N_31442);
nand U32915 (N_32915,N_31891,N_30709);
and U32916 (N_32916,N_30118,N_30286);
nor U32917 (N_32917,N_30089,N_31526);
and U32918 (N_32918,N_31927,N_31115);
nor U32919 (N_32919,N_31562,N_31932);
nand U32920 (N_32920,N_31288,N_30454);
nor U32921 (N_32921,N_31331,N_31082);
and U32922 (N_32922,N_31609,N_31757);
nor U32923 (N_32923,N_31392,N_30132);
or U32924 (N_32924,N_30832,N_30156);
nand U32925 (N_32925,N_31179,N_31426);
and U32926 (N_32926,N_31235,N_31509);
nand U32927 (N_32927,N_31784,N_31660);
and U32928 (N_32928,N_31491,N_31445);
nor U32929 (N_32929,N_30700,N_30322);
and U32930 (N_32930,N_31059,N_31659);
nand U32931 (N_32931,N_31323,N_30237);
or U32932 (N_32932,N_30342,N_30420);
nor U32933 (N_32933,N_30604,N_30919);
and U32934 (N_32934,N_30453,N_30358);
and U32935 (N_32935,N_30994,N_31333);
or U32936 (N_32936,N_30353,N_31928);
xnor U32937 (N_32937,N_30438,N_31604);
nand U32938 (N_32938,N_31564,N_31918);
or U32939 (N_32939,N_31060,N_31751);
and U32940 (N_32940,N_30381,N_30656);
nand U32941 (N_32941,N_31923,N_30893);
nand U32942 (N_32942,N_30536,N_30490);
and U32943 (N_32943,N_31606,N_31767);
or U32944 (N_32944,N_31539,N_31770);
nand U32945 (N_32945,N_30688,N_30169);
or U32946 (N_32946,N_30706,N_31915);
or U32947 (N_32947,N_31533,N_31884);
or U32948 (N_32948,N_30021,N_31447);
nand U32949 (N_32949,N_30347,N_30278);
and U32950 (N_32950,N_31796,N_31912);
nand U32951 (N_32951,N_30082,N_30666);
nand U32952 (N_32952,N_31941,N_30668);
nand U32953 (N_32953,N_30014,N_31655);
or U32954 (N_32954,N_30458,N_30633);
or U32955 (N_32955,N_31242,N_31534);
nor U32956 (N_32956,N_31024,N_31673);
and U32957 (N_32957,N_30007,N_30836);
or U32958 (N_32958,N_30530,N_30847);
nand U32959 (N_32959,N_30022,N_31209);
and U32960 (N_32960,N_31139,N_31129);
nand U32961 (N_32961,N_30971,N_30130);
nand U32962 (N_32962,N_30475,N_31414);
nor U32963 (N_32963,N_31648,N_30805);
nand U32964 (N_32964,N_30928,N_30385);
or U32965 (N_32965,N_30636,N_31238);
and U32966 (N_32966,N_30340,N_31527);
xnor U32967 (N_32967,N_30435,N_31055);
xor U32968 (N_32968,N_31598,N_31542);
or U32969 (N_32969,N_31506,N_30761);
nor U32970 (N_32970,N_30752,N_30012);
nor U32971 (N_32971,N_30514,N_31994);
xnor U32972 (N_32972,N_30655,N_31763);
and U32973 (N_32973,N_30574,N_31730);
or U32974 (N_32974,N_31931,N_30159);
xor U32975 (N_32975,N_31191,N_31588);
nand U32976 (N_32976,N_30625,N_30043);
nor U32977 (N_32977,N_30160,N_30646);
nand U32978 (N_32978,N_31782,N_31008);
nand U32979 (N_32979,N_30888,N_30102);
nand U32980 (N_32980,N_30307,N_30073);
or U32981 (N_32981,N_30719,N_30783);
and U32982 (N_32982,N_30608,N_30072);
and U32983 (N_32983,N_31398,N_30291);
or U32984 (N_32984,N_31965,N_30324);
and U32985 (N_32985,N_31061,N_31435);
or U32986 (N_32986,N_30079,N_31033);
xnor U32987 (N_32987,N_30641,N_31675);
nand U32988 (N_32988,N_31285,N_30565);
or U32989 (N_32989,N_31814,N_30659);
nand U32990 (N_32990,N_30091,N_31401);
nor U32991 (N_32991,N_30509,N_30344);
nor U32992 (N_32992,N_30684,N_30726);
nor U32993 (N_32993,N_30401,N_30584);
nand U32994 (N_32994,N_30008,N_30294);
or U32995 (N_32995,N_30293,N_30087);
nor U32996 (N_32996,N_30154,N_31505);
and U32997 (N_32997,N_30049,N_31754);
or U32998 (N_32998,N_30804,N_31461);
nand U32999 (N_32999,N_31408,N_31074);
nor U33000 (N_33000,N_30081,N_30235);
and U33001 (N_33001,N_30762,N_31104);
and U33002 (N_33002,N_31740,N_30062);
nand U33003 (N_33003,N_30501,N_31222);
xor U33004 (N_33004,N_30102,N_30077);
or U33005 (N_33005,N_31154,N_31286);
or U33006 (N_33006,N_30422,N_31320);
nor U33007 (N_33007,N_30178,N_31660);
nand U33008 (N_33008,N_30578,N_30647);
xor U33009 (N_33009,N_30292,N_30976);
xnor U33010 (N_33010,N_31779,N_30184);
xor U33011 (N_33011,N_31807,N_30659);
or U33012 (N_33012,N_31205,N_31802);
nand U33013 (N_33013,N_31210,N_30898);
xor U33014 (N_33014,N_30557,N_30330);
xnor U33015 (N_33015,N_31622,N_31793);
nor U33016 (N_33016,N_31784,N_31997);
or U33017 (N_33017,N_31644,N_31525);
and U33018 (N_33018,N_31170,N_31611);
nor U33019 (N_33019,N_30799,N_30443);
nand U33020 (N_33020,N_30192,N_30726);
xnor U33021 (N_33021,N_31342,N_30395);
xnor U33022 (N_33022,N_30415,N_30090);
nand U33023 (N_33023,N_30439,N_30400);
and U33024 (N_33024,N_30704,N_31939);
nand U33025 (N_33025,N_31377,N_31509);
and U33026 (N_33026,N_30074,N_31628);
xor U33027 (N_33027,N_31225,N_30036);
nand U33028 (N_33028,N_30079,N_31972);
nor U33029 (N_33029,N_30933,N_31629);
nor U33030 (N_33030,N_30870,N_31641);
nor U33031 (N_33031,N_31453,N_31928);
or U33032 (N_33032,N_30978,N_30367);
nor U33033 (N_33033,N_30284,N_30840);
or U33034 (N_33034,N_31724,N_31289);
or U33035 (N_33035,N_30957,N_30730);
and U33036 (N_33036,N_30708,N_30990);
and U33037 (N_33037,N_30074,N_30659);
nor U33038 (N_33038,N_31888,N_30159);
or U33039 (N_33039,N_30526,N_30864);
nor U33040 (N_33040,N_31399,N_31868);
or U33041 (N_33041,N_31704,N_30732);
nor U33042 (N_33042,N_31171,N_31447);
nor U33043 (N_33043,N_31221,N_30244);
xnor U33044 (N_33044,N_30882,N_30894);
xnor U33045 (N_33045,N_31462,N_30853);
nand U33046 (N_33046,N_31990,N_31185);
nor U33047 (N_33047,N_30277,N_30034);
or U33048 (N_33048,N_31708,N_30889);
and U33049 (N_33049,N_31331,N_31438);
nand U33050 (N_33050,N_31165,N_31475);
or U33051 (N_33051,N_30118,N_30730);
and U33052 (N_33052,N_30103,N_31946);
xor U33053 (N_33053,N_31673,N_30224);
and U33054 (N_33054,N_31939,N_31058);
and U33055 (N_33055,N_31199,N_30932);
nor U33056 (N_33056,N_30073,N_30171);
nor U33057 (N_33057,N_30540,N_31016);
or U33058 (N_33058,N_31337,N_31465);
or U33059 (N_33059,N_31096,N_30775);
xor U33060 (N_33060,N_30031,N_31376);
xor U33061 (N_33061,N_31310,N_30973);
nor U33062 (N_33062,N_30992,N_31227);
or U33063 (N_33063,N_30409,N_31564);
or U33064 (N_33064,N_30557,N_30545);
nor U33065 (N_33065,N_30374,N_31965);
or U33066 (N_33066,N_31521,N_31448);
nor U33067 (N_33067,N_30330,N_30912);
xor U33068 (N_33068,N_31202,N_30604);
and U33069 (N_33069,N_31870,N_31493);
nand U33070 (N_33070,N_30381,N_30804);
and U33071 (N_33071,N_31389,N_31181);
xnor U33072 (N_33072,N_31190,N_31502);
or U33073 (N_33073,N_30824,N_30886);
nor U33074 (N_33074,N_30945,N_31241);
nand U33075 (N_33075,N_30322,N_31384);
nand U33076 (N_33076,N_30611,N_31262);
xnor U33077 (N_33077,N_30802,N_30884);
nand U33078 (N_33078,N_30893,N_31137);
nand U33079 (N_33079,N_31605,N_31168);
and U33080 (N_33080,N_31813,N_31566);
or U33081 (N_33081,N_30206,N_31363);
nand U33082 (N_33082,N_30025,N_30299);
xnor U33083 (N_33083,N_31865,N_30075);
and U33084 (N_33084,N_31790,N_30405);
or U33085 (N_33085,N_30805,N_30631);
xnor U33086 (N_33086,N_31170,N_31972);
and U33087 (N_33087,N_31638,N_30072);
or U33088 (N_33088,N_30008,N_31030);
or U33089 (N_33089,N_31716,N_30835);
and U33090 (N_33090,N_31357,N_31909);
nor U33091 (N_33091,N_30813,N_31019);
or U33092 (N_33092,N_31007,N_31133);
nor U33093 (N_33093,N_30764,N_31705);
xor U33094 (N_33094,N_30292,N_30987);
or U33095 (N_33095,N_30166,N_31643);
nand U33096 (N_33096,N_31580,N_30095);
xnor U33097 (N_33097,N_30124,N_30099);
xnor U33098 (N_33098,N_30723,N_30164);
nand U33099 (N_33099,N_30851,N_30883);
or U33100 (N_33100,N_30670,N_31711);
or U33101 (N_33101,N_30514,N_30426);
nor U33102 (N_33102,N_31712,N_31095);
nand U33103 (N_33103,N_31226,N_31549);
xor U33104 (N_33104,N_30091,N_30037);
or U33105 (N_33105,N_31587,N_31160);
xor U33106 (N_33106,N_31194,N_31240);
nand U33107 (N_33107,N_30174,N_31026);
nand U33108 (N_33108,N_30976,N_30822);
nand U33109 (N_33109,N_31412,N_30680);
and U33110 (N_33110,N_30571,N_31050);
nand U33111 (N_33111,N_31168,N_30444);
nor U33112 (N_33112,N_31058,N_30497);
and U33113 (N_33113,N_30524,N_30087);
nor U33114 (N_33114,N_30444,N_30166);
nor U33115 (N_33115,N_31574,N_31856);
or U33116 (N_33116,N_31327,N_30272);
nand U33117 (N_33117,N_31318,N_30592);
xor U33118 (N_33118,N_30878,N_31214);
nor U33119 (N_33119,N_30371,N_31848);
and U33120 (N_33120,N_31201,N_30355);
or U33121 (N_33121,N_30643,N_31837);
nor U33122 (N_33122,N_30252,N_30079);
xor U33123 (N_33123,N_31134,N_31175);
nor U33124 (N_33124,N_30235,N_31861);
and U33125 (N_33125,N_30817,N_30006);
nor U33126 (N_33126,N_30809,N_31261);
nor U33127 (N_33127,N_30399,N_30374);
and U33128 (N_33128,N_30689,N_30731);
xor U33129 (N_33129,N_30429,N_31129);
and U33130 (N_33130,N_30629,N_30831);
xor U33131 (N_33131,N_31346,N_31603);
nand U33132 (N_33132,N_30383,N_31000);
or U33133 (N_33133,N_31770,N_30961);
or U33134 (N_33134,N_31596,N_31665);
nor U33135 (N_33135,N_30739,N_31211);
nand U33136 (N_33136,N_30152,N_31050);
nor U33137 (N_33137,N_30960,N_31583);
or U33138 (N_33138,N_31729,N_31402);
nand U33139 (N_33139,N_30459,N_31717);
xnor U33140 (N_33140,N_31132,N_30165);
xnor U33141 (N_33141,N_30078,N_31327);
nor U33142 (N_33142,N_30133,N_31048);
nor U33143 (N_33143,N_30748,N_31531);
and U33144 (N_33144,N_31072,N_31561);
nor U33145 (N_33145,N_30324,N_30588);
and U33146 (N_33146,N_31330,N_31524);
xor U33147 (N_33147,N_30997,N_31767);
or U33148 (N_33148,N_31587,N_30115);
nand U33149 (N_33149,N_30884,N_31129);
or U33150 (N_33150,N_31498,N_31035);
and U33151 (N_33151,N_31691,N_30900);
and U33152 (N_33152,N_30946,N_31435);
nand U33153 (N_33153,N_30529,N_30285);
or U33154 (N_33154,N_31226,N_30995);
nand U33155 (N_33155,N_30116,N_31893);
nor U33156 (N_33156,N_30026,N_30982);
xor U33157 (N_33157,N_31363,N_31349);
or U33158 (N_33158,N_31489,N_31206);
xor U33159 (N_33159,N_30611,N_31530);
xnor U33160 (N_33160,N_30080,N_30667);
xnor U33161 (N_33161,N_30771,N_30914);
and U33162 (N_33162,N_31086,N_30205);
nor U33163 (N_33163,N_31438,N_31355);
nand U33164 (N_33164,N_30220,N_31973);
nand U33165 (N_33165,N_30918,N_30646);
nor U33166 (N_33166,N_31452,N_31306);
nand U33167 (N_33167,N_31399,N_31369);
and U33168 (N_33168,N_31745,N_31478);
nor U33169 (N_33169,N_30128,N_30167);
and U33170 (N_33170,N_31714,N_31925);
or U33171 (N_33171,N_30687,N_31359);
xnor U33172 (N_33172,N_31059,N_31406);
and U33173 (N_33173,N_30094,N_30273);
xnor U33174 (N_33174,N_30871,N_31889);
and U33175 (N_33175,N_30532,N_31620);
xnor U33176 (N_33176,N_30968,N_30366);
and U33177 (N_33177,N_30167,N_31767);
xnor U33178 (N_33178,N_30240,N_30629);
xor U33179 (N_33179,N_30094,N_31668);
and U33180 (N_33180,N_30940,N_31000);
or U33181 (N_33181,N_30948,N_31053);
nand U33182 (N_33182,N_30812,N_30401);
and U33183 (N_33183,N_31973,N_30300);
xor U33184 (N_33184,N_31367,N_30077);
xnor U33185 (N_33185,N_31114,N_30097);
xor U33186 (N_33186,N_30950,N_30605);
xor U33187 (N_33187,N_31832,N_30185);
nand U33188 (N_33188,N_30088,N_31981);
nor U33189 (N_33189,N_30261,N_30058);
xor U33190 (N_33190,N_31709,N_30487);
xor U33191 (N_33191,N_30861,N_30488);
and U33192 (N_33192,N_31722,N_31829);
or U33193 (N_33193,N_31032,N_30323);
or U33194 (N_33194,N_31804,N_31728);
nor U33195 (N_33195,N_31809,N_31153);
nand U33196 (N_33196,N_30697,N_31552);
and U33197 (N_33197,N_30639,N_31335);
nor U33198 (N_33198,N_31003,N_30316);
or U33199 (N_33199,N_30992,N_30609);
nor U33200 (N_33200,N_30622,N_31815);
or U33201 (N_33201,N_30789,N_30517);
nor U33202 (N_33202,N_31656,N_30197);
and U33203 (N_33203,N_30117,N_31776);
nor U33204 (N_33204,N_30999,N_30799);
and U33205 (N_33205,N_31516,N_31406);
xor U33206 (N_33206,N_31796,N_30928);
nor U33207 (N_33207,N_31188,N_30609);
nand U33208 (N_33208,N_31277,N_30418);
and U33209 (N_33209,N_31698,N_31772);
and U33210 (N_33210,N_31019,N_31762);
nor U33211 (N_33211,N_31348,N_31758);
and U33212 (N_33212,N_30706,N_30263);
xnor U33213 (N_33213,N_31389,N_31230);
or U33214 (N_33214,N_31632,N_30162);
and U33215 (N_33215,N_30867,N_30364);
or U33216 (N_33216,N_31608,N_30008);
xnor U33217 (N_33217,N_30508,N_30411);
or U33218 (N_33218,N_30719,N_30704);
nand U33219 (N_33219,N_31728,N_31300);
or U33220 (N_33220,N_30614,N_31311);
nand U33221 (N_33221,N_31960,N_31598);
xor U33222 (N_33222,N_30510,N_30544);
nor U33223 (N_33223,N_30383,N_30869);
or U33224 (N_33224,N_31171,N_31286);
xnor U33225 (N_33225,N_30841,N_31199);
and U33226 (N_33226,N_31801,N_31280);
nand U33227 (N_33227,N_30816,N_30076);
xor U33228 (N_33228,N_30484,N_30456);
and U33229 (N_33229,N_31122,N_30218);
xnor U33230 (N_33230,N_30482,N_30042);
xor U33231 (N_33231,N_30989,N_30813);
nor U33232 (N_33232,N_30515,N_30755);
and U33233 (N_33233,N_30248,N_30849);
nor U33234 (N_33234,N_31852,N_30056);
nand U33235 (N_33235,N_30358,N_31428);
nor U33236 (N_33236,N_31680,N_30814);
nor U33237 (N_33237,N_30623,N_31327);
nand U33238 (N_33238,N_31356,N_30946);
and U33239 (N_33239,N_30847,N_30495);
xnor U33240 (N_33240,N_30769,N_30443);
nor U33241 (N_33241,N_30454,N_31943);
nor U33242 (N_33242,N_30746,N_31443);
xor U33243 (N_33243,N_30201,N_31895);
xor U33244 (N_33244,N_30567,N_30108);
nor U33245 (N_33245,N_31415,N_31707);
and U33246 (N_33246,N_31744,N_30040);
or U33247 (N_33247,N_31079,N_31911);
nand U33248 (N_33248,N_30428,N_31429);
xnor U33249 (N_33249,N_31217,N_30874);
xnor U33250 (N_33250,N_31212,N_30108);
nor U33251 (N_33251,N_31171,N_30939);
or U33252 (N_33252,N_30707,N_31306);
nor U33253 (N_33253,N_31735,N_31403);
xnor U33254 (N_33254,N_31118,N_30488);
or U33255 (N_33255,N_30341,N_31407);
and U33256 (N_33256,N_30826,N_30655);
xor U33257 (N_33257,N_30156,N_31971);
or U33258 (N_33258,N_30388,N_30323);
nor U33259 (N_33259,N_31309,N_31116);
or U33260 (N_33260,N_30122,N_31410);
nor U33261 (N_33261,N_30152,N_30322);
nor U33262 (N_33262,N_31833,N_31722);
or U33263 (N_33263,N_30437,N_30240);
xnor U33264 (N_33264,N_31976,N_30233);
or U33265 (N_33265,N_31221,N_30824);
nand U33266 (N_33266,N_30729,N_31843);
nor U33267 (N_33267,N_30415,N_30439);
nor U33268 (N_33268,N_30923,N_30649);
nor U33269 (N_33269,N_31502,N_30345);
and U33270 (N_33270,N_30960,N_30907);
and U33271 (N_33271,N_31343,N_30093);
and U33272 (N_33272,N_30218,N_31350);
and U33273 (N_33273,N_30794,N_30515);
or U33274 (N_33274,N_30114,N_31995);
or U33275 (N_33275,N_30218,N_30482);
and U33276 (N_33276,N_30905,N_30014);
nand U33277 (N_33277,N_31576,N_31205);
xnor U33278 (N_33278,N_31795,N_30021);
or U33279 (N_33279,N_30306,N_31984);
nor U33280 (N_33280,N_31639,N_30962);
nand U33281 (N_33281,N_30577,N_31475);
nor U33282 (N_33282,N_30725,N_30836);
nand U33283 (N_33283,N_30086,N_31857);
and U33284 (N_33284,N_31193,N_30861);
nand U33285 (N_33285,N_31736,N_31429);
and U33286 (N_33286,N_30687,N_31813);
xor U33287 (N_33287,N_30326,N_31959);
or U33288 (N_33288,N_31339,N_31601);
nand U33289 (N_33289,N_30657,N_30759);
nand U33290 (N_33290,N_30498,N_31829);
and U33291 (N_33291,N_31633,N_31244);
and U33292 (N_33292,N_30306,N_31463);
and U33293 (N_33293,N_31055,N_30366);
nand U33294 (N_33294,N_30309,N_31366);
xor U33295 (N_33295,N_31877,N_30231);
or U33296 (N_33296,N_30509,N_31330);
and U33297 (N_33297,N_30823,N_30169);
and U33298 (N_33298,N_30437,N_31134);
or U33299 (N_33299,N_31529,N_31238);
or U33300 (N_33300,N_31569,N_30215);
or U33301 (N_33301,N_30828,N_30610);
and U33302 (N_33302,N_31126,N_31427);
and U33303 (N_33303,N_30151,N_30430);
or U33304 (N_33304,N_31008,N_30918);
and U33305 (N_33305,N_31892,N_31296);
nor U33306 (N_33306,N_31699,N_30023);
or U33307 (N_33307,N_30809,N_31558);
or U33308 (N_33308,N_30724,N_30001);
xnor U33309 (N_33309,N_31916,N_30569);
or U33310 (N_33310,N_31681,N_31139);
xor U33311 (N_33311,N_30066,N_30959);
and U33312 (N_33312,N_31881,N_30999);
xor U33313 (N_33313,N_31355,N_30159);
nor U33314 (N_33314,N_31706,N_31020);
nor U33315 (N_33315,N_31287,N_30235);
or U33316 (N_33316,N_30714,N_30177);
nand U33317 (N_33317,N_30252,N_31188);
or U33318 (N_33318,N_31584,N_30380);
nor U33319 (N_33319,N_30782,N_30619);
and U33320 (N_33320,N_31424,N_30149);
nand U33321 (N_33321,N_30588,N_31147);
nor U33322 (N_33322,N_31827,N_30263);
nor U33323 (N_33323,N_30014,N_30517);
nand U33324 (N_33324,N_30413,N_30289);
xor U33325 (N_33325,N_31762,N_31142);
nor U33326 (N_33326,N_30038,N_31223);
nand U33327 (N_33327,N_31992,N_31386);
or U33328 (N_33328,N_30480,N_31539);
or U33329 (N_33329,N_30645,N_30611);
nand U33330 (N_33330,N_30961,N_30139);
xor U33331 (N_33331,N_31587,N_31109);
or U33332 (N_33332,N_31268,N_31609);
xnor U33333 (N_33333,N_31088,N_31442);
xor U33334 (N_33334,N_30161,N_30167);
nor U33335 (N_33335,N_30636,N_30032);
and U33336 (N_33336,N_31340,N_30267);
and U33337 (N_33337,N_30935,N_30713);
nor U33338 (N_33338,N_31991,N_30037);
xor U33339 (N_33339,N_30833,N_31985);
and U33340 (N_33340,N_30725,N_30336);
nor U33341 (N_33341,N_30873,N_30751);
nor U33342 (N_33342,N_30270,N_31120);
or U33343 (N_33343,N_30226,N_30683);
nor U33344 (N_33344,N_30453,N_31411);
nor U33345 (N_33345,N_31478,N_30278);
or U33346 (N_33346,N_30544,N_30166);
nor U33347 (N_33347,N_31185,N_30136);
nor U33348 (N_33348,N_30677,N_30313);
nor U33349 (N_33349,N_31602,N_30204);
nand U33350 (N_33350,N_31124,N_31133);
or U33351 (N_33351,N_30038,N_31170);
nand U33352 (N_33352,N_30192,N_30361);
or U33353 (N_33353,N_30811,N_30108);
nand U33354 (N_33354,N_31528,N_31544);
and U33355 (N_33355,N_31862,N_31059);
nor U33356 (N_33356,N_30036,N_30668);
nand U33357 (N_33357,N_31683,N_31228);
nand U33358 (N_33358,N_31659,N_31870);
nor U33359 (N_33359,N_31446,N_31940);
or U33360 (N_33360,N_30285,N_31777);
nand U33361 (N_33361,N_30128,N_31081);
nand U33362 (N_33362,N_31910,N_31960);
and U33363 (N_33363,N_30516,N_31363);
nor U33364 (N_33364,N_30614,N_31541);
nand U33365 (N_33365,N_30234,N_30778);
or U33366 (N_33366,N_31661,N_31743);
nand U33367 (N_33367,N_30117,N_30129);
or U33368 (N_33368,N_31162,N_30976);
nand U33369 (N_33369,N_30223,N_31643);
nand U33370 (N_33370,N_31346,N_30326);
xor U33371 (N_33371,N_31159,N_31183);
and U33372 (N_33372,N_30670,N_31736);
nor U33373 (N_33373,N_30544,N_31547);
xor U33374 (N_33374,N_31049,N_31893);
nor U33375 (N_33375,N_31952,N_30408);
nor U33376 (N_33376,N_30434,N_30891);
and U33377 (N_33377,N_31540,N_30597);
nor U33378 (N_33378,N_30193,N_31630);
and U33379 (N_33379,N_31594,N_30748);
and U33380 (N_33380,N_30104,N_31125);
xor U33381 (N_33381,N_30990,N_31846);
nand U33382 (N_33382,N_31866,N_31115);
nand U33383 (N_33383,N_30649,N_30862);
xor U33384 (N_33384,N_30647,N_31601);
or U33385 (N_33385,N_31436,N_30143);
xor U33386 (N_33386,N_30743,N_31479);
or U33387 (N_33387,N_31036,N_31477);
xor U33388 (N_33388,N_30787,N_30341);
or U33389 (N_33389,N_30738,N_31311);
nor U33390 (N_33390,N_31390,N_30800);
nand U33391 (N_33391,N_31155,N_31156);
nor U33392 (N_33392,N_31234,N_30650);
and U33393 (N_33393,N_30583,N_31228);
and U33394 (N_33394,N_31779,N_30757);
nor U33395 (N_33395,N_31576,N_30879);
xor U33396 (N_33396,N_31254,N_31552);
nand U33397 (N_33397,N_30426,N_30238);
nor U33398 (N_33398,N_31466,N_31981);
xnor U33399 (N_33399,N_31973,N_31662);
and U33400 (N_33400,N_30938,N_30765);
nor U33401 (N_33401,N_30264,N_31540);
nand U33402 (N_33402,N_30599,N_30885);
nor U33403 (N_33403,N_31996,N_31616);
xnor U33404 (N_33404,N_30646,N_31544);
or U33405 (N_33405,N_31158,N_31719);
and U33406 (N_33406,N_30500,N_31089);
and U33407 (N_33407,N_31426,N_30472);
xnor U33408 (N_33408,N_30540,N_30832);
nor U33409 (N_33409,N_30891,N_30981);
nor U33410 (N_33410,N_31553,N_30807);
nor U33411 (N_33411,N_31168,N_31284);
nor U33412 (N_33412,N_31316,N_30041);
xnor U33413 (N_33413,N_30856,N_31523);
and U33414 (N_33414,N_30284,N_30956);
nor U33415 (N_33415,N_30006,N_30586);
nand U33416 (N_33416,N_30348,N_30696);
and U33417 (N_33417,N_30570,N_31220);
or U33418 (N_33418,N_30157,N_30742);
xor U33419 (N_33419,N_30944,N_30785);
and U33420 (N_33420,N_31566,N_31946);
nand U33421 (N_33421,N_30303,N_30710);
or U33422 (N_33422,N_30435,N_30510);
and U33423 (N_33423,N_31177,N_31481);
xnor U33424 (N_33424,N_30766,N_30956);
xnor U33425 (N_33425,N_31011,N_31690);
nor U33426 (N_33426,N_31153,N_31445);
and U33427 (N_33427,N_31836,N_30356);
or U33428 (N_33428,N_30181,N_31564);
nor U33429 (N_33429,N_30539,N_31280);
nand U33430 (N_33430,N_31342,N_30326);
xor U33431 (N_33431,N_31933,N_30205);
and U33432 (N_33432,N_31878,N_30320);
and U33433 (N_33433,N_30356,N_30223);
nor U33434 (N_33434,N_31859,N_31053);
nor U33435 (N_33435,N_30941,N_30038);
nand U33436 (N_33436,N_31515,N_31766);
xnor U33437 (N_33437,N_31096,N_30479);
nor U33438 (N_33438,N_30755,N_30914);
xnor U33439 (N_33439,N_31226,N_30417);
nand U33440 (N_33440,N_31602,N_30330);
xnor U33441 (N_33441,N_30612,N_30683);
or U33442 (N_33442,N_31738,N_31826);
nor U33443 (N_33443,N_30132,N_30605);
and U33444 (N_33444,N_30878,N_30115);
and U33445 (N_33445,N_30543,N_31251);
or U33446 (N_33446,N_31080,N_30546);
xor U33447 (N_33447,N_31106,N_30234);
xor U33448 (N_33448,N_31503,N_30601);
nand U33449 (N_33449,N_30150,N_30312);
xnor U33450 (N_33450,N_31840,N_30408);
nand U33451 (N_33451,N_30991,N_31452);
nand U33452 (N_33452,N_31644,N_30780);
nor U33453 (N_33453,N_31958,N_30663);
nor U33454 (N_33454,N_30883,N_30325);
nand U33455 (N_33455,N_30230,N_30712);
nand U33456 (N_33456,N_30143,N_31788);
nand U33457 (N_33457,N_30352,N_30678);
xnor U33458 (N_33458,N_30141,N_31392);
xnor U33459 (N_33459,N_31476,N_30371);
xnor U33460 (N_33460,N_31238,N_31025);
xor U33461 (N_33461,N_30632,N_30020);
or U33462 (N_33462,N_31481,N_31809);
nor U33463 (N_33463,N_30902,N_30749);
nand U33464 (N_33464,N_31734,N_31374);
nand U33465 (N_33465,N_30703,N_30259);
and U33466 (N_33466,N_30149,N_30662);
or U33467 (N_33467,N_30382,N_30963);
xnor U33468 (N_33468,N_31870,N_30377);
and U33469 (N_33469,N_31012,N_31612);
and U33470 (N_33470,N_30789,N_30877);
and U33471 (N_33471,N_30445,N_30987);
nor U33472 (N_33472,N_31136,N_31744);
or U33473 (N_33473,N_31707,N_31809);
or U33474 (N_33474,N_30402,N_31331);
xnor U33475 (N_33475,N_31072,N_31662);
xor U33476 (N_33476,N_30600,N_31336);
nor U33477 (N_33477,N_31766,N_30816);
xor U33478 (N_33478,N_31193,N_31248);
nor U33479 (N_33479,N_30706,N_31650);
nand U33480 (N_33480,N_30197,N_31530);
or U33481 (N_33481,N_30190,N_30217);
and U33482 (N_33482,N_30963,N_31328);
xnor U33483 (N_33483,N_30518,N_30804);
and U33484 (N_33484,N_31208,N_30118);
and U33485 (N_33485,N_30463,N_31339);
xnor U33486 (N_33486,N_30253,N_31119);
and U33487 (N_33487,N_31096,N_31137);
nand U33488 (N_33488,N_30450,N_30399);
nor U33489 (N_33489,N_31450,N_31550);
nand U33490 (N_33490,N_30348,N_30287);
nand U33491 (N_33491,N_31343,N_31548);
nor U33492 (N_33492,N_31963,N_30914);
xor U33493 (N_33493,N_31525,N_30592);
xor U33494 (N_33494,N_30817,N_31209);
or U33495 (N_33495,N_31760,N_31714);
nand U33496 (N_33496,N_30732,N_30918);
or U33497 (N_33497,N_30157,N_30678);
nand U33498 (N_33498,N_30963,N_31627);
nor U33499 (N_33499,N_30367,N_30101);
nand U33500 (N_33500,N_30652,N_30227);
and U33501 (N_33501,N_30696,N_31099);
and U33502 (N_33502,N_30164,N_31376);
nand U33503 (N_33503,N_31997,N_30461);
and U33504 (N_33504,N_30243,N_31201);
and U33505 (N_33505,N_31979,N_30596);
xnor U33506 (N_33506,N_31803,N_31862);
and U33507 (N_33507,N_31398,N_30874);
nor U33508 (N_33508,N_31593,N_31156);
and U33509 (N_33509,N_30465,N_31099);
nor U33510 (N_33510,N_31574,N_30740);
or U33511 (N_33511,N_30381,N_30171);
and U33512 (N_33512,N_31970,N_30362);
nor U33513 (N_33513,N_31040,N_31091);
xnor U33514 (N_33514,N_31490,N_31856);
and U33515 (N_33515,N_30407,N_30256);
nor U33516 (N_33516,N_31882,N_31533);
nand U33517 (N_33517,N_31105,N_30818);
or U33518 (N_33518,N_31734,N_31727);
xor U33519 (N_33519,N_30258,N_30767);
xor U33520 (N_33520,N_31996,N_30652);
xnor U33521 (N_33521,N_31729,N_31239);
nand U33522 (N_33522,N_30325,N_31098);
or U33523 (N_33523,N_31248,N_30199);
or U33524 (N_33524,N_30772,N_31138);
nor U33525 (N_33525,N_31051,N_31338);
nand U33526 (N_33526,N_31209,N_30413);
nor U33527 (N_33527,N_31864,N_30688);
nand U33528 (N_33528,N_30021,N_30412);
nor U33529 (N_33529,N_30463,N_31288);
xnor U33530 (N_33530,N_31980,N_31142);
nand U33531 (N_33531,N_31167,N_30486);
xor U33532 (N_33532,N_30074,N_31143);
or U33533 (N_33533,N_30047,N_30690);
and U33534 (N_33534,N_30346,N_31291);
or U33535 (N_33535,N_31596,N_30906);
and U33536 (N_33536,N_31220,N_30025);
or U33537 (N_33537,N_31647,N_31428);
and U33538 (N_33538,N_30081,N_31977);
nor U33539 (N_33539,N_31819,N_31028);
nand U33540 (N_33540,N_30308,N_30900);
or U33541 (N_33541,N_31720,N_31370);
nand U33542 (N_33542,N_30329,N_30168);
or U33543 (N_33543,N_30577,N_30819);
or U33544 (N_33544,N_31945,N_31962);
and U33545 (N_33545,N_31750,N_31742);
nand U33546 (N_33546,N_30052,N_31636);
and U33547 (N_33547,N_30759,N_31280);
or U33548 (N_33548,N_30029,N_31078);
or U33549 (N_33549,N_31850,N_30947);
nor U33550 (N_33550,N_30379,N_31036);
nor U33551 (N_33551,N_30120,N_30277);
nand U33552 (N_33552,N_31631,N_30261);
or U33553 (N_33553,N_30833,N_31423);
or U33554 (N_33554,N_31637,N_31111);
xor U33555 (N_33555,N_31143,N_30621);
xnor U33556 (N_33556,N_30653,N_31811);
xnor U33557 (N_33557,N_30059,N_30323);
nand U33558 (N_33558,N_31327,N_31582);
and U33559 (N_33559,N_31168,N_30431);
nor U33560 (N_33560,N_31273,N_30301);
or U33561 (N_33561,N_31763,N_30198);
and U33562 (N_33562,N_30314,N_30552);
nor U33563 (N_33563,N_31380,N_31960);
nand U33564 (N_33564,N_30879,N_30659);
nor U33565 (N_33565,N_30531,N_31113);
and U33566 (N_33566,N_31717,N_31313);
and U33567 (N_33567,N_30127,N_30977);
or U33568 (N_33568,N_30502,N_31928);
and U33569 (N_33569,N_31492,N_31784);
nor U33570 (N_33570,N_30884,N_31941);
nor U33571 (N_33571,N_30918,N_31757);
xnor U33572 (N_33572,N_31989,N_31198);
or U33573 (N_33573,N_30115,N_31429);
or U33574 (N_33574,N_30068,N_31305);
or U33575 (N_33575,N_30514,N_31477);
nand U33576 (N_33576,N_30811,N_31030);
nand U33577 (N_33577,N_30231,N_30892);
and U33578 (N_33578,N_30015,N_31758);
or U33579 (N_33579,N_31759,N_31432);
or U33580 (N_33580,N_30148,N_30904);
nand U33581 (N_33581,N_30279,N_31777);
nor U33582 (N_33582,N_30247,N_30109);
and U33583 (N_33583,N_30166,N_30226);
and U33584 (N_33584,N_31838,N_31412);
and U33585 (N_33585,N_31164,N_30588);
nand U33586 (N_33586,N_31956,N_31971);
nand U33587 (N_33587,N_30271,N_31392);
and U33588 (N_33588,N_31447,N_30262);
nand U33589 (N_33589,N_31811,N_31551);
xnor U33590 (N_33590,N_31390,N_31133);
xnor U33591 (N_33591,N_30014,N_31485);
and U33592 (N_33592,N_31120,N_30240);
nor U33593 (N_33593,N_30222,N_30386);
nor U33594 (N_33594,N_31433,N_31890);
and U33595 (N_33595,N_30669,N_30728);
nand U33596 (N_33596,N_31868,N_31071);
nor U33597 (N_33597,N_31703,N_31951);
and U33598 (N_33598,N_31697,N_31318);
and U33599 (N_33599,N_30822,N_31411);
or U33600 (N_33600,N_31377,N_30439);
xnor U33601 (N_33601,N_30451,N_30885);
nor U33602 (N_33602,N_31787,N_31049);
or U33603 (N_33603,N_30624,N_31719);
nor U33604 (N_33604,N_30924,N_31764);
and U33605 (N_33605,N_30838,N_31714);
nor U33606 (N_33606,N_30864,N_31287);
nor U33607 (N_33607,N_31499,N_31325);
nor U33608 (N_33608,N_31367,N_30904);
and U33609 (N_33609,N_31230,N_31608);
nand U33610 (N_33610,N_30907,N_30804);
xor U33611 (N_33611,N_30194,N_30389);
and U33612 (N_33612,N_31313,N_31954);
nand U33613 (N_33613,N_30223,N_30044);
and U33614 (N_33614,N_31950,N_31662);
and U33615 (N_33615,N_31184,N_31531);
nor U33616 (N_33616,N_31779,N_31125);
nor U33617 (N_33617,N_30818,N_30492);
and U33618 (N_33618,N_30740,N_31999);
or U33619 (N_33619,N_30192,N_30204);
or U33620 (N_33620,N_30230,N_30550);
nor U33621 (N_33621,N_30959,N_31282);
and U33622 (N_33622,N_31421,N_30315);
nor U33623 (N_33623,N_31422,N_31947);
nor U33624 (N_33624,N_31254,N_30398);
nand U33625 (N_33625,N_30402,N_30853);
and U33626 (N_33626,N_31771,N_31283);
nand U33627 (N_33627,N_31112,N_30610);
xnor U33628 (N_33628,N_31162,N_31843);
or U33629 (N_33629,N_31854,N_31930);
nor U33630 (N_33630,N_31675,N_30844);
xnor U33631 (N_33631,N_30269,N_31718);
nor U33632 (N_33632,N_30083,N_30916);
xor U33633 (N_33633,N_31399,N_30107);
and U33634 (N_33634,N_30989,N_30872);
or U33635 (N_33635,N_30742,N_31054);
and U33636 (N_33636,N_31522,N_31250);
or U33637 (N_33637,N_30434,N_30884);
or U33638 (N_33638,N_31058,N_31318);
nor U33639 (N_33639,N_31840,N_31932);
nor U33640 (N_33640,N_31692,N_30913);
and U33641 (N_33641,N_31571,N_31858);
nor U33642 (N_33642,N_31735,N_30160);
and U33643 (N_33643,N_31410,N_31088);
nand U33644 (N_33644,N_30580,N_31503);
nor U33645 (N_33645,N_31172,N_31862);
xor U33646 (N_33646,N_30384,N_30899);
nor U33647 (N_33647,N_31521,N_30451);
nand U33648 (N_33648,N_31790,N_30399);
nor U33649 (N_33649,N_30104,N_31645);
nor U33650 (N_33650,N_30068,N_30038);
xnor U33651 (N_33651,N_31663,N_31096);
xnor U33652 (N_33652,N_30478,N_30596);
and U33653 (N_33653,N_30857,N_31910);
nand U33654 (N_33654,N_31908,N_30966);
nor U33655 (N_33655,N_30579,N_31929);
nor U33656 (N_33656,N_30992,N_30874);
nand U33657 (N_33657,N_31913,N_30727);
and U33658 (N_33658,N_31404,N_31715);
or U33659 (N_33659,N_30890,N_31805);
or U33660 (N_33660,N_30827,N_31046);
and U33661 (N_33661,N_30669,N_31860);
nor U33662 (N_33662,N_30322,N_31607);
nand U33663 (N_33663,N_30766,N_31110);
or U33664 (N_33664,N_31614,N_31971);
xnor U33665 (N_33665,N_30824,N_30795);
and U33666 (N_33666,N_31198,N_30423);
nor U33667 (N_33667,N_31458,N_30019);
or U33668 (N_33668,N_31397,N_30553);
nor U33669 (N_33669,N_30127,N_30173);
xnor U33670 (N_33670,N_30820,N_30826);
and U33671 (N_33671,N_30766,N_31083);
nand U33672 (N_33672,N_31193,N_31319);
nand U33673 (N_33673,N_30909,N_30123);
or U33674 (N_33674,N_30212,N_31782);
or U33675 (N_33675,N_31143,N_31312);
nor U33676 (N_33676,N_30878,N_30069);
and U33677 (N_33677,N_31200,N_31941);
and U33678 (N_33678,N_31155,N_30139);
or U33679 (N_33679,N_31113,N_30992);
xor U33680 (N_33680,N_30539,N_31438);
or U33681 (N_33681,N_30734,N_30865);
nand U33682 (N_33682,N_30339,N_30236);
nor U33683 (N_33683,N_31955,N_30061);
and U33684 (N_33684,N_30427,N_31150);
nor U33685 (N_33685,N_31579,N_31843);
and U33686 (N_33686,N_31247,N_30331);
nor U33687 (N_33687,N_30218,N_30644);
xor U33688 (N_33688,N_31934,N_31101);
or U33689 (N_33689,N_30863,N_31662);
nor U33690 (N_33690,N_31877,N_30593);
nand U33691 (N_33691,N_30886,N_31908);
nor U33692 (N_33692,N_30958,N_30413);
nor U33693 (N_33693,N_31576,N_31453);
nand U33694 (N_33694,N_30240,N_30779);
or U33695 (N_33695,N_31920,N_30001);
and U33696 (N_33696,N_30785,N_31758);
nand U33697 (N_33697,N_31395,N_31545);
and U33698 (N_33698,N_30710,N_30831);
xnor U33699 (N_33699,N_30663,N_30197);
xnor U33700 (N_33700,N_30193,N_31527);
and U33701 (N_33701,N_30923,N_30014);
and U33702 (N_33702,N_30333,N_30966);
nor U33703 (N_33703,N_30233,N_31183);
or U33704 (N_33704,N_30444,N_31724);
or U33705 (N_33705,N_30385,N_30740);
nand U33706 (N_33706,N_30224,N_31786);
or U33707 (N_33707,N_31654,N_30707);
nand U33708 (N_33708,N_30148,N_30334);
nand U33709 (N_33709,N_31646,N_30884);
xor U33710 (N_33710,N_30833,N_30602);
and U33711 (N_33711,N_30997,N_31882);
xnor U33712 (N_33712,N_30324,N_30420);
nand U33713 (N_33713,N_31516,N_31648);
and U33714 (N_33714,N_30312,N_31662);
nand U33715 (N_33715,N_30087,N_30464);
xnor U33716 (N_33716,N_30491,N_31470);
or U33717 (N_33717,N_31135,N_30266);
or U33718 (N_33718,N_31559,N_31873);
or U33719 (N_33719,N_31041,N_31052);
nor U33720 (N_33720,N_30564,N_30448);
and U33721 (N_33721,N_31946,N_30388);
or U33722 (N_33722,N_30467,N_31732);
and U33723 (N_33723,N_30812,N_30599);
xor U33724 (N_33724,N_30245,N_31776);
or U33725 (N_33725,N_30231,N_31718);
nand U33726 (N_33726,N_30788,N_31659);
and U33727 (N_33727,N_31942,N_30561);
nand U33728 (N_33728,N_30633,N_30267);
xnor U33729 (N_33729,N_31307,N_30368);
and U33730 (N_33730,N_30101,N_31593);
or U33731 (N_33731,N_31358,N_30265);
and U33732 (N_33732,N_30653,N_31932);
nor U33733 (N_33733,N_31491,N_31166);
nand U33734 (N_33734,N_30641,N_31853);
xnor U33735 (N_33735,N_30024,N_30730);
and U33736 (N_33736,N_31635,N_30194);
and U33737 (N_33737,N_31264,N_30156);
or U33738 (N_33738,N_31923,N_31117);
or U33739 (N_33739,N_31178,N_31370);
nand U33740 (N_33740,N_31429,N_31144);
xnor U33741 (N_33741,N_31616,N_30244);
nor U33742 (N_33742,N_31392,N_31535);
xor U33743 (N_33743,N_30423,N_30548);
nor U33744 (N_33744,N_30094,N_31004);
xor U33745 (N_33745,N_30923,N_30189);
nor U33746 (N_33746,N_30759,N_31141);
nor U33747 (N_33747,N_30011,N_30827);
xor U33748 (N_33748,N_31340,N_30586);
xor U33749 (N_33749,N_30832,N_31859);
nand U33750 (N_33750,N_30409,N_31685);
xnor U33751 (N_33751,N_30521,N_30060);
nor U33752 (N_33752,N_30584,N_31276);
nor U33753 (N_33753,N_31075,N_30616);
and U33754 (N_33754,N_31322,N_31798);
and U33755 (N_33755,N_30048,N_30655);
or U33756 (N_33756,N_30147,N_30077);
and U33757 (N_33757,N_31472,N_30970);
nor U33758 (N_33758,N_31318,N_30694);
nor U33759 (N_33759,N_31308,N_30255);
and U33760 (N_33760,N_31338,N_31143);
nor U33761 (N_33761,N_31936,N_30776);
nand U33762 (N_33762,N_31749,N_30165);
xnor U33763 (N_33763,N_31986,N_31791);
nor U33764 (N_33764,N_30692,N_30153);
and U33765 (N_33765,N_30166,N_30000);
xor U33766 (N_33766,N_30054,N_31044);
or U33767 (N_33767,N_30009,N_30994);
nor U33768 (N_33768,N_30079,N_30634);
nor U33769 (N_33769,N_30893,N_31207);
and U33770 (N_33770,N_30121,N_31766);
and U33771 (N_33771,N_30735,N_30149);
or U33772 (N_33772,N_30937,N_30841);
nor U33773 (N_33773,N_30777,N_30442);
xnor U33774 (N_33774,N_30025,N_31623);
and U33775 (N_33775,N_30869,N_31566);
and U33776 (N_33776,N_30066,N_31991);
nand U33777 (N_33777,N_30151,N_30854);
nand U33778 (N_33778,N_31102,N_30811);
or U33779 (N_33779,N_30148,N_31491);
nor U33780 (N_33780,N_30930,N_31016);
or U33781 (N_33781,N_30490,N_30983);
xor U33782 (N_33782,N_30596,N_31576);
or U33783 (N_33783,N_31108,N_30514);
or U33784 (N_33784,N_30010,N_31944);
and U33785 (N_33785,N_30583,N_31409);
and U33786 (N_33786,N_30181,N_30596);
xnor U33787 (N_33787,N_31917,N_31047);
or U33788 (N_33788,N_30058,N_30695);
or U33789 (N_33789,N_31739,N_31904);
nor U33790 (N_33790,N_30292,N_30270);
or U33791 (N_33791,N_31338,N_31479);
and U33792 (N_33792,N_31255,N_30647);
or U33793 (N_33793,N_31231,N_30916);
xor U33794 (N_33794,N_30686,N_30647);
xnor U33795 (N_33795,N_30884,N_31572);
and U33796 (N_33796,N_30979,N_31436);
or U33797 (N_33797,N_30792,N_30742);
and U33798 (N_33798,N_31813,N_30005);
xor U33799 (N_33799,N_30604,N_31950);
nor U33800 (N_33800,N_30389,N_30043);
and U33801 (N_33801,N_30469,N_30058);
nor U33802 (N_33802,N_31155,N_30250);
and U33803 (N_33803,N_30346,N_31116);
or U33804 (N_33804,N_31555,N_31378);
nand U33805 (N_33805,N_31997,N_31167);
and U33806 (N_33806,N_30995,N_30245);
nor U33807 (N_33807,N_30899,N_30372);
nor U33808 (N_33808,N_30721,N_31960);
xor U33809 (N_33809,N_30600,N_31234);
and U33810 (N_33810,N_30800,N_30255);
and U33811 (N_33811,N_31278,N_30045);
nand U33812 (N_33812,N_31632,N_30263);
and U33813 (N_33813,N_31719,N_30209);
or U33814 (N_33814,N_30838,N_31425);
nor U33815 (N_33815,N_31589,N_31657);
and U33816 (N_33816,N_31977,N_30827);
or U33817 (N_33817,N_31684,N_31887);
xor U33818 (N_33818,N_31367,N_31132);
nand U33819 (N_33819,N_31963,N_30824);
nand U33820 (N_33820,N_30741,N_31115);
and U33821 (N_33821,N_31582,N_31667);
nor U33822 (N_33822,N_30270,N_31480);
and U33823 (N_33823,N_30368,N_30931);
nor U33824 (N_33824,N_31505,N_30408);
or U33825 (N_33825,N_31683,N_31348);
xor U33826 (N_33826,N_31191,N_30786);
or U33827 (N_33827,N_30169,N_31250);
and U33828 (N_33828,N_31208,N_30973);
xor U33829 (N_33829,N_30280,N_30465);
or U33830 (N_33830,N_30646,N_30364);
nand U33831 (N_33831,N_30402,N_31052);
and U33832 (N_33832,N_31664,N_30478);
or U33833 (N_33833,N_30145,N_30094);
nor U33834 (N_33834,N_31720,N_31472);
and U33835 (N_33835,N_30227,N_31420);
xor U33836 (N_33836,N_30410,N_30175);
or U33837 (N_33837,N_30944,N_31410);
xor U33838 (N_33838,N_31562,N_31963);
nand U33839 (N_33839,N_31539,N_31155);
nor U33840 (N_33840,N_31491,N_30146);
nor U33841 (N_33841,N_30988,N_31730);
or U33842 (N_33842,N_31747,N_31117);
xnor U33843 (N_33843,N_31567,N_30645);
nand U33844 (N_33844,N_31012,N_30470);
and U33845 (N_33845,N_30011,N_30054);
nand U33846 (N_33846,N_31909,N_30813);
nor U33847 (N_33847,N_30532,N_30566);
xnor U33848 (N_33848,N_31620,N_31141);
and U33849 (N_33849,N_31146,N_31202);
nor U33850 (N_33850,N_31138,N_31990);
or U33851 (N_33851,N_30839,N_30692);
nand U33852 (N_33852,N_30116,N_31369);
nor U33853 (N_33853,N_30328,N_30986);
or U33854 (N_33854,N_30728,N_30107);
nand U33855 (N_33855,N_31284,N_30805);
and U33856 (N_33856,N_31582,N_30554);
xor U33857 (N_33857,N_30879,N_31261);
or U33858 (N_33858,N_31247,N_31318);
nor U33859 (N_33859,N_30523,N_31048);
nor U33860 (N_33860,N_30088,N_31643);
and U33861 (N_33861,N_31054,N_30894);
xor U33862 (N_33862,N_30328,N_31708);
nor U33863 (N_33863,N_31144,N_31375);
nand U33864 (N_33864,N_31949,N_31234);
xor U33865 (N_33865,N_30047,N_30604);
and U33866 (N_33866,N_31310,N_31715);
xnor U33867 (N_33867,N_30079,N_30467);
and U33868 (N_33868,N_31385,N_31822);
xnor U33869 (N_33869,N_31014,N_31901);
or U33870 (N_33870,N_31239,N_31201);
nor U33871 (N_33871,N_30726,N_31628);
nand U33872 (N_33872,N_30838,N_30122);
xnor U33873 (N_33873,N_30032,N_31611);
nand U33874 (N_33874,N_31985,N_30687);
nor U33875 (N_33875,N_31488,N_30221);
or U33876 (N_33876,N_30639,N_31666);
nand U33877 (N_33877,N_30606,N_30444);
and U33878 (N_33878,N_31481,N_30179);
nor U33879 (N_33879,N_31609,N_31880);
or U33880 (N_33880,N_31207,N_30131);
nand U33881 (N_33881,N_31270,N_31796);
or U33882 (N_33882,N_31080,N_30859);
nand U33883 (N_33883,N_30907,N_30179);
xor U33884 (N_33884,N_30913,N_30302);
or U33885 (N_33885,N_30178,N_30333);
or U33886 (N_33886,N_31268,N_31651);
xor U33887 (N_33887,N_30694,N_31528);
xnor U33888 (N_33888,N_31208,N_31847);
nand U33889 (N_33889,N_30528,N_30471);
and U33890 (N_33890,N_31731,N_31989);
nand U33891 (N_33891,N_30206,N_31967);
nand U33892 (N_33892,N_31782,N_31387);
and U33893 (N_33893,N_31489,N_30522);
and U33894 (N_33894,N_31687,N_31443);
nand U33895 (N_33895,N_30409,N_30545);
xor U33896 (N_33896,N_30650,N_31632);
nor U33897 (N_33897,N_30611,N_31412);
or U33898 (N_33898,N_30857,N_30885);
nor U33899 (N_33899,N_30688,N_31003);
xnor U33900 (N_33900,N_31214,N_30961);
or U33901 (N_33901,N_31272,N_31500);
nand U33902 (N_33902,N_30067,N_31518);
nand U33903 (N_33903,N_30189,N_30171);
nor U33904 (N_33904,N_30854,N_30186);
and U33905 (N_33905,N_30792,N_30994);
xor U33906 (N_33906,N_31765,N_30948);
or U33907 (N_33907,N_31122,N_31615);
nor U33908 (N_33908,N_31684,N_30446);
xnor U33909 (N_33909,N_30364,N_30918);
xnor U33910 (N_33910,N_30061,N_30980);
nor U33911 (N_33911,N_30225,N_30172);
or U33912 (N_33912,N_30816,N_30866);
nand U33913 (N_33913,N_31964,N_31083);
xor U33914 (N_33914,N_30252,N_30404);
nor U33915 (N_33915,N_31444,N_31756);
xor U33916 (N_33916,N_31519,N_30974);
nand U33917 (N_33917,N_30853,N_30073);
nand U33918 (N_33918,N_31292,N_30540);
nor U33919 (N_33919,N_31227,N_31393);
or U33920 (N_33920,N_31359,N_31274);
xnor U33921 (N_33921,N_31199,N_30634);
nand U33922 (N_33922,N_31896,N_30273);
nand U33923 (N_33923,N_31242,N_30553);
xnor U33924 (N_33924,N_31202,N_30187);
and U33925 (N_33925,N_31697,N_31321);
and U33926 (N_33926,N_31420,N_30419);
and U33927 (N_33927,N_30286,N_31983);
nand U33928 (N_33928,N_31354,N_30214);
or U33929 (N_33929,N_30535,N_31510);
or U33930 (N_33930,N_31509,N_30901);
and U33931 (N_33931,N_30273,N_30675);
nand U33932 (N_33932,N_30959,N_30679);
nor U33933 (N_33933,N_31046,N_30025);
nand U33934 (N_33934,N_31239,N_31545);
or U33935 (N_33935,N_31260,N_30022);
nor U33936 (N_33936,N_30987,N_31928);
xor U33937 (N_33937,N_31812,N_30154);
xor U33938 (N_33938,N_30019,N_30083);
xor U33939 (N_33939,N_31085,N_31656);
nor U33940 (N_33940,N_31213,N_31027);
nand U33941 (N_33941,N_30333,N_31148);
and U33942 (N_33942,N_30407,N_31202);
nor U33943 (N_33943,N_30661,N_30305);
nand U33944 (N_33944,N_30596,N_30137);
or U33945 (N_33945,N_31061,N_31026);
xnor U33946 (N_33946,N_31178,N_30749);
nand U33947 (N_33947,N_30445,N_30012);
and U33948 (N_33948,N_31525,N_30933);
xor U33949 (N_33949,N_30613,N_31691);
nand U33950 (N_33950,N_30078,N_30164);
xnor U33951 (N_33951,N_30497,N_30806);
nand U33952 (N_33952,N_30997,N_30271);
nand U33953 (N_33953,N_30912,N_31302);
or U33954 (N_33954,N_30767,N_31621);
xnor U33955 (N_33955,N_30855,N_31008);
or U33956 (N_33956,N_30730,N_31993);
nand U33957 (N_33957,N_30174,N_31262);
nand U33958 (N_33958,N_30958,N_30194);
nor U33959 (N_33959,N_31574,N_30928);
nor U33960 (N_33960,N_31749,N_30015);
and U33961 (N_33961,N_31512,N_31987);
nand U33962 (N_33962,N_30612,N_31872);
or U33963 (N_33963,N_31306,N_30064);
nor U33964 (N_33964,N_31848,N_30800);
or U33965 (N_33965,N_30107,N_30236);
and U33966 (N_33966,N_30624,N_30056);
nand U33967 (N_33967,N_30436,N_30002);
nand U33968 (N_33968,N_30734,N_30461);
nand U33969 (N_33969,N_30924,N_30122);
or U33970 (N_33970,N_30593,N_31966);
or U33971 (N_33971,N_30507,N_30781);
nor U33972 (N_33972,N_30990,N_31038);
nand U33973 (N_33973,N_31985,N_30752);
or U33974 (N_33974,N_31131,N_31032);
or U33975 (N_33975,N_30378,N_30286);
nor U33976 (N_33976,N_30290,N_31896);
nor U33977 (N_33977,N_30348,N_31641);
or U33978 (N_33978,N_31833,N_30079);
nand U33979 (N_33979,N_31267,N_31199);
or U33980 (N_33980,N_30639,N_30722);
nor U33981 (N_33981,N_30890,N_31609);
or U33982 (N_33982,N_30846,N_30443);
xnor U33983 (N_33983,N_31824,N_31762);
xnor U33984 (N_33984,N_30824,N_30117);
nor U33985 (N_33985,N_30442,N_30175);
or U33986 (N_33986,N_31798,N_31515);
and U33987 (N_33987,N_30290,N_31227);
or U33988 (N_33988,N_30276,N_31573);
nor U33989 (N_33989,N_30920,N_30725);
and U33990 (N_33990,N_30461,N_30688);
nand U33991 (N_33991,N_30799,N_31483);
xnor U33992 (N_33992,N_30470,N_31243);
xnor U33993 (N_33993,N_30809,N_31291);
xnor U33994 (N_33994,N_31182,N_30574);
and U33995 (N_33995,N_31892,N_31752);
and U33996 (N_33996,N_30860,N_31171);
or U33997 (N_33997,N_30625,N_30455);
nor U33998 (N_33998,N_31704,N_30332);
nor U33999 (N_33999,N_31423,N_30384);
nand U34000 (N_34000,N_32846,N_33068);
or U34001 (N_34001,N_32752,N_32528);
or U34002 (N_34002,N_33059,N_33661);
nor U34003 (N_34003,N_32884,N_32907);
nor U34004 (N_34004,N_32784,N_33119);
xor U34005 (N_34005,N_32627,N_33213);
or U34006 (N_34006,N_33132,N_33184);
nand U34007 (N_34007,N_33032,N_33796);
xor U34008 (N_34008,N_33070,N_33621);
xor U34009 (N_34009,N_32161,N_33260);
and U34010 (N_34010,N_33920,N_33695);
xnor U34011 (N_34011,N_33690,N_32654);
or U34012 (N_34012,N_33396,N_32670);
or U34013 (N_34013,N_32325,N_32480);
xnor U34014 (N_34014,N_32115,N_33537);
xnor U34015 (N_34015,N_33265,N_32394);
nor U34016 (N_34016,N_33423,N_32416);
nand U34017 (N_34017,N_32247,N_33089);
xnor U34018 (N_34018,N_33408,N_32045);
xor U34019 (N_34019,N_32717,N_32097);
or U34020 (N_34020,N_33222,N_33468);
nand U34021 (N_34021,N_32366,N_32707);
and U34022 (N_34022,N_33606,N_33155);
and U34023 (N_34023,N_32007,N_33307);
and U34024 (N_34024,N_32993,N_32979);
xnor U34025 (N_34025,N_32960,N_32399);
nand U34026 (N_34026,N_33977,N_33648);
nor U34027 (N_34027,N_33157,N_33512);
xnor U34028 (N_34028,N_32905,N_32684);
or U34029 (N_34029,N_33789,N_33652);
xnor U34030 (N_34030,N_33334,N_32350);
nor U34031 (N_34031,N_32167,N_33285);
and U34032 (N_34032,N_32203,N_32982);
nor U34033 (N_34033,N_33469,N_32421);
and U34034 (N_34034,N_32484,N_33017);
or U34035 (N_34035,N_33025,N_32265);
nand U34036 (N_34036,N_32499,N_33287);
xnor U34037 (N_34037,N_32780,N_33430);
or U34038 (N_34038,N_32311,N_32236);
nor U34039 (N_34039,N_33041,N_33777);
or U34040 (N_34040,N_32699,N_32648);
nand U34041 (N_34041,N_33962,N_32343);
nor U34042 (N_34042,N_33565,N_32693);
nor U34043 (N_34043,N_33060,N_33786);
nor U34044 (N_34044,N_33341,N_33769);
and U34045 (N_34045,N_32908,N_32550);
nand U34046 (N_34046,N_32296,N_33524);
nand U34047 (N_34047,N_32571,N_32331);
nor U34048 (N_34048,N_32711,N_32054);
nand U34049 (N_34049,N_33317,N_33049);
nand U34050 (N_34050,N_33475,N_33278);
or U34051 (N_34051,N_33732,N_33484);
nand U34052 (N_34052,N_32864,N_32209);
or U34053 (N_34053,N_32251,N_33206);
and U34054 (N_34054,N_33988,N_32814);
nor U34055 (N_34055,N_32577,N_32049);
nor U34056 (N_34056,N_32436,N_32113);
nand U34057 (N_34057,N_33848,N_33033);
nand U34058 (N_34058,N_32808,N_33785);
nor U34059 (N_34059,N_32603,N_32362);
xor U34060 (N_34060,N_33601,N_32047);
and U34061 (N_34061,N_33639,N_32363);
and U34062 (N_34062,N_33111,N_32815);
and U34063 (N_34063,N_33061,N_33488);
nor U34064 (N_34064,N_33584,N_33706);
and U34065 (N_34065,N_32492,N_32051);
xor U34066 (N_34066,N_32625,N_32494);
xnor U34067 (N_34067,N_33106,N_32498);
nor U34068 (N_34068,N_32156,N_33623);
and U34069 (N_34069,N_32318,N_32788);
or U34070 (N_34070,N_33841,N_32017);
xor U34071 (N_34071,N_33793,N_32244);
nor U34072 (N_34072,N_32596,N_32310);
or U34073 (N_34073,N_33139,N_33521);
xor U34074 (N_34074,N_33347,N_33442);
and U34075 (N_34075,N_33619,N_32669);
or U34076 (N_34076,N_32923,N_33831);
nand U34077 (N_34077,N_32359,N_33397);
xor U34078 (N_34078,N_32234,N_32219);
nand U34079 (N_34079,N_32730,N_32736);
xor U34080 (N_34080,N_33403,N_32664);
and U34081 (N_34081,N_33491,N_32149);
xor U34082 (N_34082,N_33216,N_32869);
nor U34083 (N_34083,N_32355,N_32823);
or U34084 (N_34084,N_32924,N_32753);
and U34085 (N_34085,N_33813,N_32691);
nor U34086 (N_34086,N_32977,N_33372);
and U34087 (N_34087,N_33338,N_32069);
xor U34088 (N_34088,N_33241,N_32061);
or U34089 (N_34089,N_32142,N_33044);
or U34090 (N_34090,N_33178,N_32866);
or U34091 (N_34091,N_32256,N_33214);
or U34092 (N_34092,N_33180,N_33507);
or U34093 (N_34093,N_32641,N_32885);
nand U34094 (N_34094,N_33913,N_33914);
xor U34095 (N_34095,N_32019,N_32677);
or U34096 (N_34096,N_32685,N_33703);
xnor U34097 (N_34097,N_33596,N_33360);
nor U34098 (N_34098,N_32062,N_32268);
or U34099 (N_34099,N_32294,N_33439);
and U34100 (N_34100,N_33083,N_32380);
xnor U34101 (N_34101,N_32606,N_33392);
and U34102 (N_34102,N_32969,N_32041);
or U34103 (N_34103,N_32879,N_32833);
nand U34104 (N_34104,N_33663,N_33683);
xnor U34105 (N_34105,N_33143,N_33603);
and U34106 (N_34106,N_32639,N_32941);
or U34107 (N_34107,N_32277,N_33928);
nor U34108 (N_34108,N_32412,N_33699);
nand U34109 (N_34109,N_33911,N_32150);
and U34110 (N_34110,N_33881,N_32280);
nor U34111 (N_34111,N_32315,N_32360);
or U34112 (N_34112,N_33868,N_33806);
and U34113 (N_34113,N_33221,N_32934);
and U34114 (N_34114,N_32887,N_33495);
or U34115 (N_34115,N_32002,N_33811);
or U34116 (N_34116,N_32594,N_32227);
nor U34117 (N_34117,N_33530,N_33934);
and U34118 (N_34118,N_33210,N_33335);
nand U34119 (N_34119,N_32369,N_32652);
or U34120 (N_34120,N_32217,N_32295);
or U34121 (N_34121,N_33199,N_33116);
nand U34122 (N_34122,N_32301,N_33664);
nand U34123 (N_34123,N_32996,N_33467);
nor U34124 (N_34124,N_32640,N_33574);
nand U34125 (N_34125,N_33926,N_33496);
and U34126 (N_34126,N_32526,N_33205);
nand U34127 (N_34127,N_32533,N_32601);
xor U34128 (N_34128,N_32012,N_33190);
or U34129 (N_34129,N_33725,N_33929);
nand U34130 (N_34130,N_32454,N_32023);
and U34131 (N_34131,N_32508,N_33906);
nand U34132 (N_34132,N_33879,N_32862);
nand U34133 (N_34133,N_33739,N_33151);
nor U34134 (N_34134,N_32581,N_32048);
or U34135 (N_34135,N_32863,N_32881);
nand U34136 (N_34136,N_33003,N_33692);
nand U34137 (N_34137,N_33932,N_32942);
nor U34138 (N_34138,N_33035,N_32290);
nand U34139 (N_34139,N_33472,N_32099);
nand U34140 (N_34140,N_33516,N_32511);
and U34141 (N_34141,N_33183,N_33972);
nand U34142 (N_34142,N_33978,N_33688);
and U34143 (N_34143,N_33961,N_33380);
xor U34144 (N_34144,N_33478,N_33994);
nor U34145 (N_34145,N_32618,N_33144);
xor U34146 (N_34146,N_32595,N_33923);
and U34147 (N_34147,N_33306,N_33544);
xor U34148 (N_34148,N_33931,N_33531);
xnor U34149 (N_34149,N_33228,N_32091);
and U34150 (N_34150,N_33646,N_33901);
and U34151 (N_34151,N_33520,N_32003);
xnor U34152 (N_34152,N_33947,N_32915);
or U34153 (N_34153,N_33254,N_32789);
and U34154 (N_34154,N_33707,N_33883);
nor U34155 (N_34155,N_32937,N_32738);
xor U34156 (N_34156,N_33607,N_32309);
or U34157 (N_34157,N_33778,N_32082);
xor U34158 (N_34158,N_32836,N_32763);
nor U34159 (N_34159,N_32672,N_33440);
or U34160 (N_34160,N_33251,N_32910);
xnor U34161 (N_34161,N_33443,N_32667);
and U34162 (N_34162,N_33450,N_32706);
nor U34163 (N_34163,N_32453,N_32218);
nand U34164 (N_34164,N_32402,N_33554);
xnor U34165 (N_34165,N_33808,N_32276);
and U34166 (N_34166,N_33721,N_33997);
nor U34167 (N_34167,N_33723,N_32258);
nor U34168 (N_34168,N_32518,N_33567);
xnor U34169 (N_34169,N_32802,N_33028);
or U34170 (N_34170,N_32133,N_33958);
nand U34171 (N_34171,N_33308,N_32348);
or U34172 (N_34172,N_32758,N_32100);
xnor U34173 (N_34173,N_33005,N_33925);
nor U34174 (N_34174,N_32678,N_33168);
nor U34175 (N_34175,N_33499,N_32774);
xnor U34176 (N_34176,N_32822,N_33342);
nor U34177 (N_34177,N_33007,N_33253);
nand U34178 (N_34178,N_32177,N_33799);
or U34179 (N_34179,N_33011,N_33055);
nand U34180 (N_34180,N_33158,N_33687);
and U34181 (N_34181,N_33289,N_32779);
xnor U34182 (N_34182,N_33724,N_32192);
nand U34183 (N_34183,N_32743,N_33800);
nor U34184 (N_34184,N_32471,N_33889);
and U34185 (N_34185,N_33192,N_33751);
and U34186 (N_34186,N_32078,N_32883);
nor U34187 (N_34187,N_33239,N_33485);
or U34188 (N_34188,N_32940,N_32810);
nand U34189 (N_34189,N_32446,N_33429);
nand U34190 (N_34190,N_32129,N_33571);
nand U34191 (N_34191,N_33627,N_33750);
xnor U34192 (N_34192,N_33252,N_32955);
xor U34193 (N_34193,N_33109,N_32169);
nor U34194 (N_34194,N_32716,N_33189);
xnor U34195 (N_34195,N_32053,N_32651);
nand U34196 (N_34196,N_33866,N_33318);
and U34197 (N_34197,N_32376,N_33402);
nand U34198 (N_34198,N_32653,N_33425);
and U34199 (N_34199,N_33676,N_33708);
xor U34200 (N_34200,N_32316,N_32722);
xor U34201 (N_34201,N_32342,N_32539);
xor U34202 (N_34202,N_33464,N_32851);
nand U34203 (N_34203,N_33263,N_33042);
or U34204 (N_34204,N_33733,N_33227);
nor U34205 (N_34205,N_33691,N_33702);
nor U34206 (N_34206,N_32103,N_32491);
xnor U34207 (N_34207,N_33212,N_32919);
or U34208 (N_34208,N_32853,N_32948);
or U34209 (N_34209,N_33629,N_32668);
xor U34210 (N_34210,N_32063,N_32897);
nor U34211 (N_34211,N_33389,N_32422);
and U34212 (N_34212,N_33066,N_32874);
and U34213 (N_34213,N_32337,N_33736);
xor U34214 (N_34214,N_32485,N_33457);
nand U34215 (N_34215,N_33744,N_32431);
nand U34216 (N_34216,N_33054,N_33470);
and U34217 (N_34217,N_33833,N_33991);
nand U34218 (N_34218,N_32336,N_33062);
xnor U34219 (N_34219,N_32478,N_32329);
xor U34220 (N_34220,N_33364,N_32189);
nor U34221 (N_34221,N_33259,N_33264);
nand U34222 (N_34222,N_32401,N_32951);
xor U34223 (N_34223,N_33427,N_33720);
nor U34224 (N_34224,N_33614,N_33453);
or U34225 (N_34225,N_33257,N_33762);
xor U34226 (N_34226,N_32524,N_33938);
nor U34227 (N_34227,N_32178,N_32661);
xnor U34228 (N_34228,N_33058,N_33486);
nand U34229 (N_34229,N_33630,N_33551);
or U34230 (N_34230,N_33505,N_33405);
xnor U34231 (N_34231,N_33741,N_32882);
nor U34232 (N_34232,N_33368,N_32503);
and U34233 (N_34233,N_32552,N_33532);
nor U34234 (N_34234,N_33581,N_33998);
or U34235 (N_34235,N_33899,N_32111);
and U34236 (N_34236,N_33477,N_33479);
nor U34237 (N_34237,N_33245,N_33247);
or U34238 (N_34238,N_33782,N_32430);
nor U34239 (N_34239,N_33127,N_33992);
or U34240 (N_34240,N_33814,N_32347);
and U34241 (N_34241,N_33550,N_32497);
nand U34242 (N_34242,N_32636,N_32395);
nor U34243 (N_34243,N_32459,N_32243);
nand U34244 (N_34244,N_33063,N_33842);
nand U34245 (N_34245,N_33710,N_33074);
nor U34246 (N_34246,N_33705,N_32614);
nand U34247 (N_34247,N_32748,N_33609);
xor U34248 (N_34248,N_33783,N_32886);
xor U34249 (N_34249,N_33594,N_32631);
nand U34250 (N_34250,N_32842,N_32573);
or U34251 (N_34251,N_32285,N_33379);
and U34252 (N_34252,N_32059,N_32899);
nor U34253 (N_34253,N_33490,N_32075);
xnor U34254 (N_34254,N_32745,N_33644);
xor U34255 (N_34255,N_33175,N_32143);
xnor U34256 (N_34256,N_32014,N_32961);
or U34257 (N_34257,N_33413,N_32119);
xnor U34258 (N_34258,N_33529,N_33193);
and U34259 (N_34259,N_33147,N_32512);
or U34260 (N_34260,N_32392,N_33501);
nand U34261 (N_34261,N_32457,N_33354);
xor U34262 (N_34262,N_33303,N_33896);
or U34263 (N_34263,N_33316,N_33164);
nor U34264 (N_34264,N_33098,N_33185);
xnor U34265 (N_34265,N_32289,N_32932);
and U34266 (N_34266,N_33828,N_33555);
nor U34267 (N_34267,N_33187,N_32997);
or U34268 (N_34268,N_33220,N_33124);
and U34269 (N_34269,N_32155,N_32957);
and U34270 (N_34270,N_32202,N_32893);
xnor U34271 (N_34271,N_32093,N_33020);
and U34272 (N_34272,N_32740,N_33492);
xnor U34273 (N_34273,N_32830,N_32544);
xor U34274 (N_34274,N_32212,N_32876);
xnor U34275 (N_34275,N_32624,N_32474);
or U34276 (N_34276,N_32643,N_33330);
xor U34277 (N_34277,N_33838,N_32770);
nor U34278 (N_34278,N_32811,N_33233);
and U34279 (N_34279,N_33951,N_33986);
xnor U34280 (N_34280,N_32757,N_33867);
xor U34281 (N_34281,N_32353,N_33023);
or U34282 (N_34282,N_32719,N_33130);
xor U34283 (N_34283,N_33355,N_32116);
and U34284 (N_34284,N_33202,N_32070);
nor U34285 (N_34285,N_32313,N_32755);
and U34286 (N_34286,N_33944,N_33314);
and U34287 (N_34287,N_32171,N_32123);
xnor U34288 (N_34288,N_33909,N_32034);
nor U34289 (N_34289,N_33846,N_33543);
nor U34290 (N_34290,N_32462,N_32279);
nor U34291 (N_34291,N_32619,N_32938);
nand U34292 (N_34292,N_32400,N_32521);
xor U34293 (N_34293,N_32267,N_33804);
nand U34294 (N_34294,N_32613,N_33323);
nand U34295 (N_34295,N_32306,N_32326);
and U34296 (N_34296,N_33506,N_33825);
or U34297 (N_34297,N_32794,N_32162);
nand U34298 (N_34298,N_32042,N_32127);
nor U34299 (N_34299,N_32859,N_32393);
xnor U34300 (N_34300,N_33784,N_33345);
nand U34301 (N_34301,N_32083,N_33340);
nor U34302 (N_34302,N_33348,N_33385);
and U34303 (N_34303,N_33517,N_32906);
or U34304 (N_34304,N_33903,N_33534);
nand U34305 (N_34305,N_33805,N_32435);
nand U34306 (N_34306,N_33001,N_32540);
nand U34307 (N_34307,N_33320,N_32819);
xor U34308 (N_34308,N_33008,N_33839);
nor U34309 (N_34309,N_32720,N_32482);
or U34310 (N_34310,N_32324,N_33471);
nor U34311 (N_34311,N_32396,N_32428);
or U34312 (N_34312,N_33311,N_33985);
nand U34313 (N_34313,N_33292,N_33709);
xnor U34314 (N_34314,N_32913,N_33526);
or U34315 (N_34315,N_33533,N_32575);
nor U34316 (N_34316,N_32662,N_32909);
and U34317 (N_34317,N_33258,N_32060);
nor U34318 (N_34318,N_32732,N_32389);
xnor U34319 (N_34319,N_33684,N_33580);
nand U34320 (N_34320,N_32989,N_32623);
or U34321 (N_34321,N_32843,N_33847);
nand U34322 (N_34322,N_32121,N_32986);
or U34323 (N_34323,N_32611,N_33309);
nand U34324 (N_34324,N_33743,N_33272);
nand U34325 (N_34325,N_33047,N_33832);
xnor U34326 (N_34326,N_32675,N_32292);
nand U34327 (N_34327,N_33641,N_32229);
nor U34328 (N_34328,N_33043,N_32010);
and U34329 (N_34329,N_32378,N_33875);
nand U34330 (N_34330,N_33394,N_33122);
xor U34331 (N_34331,N_32288,N_32172);
and U34332 (N_34332,N_32607,N_33432);
nor U34333 (N_34333,N_33820,N_33870);
and U34334 (N_34334,N_32844,N_33294);
and U34335 (N_34335,N_33624,N_32921);
and U34336 (N_34336,N_33764,N_33797);
nand U34337 (N_34337,N_33787,N_32697);
nand U34338 (N_34338,N_33416,N_32444);
nand U34339 (N_34339,N_32522,N_32184);
or U34340 (N_34340,N_32001,N_32867);
or U34341 (N_34341,N_33095,N_32074);
or U34342 (N_34342,N_33225,N_33597);
xnor U34343 (N_34343,N_32688,N_32852);
nand U34344 (N_34344,N_33036,N_33386);
nor U34345 (N_34345,N_32696,N_32663);
nor U34346 (N_34346,N_32228,N_33912);
xnor U34347 (N_34347,N_32551,N_33742);
nand U34348 (N_34348,N_32375,N_32644);
or U34349 (N_34349,N_32515,N_32320);
and U34350 (N_34350,N_33215,N_32174);
nand U34351 (N_34351,N_33395,N_33884);
xnor U34352 (N_34352,N_32242,N_33585);
and U34353 (N_34353,N_32673,N_33204);
nand U34354 (N_34354,N_32737,N_33090);
and U34355 (N_34355,N_32764,N_33288);
xor U34356 (N_34356,N_32094,N_32772);
xor U34357 (N_34357,N_32579,N_33487);
xor U34358 (N_34358,N_33296,N_33255);
or U34359 (N_34359,N_32109,N_32704);
xor U34360 (N_34360,N_33738,N_32240);
or U34361 (N_34361,N_33256,N_32441);
nor U34362 (N_34362,N_32255,N_33181);
and U34363 (N_34363,N_33924,N_32370);
or U34364 (N_34364,N_33091,N_33539);
nor U34365 (N_34365,N_32735,N_33324);
or U34366 (N_34366,N_32769,N_32469);
xnor U34367 (N_34367,N_32496,N_33758);
nand U34368 (N_34368,N_33611,N_32163);
and U34369 (N_34369,N_33541,N_33328);
nand U34370 (N_34370,N_32703,N_33411);
or U34371 (N_34371,N_32798,N_32125);
xor U34372 (N_34372,N_32175,N_32557);
nor U34373 (N_34373,N_33493,N_33933);
xnor U34374 (N_34374,N_33246,N_32504);
xor U34375 (N_34375,N_32414,N_33608);
xnor U34376 (N_34376,N_33810,N_32845);
nor U34377 (N_34377,N_33569,N_33337);
or U34378 (N_34378,N_32826,N_32965);
or U34379 (N_34379,N_32825,N_33669);
nand U34380 (N_34380,N_32341,N_32286);
xnor U34381 (N_34381,N_33547,N_33086);
nand U34382 (N_34382,N_33575,N_32009);
xnor U34383 (N_34383,N_33618,N_32762);
xor U34384 (N_34384,N_33363,N_33211);
nor U34385 (N_34385,N_32984,N_33850);
xor U34386 (N_34386,N_32413,N_32044);
nor U34387 (N_34387,N_33882,N_33999);
or U34388 (N_34388,N_32878,N_33941);
nand U34389 (N_34389,N_33862,N_33024);
nand U34390 (N_34390,N_33293,N_32966);
and U34391 (N_34391,N_33942,N_32615);
nand U34392 (N_34392,N_33350,N_32796);
xnor U34393 (N_34393,N_32807,N_32204);
nor U34394 (N_34394,N_33658,N_32210);
or U34395 (N_34395,N_32629,N_32220);
and U34396 (N_34396,N_32367,N_33231);
nand U34397 (N_34397,N_32970,N_32634);
and U34398 (N_34398,N_32781,N_33141);
and U34399 (N_34399,N_33854,N_33118);
nor U34400 (N_34400,N_32445,N_32635);
xnor U34401 (N_34401,N_33801,N_33142);
or U34402 (N_34402,N_33504,N_33818);
nand U34403 (N_34403,N_32090,N_32461);
nand U34404 (N_34404,N_32837,N_32564);
nor U34405 (N_34405,N_33374,N_32976);
or U34406 (N_34406,N_32985,N_33599);
nor U34407 (N_34407,N_33887,N_33188);
and U34408 (N_34408,N_33670,N_33349);
xor U34409 (N_34409,N_32006,N_33817);
nor U34410 (N_34410,N_33542,N_33170);
and U34411 (N_34411,N_32792,N_33081);
xor U34412 (N_34412,N_33038,N_33651);
nor U34413 (N_34413,N_32742,N_33045);
and U34414 (N_34414,N_33186,N_33895);
xnor U34415 (N_34415,N_33678,N_32777);
or U34416 (N_34416,N_32188,N_32857);
nor U34417 (N_34417,N_32364,N_33902);
xor U34418 (N_34418,N_33434,N_32804);
or U34419 (N_34419,N_32994,N_33568);
or U34420 (N_34420,N_33234,N_33726);
xnor U34421 (N_34421,N_33950,N_32397);
xnor U34422 (N_34422,N_33659,N_32532);
and U34423 (N_34423,N_33774,N_33946);
nor U34424 (N_34424,N_33084,N_33680);
and U34425 (N_34425,N_32962,N_32858);
or U34426 (N_34426,N_32566,N_33824);
nand U34427 (N_34427,N_33237,N_33390);
or U34428 (N_34428,N_33686,N_33698);
xor U34429 (N_34429,N_33050,N_32817);
xnor U34430 (N_34430,N_32795,N_32197);
or U34431 (N_34431,N_32556,N_32734);
xor U34432 (N_34432,N_32084,N_32847);
and U34433 (N_34433,N_32153,N_32968);
nand U34434 (N_34434,N_32873,N_32464);
nor U34435 (N_34435,N_32087,N_33770);
nand U34436 (N_34436,N_33983,N_33677);
nand U34437 (N_34437,N_33268,N_32750);
xnor U34438 (N_34438,N_32590,N_32000);
or U34439 (N_34439,N_33310,N_32621);
or U34440 (N_34440,N_32487,N_32447);
nor U34441 (N_34441,N_32647,N_33885);
xnor U34442 (N_34442,N_32633,N_33069);
nor U34443 (N_34443,N_33863,N_32110);
or U34444 (N_34444,N_32253,N_32233);
and U34445 (N_34445,N_32563,N_33057);
and U34446 (N_34446,N_32180,N_32191);
and U34447 (N_34447,N_33948,N_33954);
and U34448 (N_34448,N_33696,N_32281);
nand U34449 (N_34449,N_32956,N_32144);
nand U34450 (N_34450,N_33099,N_33040);
nor U34451 (N_34451,N_33734,N_33305);
nand U34452 (N_34452,N_33715,N_33152);
and U34453 (N_34453,N_33088,N_32283);
or U34454 (N_34454,N_33382,N_32535);
or U34455 (N_34455,N_33518,N_32071);
xnor U34456 (N_34456,N_33714,N_32429);
xnor U34457 (N_34457,N_33149,N_33626);
xor U34458 (N_34458,N_33240,N_33916);
and U34459 (N_34459,N_32426,N_32305);
nand U34460 (N_34460,N_32194,N_33417);
xor U34461 (N_34461,N_32818,N_32358);
nand U34462 (N_34462,N_33421,N_33788);
nor U34463 (N_34463,N_32254,N_32050);
nor U34464 (N_34464,N_32008,N_32759);
or U34465 (N_34465,N_32160,N_33339);
xor U34466 (N_34466,N_32284,N_33752);
nand U34467 (N_34467,N_33052,N_32200);
xor U34468 (N_34468,N_32850,N_33367);
nor U34469 (N_34469,N_32803,N_33344);
nor U34470 (N_34470,N_32046,N_33675);
or U34471 (N_34471,N_32458,N_32221);
or U34472 (N_34472,N_33860,N_32245);
xor U34473 (N_34473,N_32558,N_33121);
nand U34474 (N_34474,N_33995,N_33431);
xnor U34475 (N_34475,N_33500,N_33625);
and U34476 (N_34476,N_33002,N_33087);
nor U34477 (N_34477,N_32870,N_33969);
xor U34478 (N_34478,N_33325,N_33409);
nand U34479 (N_34479,N_33276,N_32592);
or U34480 (N_34480,N_33987,N_33704);
nand U34481 (N_34481,N_33123,N_32134);
xor U34482 (N_34482,N_33196,N_33377);
xnor U34483 (N_34483,N_32334,N_32185);
nand U34484 (N_34484,N_32920,N_33266);
nor U34485 (N_34485,N_32179,N_33483);
and U34486 (N_34486,N_32554,N_32914);
and U34487 (N_34487,N_33856,N_33812);
xnor U34488 (N_34488,N_32671,N_32032);
nor U34489 (N_34489,N_32991,N_33097);
xnor U34490 (N_34490,N_33718,N_33772);
and U34491 (N_34491,N_33893,N_32502);
xnor U34492 (N_34492,N_33679,N_33907);
nor U34493 (N_34493,N_33238,N_32114);
xnor U34494 (N_34494,N_33859,N_33473);
nor U34495 (N_34495,N_33853,N_32786);
nor U34496 (N_34496,N_33391,N_33834);
nor U34497 (N_34497,N_33146,N_33013);
xor U34498 (N_34498,N_32058,N_32182);
or U34499 (N_34499,N_33647,N_33638);
xnor U34500 (N_34500,N_32754,N_32183);
nand U34501 (N_34501,N_32168,N_33908);
xnor U34502 (N_34502,N_32304,N_32514);
xor U34503 (N_34503,N_32787,N_33436);
nor U34504 (N_34504,N_32181,N_33996);
nor U34505 (N_34505,N_33393,N_33072);
or U34506 (N_34506,N_32527,N_33179);
nand U34507 (N_34507,N_32856,N_33120);
and U34508 (N_34508,N_33105,N_33577);
nor U34509 (N_34509,N_33438,N_33019);
and U34510 (N_34510,N_33455,N_33967);
and U34511 (N_34511,N_33353,N_32272);
xnor U34512 (N_34512,N_32785,N_33635);
nand U34513 (N_34513,N_32889,N_32068);
nor U34514 (N_34514,N_33270,N_33298);
xnor U34515 (N_34515,N_33864,N_33979);
nor U34516 (N_34516,N_32488,N_32622);
or U34517 (N_34517,N_32105,N_32990);
xor U34518 (N_34518,N_33509,N_33207);
nor U34519 (N_34519,N_32146,N_33559);
nor U34520 (N_34520,N_32333,N_33735);
and U34521 (N_34521,N_32479,N_33176);
nand U34522 (N_34522,N_33880,N_32278);
nor U34523 (N_34523,N_32196,N_33313);
or U34524 (N_34524,N_33101,N_32021);
and U34525 (N_34525,N_32476,N_32270);
and U34526 (N_34526,N_33295,N_33582);
nand U34527 (N_34527,N_32880,N_32659);
and U34528 (N_34528,N_32384,N_32335);
or U34529 (N_34529,N_33030,N_33553);
xnor U34530 (N_34530,N_32650,N_33458);
nor U34531 (N_34531,N_32783,N_32092);
xor U34532 (N_34532,N_32222,N_32425);
nor U34533 (N_34533,N_32642,N_33980);
nand U34534 (N_34534,N_32824,N_32011);
nor U34535 (N_34535,N_33527,N_32374);
nand U34536 (N_34536,N_33319,N_32848);
nand U34537 (N_34537,N_32865,N_33966);
nor U34538 (N_34538,N_32148,N_33632);
xor U34539 (N_34539,N_33474,N_32793);
xor U34540 (N_34540,N_32193,N_33156);
nand U34541 (N_34541,N_33362,N_33333);
nand U34542 (N_34542,N_33229,N_33226);
xnor U34543 (N_34543,N_33224,N_32547);
and U34544 (N_34544,N_32117,N_32410);
xnor U34545 (N_34545,N_32809,N_33356);
and U34546 (N_34546,N_33073,N_32749);
or U34547 (N_34547,N_33280,N_33219);
nand U34548 (N_34548,N_32190,N_33463);
or U34549 (N_34549,N_33114,N_32801);
or U34550 (N_34550,N_33489,N_33572);
and U34551 (N_34551,N_32967,N_32534);
or U34552 (N_34552,N_33701,N_32600);
and U34553 (N_34553,N_33930,N_33291);
nor U34554 (N_34554,N_33071,N_33990);
or U34555 (N_34555,N_32553,N_33982);
nand U34556 (N_34556,N_33267,N_33672);
xnor U34557 (N_34557,N_33894,N_32314);
xnor U34558 (N_34558,N_33829,N_32437);
xnor U34559 (N_34559,N_32587,N_32307);
nor U34560 (N_34560,N_32282,N_33297);
nand U34561 (N_34561,N_33000,N_33633);
nand U34562 (N_34562,N_33970,N_32056);
nor U34563 (N_34563,N_32259,N_33936);
nor U34564 (N_34564,N_32570,N_32567);
xor U34565 (N_34565,N_32548,N_33617);
nand U34566 (N_34566,N_33279,N_33027);
nor U34567 (N_34567,N_32427,N_33836);
or U34568 (N_34568,N_32517,N_32766);
xor U34569 (N_34569,N_33540,N_33326);
xor U34570 (N_34570,N_32460,N_33917);
and U34571 (N_34571,N_32065,N_33763);
nand U34572 (N_34572,N_33771,N_32154);
and U34573 (N_34573,N_33419,N_32036);
nand U34574 (N_34574,N_32505,N_33444);
and U34575 (N_34575,N_33148,N_33514);
nand U34576 (N_34576,N_32312,N_32139);
and U34577 (N_34577,N_32896,N_32330);
and U34578 (N_34578,N_32377,N_33163);
xnor U34579 (N_34579,N_32328,N_32201);
nand U34580 (N_34580,N_32477,N_33301);
xor U34581 (N_34581,N_32354,N_33304);
or U34582 (N_34582,N_32170,N_32064);
and U34583 (N_34583,N_33112,N_33273);
or U34584 (N_34584,N_33162,N_32790);
nand U34585 (N_34585,N_32137,N_33102);
xor U34586 (N_34586,N_32263,N_33719);
or U34587 (N_34587,N_33343,N_32186);
xnor U34588 (N_34588,N_33538,N_33921);
nand U34589 (N_34589,N_33871,N_32516);
and U34590 (N_34590,N_33643,N_33840);
and U34591 (N_34591,N_33511,N_32574);
or U34592 (N_34592,N_33243,N_32365);
nor U34593 (N_34593,N_32523,N_32892);
nand U34594 (N_34594,N_32834,N_32656);
and U34595 (N_34595,N_33283,N_32828);
and U34596 (N_34596,N_33792,N_32812);
xor U34597 (N_34597,N_33855,N_33657);
xor U34598 (N_34598,N_33502,N_33197);
and U34599 (N_34599,N_33009,N_32760);
nand U34600 (N_34600,N_32911,N_33336);
nand U34601 (N_34601,N_32291,N_32765);
nor U34602 (N_34602,N_32657,N_33857);
or U34603 (N_34603,N_32158,N_33753);
and U34604 (N_34604,N_33274,N_32352);
xnor U34605 (N_34605,N_32411,N_32686);
nor U34606 (N_34606,N_33365,N_32152);
nor U34607 (N_34607,N_32939,N_33510);
nand U34608 (N_34608,N_33956,N_33375);
xor U34609 (N_34609,N_33203,N_32266);
nor U34610 (N_34610,N_33466,N_32727);
or U34611 (N_34611,N_32088,N_33031);
xor U34612 (N_34612,N_32971,N_33731);
xor U34613 (N_34613,N_33503,N_33352);
nand U34614 (N_34614,N_33006,N_32322);
and U34615 (N_34615,N_32832,N_32560);
nor U34616 (N_34616,N_32124,N_33217);
nor U34617 (N_34617,N_32135,N_33174);
or U34618 (N_34618,N_33898,N_32925);
and U34619 (N_34619,N_33100,N_33765);
xor U34620 (N_34620,N_32569,N_33660);
nand U34621 (N_34621,N_33960,N_32321);
nor U34622 (N_34622,N_33939,N_32249);
or U34623 (N_34623,N_33384,N_32404);
and U34624 (N_34624,N_33545,N_33236);
and U34625 (N_34625,N_32854,N_32257);
nor U34626 (N_34626,N_33876,N_33634);
or U34627 (N_34627,N_33357,N_33315);
and U34628 (N_34628,N_32066,N_33636);
nor U34629 (N_34629,N_32264,N_32646);
nor U34630 (N_34630,N_33172,N_32705);
xnor U34631 (N_34631,N_32473,N_33015);
nor U34632 (N_34632,N_33681,N_32346);
xor U34633 (N_34633,N_32373,N_32871);
xnor U34634 (N_34634,N_32992,N_33113);
nor U34635 (N_34635,N_32778,N_33459);
nand U34636 (N_34636,N_32385,N_33249);
xnor U34637 (N_34637,N_33694,N_33194);
nand U34638 (N_34638,N_32026,N_33420);
nor U34639 (N_34639,N_33103,N_32718);
or U34640 (N_34640,N_33940,N_33747);
and U34641 (N_34641,N_32912,N_33195);
and U34642 (N_34642,N_32841,N_32981);
nor U34643 (N_34643,N_32945,N_32340);
nor U34644 (N_34644,N_33461,N_32875);
nor U34645 (N_34645,N_32868,N_33620);
nand U34646 (N_34646,N_33845,N_32408);
and U34647 (N_34647,N_32423,N_33437);
nand U34648 (N_34648,N_32239,N_32302);
or U34649 (N_34649,N_32261,N_32187);
nor U34650 (N_34650,N_33415,N_32043);
or U34651 (N_34651,N_33016,N_32983);
nor U34652 (N_34652,N_33277,N_32332);
and U34653 (N_34653,N_32238,N_32470);
nor U34654 (N_34654,N_32739,N_33046);
or U34655 (N_34655,N_32591,N_33685);
and U34656 (N_34656,N_33410,N_32929);
and U34657 (N_34657,N_32952,N_33414);
and U34658 (N_34658,N_33284,N_33080);
and U34659 (N_34659,N_33110,N_33079);
nor U34660 (N_34660,N_33888,N_33984);
and U34661 (N_34661,N_32954,N_32035);
nand U34662 (N_34662,N_33600,N_32608);
and U34663 (N_34663,N_32159,N_32964);
xor U34664 (N_34664,N_33760,N_33562);
or U34665 (N_34665,N_33815,N_33094);
or U34666 (N_34666,N_33673,N_32767);
or U34667 (N_34667,N_32723,N_33359);
and U34668 (N_34668,N_33613,N_32317);
or U34669 (N_34669,N_32998,N_32073);
xnor U34670 (N_34670,N_32835,N_33076);
nand U34671 (N_34671,N_33826,N_32593);
xnor U34672 (N_34672,N_33745,N_33697);
or U34673 (N_34673,N_32546,N_32645);
nand U34674 (N_34674,N_32004,N_32138);
nor U34675 (N_34675,N_32501,N_33570);
nand U34676 (N_34676,N_33656,N_32543);
nand U34677 (N_34677,N_32604,N_33631);
and U34678 (N_34678,N_33791,N_32610);
nor U34679 (N_34679,N_32274,N_32486);
nor U34680 (N_34680,N_32589,N_33067);
nor U34681 (N_34681,N_32145,N_32542);
and U34682 (N_34682,N_32205,N_32520);
nand U34683 (N_34683,N_32466,N_33564);
nand U34684 (N_34684,N_33579,N_33981);
xnor U34685 (N_34685,N_32849,N_32407);
nand U34686 (N_34686,N_33910,N_32140);
or U34687 (N_34687,N_33729,N_32132);
nand U34688 (N_34688,N_33612,N_33150);
nor U34689 (N_34689,N_32450,N_33248);
nand U34690 (N_34690,N_33232,N_33655);
and U34691 (N_34691,N_33964,N_33056);
nor U34692 (N_34692,N_32820,N_33129);
nor U34693 (N_34693,N_33802,N_32297);
and U34694 (N_34694,N_33602,N_33727);
and U34695 (N_34695,N_33053,N_33640);
and U34696 (N_34696,N_32442,N_33498);
xor U34697 (N_34697,N_33145,N_32710);
or U34698 (N_34698,N_33302,N_32415);
or U34699 (N_34699,N_32141,N_32744);
xnor U34700 (N_34700,N_33610,N_32768);
and U34701 (N_34701,N_33160,N_32361);
nor U34702 (N_34702,N_33522,N_32582);
or U34703 (N_34703,N_32588,N_32751);
xnor U34704 (N_34704,N_32096,N_32894);
nor U34705 (N_34705,N_32872,N_33989);
nor U34706 (N_34706,N_33905,N_33823);
xor U34707 (N_34707,N_33821,N_32237);
nand U34708 (N_34708,N_32199,N_33104);
xor U34709 (N_34709,N_33682,N_32687);
xnor U34710 (N_34710,N_32729,N_33756);
or U34711 (N_34711,N_32821,N_32463);
and U34712 (N_34712,N_33968,N_32947);
or U34713 (N_34713,N_32120,N_33107);
nand U34714 (N_34714,N_33892,N_33737);
and U34715 (N_34715,N_32164,N_33795);
and U34716 (N_34716,N_33401,N_32095);
or U34717 (N_34717,N_32531,N_33890);
or U34718 (N_34718,N_32612,N_32029);
nand U34719 (N_34719,N_33807,N_33587);
xor U34720 (N_34720,N_33662,N_33528);
nor U34721 (N_34721,N_33494,N_32371);
and U34722 (N_34722,N_33974,N_32695);
xnor U34723 (N_34723,N_32448,N_33849);
and U34724 (N_34724,N_32958,N_32122);
and U34725 (N_34725,N_32076,N_32419);
nand U34726 (N_34726,N_33137,N_32357);
and U34727 (N_34727,N_33412,N_33900);
or U34728 (N_34728,N_32541,N_33300);
nand U34729 (N_34729,N_32089,N_33262);
or U34730 (N_34730,N_32102,N_33452);
xnor U34731 (N_34731,N_32731,N_33667);
xnor U34732 (N_34732,N_32434,N_32805);
or U34733 (N_34733,N_33154,N_33955);
xor U34734 (N_34734,N_33388,N_32107);
and U34735 (N_34735,N_32690,N_32602);
nor U34736 (N_34736,N_32398,N_33476);
xor U34737 (N_34737,N_32465,N_33092);
nand U34738 (N_34738,N_32944,N_32901);
nand U34739 (N_34739,N_32112,N_32468);
or U34740 (N_34740,N_32987,N_33711);
nand U34741 (N_34741,N_32490,N_32128);
nand U34742 (N_34742,N_32443,N_32489);
xnor U34743 (N_34743,N_33012,N_33654);
or U34744 (N_34744,N_32287,N_33428);
nor U34745 (N_34745,N_32839,N_32922);
or U34746 (N_34746,N_32166,N_32300);
nor U34747 (N_34747,N_32549,N_32791);
or U34748 (N_34748,N_33085,N_33915);
and U34749 (N_34749,N_33604,N_33117);
nor U34750 (N_34750,N_32617,N_32231);
xor U34751 (N_34751,N_33761,N_32027);
nor U34752 (N_34752,N_32782,N_32130);
or U34753 (N_34753,N_33322,N_32269);
nor U34754 (N_34754,N_32387,N_32708);
nand U34755 (N_34755,N_33622,N_33201);
nand U34756 (N_34756,N_32356,N_33208);
nand U34757 (N_34757,N_32165,N_32386);
nand U34758 (N_34758,N_33376,N_32714);
nand U34759 (N_34759,N_33693,N_33433);
or U34760 (N_34760,N_32559,N_33358);
or U34761 (N_34761,N_33445,N_32081);
nor U34762 (N_34762,N_32630,N_32680);
xnor U34763 (N_34763,N_32455,N_32565);
or U34764 (N_34764,N_33878,N_32761);
nand U34765 (N_34765,N_32683,N_33837);
and U34766 (N_34766,N_33843,N_33637);
nand U34767 (N_34767,N_33383,N_32030);
and U34768 (N_34768,N_33767,N_33589);
nand U34769 (N_34769,N_33198,N_33776);
nand U34770 (N_34770,N_32418,N_33549);
xnor U34771 (N_34771,N_33748,N_32157);
or U34772 (N_34772,N_32701,N_33406);
xnor U34773 (N_34773,N_32495,N_32813);
nor U34774 (N_34774,N_33165,N_32679);
xnor U34775 (N_34775,N_33039,N_32224);
and U34776 (N_34776,N_32605,N_33331);
or U34777 (N_34777,N_33773,N_32946);
nor U34778 (N_34778,N_32176,N_32519);
xnor U34779 (N_34779,N_32005,N_32206);
nor U34780 (N_34780,N_32988,N_32891);
and U34781 (N_34781,N_32658,N_32085);
nor U34782 (N_34782,N_32319,N_33218);
nand U34783 (N_34783,N_33460,N_32235);
xor U34784 (N_34784,N_32260,N_32530);
or U34785 (N_34785,N_32806,N_33022);
and U34786 (N_34786,N_33586,N_33159);
and U34787 (N_34787,N_33034,N_33728);
xor U34788 (N_34788,N_33351,N_32715);
nor U34789 (N_34789,N_33713,N_32057);
nand U34790 (N_34790,N_32713,N_33381);
nor U34791 (N_34791,N_33407,N_32339);
and U34792 (N_34792,N_33242,N_33874);
xor U34793 (N_34793,N_33096,N_33523);
xnor U34794 (N_34794,N_32773,N_32475);
and U34795 (N_34795,N_33965,N_32262);
xor U34796 (N_34796,N_32079,N_32351);
or U34797 (N_34797,N_32933,N_32598);
and U34798 (N_34798,N_32323,N_32230);
nor U34799 (N_34799,N_32525,N_33418);
xnor U34800 (N_34800,N_33858,N_32022);
xor U34801 (N_34801,N_33051,N_33943);
and U34802 (N_34802,N_32537,N_32147);
and U34803 (N_34803,N_32628,N_33282);
and U34804 (N_34804,N_33605,N_33595);
nand U34805 (N_34805,N_33779,N_33014);
or U34806 (N_34806,N_33387,N_33963);
nor U34807 (N_34807,N_32118,N_33976);
nand U34808 (N_34808,N_32031,N_32198);
or U34809 (N_34809,N_33766,N_33556);
or U34810 (N_34810,N_32382,N_33497);
xor U34811 (N_34811,N_32214,N_33134);
nor U34812 (N_34812,N_32131,N_33918);
and U34813 (N_34813,N_33370,N_32626);
or U34814 (N_34814,N_32507,N_32877);
nor U34815 (N_34815,N_33535,N_33018);
or U34816 (N_34816,N_32694,N_33790);
and U34817 (N_34817,N_33583,N_32561);
nand U34818 (N_34818,N_33877,N_33588);
nor U34819 (N_34819,N_33759,N_32775);
nand U34820 (N_34820,N_33873,N_33749);
and U34821 (N_34821,N_33513,N_32344);
nand U34822 (N_34822,N_33794,N_32959);
or U34823 (N_34823,N_32741,N_32637);
xor U34824 (N_34824,N_32724,N_32223);
xor U34825 (N_34825,N_33128,N_32252);
or U34826 (N_34826,N_32973,N_33891);
or U34827 (N_34827,N_33182,N_33835);
nor U34828 (N_34828,N_32660,N_33271);
xor U34829 (N_34829,N_32888,N_32391);
nor U34830 (N_34830,N_33078,N_32308);
nor U34831 (N_34831,N_33730,N_33945);
and U34832 (N_34832,N_33757,N_32700);
nor U34833 (N_34833,N_33666,N_33021);
and U34834 (N_34834,N_33082,N_33536);
and U34835 (N_34835,N_33953,N_33844);
nand U34836 (N_34836,N_33010,N_32481);
nand U34837 (N_34837,N_33775,N_33519);
xnor U34838 (N_34838,N_33093,N_32016);
and U34839 (N_34839,N_33573,N_32298);
and U34840 (N_34840,N_33191,N_32676);
or U34841 (N_34841,N_32098,N_32345);
nor U34842 (N_34842,N_33869,N_33077);
or U34843 (N_34843,N_32712,N_33689);
xnor U34844 (N_34844,N_32493,N_32368);
and U34845 (N_34845,N_32995,N_33426);
and U34846 (N_34846,N_32725,N_33400);
nor U34847 (N_34847,N_32432,N_32609);
nor U34848 (N_34848,N_33616,N_33904);
nand U34849 (N_34849,N_33591,N_32620);
nand U34850 (N_34850,N_32928,N_33615);
nand U34851 (N_34851,N_33167,N_33798);
xor U34852 (N_34852,N_32383,N_32855);
nor U34853 (N_34853,N_33126,N_32108);
nor U34854 (N_34854,N_33645,N_32080);
nor U34855 (N_34855,N_32616,N_33593);
and U34856 (N_34856,N_33075,N_32584);
nand U34857 (N_34857,N_32902,N_33166);
nand U34858 (N_34858,N_33171,N_32578);
nand U34859 (N_34859,N_33230,N_33872);
and U34860 (N_34860,N_32072,N_32916);
xor U34861 (N_34861,N_33668,N_32900);
nor U34862 (N_34862,N_32104,N_33861);
or U34863 (N_34863,N_32250,N_33957);
nor U34864 (N_34864,N_33566,N_32963);
xor U34865 (N_34865,N_32681,N_32682);
nand U34866 (N_34866,N_33919,N_33803);
or U34867 (N_34867,N_33558,N_33446);
xor U34868 (N_34868,N_32303,N_32126);
nor U34869 (N_34869,N_33329,N_32246);
nand U34870 (N_34870,N_33004,N_33480);
nand U34871 (N_34871,N_32039,N_32173);
xor U34872 (N_34872,N_32293,N_32733);
and U34873 (N_34873,N_32585,N_33299);
and U34874 (N_34874,N_32953,N_33378);
nand U34875 (N_34875,N_33131,N_33454);
or U34876 (N_34876,N_33628,N_32545);
and U34877 (N_34877,N_33959,N_32420);
or U34878 (N_34878,N_33244,N_33700);
and U34879 (N_34879,N_32931,N_33361);
nand U34880 (N_34880,N_32632,N_32509);
nand U34881 (N_34881,N_33422,N_32483);
nand U34882 (N_34882,N_32950,N_32438);
xor U34883 (N_34883,N_33642,N_32917);
nand U34884 (N_34884,N_33740,N_32568);
and U34885 (N_34885,N_33108,N_33448);
nor U34886 (N_34886,N_32195,N_33578);
nand U34887 (N_34887,N_32038,N_33590);
nand U34888 (N_34888,N_32037,N_32456);
nor U34889 (N_34889,N_33937,N_32299);
and U34890 (N_34890,N_33717,N_33561);
xor U34891 (N_34891,N_32927,N_33441);
and U34892 (N_34892,N_32439,N_32055);
and U34893 (N_34893,N_32271,N_33161);
xor U34894 (N_34894,N_32213,N_33140);
or U34895 (N_34895,N_32013,N_33852);
nand U34896 (N_34896,N_32726,N_32215);
xor U34897 (N_34897,N_32379,N_32513);
nand U34898 (N_34898,N_32020,N_33665);
or U34899 (N_34899,N_33971,N_33133);
nor U34900 (N_34900,N_32417,N_32225);
and U34901 (N_34901,N_32086,N_33592);
nand U34902 (N_34902,N_32838,N_33281);
nand U34903 (N_34903,N_33153,N_32918);
or U34904 (N_34904,N_32943,N_33462);
nor U34905 (N_34905,N_33327,N_32248);
nand U34906 (N_34906,N_32067,N_32207);
nand U34907 (N_34907,N_32472,N_33138);
or U34908 (N_34908,N_32433,N_32776);
and U34909 (N_34909,N_32151,N_32033);
nand U34910 (N_34910,N_33286,N_32975);
or U34911 (N_34911,N_32538,N_33366);
nand U34912 (N_34912,N_32800,N_33275);
and U34913 (N_34913,N_32452,N_33809);
xor U34914 (N_34914,N_33922,N_32241);
and U34915 (N_34915,N_32077,N_32978);
xor U34916 (N_34916,N_33321,N_32136);
or U34917 (N_34917,N_33935,N_32529);
xnor U34918 (N_34918,N_32403,N_32052);
and U34919 (N_34919,N_32327,N_32572);
or U34920 (N_34920,N_33952,N_33754);
nor U34921 (N_34921,N_33674,N_33404);
nor U34922 (N_34922,N_33398,N_33482);
nand U34923 (N_34923,N_32583,N_33649);
and U34924 (N_34924,N_33373,N_33449);
xnor U34925 (N_34925,N_32449,N_33781);
nand U34926 (N_34926,N_33235,N_32655);
or U34927 (N_34927,N_33822,N_32816);
and U34928 (N_34928,N_32500,N_32599);
nand U34929 (N_34929,N_32015,N_32440);
xnor U34930 (N_34930,N_32840,N_32349);
nand U34931 (N_34931,N_33546,N_33200);
or U34932 (N_34932,N_32898,N_32972);
xnor U34933 (N_34933,N_32424,N_33816);
nand U34934 (N_34934,N_32211,N_33886);
or U34935 (N_34935,N_33780,N_33949);
nor U34936 (N_34936,N_33515,N_32756);
and U34937 (N_34937,N_33576,N_33026);
nand U34938 (N_34938,N_33819,N_33975);
nor U34939 (N_34939,N_33048,N_32372);
xnor U34940 (N_34940,N_33973,N_32405);
nand U34941 (N_34941,N_33768,N_32861);
and U34942 (N_34942,N_32106,N_32451);
and U34943 (N_34943,N_32536,N_32388);
xnor U34944 (N_34944,N_33851,N_33563);
or U34945 (N_34945,N_33346,N_33830);
nor U34946 (N_34946,N_32226,N_33223);
or U34947 (N_34947,N_32974,N_32692);
nand U34948 (N_34948,N_33508,N_32728);
nor U34949 (N_34949,N_32935,N_32797);
nand U34950 (N_34950,N_33712,N_32930);
nor U34951 (N_34951,N_32024,N_32665);
xor U34952 (N_34952,N_33290,N_33173);
nand U34953 (N_34953,N_32890,N_32040);
xor U34954 (N_34954,N_32028,N_32409);
nor U34955 (N_34955,N_32025,N_32666);
xnor U34956 (N_34956,N_32510,N_32926);
or U34957 (N_34957,N_33456,N_33557);
or U34958 (N_34958,N_33037,N_33371);
nor U34959 (N_34959,N_33525,N_32831);
xor U34960 (N_34960,N_33250,N_32638);
xor U34961 (N_34961,N_32829,N_32799);
and U34962 (N_34962,N_32381,N_33332);
nand U34963 (N_34963,N_32216,N_33465);
and U34964 (N_34964,N_32771,N_33653);
and U34965 (N_34965,N_33125,N_33746);
xnor U34966 (N_34966,N_33481,N_32746);
xnor U34967 (N_34967,N_32674,N_32101);
xnor U34968 (N_34968,N_33827,N_32721);
nor U34969 (N_34969,N_32904,N_32338);
nor U34970 (N_34970,N_32390,N_33927);
xor U34971 (N_34971,N_32580,N_32980);
xnor U34972 (N_34972,N_33369,N_32709);
nor U34973 (N_34973,N_32949,N_33064);
nor U34974 (N_34974,N_33065,N_32018);
xnor U34975 (N_34975,N_32649,N_32860);
xor U34976 (N_34976,N_32275,N_33135);
xnor U34977 (N_34977,N_32467,N_33312);
xor U34978 (N_34978,N_33897,N_33548);
nor U34979 (N_34979,N_33552,N_32576);
or U34980 (N_34980,N_33169,N_32999);
or U34981 (N_34981,N_32597,N_33755);
nand U34982 (N_34982,N_33209,N_32698);
nand U34983 (N_34983,N_32506,N_33993);
xnor U34984 (N_34984,N_32273,N_32903);
nor U34985 (N_34985,N_32586,N_33029);
xor U34986 (N_34986,N_32895,N_33115);
or U34987 (N_34987,N_33650,N_33716);
nand U34988 (N_34988,N_32689,N_32936);
nand U34989 (N_34989,N_33424,N_32562);
or U34990 (N_34990,N_32232,N_33435);
nor U34991 (N_34991,N_32747,N_33598);
nor U34992 (N_34992,N_32555,N_33177);
nor U34993 (N_34993,N_32208,N_33261);
nand U34994 (N_34994,N_32827,N_33269);
xnor U34995 (N_34995,N_32702,N_33671);
and U34996 (N_34996,N_33136,N_33447);
xnor U34997 (N_34997,N_33865,N_33560);
and U34998 (N_34998,N_33399,N_33451);
and U34999 (N_34999,N_32406,N_33722);
xnor U35000 (N_35000,N_32615,N_32370);
or U35001 (N_35001,N_32666,N_32611);
or U35002 (N_35002,N_33820,N_32744);
or U35003 (N_35003,N_33279,N_32876);
nor U35004 (N_35004,N_33238,N_33233);
and U35005 (N_35005,N_33835,N_32313);
and U35006 (N_35006,N_33244,N_32625);
nand U35007 (N_35007,N_32900,N_33601);
and U35008 (N_35008,N_32572,N_33573);
and U35009 (N_35009,N_32399,N_32567);
xor U35010 (N_35010,N_33094,N_32228);
nor U35011 (N_35011,N_33158,N_32139);
and U35012 (N_35012,N_33204,N_33561);
nor U35013 (N_35013,N_32453,N_32720);
and U35014 (N_35014,N_32165,N_33993);
or U35015 (N_35015,N_32299,N_32448);
or U35016 (N_35016,N_33782,N_32967);
or U35017 (N_35017,N_32266,N_33189);
or U35018 (N_35018,N_33365,N_32319);
and U35019 (N_35019,N_33291,N_33808);
xnor U35020 (N_35020,N_32470,N_32979);
or U35021 (N_35021,N_33307,N_32936);
xor U35022 (N_35022,N_32446,N_33587);
and U35023 (N_35023,N_33958,N_33633);
nor U35024 (N_35024,N_33939,N_33623);
and U35025 (N_35025,N_33829,N_33577);
nor U35026 (N_35026,N_32596,N_33907);
and U35027 (N_35027,N_32093,N_32205);
nor U35028 (N_35028,N_32079,N_32340);
and U35029 (N_35029,N_33676,N_33045);
or U35030 (N_35030,N_33550,N_33536);
nand U35031 (N_35031,N_33003,N_32546);
and U35032 (N_35032,N_32639,N_32238);
nor U35033 (N_35033,N_32633,N_32409);
xor U35034 (N_35034,N_33512,N_33791);
or U35035 (N_35035,N_32217,N_32141);
or U35036 (N_35036,N_33882,N_33630);
and U35037 (N_35037,N_33606,N_32834);
nor U35038 (N_35038,N_33922,N_33831);
and U35039 (N_35039,N_33009,N_32348);
or U35040 (N_35040,N_32312,N_33417);
and U35041 (N_35041,N_32202,N_32776);
nor U35042 (N_35042,N_33577,N_32748);
xnor U35043 (N_35043,N_32962,N_32010);
and U35044 (N_35044,N_33882,N_33581);
and U35045 (N_35045,N_33469,N_32646);
nor U35046 (N_35046,N_33157,N_32063);
or U35047 (N_35047,N_33523,N_33008);
nor U35048 (N_35048,N_32350,N_33757);
or U35049 (N_35049,N_33293,N_33757);
nand U35050 (N_35050,N_33742,N_32826);
nor U35051 (N_35051,N_33613,N_33506);
nand U35052 (N_35052,N_32050,N_32804);
or U35053 (N_35053,N_32225,N_32271);
xnor U35054 (N_35054,N_32720,N_32035);
nor U35055 (N_35055,N_33905,N_32729);
xnor U35056 (N_35056,N_33304,N_32746);
xnor U35057 (N_35057,N_33277,N_33073);
nor U35058 (N_35058,N_33514,N_32399);
or U35059 (N_35059,N_32154,N_33384);
and U35060 (N_35060,N_32486,N_32818);
and U35061 (N_35061,N_33930,N_32137);
xnor U35062 (N_35062,N_32800,N_33658);
xnor U35063 (N_35063,N_32012,N_33382);
xnor U35064 (N_35064,N_32986,N_32193);
xor U35065 (N_35065,N_33700,N_33935);
or U35066 (N_35066,N_32848,N_32335);
or U35067 (N_35067,N_33727,N_33121);
nand U35068 (N_35068,N_33167,N_33273);
or U35069 (N_35069,N_32705,N_33934);
nor U35070 (N_35070,N_33969,N_33248);
xor U35071 (N_35071,N_33998,N_33495);
or U35072 (N_35072,N_32174,N_33360);
and U35073 (N_35073,N_33603,N_33851);
xor U35074 (N_35074,N_33612,N_32171);
nor U35075 (N_35075,N_33689,N_33859);
or U35076 (N_35076,N_33669,N_33576);
xnor U35077 (N_35077,N_32498,N_33402);
nor U35078 (N_35078,N_32103,N_33442);
nand U35079 (N_35079,N_33201,N_33375);
and U35080 (N_35080,N_33120,N_33001);
or U35081 (N_35081,N_32102,N_32465);
nor U35082 (N_35082,N_33913,N_32958);
nor U35083 (N_35083,N_33421,N_33116);
and U35084 (N_35084,N_33013,N_33752);
nand U35085 (N_35085,N_33576,N_33637);
xnor U35086 (N_35086,N_32680,N_33909);
nand U35087 (N_35087,N_33026,N_33224);
nand U35088 (N_35088,N_32789,N_32644);
or U35089 (N_35089,N_33297,N_32646);
nor U35090 (N_35090,N_32438,N_32543);
xor U35091 (N_35091,N_33915,N_33780);
xor U35092 (N_35092,N_33483,N_32805);
or U35093 (N_35093,N_33113,N_32162);
nand U35094 (N_35094,N_33003,N_32272);
nand U35095 (N_35095,N_32330,N_32331);
nand U35096 (N_35096,N_33406,N_32782);
or U35097 (N_35097,N_33096,N_33931);
and U35098 (N_35098,N_32656,N_32638);
nor U35099 (N_35099,N_32698,N_33365);
nand U35100 (N_35100,N_33453,N_33997);
xor U35101 (N_35101,N_33794,N_33751);
and U35102 (N_35102,N_33274,N_33317);
or U35103 (N_35103,N_33871,N_33113);
nor U35104 (N_35104,N_33217,N_32482);
and U35105 (N_35105,N_32267,N_33375);
nand U35106 (N_35106,N_32514,N_32152);
or U35107 (N_35107,N_33382,N_32609);
or U35108 (N_35108,N_32466,N_32190);
xnor U35109 (N_35109,N_33222,N_32113);
nor U35110 (N_35110,N_33071,N_33802);
and U35111 (N_35111,N_33944,N_32943);
nand U35112 (N_35112,N_32431,N_32689);
and U35113 (N_35113,N_33000,N_33404);
xnor U35114 (N_35114,N_33322,N_32775);
and U35115 (N_35115,N_32642,N_33750);
or U35116 (N_35116,N_33252,N_32260);
or U35117 (N_35117,N_33610,N_33189);
or U35118 (N_35118,N_32679,N_32498);
nand U35119 (N_35119,N_32160,N_32392);
nand U35120 (N_35120,N_32323,N_32689);
xor U35121 (N_35121,N_33566,N_33303);
or U35122 (N_35122,N_32736,N_32240);
nand U35123 (N_35123,N_33304,N_32601);
or U35124 (N_35124,N_32446,N_33186);
and U35125 (N_35125,N_33352,N_32559);
xor U35126 (N_35126,N_32518,N_32365);
and U35127 (N_35127,N_32822,N_32046);
and U35128 (N_35128,N_33486,N_32066);
nand U35129 (N_35129,N_32706,N_33220);
nand U35130 (N_35130,N_32521,N_32401);
and U35131 (N_35131,N_32698,N_32371);
nor U35132 (N_35132,N_32477,N_33181);
or U35133 (N_35133,N_32552,N_33693);
nor U35134 (N_35134,N_33599,N_33485);
xnor U35135 (N_35135,N_32854,N_32452);
or U35136 (N_35136,N_33495,N_33726);
xor U35137 (N_35137,N_32758,N_33585);
or U35138 (N_35138,N_32087,N_32372);
or U35139 (N_35139,N_32495,N_33119);
nand U35140 (N_35140,N_32015,N_33825);
xor U35141 (N_35141,N_33010,N_33097);
and U35142 (N_35142,N_32228,N_32545);
and U35143 (N_35143,N_33869,N_32347);
nand U35144 (N_35144,N_32658,N_32899);
xor U35145 (N_35145,N_33045,N_32367);
nor U35146 (N_35146,N_33064,N_33373);
nor U35147 (N_35147,N_32216,N_32325);
xor U35148 (N_35148,N_32590,N_32469);
or U35149 (N_35149,N_32696,N_32550);
nand U35150 (N_35150,N_32065,N_32237);
xnor U35151 (N_35151,N_32130,N_33757);
nand U35152 (N_35152,N_32081,N_32340);
nand U35153 (N_35153,N_33990,N_32898);
or U35154 (N_35154,N_32513,N_33360);
and U35155 (N_35155,N_32856,N_33541);
nand U35156 (N_35156,N_32361,N_33240);
nor U35157 (N_35157,N_32182,N_33151);
xnor U35158 (N_35158,N_32658,N_33829);
and U35159 (N_35159,N_33492,N_33160);
and U35160 (N_35160,N_32999,N_33615);
or U35161 (N_35161,N_33909,N_32329);
or U35162 (N_35162,N_32130,N_33715);
or U35163 (N_35163,N_32671,N_33932);
xnor U35164 (N_35164,N_32196,N_32518);
nand U35165 (N_35165,N_32481,N_33077);
nand U35166 (N_35166,N_33642,N_33512);
nor U35167 (N_35167,N_32854,N_33196);
and U35168 (N_35168,N_33829,N_32888);
nor U35169 (N_35169,N_33089,N_32810);
xnor U35170 (N_35170,N_33807,N_33833);
xnor U35171 (N_35171,N_32192,N_33894);
nor U35172 (N_35172,N_33618,N_33202);
or U35173 (N_35173,N_33192,N_33857);
xor U35174 (N_35174,N_32062,N_32379);
nand U35175 (N_35175,N_32299,N_33355);
or U35176 (N_35176,N_32944,N_32306);
or U35177 (N_35177,N_32485,N_33674);
xor U35178 (N_35178,N_32753,N_33743);
xnor U35179 (N_35179,N_32467,N_33683);
or U35180 (N_35180,N_33682,N_32006);
and U35181 (N_35181,N_33971,N_33266);
xnor U35182 (N_35182,N_32001,N_32312);
and U35183 (N_35183,N_32823,N_33512);
nor U35184 (N_35184,N_32292,N_33049);
xnor U35185 (N_35185,N_32052,N_32747);
xnor U35186 (N_35186,N_33898,N_33943);
nor U35187 (N_35187,N_33408,N_33713);
and U35188 (N_35188,N_32513,N_32007);
or U35189 (N_35189,N_32651,N_33247);
xor U35190 (N_35190,N_32054,N_32997);
and U35191 (N_35191,N_32226,N_33491);
nor U35192 (N_35192,N_32403,N_33388);
or U35193 (N_35193,N_32063,N_32112);
or U35194 (N_35194,N_32929,N_33458);
and U35195 (N_35195,N_32372,N_33581);
or U35196 (N_35196,N_33741,N_32494);
xor U35197 (N_35197,N_32810,N_32019);
xor U35198 (N_35198,N_33032,N_33752);
and U35199 (N_35199,N_32057,N_33672);
xor U35200 (N_35200,N_33402,N_33178);
nand U35201 (N_35201,N_32253,N_32643);
and U35202 (N_35202,N_32856,N_33494);
nor U35203 (N_35203,N_33487,N_32633);
nand U35204 (N_35204,N_33421,N_33706);
nor U35205 (N_35205,N_33335,N_32225);
and U35206 (N_35206,N_33196,N_32622);
nand U35207 (N_35207,N_33113,N_32443);
nor U35208 (N_35208,N_32280,N_32806);
and U35209 (N_35209,N_32985,N_33143);
nor U35210 (N_35210,N_33763,N_32684);
nor U35211 (N_35211,N_33649,N_32391);
nand U35212 (N_35212,N_32300,N_32564);
xor U35213 (N_35213,N_33215,N_32540);
or U35214 (N_35214,N_33911,N_32324);
and U35215 (N_35215,N_32962,N_32109);
and U35216 (N_35216,N_32121,N_33364);
nand U35217 (N_35217,N_33888,N_32987);
xor U35218 (N_35218,N_32977,N_32136);
nand U35219 (N_35219,N_32461,N_32081);
nor U35220 (N_35220,N_32482,N_32722);
and U35221 (N_35221,N_33164,N_33052);
nor U35222 (N_35222,N_33996,N_32091);
nand U35223 (N_35223,N_32031,N_32513);
nor U35224 (N_35224,N_32827,N_33643);
xnor U35225 (N_35225,N_33005,N_33467);
nand U35226 (N_35226,N_32540,N_32448);
nand U35227 (N_35227,N_33178,N_32763);
xnor U35228 (N_35228,N_32396,N_32012);
or U35229 (N_35229,N_32373,N_33594);
nand U35230 (N_35230,N_33520,N_32350);
xor U35231 (N_35231,N_33067,N_32053);
nand U35232 (N_35232,N_33190,N_33502);
xor U35233 (N_35233,N_32958,N_33088);
and U35234 (N_35234,N_33822,N_32294);
nand U35235 (N_35235,N_32277,N_33767);
xnor U35236 (N_35236,N_32285,N_33382);
nor U35237 (N_35237,N_33058,N_33545);
or U35238 (N_35238,N_32330,N_33256);
xor U35239 (N_35239,N_32661,N_32576);
nand U35240 (N_35240,N_32106,N_33004);
xor U35241 (N_35241,N_32523,N_33732);
or U35242 (N_35242,N_32488,N_33156);
xnor U35243 (N_35243,N_32760,N_32183);
nand U35244 (N_35244,N_33342,N_33747);
or U35245 (N_35245,N_33593,N_32689);
or U35246 (N_35246,N_33127,N_33122);
xnor U35247 (N_35247,N_32832,N_33838);
and U35248 (N_35248,N_33765,N_32943);
or U35249 (N_35249,N_32565,N_33489);
nand U35250 (N_35250,N_33778,N_32796);
nor U35251 (N_35251,N_33003,N_32764);
nand U35252 (N_35252,N_33717,N_32966);
xor U35253 (N_35253,N_32383,N_32417);
xor U35254 (N_35254,N_33137,N_33689);
and U35255 (N_35255,N_33867,N_32108);
nand U35256 (N_35256,N_32569,N_33220);
nor U35257 (N_35257,N_32933,N_32688);
xnor U35258 (N_35258,N_32006,N_32844);
and U35259 (N_35259,N_33091,N_33010);
nor U35260 (N_35260,N_32281,N_32013);
xnor U35261 (N_35261,N_32819,N_32900);
xnor U35262 (N_35262,N_33451,N_32468);
nand U35263 (N_35263,N_32876,N_33506);
and U35264 (N_35264,N_32678,N_33863);
and U35265 (N_35265,N_32207,N_32363);
nor U35266 (N_35266,N_33702,N_33822);
or U35267 (N_35267,N_33579,N_33890);
nor U35268 (N_35268,N_32721,N_33758);
nor U35269 (N_35269,N_33316,N_33429);
nand U35270 (N_35270,N_33083,N_33475);
and U35271 (N_35271,N_33959,N_32278);
nor U35272 (N_35272,N_32384,N_33402);
and U35273 (N_35273,N_33724,N_33344);
nor U35274 (N_35274,N_32432,N_33241);
and U35275 (N_35275,N_33262,N_33839);
and U35276 (N_35276,N_33463,N_33487);
xnor U35277 (N_35277,N_33084,N_32391);
xnor U35278 (N_35278,N_33478,N_32834);
or U35279 (N_35279,N_33179,N_32193);
nand U35280 (N_35280,N_32704,N_33255);
nand U35281 (N_35281,N_32699,N_32497);
xnor U35282 (N_35282,N_33587,N_32530);
xnor U35283 (N_35283,N_32825,N_33916);
or U35284 (N_35284,N_32171,N_33250);
and U35285 (N_35285,N_32704,N_32619);
or U35286 (N_35286,N_32709,N_32495);
nor U35287 (N_35287,N_32225,N_33736);
nand U35288 (N_35288,N_33222,N_32700);
and U35289 (N_35289,N_33877,N_33701);
nor U35290 (N_35290,N_33251,N_33655);
nor U35291 (N_35291,N_32759,N_33007);
nand U35292 (N_35292,N_33486,N_33442);
xnor U35293 (N_35293,N_33243,N_32792);
nand U35294 (N_35294,N_32132,N_33324);
and U35295 (N_35295,N_33579,N_33548);
xor U35296 (N_35296,N_32166,N_33208);
nand U35297 (N_35297,N_33829,N_33417);
xor U35298 (N_35298,N_33007,N_32923);
nor U35299 (N_35299,N_33419,N_33477);
or U35300 (N_35300,N_32662,N_33556);
or U35301 (N_35301,N_33402,N_32355);
xor U35302 (N_35302,N_32673,N_32490);
and U35303 (N_35303,N_33859,N_33349);
and U35304 (N_35304,N_32626,N_32008);
nand U35305 (N_35305,N_32317,N_32856);
or U35306 (N_35306,N_33609,N_33517);
xnor U35307 (N_35307,N_32263,N_32608);
xnor U35308 (N_35308,N_32455,N_33732);
xnor U35309 (N_35309,N_33037,N_32125);
nor U35310 (N_35310,N_33276,N_32932);
xor U35311 (N_35311,N_33717,N_32742);
nand U35312 (N_35312,N_32594,N_33346);
and U35313 (N_35313,N_33131,N_33636);
nand U35314 (N_35314,N_33037,N_32467);
and U35315 (N_35315,N_32402,N_33313);
nor U35316 (N_35316,N_32408,N_32090);
nor U35317 (N_35317,N_32695,N_33852);
nor U35318 (N_35318,N_33601,N_33034);
xnor U35319 (N_35319,N_32319,N_32039);
or U35320 (N_35320,N_33417,N_33078);
or U35321 (N_35321,N_32050,N_32202);
and U35322 (N_35322,N_33396,N_32744);
or U35323 (N_35323,N_33904,N_32794);
or U35324 (N_35324,N_32947,N_32615);
nand U35325 (N_35325,N_33132,N_33677);
nand U35326 (N_35326,N_33420,N_33526);
nand U35327 (N_35327,N_33478,N_32716);
and U35328 (N_35328,N_33989,N_32652);
nand U35329 (N_35329,N_32228,N_33626);
and U35330 (N_35330,N_33829,N_33308);
nor U35331 (N_35331,N_32299,N_32348);
xnor U35332 (N_35332,N_32180,N_33107);
or U35333 (N_35333,N_32043,N_32051);
nor U35334 (N_35334,N_33087,N_33553);
and U35335 (N_35335,N_32691,N_32951);
nor U35336 (N_35336,N_33671,N_33747);
xor U35337 (N_35337,N_32536,N_32191);
xnor U35338 (N_35338,N_33215,N_33695);
or U35339 (N_35339,N_32750,N_33788);
nor U35340 (N_35340,N_32767,N_32259);
nand U35341 (N_35341,N_32294,N_33944);
nand U35342 (N_35342,N_32441,N_32599);
nor U35343 (N_35343,N_32004,N_32933);
nor U35344 (N_35344,N_32725,N_32194);
nand U35345 (N_35345,N_33286,N_33266);
xnor U35346 (N_35346,N_33485,N_33346);
nor U35347 (N_35347,N_32536,N_32263);
nand U35348 (N_35348,N_33842,N_32603);
xnor U35349 (N_35349,N_33817,N_33776);
and U35350 (N_35350,N_33316,N_32041);
nand U35351 (N_35351,N_33241,N_32518);
xnor U35352 (N_35352,N_33236,N_32577);
nor U35353 (N_35353,N_33716,N_33549);
nand U35354 (N_35354,N_32073,N_32707);
or U35355 (N_35355,N_32000,N_32097);
and U35356 (N_35356,N_32259,N_32806);
and U35357 (N_35357,N_33402,N_32837);
and U35358 (N_35358,N_33000,N_33588);
nand U35359 (N_35359,N_32618,N_33917);
nor U35360 (N_35360,N_33623,N_32060);
nor U35361 (N_35361,N_33246,N_32407);
xor U35362 (N_35362,N_32155,N_32086);
or U35363 (N_35363,N_33124,N_33591);
nor U35364 (N_35364,N_32001,N_32220);
and U35365 (N_35365,N_32960,N_33339);
nand U35366 (N_35366,N_32524,N_33272);
and U35367 (N_35367,N_33876,N_32755);
nor U35368 (N_35368,N_32286,N_32613);
and U35369 (N_35369,N_33004,N_32679);
xnor U35370 (N_35370,N_33810,N_32151);
nand U35371 (N_35371,N_32907,N_32633);
and U35372 (N_35372,N_32389,N_32271);
nand U35373 (N_35373,N_33782,N_33064);
and U35374 (N_35374,N_32968,N_32277);
xnor U35375 (N_35375,N_32983,N_33339);
xnor U35376 (N_35376,N_33935,N_33615);
xor U35377 (N_35377,N_32205,N_32999);
or U35378 (N_35378,N_33779,N_33513);
or U35379 (N_35379,N_32016,N_32798);
or U35380 (N_35380,N_33837,N_32768);
or U35381 (N_35381,N_33935,N_33523);
nand U35382 (N_35382,N_32144,N_33654);
nor U35383 (N_35383,N_32778,N_33426);
nand U35384 (N_35384,N_33481,N_33755);
and U35385 (N_35385,N_32109,N_33655);
nand U35386 (N_35386,N_33076,N_33831);
nand U35387 (N_35387,N_32294,N_33212);
or U35388 (N_35388,N_32340,N_33161);
xor U35389 (N_35389,N_32042,N_33680);
xnor U35390 (N_35390,N_33474,N_32018);
nor U35391 (N_35391,N_32885,N_32267);
xnor U35392 (N_35392,N_33191,N_32388);
nor U35393 (N_35393,N_32766,N_32165);
and U35394 (N_35394,N_32811,N_33410);
or U35395 (N_35395,N_32805,N_32349);
and U35396 (N_35396,N_32887,N_32368);
nand U35397 (N_35397,N_33598,N_33920);
nand U35398 (N_35398,N_32799,N_32865);
and U35399 (N_35399,N_32729,N_33827);
and U35400 (N_35400,N_32717,N_32434);
nand U35401 (N_35401,N_32076,N_33882);
nand U35402 (N_35402,N_32222,N_32515);
nand U35403 (N_35403,N_33717,N_33013);
xor U35404 (N_35404,N_33355,N_32628);
or U35405 (N_35405,N_32930,N_33914);
nand U35406 (N_35406,N_32792,N_32154);
nor U35407 (N_35407,N_32442,N_33164);
xor U35408 (N_35408,N_33470,N_33223);
and U35409 (N_35409,N_32269,N_33336);
nor U35410 (N_35410,N_32736,N_32299);
nand U35411 (N_35411,N_32975,N_33403);
xor U35412 (N_35412,N_32961,N_33337);
nor U35413 (N_35413,N_33833,N_33519);
and U35414 (N_35414,N_32631,N_32093);
and U35415 (N_35415,N_33206,N_32668);
or U35416 (N_35416,N_33504,N_33688);
or U35417 (N_35417,N_32430,N_32617);
or U35418 (N_35418,N_32246,N_33474);
nand U35419 (N_35419,N_32453,N_33823);
or U35420 (N_35420,N_33493,N_32620);
or U35421 (N_35421,N_32438,N_33313);
nor U35422 (N_35422,N_32453,N_33624);
xor U35423 (N_35423,N_32601,N_32491);
nand U35424 (N_35424,N_32654,N_33641);
nor U35425 (N_35425,N_32542,N_33755);
and U35426 (N_35426,N_33473,N_33655);
nand U35427 (N_35427,N_33964,N_32516);
and U35428 (N_35428,N_33488,N_32795);
or U35429 (N_35429,N_32920,N_33673);
nor U35430 (N_35430,N_33225,N_32656);
or U35431 (N_35431,N_33506,N_32246);
or U35432 (N_35432,N_32328,N_32535);
and U35433 (N_35433,N_32319,N_32646);
and U35434 (N_35434,N_32074,N_33928);
nand U35435 (N_35435,N_33899,N_32805);
xor U35436 (N_35436,N_32431,N_33447);
nand U35437 (N_35437,N_33884,N_33739);
and U35438 (N_35438,N_32766,N_32236);
nor U35439 (N_35439,N_32366,N_32462);
nand U35440 (N_35440,N_32026,N_33346);
xnor U35441 (N_35441,N_32686,N_33426);
or U35442 (N_35442,N_32929,N_32435);
or U35443 (N_35443,N_32201,N_33538);
xor U35444 (N_35444,N_32339,N_32404);
nor U35445 (N_35445,N_33868,N_32945);
xor U35446 (N_35446,N_32986,N_32451);
and U35447 (N_35447,N_32587,N_33060);
xnor U35448 (N_35448,N_33236,N_32535);
or U35449 (N_35449,N_32756,N_33683);
nand U35450 (N_35450,N_32720,N_32061);
nor U35451 (N_35451,N_32906,N_33935);
or U35452 (N_35452,N_33878,N_32055);
xor U35453 (N_35453,N_32017,N_33382);
or U35454 (N_35454,N_32187,N_32133);
nor U35455 (N_35455,N_33657,N_32208);
nand U35456 (N_35456,N_32978,N_33903);
xor U35457 (N_35457,N_32538,N_33110);
nand U35458 (N_35458,N_32397,N_33344);
and U35459 (N_35459,N_33468,N_32203);
nor U35460 (N_35460,N_32140,N_32008);
or U35461 (N_35461,N_32630,N_32985);
and U35462 (N_35462,N_33634,N_33118);
or U35463 (N_35463,N_32672,N_33159);
xnor U35464 (N_35464,N_32928,N_33040);
nor U35465 (N_35465,N_33093,N_33010);
and U35466 (N_35466,N_32105,N_32770);
nor U35467 (N_35467,N_33439,N_32980);
or U35468 (N_35468,N_33996,N_33924);
nor U35469 (N_35469,N_33992,N_33128);
nor U35470 (N_35470,N_32165,N_33173);
nor U35471 (N_35471,N_33052,N_33559);
nand U35472 (N_35472,N_33993,N_33606);
or U35473 (N_35473,N_32141,N_32591);
nand U35474 (N_35474,N_33056,N_32486);
nand U35475 (N_35475,N_33272,N_32957);
and U35476 (N_35476,N_32114,N_33993);
nand U35477 (N_35477,N_33036,N_33704);
xnor U35478 (N_35478,N_32294,N_32468);
nand U35479 (N_35479,N_33300,N_33164);
xnor U35480 (N_35480,N_32308,N_32115);
xor U35481 (N_35481,N_32765,N_33317);
or U35482 (N_35482,N_33509,N_33220);
nor U35483 (N_35483,N_33195,N_32832);
nand U35484 (N_35484,N_33619,N_33741);
xor U35485 (N_35485,N_32081,N_33628);
nand U35486 (N_35486,N_32321,N_32744);
nor U35487 (N_35487,N_32545,N_33237);
and U35488 (N_35488,N_33981,N_33506);
and U35489 (N_35489,N_33541,N_33391);
or U35490 (N_35490,N_32123,N_33657);
or U35491 (N_35491,N_33246,N_33820);
nor U35492 (N_35492,N_33826,N_32176);
nand U35493 (N_35493,N_33370,N_32768);
xnor U35494 (N_35494,N_33658,N_32583);
or U35495 (N_35495,N_32091,N_33832);
and U35496 (N_35496,N_33224,N_33612);
or U35497 (N_35497,N_32401,N_33145);
xnor U35498 (N_35498,N_33022,N_32431);
nand U35499 (N_35499,N_32869,N_32502);
nor U35500 (N_35500,N_33935,N_32332);
xnor U35501 (N_35501,N_33255,N_32056);
nor U35502 (N_35502,N_32827,N_32455);
nand U35503 (N_35503,N_33305,N_33827);
and U35504 (N_35504,N_33073,N_32526);
nor U35505 (N_35505,N_33184,N_33765);
nand U35506 (N_35506,N_33394,N_32628);
nor U35507 (N_35507,N_33737,N_33729);
xnor U35508 (N_35508,N_32802,N_33158);
xnor U35509 (N_35509,N_32834,N_33898);
and U35510 (N_35510,N_32511,N_33488);
nor U35511 (N_35511,N_32042,N_33253);
nand U35512 (N_35512,N_32665,N_32213);
and U35513 (N_35513,N_33115,N_32818);
nor U35514 (N_35514,N_33103,N_33234);
xnor U35515 (N_35515,N_32490,N_32124);
xnor U35516 (N_35516,N_33802,N_32307);
xor U35517 (N_35517,N_33189,N_33613);
xor U35518 (N_35518,N_33834,N_32829);
or U35519 (N_35519,N_33627,N_33666);
xnor U35520 (N_35520,N_32259,N_32454);
or U35521 (N_35521,N_32947,N_33270);
nand U35522 (N_35522,N_33016,N_32114);
xnor U35523 (N_35523,N_33588,N_32514);
xnor U35524 (N_35524,N_32412,N_32368);
xor U35525 (N_35525,N_32424,N_32997);
nor U35526 (N_35526,N_32323,N_32500);
or U35527 (N_35527,N_33510,N_33325);
nor U35528 (N_35528,N_32626,N_33559);
or U35529 (N_35529,N_32111,N_32258);
or U35530 (N_35530,N_32408,N_32570);
or U35531 (N_35531,N_33399,N_32605);
xnor U35532 (N_35532,N_33334,N_32634);
or U35533 (N_35533,N_33395,N_33074);
nor U35534 (N_35534,N_33670,N_32373);
or U35535 (N_35535,N_32091,N_33631);
nand U35536 (N_35536,N_32552,N_32529);
nand U35537 (N_35537,N_32023,N_33594);
xor U35538 (N_35538,N_33719,N_33186);
nand U35539 (N_35539,N_32726,N_33877);
xnor U35540 (N_35540,N_33374,N_32532);
xor U35541 (N_35541,N_32552,N_32912);
nor U35542 (N_35542,N_33019,N_33282);
nand U35543 (N_35543,N_32843,N_33382);
or U35544 (N_35544,N_32659,N_32102);
nand U35545 (N_35545,N_33003,N_33951);
nor U35546 (N_35546,N_32202,N_32189);
xnor U35547 (N_35547,N_33009,N_32973);
xor U35548 (N_35548,N_33502,N_32775);
or U35549 (N_35549,N_33335,N_33181);
xor U35550 (N_35550,N_33015,N_33006);
and U35551 (N_35551,N_33218,N_32662);
or U35552 (N_35552,N_32650,N_33221);
or U35553 (N_35553,N_33655,N_32641);
nor U35554 (N_35554,N_32136,N_33088);
nand U35555 (N_35555,N_33503,N_32701);
nand U35556 (N_35556,N_32779,N_32412);
nor U35557 (N_35557,N_33299,N_33115);
nand U35558 (N_35558,N_32890,N_32503);
nor U35559 (N_35559,N_32960,N_33580);
and U35560 (N_35560,N_32939,N_32735);
nand U35561 (N_35561,N_32126,N_33336);
nand U35562 (N_35562,N_32805,N_32373);
nand U35563 (N_35563,N_32953,N_32119);
nor U35564 (N_35564,N_33594,N_32722);
and U35565 (N_35565,N_32477,N_32302);
nand U35566 (N_35566,N_32444,N_33486);
nor U35567 (N_35567,N_32965,N_32603);
and U35568 (N_35568,N_32341,N_33198);
xor U35569 (N_35569,N_32365,N_32458);
nand U35570 (N_35570,N_33860,N_33742);
nand U35571 (N_35571,N_33778,N_33195);
and U35572 (N_35572,N_32966,N_32386);
xor U35573 (N_35573,N_32293,N_33462);
xnor U35574 (N_35574,N_33865,N_33641);
nand U35575 (N_35575,N_33706,N_32662);
or U35576 (N_35576,N_33041,N_32615);
xor U35577 (N_35577,N_33946,N_33404);
or U35578 (N_35578,N_32925,N_33230);
xnor U35579 (N_35579,N_32489,N_32701);
nor U35580 (N_35580,N_33655,N_33793);
nand U35581 (N_35581,N_32364,N_33203);
and U35582 (N_35582,N_32849,N_32221);
nand U35583 (N_35583,N_32123,N_32958);
xnor U35584 (N_35584,N_32315,N_32601);
nand U35585 (N_35585,N_33569,N_33587);
or U35586 (N_35586,N_32397,N_33202);
nor U35587 (N_35587,N_32936,N_33958);
or U35588 (N_35588,N_33930,N_33816);
nor U35589 (N_35589,N_33235,N_32691);
nand U35590 (N_35590,N_32682,N_33342);
nor U35591 (N_35591,N_33257,N_32626);
and U35592 (N_35592,N_33270,N_32136);
or U35593 (N_35593,N_33711,N_33463);
or U35594 (N_35594,N_33490,N_32652);
or U35595 (N_35595,N_32601,N_32084);
nor U35596 (N_35596,N_32039,N_32995);
nor U35597 (N_35597,N_32620,N_33488);
nor U35598 (N_35598,N_33506,N_32990);
and U35599 (N_35599,N_33956,N_32041);
xnor U35600 (N_35600,N_32656,N_32139);
or U35601 (N_35601,N_33273,N_33035);
nor U35602 (N_35602,N_33845,N_33610);
nand U35603 (N_35603,N_32081,N_32045);
nor U35604 (N_35604,N_32126,N_32282);
or U35605 (N_35605,N_33484,N_32945);
xnor U35606 (N_35606,N_33810,N_33947);
nand U35607 (N_35607,N_33408,N_32068);
nor U35608 (N_35608,N_32056,N_33007);
xnor U35609 (N_35609,N_33739,N_33953);
nor U35610 (N_35610,N_33013,N_33980);
nand U35611 (N_35611,N_32031,N_32004);
nand U35612 (N_35612,N_32398,N_33662);
nand U35613 (N_35613,N_33354,N_33835);
nand U35614 (N_35614,N_32055,N_32928);
and U35615 (N_35615,N_33063,N_32502);
and U35616 (N_35616,N_33435,N_32457);
nor U35617 (N_35617,N_32631,N_33054);
or U35618 (N_35618,N_32664,N_32216);
xnor U35619 (N_35619,N_33173,N_33986);
nor U35620 (N_35620,N_33772,N_33587);
nand U35621 (N_35621,N_33153,N_33166);
and U35622 (N_35622,N_32242,N_33912);
and U35623 (N_35623,N_32317,N_33639);
and U35624 (N_35624,N_32841,N_32642);
and U35625 (N_35625,N_32787,N_33356);
xor U35626 (N_35626,N_33196,N_32226);
and U35627 (N_35627,N_33603,N_33841);
xor U35628 (N_35628,N_33360,N_33426);
nor U35629 (N_35629,N_32266,N_33169);
nor U35630 (N_35630,N_33287,N_33277);
and U35631 (N_35631,N_33030,N_32455);
xor U35632 (N_35632,N_33129,N_33358);
nand U35633 (N_35633,N_32388,N_32385);
nor U35634 (N_35634,N_32230,N_32629);
xor U35635 (N_35635,N_32528,N_33601);
and U35636 (N_35636,N_32817,N_32660);
and U35637 (N_35637,N_33231,N_33567);
or U35638 (N_35638,N_33620,N_33819);
nand U35639 (N_35639,N_33769,N_33718);
nor U35640 (N_35640,N_33476,N_33345);
nor U35641 (N_35641,N_32969,N_32036);
nor U35642 (N_35642,N_33733,N_32828);
or U35643 (N_35643,N_32711,N_32854);
xor U35644 (N_35644,N_32130,N_33875);
xnor U35645 (N_35645,N_33906,N_33819);
nor U35646 (N_35646,N_32741,N_32236);
nor U35647 (N_35647,N_32680,N_33803);
nand U35648 (N_35648,N_33844,N_32266);
or U35649 (N_35649,N_33018,N_33144);
nand U35650 (N_35650,N_33260,N_32636);
nand U35651 (N_35651,N_33049,N_33370);
xnor U35652 (N_35652,N_33336,N_32084);
nand U35653 (N_35653,N_32724,N_32836);
xor U35654 (N_35654,N_32251,N_33931);
and U35655 (N_35655,N_33009,N_32332);
or U35656 (N_35656,N_33104,N_33949);
nor U35657 (N_35657,N_32199,N_33785);
or U35658 (N_35658,N_32918,N_33727);
or U35659 (N_35659,N_32798,N_32573);
or U35660 (N_35660,N_33432,N_33823);
or U35661 (N_35661,N_33302,N_32362);
or U35662 (N_35662,N_33817,N_32834);
nor U35663 (N_35663,N_32547,N_33369);
or U35664 (N_35664,N_33173,N_33978);
xor U35665 (N_35665,N_33124,N_33755);
nor U35666 (N_35666,N_32632,N_32000);
xnor U35667 (N_35667,N_32040,N_32299);
and U35668 (N_35668,N_33074,N_33143);
xor U35669 (N_35669,N_33513,N_32945);
or U35670 (N_35670,N_33507,N_33795);
and U35671 (N_35671,N_33638,N_32284);
nand U35672 (N_35672,N_33036,N_33579);
nor U35673 (N_35673,N_33962,N_32953);
nand U35674 (N_35674,N_33169,N_32137);
or U35675 (N_35675,N_32936,N_33272);
or U35676 (N_35676,N_33832,N_33872);
nor U35677 (N_35677,N_32058,N_33999);
nand U35678 (N_35678,N_32934,N_32675);
nor U35679 (N_35679,N_33969,N_32610);
nor U35680 (N_35680,N_32699,N_32377);
or U35681 (N_35681,N_32351,N_32541);
or U35682 (N_35682,N_33698,N_33165);
or U35683 (N_35683,N_33464,N_32280);
and U35684 (N_35684,N_32783,N_33421);
nand U35685 (N_35685,N_32725,N_33080);
xor U35686 (N_35686,N_32274,N_32603);
or U35687 (N_35687,N_32515,N_33224);
and U35688 (N_35688,N_33166,N_33600);
and U35689 (N_35689,N_33931,N_32753);
nand U35690 (N_35690,N_32592,N_32951);
xor U35691 (N_35691,N_32071,N_33922);
xor U35692 (N_35692,N_32274,N_33853);
and U35693 (N_35693,N_33979,N_33225);
or U35694 (N_35694,N_32646,N_32743);
nand U35695 (N_35695,N_32332,N_32224);
or U35696 (N_35696,N_32445,N_33644);
xnor U35697 (N_35697,N_33374,N_32575);
or U35698 (N_35698,N_32159,N_32101);
xnor U35699 (N_35699,N_32382,N_33561);
nor U35700 (N_35700,N_32332,N_32862);
xnor U35701 (N_35701,N_32653,N_33816);
xor U35702 (N_35702,N_33525,N_32323);
nor U35703 (N_35703,N_32600,N_32881);
nand U35704 (N_35704,N_32641,N_33238);
and U35705 (N_35705,N_33230,N_32942);
xnor U35706 (N_35706,N_32139,N_32354);
nor U35707 (N_35707,N_32010,N_32953);
and U35708 (N_35708,N_33992,N_33848);
or U35709 (N_35709,N_33521,N_32136);
nor U35710 (N_35710,N_33163,N_32285);
xnor U35711 (N_35711,N_32734,N_33949);
nand U35712 (N_35712,N_32794,N_33798);
nand U35713 (N_35713,N_32375,N_33034);
nand U35714 (N_35714,N_33962,N_32776);
nor U35715 (N_35715,N_32740,N_33933);
and U35716 (N_35716,N_32899,N_33961);
xor U35717 (N_35717,N_33515,N_33067);
xnor U35718 (N_35718,N_33358,N_33244);
and U35719 (N_35719,N_32514,N_32449);
and U35720 (N_35720,N_32419,N_32134);
or U35721 (N_35721,N_33923,N_33710);
nor U35722 (N_35722,N_33952,N_33336);
and U35723 (N_35723,N_33157,N_32248);
xnor U35724 (N_35724,N_32025,N_33358);
xor U35725 (N_35725,N_32236,N_33410);
nor U35726 (N_35726,N_33928,N_33884);
or U35727 (N_35727,N_33776,N_32044);
nor U35728 (N_35728,N_33370,N_32128);
nor U35729 (N_35729,N_33183,N_32528);
or U35730 (N_35730,N_33035,N_33482);
or U35731 (N_35731,N_32204,N_32203);
xor U35732 (N_35732,N_32372,N_32661);
nand U35733 (N_35733,N_32159,N_33441);
and U35734 (N_35734,N_33270,N_32182);
and U35735 (N_35735,N_33638,N_32341);
and U35736 (N_35736,N_32590,N_33579);
nand U35737 (N_35737,N_33189,N_32821);
or U35738 (N_35738,N_33262,N_33773);
and U35739 (N_35739,N_32900,N_32625);
nand U35740 (N_35740,N_32541,N_32189);
or U35741 (N_35741,N_33188,N_33614);
and U35742 (N_35742,N_33603,N_32549);
xnor U35743 (N_35743,N_32594,N_33873);
or U35744 (N_35744,N_32049,N_33193);
and U35745 (N_35745,N_33052,N_33127);
nor U35746 (N_35746,N_32671,N_32805);
or U35747 (N_35747,N_33744,N_32042);
nand U35748 (N_35748,N_32456,N_32511);
nor U35749 (N_35749,N_33015,N_33433);
and U35750 (N_35750,N_32506,N_32383);
nor U35751 (N_35751,N_33478,N_32925);
or U35752 (N_35752,N_33094,N_33024);
xnor U35753 (N_35753,N_32720,N_32233);
nand U35754 (N_35754,N_33735,N_32779);
or U35755 (N_35755,N_33386,N_32340);
xor U35756 (N_35756,N_33122,N_32450);
or U35757 (N_35757,N_32526,N_32316);
nor U35758 (N_35758,N_32872,N_33631);
and U35759 (N_35759,N_32797,N_33888);
and U35760 (N_35760,N_33229,N_33901);
xor U35761 (N_35761,N_33459,N_33805);
xor U35762 (N_35762,N_33804,N_33136);
or U35763 (N_35763,N_32355,N_33248);
or U35764 (N_35764,N_32924,N_32099);
xor U35765 (N_35765,N_32851,N_32982);
nor U35766 (N_35766,N_33010,N_33942);
nor U35767 (N_35767,N_32161,N_32791);
nor U35768 (N_35768,N_33652,N_32202);
and U35769 (N_35769,N_32651,N_33598);
and U35770 (N_35770,N_33501,N_32001);
or U35771 (N_35771,N_32176,N_32070);
nand U35772 (N_35772,N_32781,N_33807);
and U35773 (N_35773,N_33697,N_33906);
or U35774 (N_35774,N_32922,N_33355);
nand U35775 (N_35775,N_32505,N_33282);
xnor U35776 (N_35776,N_33428,N_32272);
and U35777 (N_35777,N_32448,N_33212);
nor U35778 (N_35778,N_33853,N_32785);
xor U35779 (N_35779,N_33729,N_32212);
xnor U35780 (N_35780,N_33260,N_33259);
or U35781 (N_35781,N_32277,N_33887);
or U35782 (N_35782,N_32522,N_32840);
and U35783 (N_35783,N_32784,N_33677);
xnor U35784 (N_35784,N_32963,N_32795);
nor U35785 (N_35785,N_33479,N_33652);
nor U35786 (N_35786,N_33105,N_32809);
nor U35787 (N_35787,N_33325,N_33020);
xor U35788 (N_35788,N_33184,N_32564);
nor U35789 (N_35789,N_33704,N_33098);
xor U35790 (N_35790,N_32263,N_33804);
or U35791 (N_35791,N_32833,N_33798);
or U35792 (N_35792,N_33848,N_32999);
xnor U35793 (N_35793,N_33293,N_33993);
nand U35794 (N_35794,N_33516,N_33451);
xor U35795 (N_35795,N_32134,N_32922);
nor U35796 (N_35796,N_33900,N_32735);
and U35797 (N_35797,N_33573,N_33022);
xor U35798 (N_35798,N_32581,N_32315);
or U35799 (N_35799,N_32587,N_33403);
or U35800 (N_35800,N_33842,N_33918);
and U35801 (N_35801,N_32272,N_33725);
nor U35802 (N_35802,N_32091,N_32303);
and U35803 (N_35803,N_32281,N_32173);
nand U35804 (N_35804,N_33411,N_32584);
nor U35805 (N_35805,N_33504,N_32350);
and U35806 (N_35806,N_33365,N_32889);
or U35807 (N_35807,N_32503,N_33264);
or U35808 (N_35808,N_32077,N_32766);
xnor U35809 (N_35809,N_32534,N_33187);
and U35810 (N_35810,N_33415,N_32435);
or U35811 (N_35811,N_33116,N_33399);
nor U35812 (N_35812,N_33987,N_32162);
nand U35813 (N_35813,N_32610,N_33630);
xnor U35814 (N_35814,N_33184,N_32536);
nand U35815 (N_35815,N_32130,N_33772);
or U35816 (N_35816,N_33945,N_32257);
and U35817 (N_35817,N_33875,N_33766);
nor U35818 (N_35818,N_33371,N_33957);
nand U35819 (N_35819,N_32683,N_33335);
nand U35820 (N_35820,N_33287,N_33936);
nor U35821 (N_35821,N_32011,N_32502);
or U35822 (N_35822,N_32455,N_32268);
xor U35823 (N_35823,N_32971,N_32346);
xnor U35824 (N_35824,N_33787,N_32916);
and U35825 (N_35825,N_33429,N_32453);
or U35826 (N_35826,N_32713,N_33041);
or U35827 (N_35827,N_33179,N_32557);
nor U35828 (N_35828,N_32006,N_33815);
or U35829 (N_35829,N_33025,N_33356);
xnor U35830 (N_35830,N_33295,N_32688);
xnor U35831 (N_35831,N_32996,N_33441);
nand U35832 (N_35832,N_33869,N_32916);
nand U35833 (N_35833,N_33827,N_32687);
nand U35834 (N_35834,N_33817,N_32412);
and U35835 (N_35835,N_33730,N_33330);
and U35836 (N_35836,N_33414,N_32790);
nand U35837 (N_35837,N_33952,N_32044);
nand U35838 (N_35838,N_32185,N_32248);
nor U35839 (N_35839,N_32196,N_33799);
and U35840 (N_35840,N_33067,N_33637);
xnor U35841 (N_35841,N_33410,N_32798);
or U35842 (N_35842,N_32012,N_32716);
xor U35843 (N_35843,N_33219,N_32031);
xnor U35844 (N_35844,N_33117,N_32807);
and U35845 (N_35845,N_33768,N_33138);
and U35846 (N_35846,N_32105,N_33263);
and U35847 (N_35847,N_33917,N_32353);
xnor U35848 (N_35848,N_32776,N_33379);
or U35849 (N_35849,N_33739,N_33429);
xor U35850 (N_35850,N_32872,N_32803);
xnor U35851 (N_35851,N_33189,N_32918);
and U35852 (N_35852,N_33464,N_32702);
or U35853 (N_35853,N_32746,N_32520);
xor U35854 (N_35854,N_33316,N_32083);
and U35855 (N_35855,N_32178,N_32503);
or U35856 (N_35856,N_32085,N_33162);
or U35857 (N_35857,N_32239,N_33126);
and U35858 (N_35858,N_32982,N_33281);
nor U35859 (N_35859,N_33706,N_32486);
and U35860 (N_35860,N_32838,N_32057);
xnor U35861 (N_35861,N_33885,N_32977);
nor U35862 (N_35862,N_33082,N_32525);
or U35863 (N_35863,N_33759,N_33532);
or U35864 (N_35864,N_32423,N_32401);
nor U35865 (N_35865,N_33766,N_32452);
and U35866 (N_35866,N_33586,N_32958);
nor U35867 (N_35867,N_33443,N_32349);
nand U35868 (N_35868,N_33809,N_32779);
nand U35869 (N_35869,N_33391,N_33241);
or U35870 (N_35870,N_32766,N_33823);
and U35871 (N_35871,N_33937,N_32680);
nor U35872 (N_35872,N_32521,N_32919);
nor U35873 (N_35873,N_33037,N_33679);
and U35874 (N_35874,N_32614,N_32900);
or U35875 (N_35875,N_32214,N_33473);
nor U35876 (N_35876,N_32215,N_33300);
xnor U35877 (N_35877,N_33341,N_32558);
nor U35878 (N_35878,N_33842,N_33678);
nand U35879 (N_35879,N_32624,N_32838);
or U35880 (N_35880,N_32664,N_33711);
nand U35881 (N_35881,N_33518,N_33656);
and U35882 (N_35882,N_33570,N_33886);
and U35883 (N_35883,N_32375,N_32399);
and U35884 (N_35884,N_33087,N_32073);
and U35885 (N_35885,N_32223,N_33580);
xnor U35886 (N_35886,N_32640,N_32845);
xnor U35887 (N_35887,N_33067,N_33498);
xor U35888 (N_35888,N_32455,N_32198);
and U35889 (N_35889,N_32479,N_33074);
and U35890 (N_35890,N_33225,N_32294);
and U35891 (N_35891,N_32660,N_32664);
nor U35892 (N_35892,N_33733,N_32662);
or U35893 (N_35893,N_33545,N_32974);
xnor U35894 (N_35894,N_33030,N_33569);
and U35895 (N_35895,N_32742,N_32858);
xor U35896 (N_35896,N_33753,N_33965);
and U35897 (N_35897,N_33732,N_32640);
nor U35898 (N_35898,N_32691,N_32064);
xor U35899 (N_35899,N_32151,N_33059);
nor U35900 (N_35900,N_32865,N_32784);
xnor U35901 (N_35901,N_33482,N_32200);
and U35902 (N_35902,N_33992,N_33647);
nand U35903 (N_35903,N_33222,N_33905);
nand U35904 (N_35904,N_33834,N_33357);
nand U35905 (N_35905,N_32114,N_32203);
or U35906 (N_35906,N_33686,N_32023);
nor U35907 (N_35907,N_33989,N_32006);
and U35908 (N_35908,N_33094,N_33756);
or U35909 (N_35909,N_32480,N_32759);
and U35910 (N_35910,N_33172,N_32073);
nor U35911 (N_35911,N_33125,N_33861);
nor U35912 (N_35912,N_32562,N_32045);
xnor U35913 (N_35913,N_33157,N_33986);
nor U35914 (N_35914,N_32962,N_33958);
or U35915 (N_35915,N_32853,N_32572);
and U35916 (N_35916,N_33603,N_32757);
nand U35917 (N_35917,N_33850,N_32349);
xor U35918 (N_35918,N_32558,N_32721);
or U35919 (N_35919,N_32496,N_32566);
or U35920 (N_35920,N_32938,N_33764);
nor U35921 (N_35921,N_33554,N_32292);
and U35922 (N_35922,N_32371,N_33588);
or U35923 (N_35923,N_33128,N_33304);
nand U35924 (N_35924,N_33431,N_33084);
and U35925 (N_35925,N_33939,N_32592);
nand U35926 (N_35926,N_33829,N_32553);
xor U35927 (N_35927,N_33708,N_33526);
or U35928 (N_35928,N_32911,N_32584);
and U35929 (N_35929,N_33050,N_33887);
nor U35930 (N_35930,N_33117,N_33342);
and U35931 (N_35931,N_32544,N_32368);
nor U35932 (N_35932,N_33338,N_33128);
xnor U35933 (N_35933,N_33733,N_33161);
or U35934 (N_35934,N_33820,N_32132);
or U35935 (N_35935,N_33782,N_33423);
and U35936 (N_35936,N_33726,N_33557);
and U35937 (N_35937,N_32601,N_33829);
xnor U35938 (N_35938,N_33218,N_32325);
nand U35939 (N_35939,N_33399,N_33286);
and U35940 (N_35940,N_32082,N_32984);
nor U35941 (N_35941,N_32367,N_32402);
nand U35942 (N_35942,N_32193,N_33098);
or U35943 (N_35943,N_32129,N_32352);
nor U35944 (N_35944,N_33945,N_33428);
xnor U35945 (N_35945,N_32262,N_32342);
nor U35946 (N_35946,N_33703,N_32074);
or U35947 (N_35947,N_33284,N_33618);
or U35948 (N_35948,N_33348,N_32948);
and U35949 (N_35949,N_32174,N_33264);
and U35950 (N_35950,N_33314,N_33622);
and U35951 (N_35951,N_33783,N_32666);
xor U35952 (N_35952,N_33070,N_32957);
xor U35953 (N_35953,N_32494,N_32567);
nor U35954 (N_35954,N_32059,N_32357);
or U35955 (N_35955,N_32247,N_32081);
nor U35956 (N_35956,N_32726,N_33642);
xnor U35957 (N_35957,N_33016,N_32199);
and U35958 (N_35958,N_33001,N_33296);
or U35959 (N_35959,N_33073,N_32140);
or U35960 (N_35960,N_32991,N_33445);
xnor U35961 (N_35961,N_32380,N_32184);
or U35962 (N_35962,N_33794,N_32638);
nor U35963 (N_35963,N_33620,N_32225);
or U35964 (N_35964,N_33942,N_32147);
and U35965 (N_35965,N_32734,N_33508);
xor U35966 (N_35966,N_33159,N_32361);
and U35967 (N_35967,N_33408,N_32259);
or U35968 (N_35968,N_32415,N_33661);
or U35969 (N_35969,N_33323,N_32626);
nand U35970 (N_35970,N_32494,N_32632);
nor U35971 (N_35971,N_32886,N_33711);
or U35972 (N_35972,N_33007,N_32206);
or U35973 (N_35973,N_32419,N_32991);
nor U35974 (N_35974,N_33382,N_32309);
xor U35975 (N_35975,N_33798,N_33548);
nand U35976 (N_35976,N_32564,N_33835);
and U35977 (N_35977,N_32067,N_33150);
xor U35978 (N_35978,N_33116,N_32705);
xnor U35979 (N_35979,N_33004,N_32116);
nand U35980 (N_35980,N_32634,N_33393);
xor U35981 (N_35981,N_33138,N_32195);
nand U35982 (N_35982,N_33779,N_32027);
xnor U35983 (N_35983,N_32980,N_32797);
or U35984 (N_35984,N_32087,N_32909);
nand U35985 (N_35985,N_33492,N_32936);
nor U35986 (N_35986,N_32369,N_33857);
xnor U35987 (N_35987,N_32214,N_32134);
nor U35988 (N_35988,N_32672,N_32328);
nand U35989 (N_35989,N_32622,N_33215);
nand U35990 (N_35990,N_33862,N_33538);
or U35991 (N_35991,N_33484,N_32900);
or U35992 (N_35992,N_33037,N_33116);
nand U35993 (N_35993,N_33071,N_33418);
or U35994 (N_35994,N_32133,N_33154);
and U35995 (N_35995,N_32156,N_33171);
nor U35996 (N_35996,N_33106,N_33038);
xnor U35997 (N_35997,N_33894,N_32558);
nand U35998 (N_35998,N_32862,N_33274);
or U35999 (N_35999,N_32274,N_33331);
or U36000 (N_36000,N_35387,N_34894);
xor U36001 (N_36001,N_34843,N_35527);
nor U36002 (N_36002,N_34483,N_34424);
or U36003 (N_36003,N_34592,N_35436);
nand U36004 (N_36004,N_34718,N_34697);
or U36005 (N_36005,N_34480,N_34759);
and U36006 (N_36006,N_35694,N_35965);
xnor U36007 (N_36007,N_34425,N_34521);
or U36008 (N_36008,N_35792,N_35117);
xnor U36009 (N_36009,N_34048,N_35307);
and U36010 (N_36010,N_35973,N_34498);
or U36011 (N_36011,N_34310,N_34403);
nand U36012 (N_36012,N_34947,N_35464);
xnor U36013 (N_36013,N_34998,N_35507);
nand U36014 (N_36014,N_34524,N_34172);
or U36015 (N_36015,N_34383,N_35429);
xor U36016 (N_36016,N_34852,N_34451);
nand U36017 (N_36017,N_35584,N_35373);
or U36018 (N_36018,N_35636,N_35946);
and U36019 (N_36019,N_34262,N_35615);
nand U36020 (N_36020,N_34788,N_34247);
nor U36021 (N_36021,N_34157,N_34146);
nand U36022 (N_36022,N_34201,N_35342);
xor U36023 (N_36023,N_34740,N_35693);
or U36024 (N_36024,N_34409,N_34064);
nand U36025 (N_36025,N_34095,N_35617);
nand U36026 (N_36026,N_35660,N_35348);
nor U36027 (N_36027,N_35828,N_34765);
or U36028 (N_36028,N_34362,N_34946);
nor U36029 (N_36029,N_35169,N_34537);
nand U36030 (N_36030,N_34151,N_34804);
nand U36031 (N_36031,N_35673,N_34630);
or U36032 (N_36032,N_35824,N_34319);
nor U36033 (N_36033,N_34924,N_34639);
nor U36034 (N_36034,N_35729,N_34550);
xor U36035 (N_36035,N_34527,N_34265);
nor U36036 (N_36036,N_35960,N_34976);
nor U36037 (N_36037,N_35504,N_34066);
nor U36038 (N_36038,N_34100,N_34254);
and U36039 (N_36039,N_35780,N_34823);
nor U36040 (N_36040,N_34887,N_34563);
nor U36041 (N_36041,N_35880,N_35081);
and U36042 (N_36042,N_35772,N_34034);
and U36043 (N_36043,N_35893,N_34241);
xnor U36044 (N_36044,N_34667,N_35460);
or U36045 (N_36045,N_35874,N_34210);
xnor U36046 (N_36046,N_35392,N_35417);
or U36047 (N_36047,N_35346,N_35817);
and U36048 (N_36048,N_34054,N_35931);
and U36049 (N_36049,N_34567,N_35606);
or U36050 (N_36050,N_34845,N_34952);
nor U36051 (N_36051,N_34678,N_35740);
nand U36052 (N_36052,N_35732,N_35811);
xor U36053 (N_36053,N_35399,N_35895);
xnor U36054 (N_36054,N_34077,N_35843);
nand U36055 (N_36055,N_35754,N_34159);
or U36056 (N_36056,N_35784,N_35067);
and U36057 (N_36057,N_35790,N_34906);
nand U36058 (N_36058,N_34990,N_34553);
and U36059 (N_36059,N_35009,N_34123);
xnor U36060 (N_36060,N_35863,N_34420);
nand U36061 (N_36061,N_34945,N_34781);
and U36062 (N_36062,N_34074,N_34986);
xor U36063 (N_36063,N_35188,N_34437);
nand U36064 (N_36064,N_35333,N_34369);
nor U36065 (N_36065,N_34596,N_35461);
xnor U36066 (N_36066,N_34520,N_34880);
and U36067 (N_36067,N_34087,N_34791);
nor U36068 (N_36068,N_34711,N_35583);
xnor U36069 (N_36069,N_34436,N_35289);
nor U36070 (N_36070,N_34354,N_35968);
and U36071 (N_36071,N_34111,N_34811);
nor U36072 (N_36072,N_35275,N_35034);
xor U36073 (N_36073,N_34875,N_34899);
nand U36074 (N_36074,N_34005,N_35291);
xor U36075 (N_36075,N_34604,N_35924);
xnor U36076 (N_36076,N_35761,N_35263);
or U36077 (N_36077,N_35126,N_35697);
nand U36078 (N_36078,N_34488,N_34370);
nor U36079 (N_36079,N_34477,N_35538);
nor U36080 (N_36080,N_34091,N_34031);
xor U36081 (N_36081,N_34421,N_35325);
and U36082 (N_36082,N_34876,N_35410);
and U36083 (N_36083,N_35783,N_34546);
xor U36084 (N_36084,N_35500,N_34251);
or U36085 (N_36085,N_34794,N_35975);
xor U36086 (N_36086,N_34399,N_35032);
nor U36087 (N_36087,N_35757,N_34522);
nor U36088 (N_36088,N_35119,N_35727);
nor U36089 (N_36089,N_35554,N_34979);
and U36090 (N_36090,N_34859,N_34284);
nor U36091 (N_36091,N_34106,N_35206);
or U36092 (N_36092,N_34191,N_35198);
nor U36093 (N_36093,N_35233,N_35349);
or U36094 (N_36094,N_34766,N_34486);
or U36095 (N_36095,N_35962,N_34177);
and U36096 (N_36096,N_34108,N_34808);
nand U36097 (N_36097,N_34942,N_34590);
or U36098 (N_36098,N_35245,N_34043);
nand U36099 (N_36099,N_34891,N_35526);
nand U36100 (N_36100,N_34663,N_35593);
nor U36101 (N_36101,N_34067,N_35108);
xor U36102 (N_36102,N_35222,N_34308);
nor U36103 (N_36103,N_34168,N_35803);
nor U36104 (N_36104,N_35015,N_35278);
and U36105 (N_36105,N_34250,N_35488);
nand U36106 (N_36106,N_35293,N_35330);
xor U36107 (N_36107,N_35087,N_34286);
and U36108 (N_36108,N_35686,N_34839);
xnor U36109 (N_36109,N_35829,N_35378);
nand U36110 (N_36110,N_35989,N_34120);
nand U36111 (N_36111,N_34659,N_34838);
and U36112 (N_36112,N_34400,N_35313);
and U36113 (N_36113,N_34615,N_34001);
xor U36114 (N_36114,N_34216,N_35539);
xor U36115 (N_36115,N_34778,N_35592);
and U36116 (N_36116,N_35101,N_34490);
nor U36117 (N_36117,N_34675,N_34164);
nand U36118 (N_36118,N_35231,N_35655);
and U36119 (N_36119,N_34497,N_35285);
nor U36120 (N_36120,N_35100,N_35114);
nor U36121 (N_36121,N_34570,N_35869);
nor U36122 (N_36122,N_34294,N_34019);
nor U36123 (N_36123,N_34135,N_35282);
nor U36124 (N_36124,N_35215,N_35633);
xor U36125 (N_36125,N_34082,N_35243);
nand U36126 (N_36126,N_34229,N_34605);
xnor U36127 (N_36127,N_35659,N_35745);
nor U36128 (N_36128,N_34652,N_35758);
or U36129 (N_36129,N_34050,N_35048);
nor U36130 (N_36130,N_34381,N_34461);
and U36131 (N_36131,N_35070,N_35557);
nand U36132 (N_36132,N_35455,N_34260);
nor U36133 (N_36133,N_34471,N_35176);
xnor U36134 (N_36134,N_34897,N_34637);
or U36135 (N_36135,N_34846,N_34674);
or U36136 (N_36136,N_35078,N_34346);
and U36137 (N_36137,N_34474,N_35497);
and U36138 (N_36138,N_34878,N_35855);
nor U36139 (N_36139,N_34328,N_35988);
nand U36140 (N_36140,N_35679,N_35845);
xnor U36141 (N_36141,N_34453,N_35244);
or U36142 (N_36142,N_34641,N_35457);
nand U36143 (N_36143,N_34693,N_34844);
xor U36144 (N_36144,N_35148,N_35897);
or U36145 (N_36145,N_35248,N_34248);
nand U36146 (N_36146,N_35751,N_34864);
nor U36147 (N_36147,N_35207,N_34809);
nand U36148 (N_36148,N_35260,N_34447);
xor U36149 (N_36149,N_35859,N_34355);
nor U36150 (N_36150,N_35726,N_34654);
and U36151 (N_36151,N_34452,N_35854);
or U36152 (N_36152,N_34938,N_34326);
and U36153 (N_36153,N_35664,N_35876);
or U36154 (N_36154,N_35273,N_34917);
nor U36155 (N_36155,N_35145,N_35456);
nand U36156 (N_36156,N_34016,N_35232);
xor U36157 (N_36157,N_34589,N_35577);
nor U36158 (N_36158,N_34819,N_34686);
xor U36159 (N_36159,N_35900,N_34830);
or U36160 (N_36160,N_34866,N_35086);
or U36161 (N_36161,N_35840,N_35923);
and U36162 (N_36162,N_35107,N_35193);
nor U36163 (N_36163,N_34463,N_35681);
xor U36164 (N_36164,N_35423,N_35251);
xnor U36165 (N_36165,N_34613,N_35629);
nor U36166 (N_36166,N_34330,N_34515);
or U36167 (N_36167,N_34874,N_35130);
and U36168 (N_36168,N_35985,N_35481);
and U36169 (N_36169,N_34148,N_35560);
xnor U36170 (N_36170,N_34705,N_34462);
xnor U36171 (N_36171,N_35031,N_35297);
nand U36172 (N_36172,N_34372,N_34669);
or U36173 (N_36173,N_35856,N_35344);
and U36174 (N_36174,N_34642,N_35521);
or U36175 (N_36175,N_35350,N_35345);
or U36176 (N_36176,N_35091,N_35061);
nand U36177 (N_36177,N_34293,N_35391);
and U36178 (N_36178,N_34199,N_35074);
nor U36179 (N_36179,N_35190,N_35068);
and U36180 (N_36180,N_34134,N_34015);
nand U36181 (N_36181,N_34418,N_35274);
nor U36182 (N_36182,N_35029,N_35258);
and U36183 (N_36183,N_34953,N_35548);
nand U36184 (N_36184,N_35259,N_34353);
or U36185 (N_36185,N_35738,N_34239);
nand U36186 (N_36186,N_35640,N_34832);
xnor U36187 (N_36187,N_34854,N_35885);
xnor U36188 (N_36188,N_34679,N_35062);
and U36189 (N_36189,N_35478,N_35842);
and U36190 (N_36190,N_35065,N_34777);
or U36191 (N_36191,N_35421,N_34349);
nor U36192 (N_36192,N_34607,N_35006);
or U36193 (N_36193,N_34454,N_34824);
or U36194 (N_36194,N_35050,N_35037);
and U36195 (N_36195,N_35873,N_34132);
nor U36196 (N_36196,N_34716,N_34411);
and U36197 (N_36197,N_35921,N_34807);
nand U36198 (N_36198,N_35105,N_35503);
or U36199 (N_36199,N_35103,N_34367);
nor U36200 (N_36200,N_35237,N_35762);
nand U36201 (N_36201,N_34368,N_34390);
or U36202 (N_36202,N_35935,N_34784);
and U36203 (N_36203,N_35256,N_34303);
or U36204 (N_36204,N_35699,N_34534);
nor U36205 (N_36205,N_35737,N_35360);
nor U36206 (N_36206,N_35279,N_35904);
nor U36207 (N_36207,N_35280,N_34526);
and U36208 (N_36208,N_34803,N_34327);
nor U36209 (N_36209,N_34181,N_34103);
nor U36210 (N_36210,N_34581,N_35292);
nand U36211 (N_36211,N_35127,N_34512);
nand U36212 (N_36212,N_34198,N_35498);
and U36213 (N_36213,N_35864,N_35013);
and U36214 (N_36214,N_35098,N_35099);
nor U36215 (N_36215,N_35561,N_34158);
nor U36216 (N_36216,N_34047,N_34283);
nor U36217 (N_36217,N_34279,N_35230);
xnor U36218 (N_36218,N_35299,N_35505);
xor U36219 (N_36219,N_34636,N_34309);
nand U36220 (N_36220,N_34222,N_35118);
xnor U36221 (N_36221,N_35357,N_35083);
nand U36222 (N_36222,N_34538,N_34936);
nand U36223 (N_36223,N_34528,N_35324);
and U36224 (N_36224,N_35994,N_35340);
nor U36225 (N_36225,N_34207,N_34772);
nand U36226 (N_36226,N_35722,N_34729);
xor U36227 (N_36227,N_34566,N_35702);
or U36228 (N_36228,N_34053,N_34183);
nand U36229 (N_36229,N_34236,N_35550);
nand U36230 (N_36230,N_34982,N_35690);
or U36231 (N_36231,N_34767,N_35588);
and U36232 (N_36232,N_35058,N_34227);
xor U36233 (N_36233,N_35518,N_35677);
or U36234 (N_36234,N_35156,N_35007);
nand U36235 (N_36235,N_34045,N_34506);
xor U36236 (N_36236,N_35508,N_34336);
nor U36237 (N_36237,N_34495,N_34140);
nand U36238 (N_36238,N_34881,N_34127);
and U36239 (N_36239,N_35747,N_34391);
and U36240 (N_36240,N_35870,N_34935);
nor U36241 (N_36241,N_34836,N_35925);
or U36242 (N_36242,N_35600,N_35853);
xor U36243 (N_36243,N_35992,N_34700);
and U36244 (N_36244,N_35331,N_34909);
xnor U36245 (N_36245,N_34593,N_34408);
and U36246 (N_36246,N_35332,N_34097);
nand U36247 (N_36247,N_35947,N_35578);
xnor U36248 (N_36248,N_34601,N_34775);
nand U36249 (N_36249,N_34046,N_34847);
or U36250 (N_36250,N_34918,N_34371);
nand U36251 (N_36251,N_34745,N_34292);
xnor U36252 (N_36252,N_35017,N_35908);
and U36253 (N_36253,N_35742,N_35306);
nand U36254 (N_36254,N_34757,N_35320);
xor U36255 (N_36255,N_34829,N_34196);
nand U36256 (N_36256,N_35701,N_34234);
and U36257 (N_36257,N_35838,N_35678);
or U36258 (N_36258,N_34873,N_35899);
or U36259 (N_36259,N_35140,N_35905);
or U36260 (N_36260,N_35703,N_34750);
nor U36261 (N_36261,N_35609,N_35008);
and U36262 (N_36262,N_34396,N_35490);
xor U36263 (N_36263,N_35730,N_34650);
xnor U36264 (N_36264,N_34985,N_34029);
and U36265 (N_36265,N_34802,N_34037);
nor U36266 (N_36266,N_34357,N_35005);
and U36267 (N_36267,N_34093,N_34568);
and U36268 (N_36268,N_34402,N_35163);
or U36269 (N_36269,N_35316,N_35642);
xor U36270 (N_36270,N_34114,N_34558);
nor U36271 (N_36271,N_35265,N_34184);
or U36272 (N_36272,N_34584,N_35430);
and U36273 (N_36273,N_35819,N_34442);
xnor U36274 (N_36274,N_34042,N_35705);
and U36275 (N_36275,N_34143,N_35113);
or U36276 (N_36276,N_35568,N_35513);
or U36277 (N_36277,N_35782,N_34287);
or U36278 (N_36278,N_35023,N_34541);
and U36279 (N_36279,N_34209,N_34689);
and U36280 (N_36280,N_34167,N_35733);
or U36281 (N_36281,N_34171,N_34000);
xor U36282 (N_36282,N_35653,N_35489);
xor U36283 (N_36283,N_35076,N_34943);
nor U36284 (N_36284,N_35066,N_35261);
nand U36285 (N_36285,N_34315,N_34560);
xor U36286 (N_36286,N_34748,N_34302);
nor U36287 (N_36287,N_34826,N_35494);
and U36288 (N_36288,N_35453,N_34492);
nand U36289 (N_36289,N_35860,N_35334);
nand U36290 (N_36290,N_34217,N_35090);
and U36291 (N_36291,N_35798,N_34118);
or U36292 (N_36292,N_35173,N_34124);
or U36293 (N_36293,N_34364,N_35735);
nor U36294 (N_36294,N_35403,N_34743);
and U36295 (N_36295,N_35030,N_35255);
nor U36296 (N_36296,N_35797,N_35941);
nor U36297 (N_36297,N_35416,N_34923);
nor U36298 (N_36298,N_35815,N_34244);
and U36299 (N_36299,N_35926,N_34385);
or U36300 (N_36300,N_34226,N_34569);
nor U36301 (N_36301,N_34361,N_34688);
or U36302 (N_36302,N_34602,N_34220);
and U36303 (N_36303,N_35779,N_34041);
xnor U36304 (N_36304,N_35314,N_34291);
nand U36305 (N_36305,N_35055,N_34533);
or U36306 (N_36306,N_35069,N_34722);
and U36307 (N_36307,N_35247,N_35442);
or U36308 (N_36308,N_34987,N_34083);
or U36309 (N_36309,N_34933,N_34741);
nor U36310 (N_36310,N_35418,N_34010);
and U36311 (N_36311,N_34232,N_35658);
nand U36312 (N_36312,N_35888,N_35448);
and U36313 (N_36313,N_35122,N_34896);
and U36314 (N_36314,N_35052,N_35197);
or U36315 (N_36315,N_35209,N_35638);
or U36316 (N_36316,N_34908,N_35011);
or U36317 (N_36317,N_34825,N_35525);
nand U36318 (N_36318,N_34386,N_35585);
or U36319 (N_36319,N_35810,N_34738);
xnor U36320 (N_36320,N_34395,N_34059);
nand U36321 (N_36321,N_34671,N_34511);
xor U36322 (N_36322,N_34363,N_34027);
or U36323 (N_36323,N_34009,N_35850);
xnor U36324 (N_36324,N_34187,N_35580);
nor U36325 (N_36325,N_34963,N_34467);
nor U36326 (N_36326,N_34837,N_35039);
xnor U36327 (N_36327,N_35045,N_35878);
and U36328 (N_36328,N_35915,N_34728);
or U36329 (N_36329,N_34180,N_34119);
nor U36330 (N_36330,N_34656,N_34821);
nor U36331 (N_36331,N_35650,N_34956);
or U36332 (N_36332,N_35572,N_35096);
nor U36333 (N_36333,N_35450,N_35106);
and U36334 (N_36334,N_34653,N_34306);
or U36335 (N_36335,N_34194,N_34696);
or U36336 (N_36336,N_34237,N_34094);
and U36337 (N_36337,N_34358,N_35196);
nor U36338 (N_36338,N_35945,N_35929);
or U36339 (N_36339,N_35812,N_34456);
nand U36340 (N_36340,N_35698,N_35541);
and U36341 (N_36341,N_35420,N_34182);
xnor U36342 (N_36342,N_34049,N_35555);
nor U36343 (N_36343,N_35953,N_35704);
xnor U36344 (N_36344,N_35857,N_34366);
xnor U36345 (N_36345,N_35626,N_34856);
and U36346 (N_36346,N_34410,N_35272);
or U36347 (N_36347,N_34518,N_34877);
xor U36348 (N_36348,N_35322,N_35123);
nand U36349 (N_36349,N_34692,N_35276);
or U36350 (N_36350,N_34397,N_34130);
nand U36351 (N_36351,N_34892,N_34275);
or U36352 (N_36352,N_34609,N_35928);
xor U36353 (N_36353,N_34582,N_34869);
and U36354 (N_36354,N_34282,N_35760);
nor U36355 (N_36355,N_34916,N_34508);
xor U36356 (N_36356,N_34024,N_35385);
and U36357 (N_36357,N_35903,N_35594);
nand U36358 (N_36358,N_35298,N_35672);
or U36359 (N_36359,N_35451,N_34028);
or U36360 (N_36360,N_35586,N_35789);
nand U36361 (N_36361,N_34006,N_34481);
nand U36362 (N_36362,N_34479,N_35907);
nor U36363 (N_36363,N_34070,N_34756);
and U36364 (N_36364,N_35394,N_35491);
xnor U36365 (N_36365,N_34195,N_35748);
and U36366 (N_36366,N_35157,N_34631);
nor U36367 (N_36367,N_35944,N_35717);
or U36368 (N_36368,N_34365,N_34635);
nor U36369 (N_36369,N_34989,N_34870);
and U36370 (N_36370,N_34991,N_34713);
nor U36371 (N_36371,N_35089,N_34510);
or U36372 (N_36372,N_34499,N_35001);
xnor U36373 (N_36373,N_35567,N_35250);
nand U36374 (N_36374,N_34039,N_35014);
and U36375 (N_36375,N_34071,N_35665);
and U36376 (N_36376,N_35270,N_34660);
nor U36377 (N_36377,N_34038,N_35449);
and U36378 (N_36378,N_35781,N_35472);
nor U36379 (N_36379,N_35901,N_35415);
nor U36380 (N_36380,N_34081,N_34647);
nand U36381 (N_36381,N_34968,N_35178);
or U36382 (N_36382,N_34125,N_35934);
and U36383 (N_36383,N_34221,N_35223);
nor U36384 (N_36384,N_35004,N_35361);
and U36385 (N_36385,N_34138,N_35177);
and U36386 (N_36386,N_35047,N_35830);
or U36387 (N_36387,N_34036,N_35906);
nand U36388 (N_36388,N_34380,N_34812);
nor U36389 (N_36389,N_35963,N_35604);
nand U36390 (N_36390,N_35827,N_35881);
xor U36391 (N_36391,N_35235,N_34117);
nand U36392 (N_36392,N_35506,N_34519);
or U36393 (N_36393,N_34727,N_34446);
xnor U36394 (N_36394,N_35605,N_34890);
or U36395 (N_36395,N_35796,N_35294);
nor U36396 (N_36396,N_34435,N_35184);
nand U36397 (N_36397,N_34907,N_34703);
xor U36398 (N_36398,N_34186,N_35977);
nor U36399 (N_36399,N_35930,N_34507);
nand U36400 (N_36400,N_35582,N_35386);
and U36401 (N_36401,N_35000,N_35212);
and U36402 (N_36402,N_35821,N_35407);
xor U36403 (N_36403,N_35341,N_34044);
nand U36404 (N_36404,N_35865,N_34651);
or U36405 (N_36405,N_34061,N_35200);
and U36406 (N_36406,N_35304,N_34680);
nor U36407 (N_36407,N_34640,N_34910);
xnor U36408 (N_36408,N_35111,N_35771);
xnor U36409 (N_36409,N_34433,N_35639);
nor U36410 (N_36410,N_35950,N_35847);
or U36411 (N_36411,N_35060,N_35569);
or U36412 (N_36412,N_34206,N_34324);
xor U36413 (N_36413,N_34734,N_34600);
or U36414 (N_36414,N_34281,N_35120);
or U36415 (N_36415,N_35133,N_34300);
nand U36416 (N_36416,N_34776,N_34649);
xor U36417 (N_36417,N_35902,N_35602);
or U36418 (N_36418,N_34888,N_35519);
nor U36419 (N_36419,N_34598,N_34643);
xor U36420 (N_36420,N_34954,N_34491);
nor U36421 (N_36421,N_34185,N_35326);
xnor U36422 (N_36422,N_35210,N_35918);
and U36423 (N_36423,N_35354,N_34732);
or U36424 (N_36424,N_35927,N_35452);
nor U36425 (N_36425,N_35328,N_35707);
nand U36426 (N_36426,N_34394,N_35831);
nor U36427 (N_36427,N_35401,N_35095);
xor U36428 (N_36428,N_34964,N_34141);
or U36429 (N_36429,N_34707,N_35628);
xnor U36430 (N_36430,N_35195,N_34549);
and U36431 (N_36431,N_34145,N_35142);
or U36432 (N_36432,N_34154,N_35898);
xor U36433 (N_36433,N_34202,N_35598);
nand U36434 (N_36434,N_35174,N_35581);
and U36435 (N_36435,N_35203,N_35028);
and U36436 (N_36436,N_35158,N_35180);
nand U36437 (N_36437,N_35219,N_34208);
nand U36438 (N_36438,N_35024,N_35020);
xnor U36439 (N_36439,N_34706,N_35563);
or U36440 (N_36440,N_35942,N_35434);
xnor U36441 (N_36441,N_34747,N_35110);
xnor U36442 (N_36442,N_34084,N_34966);
nor U36443 (N_36443,N_34633,N_34502);
xor U36444 (N_36444,N_34253,N_35161);
xnor U36445 (N_36445,N_35713,N_35229);
nor U36446 (N_36446,N_34088,N_34258);
and U36447 (N_36447,N_35768,N_34110);
nor U36448 (N_36448,N_35057,N_34599);
nand U36449 (N_36449,N_35366,N_35603);
nand U36450 (N_36450,N_35700,N_34090);
or U36451 (N_36451,N_35621,N_34407);
xnor U36452 (N_36452,N_35858,N_35234);
nor U36453 (N_36453,N_35301,N_35957);
nor U36454 (N_36454,N_34623,N_34967);
and U36455 (N_36455,N_34670,N_35405);
nand U36456 (N_36456,N_34035,N_35972);
xnor U36457 (N_36457,N_34311,N_34487);
or U36458 (N_36458,N_34270,N_34762);
and U36459 (N_36459,N_35021,N_35997);
nand U36460 (N_36460,N_35545,N_34928);
xnor U36461 (N_36461,N_35137,N_35082);
nor U36462 (N_36462,N_35192,N_34032);
xor U36463 (N_36463,N_34789,N_35043);
and U36464 (N_36464,N_35335,N_34941);
nand U36465 (N_36465,N_34392,N_35611);
and U36466 (N_36466,N_34344,N_34080);
xnor U36467 (N_36467,N_35509,N_34595);
or U36468 (N_36468,N_35042,N_34257);
and U36469 (N_36469,N_35573,N_35851);
nor U36470 (N_36470,N_34322,N_34949);
xor U36471 (N_36471,N_34011,N_34225);
or U36472 (N_36472,N_35971,N_34337);
nand U36473 (N_36473,N_34256,N_34969);
or U36474 (N_36474,N_35254,N_34485);
xor U36475 (N_36475,N_34545,N_34993);
xnor U36476 (N_36476,N_34708,N_35336);
nand U36477 (N_36477,N_35049,N_35599);
or U36478 (N_36478,N_35438,N_35474);
nor U36479 (N_36479,N_34542,N_34721);
xor U36480 (N_36480,N_34797,N_35752);
or U36481 (N_36481,N_35290,N_34925);
xnor U36482 (N_36482,N_35775,N_34587);
xnor U36483 (N_36483,N_35367,N_35937);
nor U36484 (N_36484,N_34579,N_35439);
nand U36485 (N_36485,N_35167,N_34988);
or U36486 (N_36486,N_35984,N_35063);
nand U36487 (N_36487,N_34002,N_35199);
or U36488 (N_36488,N_34597,N_35495);
nand U36489 (N_36489,N_35296,N_34406);
and U36490 (N_36490,N_34618,N_35287);
or U36491 (N_36491,N_34457,N_35656);
and U36492 (N_36492,N_35685,N_35868);
and U36493 (N_36493,N_34230,N_34438);
and U36494 (N_36494,N_34339,N_34144);
xor U36495 (N_36495,N_35825,N_35894);
nor U36496 (N_36496,N_34440,N_34018);
and U36497 (N_36497,N_34571,N_35022);
xnor U36498 (N_36498,N_34445,N_35684);
and U36499 (N_36499,N_35809,N_34351);
nand U36500 (N_36500,N_35832,N_34165);
nand U36501 (N_36501,N_34160,N_34153);
nor U36502 (N_36502,N_34695,N_34842);
and U36503 (N_36503,N_35266,N_34769);
xnor U36504 (N_36504,N_34213,N_35182);
nand U36505 (N_36505,N_34816,N_34724);
or U36506 (N_36506,N_34161,N_34760);
nand U36507 (N_36507,N_35277,N_35054);
and U36508 (N_36508,N_34914,N_35147);
or U36509 (N_36509,N_34974,N_35071);
or U36510 (N_36510,N_34562,N_35964);
xnor U36511 (N_36511,N_34525,N_34922);
or U36512 (N_36512,N_34464,N_35471);
or U36513 (N_36513,N_35435,N_34684);
nor U36514 (N_36514,N_34704,N_34252);
or U36515 (N_36515,N_35041,N_34263);
nor U36516 (N_36516,N_35823,N_34416);
nand U36517 (N_36517,N_34065,N_35711);
nor U36518 (N_36518,N_35959,N_34448);
nand U36519 (N_36519,N_34632,N_35470);
xnor U36520 (N_36520,N_34849,N_34810);
nand U36521 (N_36521,N_35954,N_34926);
nand U36522 (N_36522,N_35770,N_34166);
xor U36523 (N_36523,N_35224,N_34735);
or U36524 (N_36524,N_34919,N_35351);
nand U36525 (N_36525,N_34003,N_34299);
or U36526 (N_36526,N_34574,N_35121);
or U36527 (N_36527,N_35511,N_35413);
nor U36528 (N_36528,N_34867,N_35515);
nor U36529 (N_36529,N_35205,N_35844);
nand U36530 (N_36530,N_35125,N_35154);
or U36531 (N_36531,N_34648,N_35426);
nor U36532 (N_36532,N_35696,N_34503);
xor U36533 (N_36533,N_34783,N_34469);
nand U36534 (N_36534,N_35731,N_34673);
nor U36535 (N_36535,N_35645,N_34886);
xor U36536 (N_36536,N_34872,N_35766);
xnor U36537 (N_36537,N_35473,N_35689);
or U36538 (N_36538,N_34173,N_35171);
nor U36539 (N_36539,N_34350,N_34489);
or U36540 (N_36540,N_34268,N_34796);
or U36541 (N_36541,N_34298,N_35922);
or U36542 (N_36542,N_34189,N_34278);
and U36543 (N_36543,N_34192,N_35211);
nand U36544 (N_36544,N_34142,N_35932);
nand U36545 (N_36545,N_35565,N_35785);
nor U36546 (N_36546,N_35059,N_34749);
or U36547 (N_36547,N_34710,N_35531);
xnor U36548 (N_36548,N_35310,N_34580);
nand U36549 (N_36549,N_34352,N_35221);
xnor U36550 (N_36550,N_34662,N_34806);
and U36551 (N_36551,N_35590,N_35053);
or U36552 (N_36552,N_35406,N_35384);
nand U36553 (N_36553,N_35104,N_34608);
or U36554 (N_36554,N_35627,N_35651);
xnor U36555 (N_36555,N_35795,N_35532);
nand U36556 (N_36556,N_34755,N_34594);
or U36557 (N_36557,N_34007,N_34719);
nor U36558 (N_36558,N_35374,N_35818);
and U36559 (N_36559,N_34434,N_34384);
nor U36560 (N_36560,N_35358,N_34548);
nor U36561 (N_36561,N_34573,N_35618);
and U36562 (N_36562,N_34576,N_35788);
nor U36563 (N_36563,N_35343,N_34795);
xor U36564 (N_36564,N_34136,N_35533);
or U36565 (N_36565,N_34494,N_35400);
and U36566 (N_36566,N_35777,N_35485);
or U36567 (N_36567,N_34219,N_34178);
nor U36568 (N_36568,N_34617,N_34556);
nor U36569 (N_36569,N_34628,N_35914);
nor U36570 (N_36570,N_35102,N_34063);
or U36571 (N_36571,N_34860,N_35132);
nor U36572 (N_36572,N_34333,N_34901);
nand U36573 (N_36573,N_34444,N_35300);
nor U36574 (N_36574,N_34296,N_35164);
nor U36575 (N_36575,N_34962,N_35616);
nor U36576 (N_36576,N_35136,N_35970);
nand U36577 (N_36577,N_34266,N_34413);
nor U36578 (N_36578,N_34627,N_34131);
xor U36579 (N_36579,N_35591,N_34427);
nor U36580 (N_36580,N_34793,N_34021);
nand U36581 (N_36581,N_34929,N_34668);
nand U36582 (N_36582,N_35012,N_34112);
nand U36583 (N_36583,N_34122,N_34913);
xnor U36584 (N_36584,N_34297,N_35166);
and U36585 (N_36585,N_34858,N_34723);
nand U36586 (N_36586,N_34624,N_35769);
and U36587 (N_36587,N_34417,N_35072);
xnor U36588 (N_36588,N_34092,N_34551);
and U36589 (N_36589,N_34105,N_35201);
xnor U36590 (N_36590,N_34742,N_35608);
nor U36591 (N_36591,N_35267,N_35003);
nor U36592 (N_36592,N_34699,N_35402);
nand U36593 (N_36593,N_34992,N_34211);
xor U36594 (N_36594,N_35813,N_34959);
nand U36595 (N_36595,N_34712,N_34831);
or U36596 (N_36596,N_34200,N_34460);
and U36597 (N_36597,N_34977,N_34883);
and U36598 (N_36598,N_35999,N_35980);
nor U36599 (N_36599,N_34882,N_34345);
nand U36600 (N_36600,N_35750,N_35303);
and U36601 (N_36601,N_35469,N_35295);
and U36602 (N_36602,N_35033,N_34879);
or U36603 (N_36603,N_34242,N_34235);
nor U36604 (N_36604,N_35791,N_34415);
nand U36605 (N_36605,N_34687,N_34621);
xnor U36606 (N_36606,N_35139,N_34619);
nand U36607 (N_36607,N_34255,N_34033);
xnor U36608 (N_36608,N_35271,N_35816);
or U36609 (N_36609,N_34981,N_34676);
nand U36610 (N_36610,N_35619,N_35204);
and U36611 (N_36611,N_35936,N_34203);
nand U36612 (N_36612,N_35546,N_34939);
nor U36613 (N_36613,N_35317,N_35445);
nand U36614 (N_36614,N_35264,N_35444);
xnor U36615 (N_36615,N_34419,N_34426);
nand U36616 (N_36616,N_34073,N_35801);
or U36617 (N_36617,N_35479,N_35933);
or U36618 (N_36618,N_34233,N_35570);
and U36619 (N_36619,N_35804,N_35909);
xor U36620 (N_36620,N_34387,N_35875);
and U36621 (N_36621,N_35372,N_35836);
nand U36622 (N_36622,N_34799,N_35983);
nand U36623 (N_36623,N_34078,N_34149);
and U36624 (N_36624,N_34501,N_35912);
nor U36625 (N_36625,N_35643,N_35183);
nor U36626 (N_36626,N_34770,N_34318);
and U36627 (N_36627,N_35647,N_34430);
nand U36628 (N_36628,N_35607,N_35974);
xor U36629 (N_36629,N_34805,N_34482);
nand U36630 (N_36630,N_34176,N_35152);
nor U36631 (N_36631,N_34915,N_34261);
xnor U36632 (N_36632,N_35329,N_34980);
nand U36633 (N_36633,N_34958,N_34374);
xnor U36634 (N_36634,N_35806,N_34972);
nor U36635 (N_36635,N_34163,N_35637);
nor U36636 (N_36636,N_34431,N_35744);
nand U36637 (N_36637,N_34865,N_35715);
and U36638 (N_36638,N_35162,N_34338);
xnor U36639 (N_36639,N_35807,N_35356);
xnor U36640 (N_36640,N_35765,N_35431);
or U36641 (N_36641,N_35961,N_35422);
nor U36642 (N_36642,N_34398,N_35630);
nand U36643 (N_36643,N_35896,N_35996);
nand U36644 (N_36644,N_34996,N_35883);
nor U36645 (N_36645,N_34683,N_35514);
nand U36646 (N_36646,N_34025,N_35692);
xor U36647 (N_36647,N_34218,N_35522);
and U36648 (N_36648,N_35321,N_35216);
nor U36649 (N_36649,N_35670,N_34955);
and U36650 (N_36650,N_34620,N_35547);
nand U36651 (N_36651,N_34478,N_35355);
or U36652 (N_36652,N_35520,N_34376);
nand U36653 (N_36653,N_34432,N_34026);
xnor U36654 (N_36654,N_35144,N_34714);
nand U36655 (N_36655,N_35676,N_35755);
nor U36656 (N_36656,N_34030,N_35510);
or U36657 (N_36657,N_34984,N_34393);
xor U36658 (N_36658,N_34681,N_34414);
nand U36659 (N_36659,N_35663,N_35483);
and U36660 (N_36660,N_34304,N_34540);
or U36661 (N_36661,N_34665,N_34147);
or U36662 (N_36662,N_35112,N_34017);
or U36663 (N_36663,N_34661,N_35728);
or U36664 (N_36664,N_34818,N_35826);
nand U36665 (N_36665,N_35465,N_35036);
or U36666 (N_36666,N_35919,N_34062);
and U36667 (N_36667,N_35185,N_35269);
and U36668 (N_36668,N_35820,N_35044);
or U36669 (N_36669,N_34817,N_35986);
nand U36670 (N_36670,N_35708,N_35040);
nor U36671 (N_36671,N_34813,N_34193);
nor U36672 (N_36672,N_35862,N_34459);
or U36673 (N_36673,N_34329,N_34957);
xor U36674 (N_36674,N_35257,N_34725);
or U36675 (N_36675,N_34657,N_34343);
and U36676 (N_36676,N_34276,N_35793);
xnor U36677 (N_36677,N_35833,N_35077);
nor U36678 (N_36678,N_35380,N_35920);
xnor U36679 (N_36679,N_35441,N_35721);
xnor U36680 (N_36680,N_34694,N_35227);
xnor U36681 (N_36681,N_34517,N_35396);
nor U36682 (N_36682,N_35958,N_35998);
nor U36683 (N_36683,N_35982,N_35652);
or U36684 (N_36684,N_35409,N_35579);
xor U36685 (N_36685,N_35226,N_34611);
or U36686 (N_36686,N_34126,N_35871);
nor U36687 (N_36687,N_35601,N_35141);
nand U36688 (N_36688,N_34828,N_35446);
xnor U36689 (N_36689,N_35682,N_35362);
nand U36690 (N_36690,N_34137,N_35800);
nor U36691 (N_36691,N_34814,N_34382);
nor U36692 (N_36692,N_34904,N_34246);
or U36693 (N_36693,N_34932,N_35064);
xor U36694 (N_36694,N_35160,N_35674);
nand U36695 (N_36695,N_35814,N_34404);
xor U36696 (N_36696,N_35553,N_35517);
nand U36697 (N_36697,N_34840,N_35556);
nor U36698 (N_36698,N_35612,N_34267);
and U36699 (N_36699,N_35252,N_34625);
or U36700 (N_36700,N_35389,N_35337);
nand U36701 (N_36701,N_34927,N_35759);
nor U36702 (N_36702,N_35889,N_35437);
nand U36703 (N_36703,N_35440,N_34895);
nor U36704 (N_36704,N_35566,N_34764);
xor U36705 (N_36705,N_34720,N_34585);
and U36706 (N_36706,N_35208,N_35808);
nor U36707 (N_36707,N_35486,N_35886);
xor U36708 (N_36708,N_35466,N_35837);
xor U36709 (N_36709,N_34325,N_35691);
or U36710 (N_36710,N_34223,N_34583);
and U36711 (N_36711,N_34753,N_35038);
xor U36712 (N_36712,N_34133,N_35459);
or U36713 (N_36713,N_35246,N_34672);
xnor U36714 (N_36714,N_34934,N_34277);
xor U36715 (N_36715,N_35537,N_35443);
nand U36716 (N_36716,N_34072,N_35763);
and U36717 (N_36717,N_34529,N_35734);
and U36718 (N_36718,N_35534,N_35482);
or U36719 (N_36719,N_35283,N_35462);
nor U36720 (N_36720,N_34401,N_35990);
xor U36721 (N_36721,N_35116,N_34099);
and U36722 (N_36722,N_34290,N_35597);
nand U36723 (N_36723,N_35249,N_34023);
nand U36724 (N_36724,N_34544,N_35657);
and U36725 (N_36725,N_34121,N_34472);
nor U36726 (N_36726,N_34614,N_35487);
and U36727 (N_36727,N_35948,N_34572);
nand U36728 (N_36728,N_34285,N_34473);
nor U36729 (N_36729,N_34578,N_34564);
nor U36730 (N_36730,N_35536,N_35170);
nand U36731 (N_36731,N_34965,N_34575);
xor U36732 (N_36732,N_35718,N_34557);
xor U36733 (N_36733,N_34040,N_34612);
and U36734 (N_36734,N_34834,N_35146);
and U36735 (N_36735,N_35027,N_34079);
and U36736 (N_36736,N_34484,N_34150);
or U36737 (N_36737,N_34833,N_35035);
nor U36738 (N_36738,N_35787,N_34780);
nand U36739 (N_36739,N_35094,N_34944);
xnor U36740 (N_36740,N_34863,N_35225);
nand U36741 (N_36741,N_35138,N_34905);
and U36742 (N_36742,N_34348,N_34677);
nor U36743 (N_36743,N_34068,N_34340);
or U36744 (N_36744,N_35562,N_34115);
xor U36745 (N_36745,N_34626,N_35390);
nor U36746 (N_36746,N_34504,N_34634);
nor U36747 (N_36747,N_34273,N_35879);
and U36748 (N_36748,N_35724,N_35228);
xnor U36749 (N_36749,N_35085,N_34752);
or U36750 (N_36750,N_34271,N_35767);
and U36751 (N_36751,N_34975,N_34763);
nand U36752 (N_36752,N_35596,N_35395);
or U36753 (N_36753,N_35610,N_34827);
xor U36754 (N_36754,N_35218,N_35217);
nand U36755 (N_36755,N_34690,N_34884);
or U36756 (N_36756,N_35549,N_34666);
and U36757 (N_36757,N_35675,N_34312);
xor U36758 (N_36758,N_35393,N_34547);
xnor U36759 (N_36759,N_34820,N_35861);
nor U36760 (N_36760,N_35849,N_35976);
or U36761 (N_36761,N_35587,N_35432);
nor U36762 (N_36762,N_34098,N_35969);
xor U36763 (N_36763,N_34240,N_35589);
nand U36764 (N_36764,N_35736,N_34616);
nand U36765 (N_36765,N_35268,N_34898);
and U36766 (N_36766,N_34373,N_35327);
nand U36767 (N_36767,N_35529,N_34116);
xor U36768 (N_36768,N_34375,N_35741);
or U36769 (N_36769,N_35115,N_35312);
and U36770 (N_36770,N_35952,N_35363);
and U36771 (N_36771,N_34458,N_34102);
nand U36772 (N_36772,N_34475,N_35839);
or U36773 (N_36773,N_34822,N_34493);
or U36774 (N_36774,N_34378,N_35544);
xnor U36775 (N_36775,N_35025,N_35979);
or U36776 (N_36776,N_34761,N_35412);
nand U36777 (N_36777,N_35917,N_34317);
nor U36778 (N_36778,N_35214,N_34249);
xnor U36779 (N_36779,N_35706,N_34855);
and U36780 (N_36780,N_35786,N_35241);
and U36781 (N_36781,N_35613,N_35949);
or U36782 (N_36782,N_34751,N_34377);
nand U36783 (N_36783,N_34264,N_35404);
nand U36784 (N_36784,N_34014,N_35662);
nand U36785 (N_36785,N_35966,N_35552);
or U36786 (N_36786,N_34698,N_35622);
and U36787 (N_36787,N_35097,N_35625);
or U36788 (N_36788,N_35002,N_34004);
xnor U36789 (N_36789,N_35433,N_35375);
nor U36790 (N_36790,N_35262,N_35939);
xnor U36791 (N_36791,N_34179,N_35239);
nand U36792 (N_36792,N_34441,N_34020);
nand U36793 (N_36793,N_35938,N_34970);
nand U36794 (N_36794,N_35981,N_34516);
nand U36795 (N_36795,N_34188,N_35620);
xor U36796 (N_36796,N_34389,N_34175);
and U36797 (N_36797,N_34259,N_35882);
nor U36798 (N_36798,N_35213,N_34702);
or U36799 (N_36799,N_35134,N_35189);
nor U36800 (N_36800,N_35669,N_34787);
xor U36801 (N_36801,N_35370,N_34997);
or U36802 (N_36802,N_34554,N_35179);
or U36803 (N_36803,N_35109,N_35774);
xor U36804 (N_36804,N_34709,N_35347);
nand U36805 (N_36805,N_35302,N_34305);
nor U36806 (N_36806,N_34513,N_34428);
nand U36807 (N_36807,N_34245,N_35467);
and U36808 (N_36808,N_34937,N_35046);
or U36809 (N_36809,N_34342,N_35016);
and U36810 (N_36810,N_34379,N_34422);
xnor U36811 (N_36811,N_35887,N_35319);
or U36812 (N_36812,N_35940,N_34129);
nand U36813 (N_36813,N_35181,N_35654);
or U36814 (N_36814,N_35073,N_35010);
nor U36815 (N_36815,N_35502,N_35891);
nor U36816 (N_36816,N_35079,N_34801);
nor U36817 (N_36817,N_35175,N_34591);
nor U36818 (N_36818,N_34746,N_34622);
nand U36819 (N_36819,N_34505,N_35155);
or U36820 (N_36820,N_34739,N_35540);
nor U36821 (N_36821,N_34069,N_35365);
nor U36822 (N_36822,N_35026,N_34443);
or U36823 (N_36823,N_34658,N_34055);
and U36824 (N_36824,N_34912,N_35468);
nor U36825 (N_36825,N_35671,N_34664);
or U36826 (N_36826,N_34331,N_34638);
or U36827 (N_36827,N_34532,N_35835);
and U36828 (N_36828,N_34316,N_35253);
or U36829 (N_36829,N_35499,N_35595);
nor U36830 (N_36830,N_35841,N_34314);
nand U36831 (N_36831,N_34920,N_34334);
nand U36832 (N_36832,N_34555,N_34076);
or U36833 (N_36833,N_35075,N_35913);
or U36834 (N_36834,N_35383,N_35484);
xor U36835 (N_36835,N_34170,N_35680);
nand U36836 (N_36836,N_34950,N_35512);
or U36837 (N_36837,N_34857,N_35756);
nor U36838 (N_36838,N_34162,N_34655);
nand U36839 (N_36839,N_35458,N_34214);
and U36840 (N_36840,N_34280,N_34530);
and U36841 (N_36841,N_34773,N_35846);
nor U36842 (N_36842,N_35634,N_34782);
xor U36843 (N_36843,N_35720,N_34470);
and U36844 (N_36844,N_35187,N_34893);
and U36845 (N_36845,N_35773,N_34295);
nor U36846 (N_36846,N_35093,N_35371);
and U36847 (N_36847,N_34107,N_35890);
xor U36848 (N_36848,N_34012,N_35381);
xor U36849 (N_36849,N_34051,N_34726);
xnor U36850 (N_36850,N_34646,N_35159);
nor U36851 (N_36851,N_34940,N_34238);
or U36852 (N_36852,N_35151,N_35447);
and U36853 (N_36853,N_35877,N_35575);
and U36854 (N_36854,N_35242,N_34056);
and U36855 (N_36855,N_34862,N_35143);
or U36856 (N_36856,N_34771,N_35463);
xnor U36857 (N_36857,N_35088,N_35571);
or U36858 (N_36858,N_35056,N_34335);
or U36859 (N_36859,N_34961,N_35635);
nor U36860 (N_36860,N_35315,N_35866);
or U36861 (N_36861,N_34768,N_34790);
xnor U36862 (N_36862,N_35753,N_35530);
nor U36863 (N_36863,N_34190,N_34013);
xor U36864 (N_36864,N_35149,N_35501);
or U36865 (N_36865,N_34388,N_34231);
nand U36866 (N_36866,N_35995,N_34429);
nand U36867 (N_36867,N_34835,N_35339);
nand U36868 (N_36868,N_35414,N_34359);
nor U36869 (N_36869,N_35186,N_34588);
nand U36870 (N_36870,N_34754,N_34868);
and U36871 (N_36871,N_35359,N_35631);
or U36872 (N_36872,N_34691,N_35092);
and U36873 (N_36873,N_35165,N_34973);
and U36874 (N_36874,N_35746,N_35153);
or U36875 (N_36875,N_34815,N_34539);
nand U36876 (N_36876,N_35683,N_35475);
nor U36877 (N_36877,N_35764,N_35281);
nand U36878 (N_36878,N_35150,N_35688);
nor U36879 (N_36879,N_35172,N_34902);
nor U36880 (N_36880,N_34509,N_35535);
xnor U36881 (N_36881,N_35454,N_35428);
or U36882 (N_36882,N_34439,N_34465);
and U36883 (N_36883,N_34215,N_35425);
xnor U36884 (N_36884,N_34449,N_35397);
xnor U36885 (N_36885,N_34903,N_35019);
and U36886 (N_36886,N_34931,N_34008);
xor U36887 (N_36887,N_35911,N_35834);
nand U36888 (N_36888,N_35712,N_35427);
or U36889 (N_36889,N_34736,N_35951);
nor U36890 (N_36890,N_34543,N_34156);
xor U36891 (N_36891,N_35576,N_34360);
nand U36892 (N_36892,N_34786,N_35624);
xnor U36893 (N_36893,N_35318,N_35687);
nor U36894 (N_36894,N_35542,N_35623);
xnor U36895 (N_36895,N_35288,N_35018);
nor U36896 (N_36896,N_35124,N_34205);
nor U36897 (N_36897,N_35667,N_35778);
xnor U36898 (N_36898,N_34212,N_34109);
nor U36899 (N_36899,N_34552,N_35543);
xnor U36900 (N_36900,N_35476,N_34995);
nand U36901 (N_36901,N_35220,N_35379);
nand U36902 (N_36902,N_34978,N_34535);
xnor U36903 (N_36903,N_35368,N_35309);
nor U36904 (N_36904,N_34861,N_34423);
nor U36905 (N_36905,N_34096,N_35411);
nand U36906 (N_36906,N_35644,N_34057);
or U36907 (N_36907,N_34701,N_34531);
or U36908 (N_36908,N_35719,N_35710);
and U36909 (N_36909,N_35558,N_35286);
xnor U36910 (N_36910,N_34243,N_34733);
nor U36911 (N_36911,N_34871,N_34851);
nand U36912 (N_36912,N_34800,N_35564);
nor U36913 (N_36913,N_34104,N_35802);
or U36914 (N_36914,N_34744,N_35492);
nor U36915 (N_36915,N_34022,N_35646);
nand U36916 (N_36916,N_35131,N_34321);
nand U36917 (N_36917,N_35352,N_35084);
or U36918 (N_36918,N_35956,N_34779);
nand U36919 (N_36919,N_34644,N_34536);
nand U36920 (N_36920,N_34889,N_35191);
xor U36921 (N_36921,N_35051,N_35480);
nand U36922 (N_36922,N_35194,N_35382);
nand U36923 (N_36923,N_35943,N_34052);
or U36924 (N_36924,N_35714,N_34169);
nor U36925 (N_36925,N_34715,N_34994);
nand U36926 (N_36926,N_35477,N_35369);
xor U36927 (N_36927,N_34930,N_34960);
xor U36928 (N_36928,N_34885,N_35305);
or U36929 (N_36929,N_34086,N_34356);
nor U36930 (N_36930,N_34155,N_34774);
nor U36931 (N_36931,N_34951,N_35080);
nor U36932 (N_36932,N_34514,N_34561);
xnor U36933 (N_36933,N_34603,N_35661);
xor U36934 (N_36934,N_34113,N_34758);
xnor U36935 (N_36935,N_34347,N_34971);
nand U36936 (N_36936,N_35408,N_34323);
nor U36937 (N_36937,N_35419,N_34228);
nor U36938 (N_36938,N_35955,N_35559);
xnor U36939 (N_36939,N_35805,N_34455);
nor U36940 (N_36940,N_34204,N_35867);
or U36941 (N_36941,N_34785,N_35338);
nor U36942 (N_36942,N_35987,N_35284);
or U36943 (N_36943,N_35424,N_35614);
nand U36944 (N_36944,N_35311,N_34341);
and U36945 (N_36945,N_34798,N_34412);
xor U36946 (N_36946,N_34792,N_34058);
nor U36947 (N_36947,N_35129,N_35528);
and U36948 (N_36948,N_35852,N_34586);
xor U36949 (N_36949,N_34850,N_35493);
and U36950 (N_36950,N_35238,N_35749);
nor U36951 (N_36951,N_34085,N_34089);
nor U36952 (N_36952,N_35524,N_34272);
or U36953 (N_36953,N_34900,N_34288);
or U36954 (N_36954,N_34911,N_35695);
xor U36955 (N_36955,N_34848,N_34841);
or U36956 (N_36956,N_35496,N_34983);
and U36957 (N_36957,N_34999,N_35910);
or U36958 (N_36958,N_34730,N_34332);
nand U36959 (N_36959,N_35551,N_35725);
nor U36960 (N_36960,N_34610,N_34060);
or U36961 (N_36961,N_34948,N_34405);
nor U36962 (N_36962,N_34468,N_34731);
nand U36963 (N_36963,N_34224,N_35739);
nor U36964 (N_36964,N_34717,N_34559);
nor U36965 (N_36965,N_35574,N_34174);
nand U36966 (N_36966,N_35364,N_34128);
and U36967 (N_36967,N_35723,N_34307);
nand U36968 (N_36968,N_34139,N_35743);
nor U36969 (N_36969,N_34523,N_34565);
xor U36970 (N_36970,N_35822,N_35641);
or U36971 (N_36971,N_35668,N_35516);
or U36972 (N_36972,N_35398,N_35649);
xnor U36973 (N_36973,N_35632,N_34500);
nor U36974 (N_36974,N_35892,N_34685);
nand U36975 (N_36975,N_35353,N_35202);
nor U36976 (N_36976,N_35323,N_34629);
nor U36977 (N_36977,N_34269,N_34197);
xnor U36978 (N_36978,N_35236,N_34301);
xnor U36979 (N_36979,N_35128,N_35388);
and U36980 (N_36980,N_34313,N_35872);
nand U36981 (N_36981,N_35794,N_35648);
and U36982 (N_36982,N_34645,N_34496);
nand U36983 (N_36983,N_35135,N_35848);
and U36984 (N_36984,N_35168,N_34320);
and U36985 (N_36985,N_35776,N_35993);
and U36986 (N_36986,N_34289,N_35967);
and U36987 (N_36987,N_34476,N_34606);
nand U36988 (N_36988,N_35666,N_34921);
nand U36989 (N_36989,N_35308,N_34152);
nor U36990 (N_36990,N_34101,N_35716);
nor U36991 (N_36991,N_35916,N_34853);
nand U36992 (N_36992,N_34737,N_34274);
and U36993 (N_36993,N_34682,N_35523);
xor U36994 (N_36994,N_35799,N_34450);
or U36995 (N_36995,N_34466,N_35978);
or U36996 (N_36996,N_35376,N_35991);
nand U36997 (N_36997,N_35240,N_34577);
xnor U36998 (N_36998,N_35377,N_35884);
xnor U36999 (N_36999,N_34075,N_35709);
nand U37000 (N_37000,N_35496,N_35004);
and U37001 (N_37001,N_35517,N_35595);
nand U37002 (N_37002,N_35523,N_34211);
nor U37003 (N_37003,N_35172,N_34177);
or U37004 (N_37004,N_34444,N_35250);
xor U37005 (N_37005,N_34414,N_34721);
nor U37006 (N_37006,N_35078,N_35720);
and U37007 (N_37007,N_35673,N_35507);
xor U37008 (N_37008,N_35175,N_34986);
or U37009 (N_37009,N_35392,N_35639);
or U37010 (N_37010,N_35505,N_34081);
nand U37011 (N_37011,N_34421,N_34475);
nor U37012 (N_37012,N_34955,N_34566);
xnor U37013 (N_37013,N_35081,N_34372);
xor U37014 (N_37014,N_35335,N_34066);
or U37015 (N_37015,N_34891,N_35404);
nand U37016 (N_37016,N_34248,N_35209);
nand U37017 (N_37017,N_34927,N_35068);
nand U37018 (N_37018,N_34665,N_35728);
xnor U37019 (N_37019,N_34858,N_34435);
nand U37020 (N_37020,N_34969,N_34365);
nand U37021 (N_37021,N_34242,N_35474);
or U37022 (N_37022,N_34248,N_35411);
nor U37023 (N_37023,N_34737,N_35766);
xor U37024 (N_37024,N_35273,N_35020);
xor U37025 (N_37025,N_35988,N_34314);
and U37026 (N_37026,N_35284,N_34138);
and U37027 (N_37027,N_35207,N_35195);
or U37028 (N_37028,N_34310,N_34024);
nor U37029 (N_37029,N_35054,N_34172);
or U37030 (N_37030,N_34328,N_34260);
or U37031 (N_37031,N_35031,N_35494);
nand U37032 (N_37032,N_35355,N_35011);
or U37033 (N_37033,N_34652,N_35505);
and U37034 (N_37034,N_34964,N_34446);
nor U37035 (N_37035,N_34034,N_34883);
xor U37036 (N_37036,N_35144,N_34215);
or U37037 (N_37037,N_34376,N_35362);
and U37038 (N_37038,N_34696,N_35490);
nand U37039 (N_37039,N_34792,N_34546);
or U37040 (N_37040,N_34995,N_35045);
or U37041 (N_37041,N_35416,N_34503);
nand U37042 (N_37042,N_34133,N_35347);
or U37043 (N_37043,N_34034,N_35535);
and U37044 (N_37044,N_35717,N_35421);
or U37045 (N_37045,N_35189,N_35532);
nor U37046 (N_37046,N_34944,N_35803);
nand U37047 (N_37047,N_35938,N_34539);
or U37048 (N_37048,N_34814,N_34329);
or U37049 (N_37049,N_34174,N_35636);
or U37050 (N_37050,N_35333,N_35301);
or U37051 (N_37051,N_35773,N_34399);
xnor U37052 (N_37052,N_35742,N_34132);
nand U37053 (N_37053,N_35035,N_34187);
or U37054 (N_37054,N_35484,N_35369);
nand U37055 (N_37055,N_35468,N_35637);
and U37056 (N_37056,N_35364,N_34576);
nand U37057 (N_37057,N_35880,N_35984);
and U37058 (N_37058,N_35564,N_34660);
nor U37059 (N_37059,N_34046,N_34470);
nand U37060 (N_37060,N_34324,N_35986);
and U37061 (N_37061,N_34257,N_35127);
nand U37062 (N_37062,N_34092,N_35906);
and U37063 (N_37063,N_34174,N_34408);
or U37064 (N_37064,N_34533,N_35126);
xnor U37065 (N_37065,N_34203,N_34728);
or U37066 (N_37066,N_34613,N_35087);
and U37067 (N_37067,N_35690,N_35216);
nand U37068 (N_37068,N_35690,N_34964);
xnor U37069 (N_37069,N_34252,N_35789);
nand U37070 (N_37070,N_35592,N_34214);
nand U37071 (N_37071,N_35621,N_35699);
or U37072 (N_37072,N_35109,N_35038);
xnor U37073 (N_37073,N_34025,N_34149);
or U37074 (N_37074,N_34907,N_34239);
nor U37075 (N_37075,N_34310,N_34835);
xnor U37076 (N_37076,N_34995,N_35606);
nor U37077 (N_37077,N_34626,N_35900);
nor U37078 (N_37078,N_35107,N_35613);
nor U37079 (N_37079,N_34230,N_34527);
nor U37080 (N_37080,N_34656,N_35321);
or U37081 (N_37081,N_34054,N_34991);
and U37082 (N_37082,N_35873,N_35984);
nor U37083 (N_37083,N_35612,N_34225);
nand U37084 (N_37084,N_34433,N_34196);
and U37085 (N_37085,N_35155,N_34397);
nand U37086 (N_37086,N_35610,N_34618);
and U37087 (N_37087,N_34990,N_34072);
or U37088 (N_37088,N_35676,N_34799);
nor U37089 (N_37089,N_34016,N_35073);
nor U37090 (N_37090,N_34326,N_35121);
nor U37091 (N_37091,N_34477,N_35356);
and U37092 (N_37092,N_35374,N_34544);
and U37093 (N_37093,N_35427,N_35130);
xnor U37094 (N_37094,N_35624,N_34469);
and U37095 (N_37095,N_35019,N_34030);
or U37096 (N_37096,N_35687,N_35532);
or U37097 (N_37097,N_35195,N_35869);
or U37098 (N_37098,N_34239,N_35869);
nand U37099 (N_37099,N_34374,N_34992);
xor U37100 (N_37100,N_35897,N_35619);
or U37101 (N_37101,N_34455,N_35002);
nor U37102 (N_37102,N_34373,N_35907);
nand U37103 (N_37103,N_34345,N_35783);
nand U37104 (N_37104,N_35748,N_35470);
nor U37105 (N_37105,N_35203,N_35354);
nand U37106 (N_37106,N_35121,N_35317);
or U37107 (N_37107,N_35268,N_34549);
and U37108 (N_37108,N_34362,N_34749);
and U37109 (N_37109,N_35946,N_35848);
nand U37110 (N_37110,N_35508,N_35943);
and U37111 (N_37111,N_34119,N_34810);
and U37112 (N_37112,N_35983,N_34571);
nor U37113 (N_37113,N_34463,N_35441);
and U37114 (N_37114,N_35197,N_35238);
and U37115 (N_37115,N_34878,N_35707);
nand U37116 (N_37116,N_34393,N_34402);
and U37117 (N_37117,N_35352,N_34248);
and U37118 (N_37118,N_35426,N_35433);
and U37119 (N_37119,N_35772,N_35792);
nor U37120 (N_37120,N_34837,N_34010);
or U37121 (N_37121,N_34245,N_35110);
or U37122 (N_37122,N_35124,N_34308);
or U37123 (N_37123,N_34898,N_35262);
nor U37124 (N_37124,N_35366,N_34568);
and U37125 (N_37125,N_34174,N_35343);
xnor U37126 (N_37126,N_35192,N_34856);
and U37127 (N_37127,N_35469,N_34475);
nor U37128 (N_37128,N_34920,N_35556);
xor U37129 (N_37129,N_34465,N_35731);
or U37130 (N_37130,N_34030,N_34693);
and U37131 (N_37131,N_35128,N_35455);
nor U37132 (N_37132,N_34250,N_34066);
or U37133 (N_37133,N_34475,N_34241);
xor U37134 (N_37134,N_35258,N_34334);
nand U37135 (N_37135,N_34617,N_34641);
and U37136 (N_37136,N_34707,N_35787);
nand U37137 (N_37137,N_34879,N_34824);
and U37138 (N_37138,N_34013,N_35886);
xnor U37139 (N_37139,N_35181,N_35366);
xnor U37140 (N_37140,N_35108,N_34581);
and U37141 (N_37141,N_35120,N_35103);
and U37142 (N_37142,N_35784,N_34368);
or U37143 (N_37143,N_34839,N_35396);
xnor U37144 (N_37144,N_34615,N_35114);
xor U37145 (N_37145,N_34503,N_34766);
xnor U37146 (N_37146,N_35036,N_35983);
nor U37147 (N_37147,N_35401,N_34040);
nor U37148 (N_37148,N_34884,N_35840);
nor U37149 (N_37149,N_34766,N_34586);
nand U37150 (N_37150,N_35979,N_34631);
or U37151 (N_37151,N_35000,N_35879);
or U37152 (N_37152,N_35689,N_34270);
and U37153 (N_37153,N_34354,N_35704);
and U37154 (N_37154,N_35691,N_34301);
nand U37155 (N_37155,N_35582,N_34434);
and U37156 (N_37156,N_34837,N_35175);
xor U37157 (N_37157,N_34193,N_35913);
or U37158 (N_37158,N_34009,N_34526);
or U37159 (N_37159,N_35438,N_35361);
or U37160 (N_37160,N_34393,N_35602);
or U37161 (N_37161,N_34658,N_34795);
or U37162 (N_37162,N_35855,N_35912);
xor U37163 (N_37163,N_34143,N_34673);
and U37164 (N_37164,N_34640,N_35934);
and U37165 (N_37165,N_34111,N_35084);
nand U37166 (N_37166,N_35741,N_34673);
nor U37167 (N_37167,N_34699,N_34956);
xor U37168 (N_37168,N_34936,N_35717);
and U37169 (N_37169,N_34201,N_34483);
nand U37170 (N_37170,N_35642,N_35969);
and U37171 (N_37171,N_34828,N_35414);
and U37172 (N_37172,N_34638,N_35505);
nand U37173 (N_37173,N_34055,N_34346);
or U37174 (N_37174,N_34036,N_34295);
xnor U37175 (N_37175,N_34824,N_34036);
nand U37176 (N_37176,N_35312,N_34037);
nor U37177 (N_37177,N_35577,N_35687);
xnor U37178 (N_37178,N_34598,N_35087);
xnor U37179 (N_37179,N_34064,N_34750);
nor U37180 (N_37180,N_34866,N_35087);
nor U37181 (N_37181,N_34388,N_35080);
nand U37182 (N_37182,N_35519,N_35037);
nor U37183 (N_37183,N_34090,N_35558);
nand U37184 (N_37184,N_35733,N_35882);
xor U37185 (N_37185,N_34705,N_35442);
or U37186 (N_37186,N_35012,N_34788);
or U37187 (N_37187,N_34585,N_34130);
xor U37188 (N_37188,N_34995,N_34270);
xor U37189 (N_37189,N_35643,N_35923);
nor U37190 (N_37190,N_35314,N_35266);
xnor U37191 (N_37191,N_34757,N_34365);
nand U37192 (N_37192,N_35674,N_34019);
xor U37193 (N_37193,N_35636,N_35289);
or U37194 (N_37194,N_35631,N_34767);
xnor U37195 (N_37195,N_34695,N_35020);
xnor U37196 (N_37196,N_35186,N_34317);
and U37197 (N_37197,N_35117,N_35420);
xnor U37198 (N_37198,N_34320,N_35869);
nand U37199 (N_37199,N_34492,N_34920);
nand U37200 (N_37200,N_34915,N_35530);
nor U37201 (N_37201,N_34419,N_35442);
or U37202 (N_37202,N_35419,N_35839);
or U37203 (N_37203,N_35375,N_34258);
or U37204 (N_37204,N_35926,N_35150);
or U37205 (N_37205,N_35273,N_35227);
nor U37206 (N_37206,N_35930,N_35635);
nor U37207 (N_37207,N_34476,N_34686);
or U37208 (N_37208,N_35842,N_35683);
or U37209 (N_37209,N_35291,N_34530);
nor U37210 (N_37210,N_35413,N_35408);
nor U37211 (N_37211,N_35090,N_34764);
nor U37212 (N_37212,N_35229,N_35400);
and U37213 (N_37213,N_35662,N_35112);
nor U37214 (N_37214,N_34428,N_34218);
nor U37215 (N_37215,N_34216,N_35639);
nor U37216 (N_37216,N_34430,N_34583);
nand U37217 (N_37217,N_35594,N_35006);
or U37218 (N_37218,N_34303,N_34037);
and U37219 (N_37219,N_34303,N_35325);
nand U37220 (N_37220,N_34466,N_34824);
xor U37221 (N_37221,N_34750,N_35059);
nand U37222 (N_37222,N_35917,N_34683);
nor U37223 (N_37223,N_35964,N_35398);
nor U37224 (N_37224,N_34353,N_34339);
or U37225 (N_37225,N_35230,N_34893);
nor U37226 (N_37226,N_34733,N_35401);
nand U37227 (N_37227,N_34902,N_34370);
or U37228 (N_37228,N_34833,N_35706);
nand U37229 (N_37229,N_34219,N_34237);
and U37230 (N_37230,N_34450,N_34400);
nor U37231 (N_37231,N_35668,N_35910);
nor U37232 (N_37232,N_35134,N_34610);
nand U37233 (N_37233,N_35621,N_35142);
and U37234 (N_37234,N_34331,N_35370);
or U37235 (N_37235,N_34388,N_34552);
and U37236 (N_37236,N_35680,N_35183);
nor U37237 (N_37237,N_34621,N_34510);
or U37238 (N_37238,N_34820,N_35571);
xor U37239 (N_37239,N_35427,N_34700);
or U37240 (N_37240,N_34522,N_34414);
nor U37241 (N_37241,N_35528,N_35988);
nor U37242 (N_37242,N_34278,N_35591);
and U37243 (N_37243,N_34040,N_35150);
and U37244 (N_37244,N_35869,N_34460);
nor U37245 (N_37245,N_34057,N_34143);
nor U37246 (N_37246,N_34015,N_34416);
nand U37247 (N_37247,N_35420,N_34758);
or U37248 (N_37248,N_35117,N_34462);
and U37249 (N_37249,N_35066,N_34423);
and U37250 (N_37250,N_34990,N_34137);
and U37251 (N_37251,N_34427,N_35207);
or U37252 (N_37252,N_35706,N_35810);
nand U37253 (N_37253,N_34753,N_34343);
xor U37254 (N_37254,N_35726,N_35121);
nand U37255 (N_37255,N_34992,N_35741);
and U37256 (N_37256,N_34571,N_35118);
and U37257 (N_37257,N_34603,N_35002);
nand U37258 (N_37258,N_34762,N_35875);
nand U37259 (N_37259,N_35791,N_34201);
or U37260 (N_37260,N_35797,N_35503);
nand U37261 (N_37261,N_35682,N_34805);
xnor U37262 (N_37262,N_35919,N_35387);
or U37263 (N_37263,N_34680,N_35495);
or U37264 (N_37264,N_34414,N_34813);
or U37265 (N_37265,N_35277,N_35446);
or U37266 (N_37266,N_34013,N_34897);
or U37267 (N_37267,N_35519,N_35577);
xor U37268 (N_37268,N_34665,N_35923);
nand U37269 (N_37269,N_35729,N_35756);
and U37270 (N_37270,N_34421,N_35191);
nand U37271 (N_37271,N_34131,N_34923);
nand U37272 (N_37272,N_34537,N_35937);
or U37273 (N_37273,N_34029,N_34120);
nor U37274 (N_37274,N_35693,N_34361);
nand U37275 (N_37275,N_35586,N_34205);
or U37276 (N_37276,N_35071,N_35911);
or U37277 (N_37277,N_35263,N_35182);
xnor U37278 (N_37278,N_35085,N_35412);
xnor U37279 (N_37279,N_35793,N_35762);
or U37280 (N_37280,N_34902,N_35439);
xor U37281 (N_37281,N_34113,N_34130);
xnor U37282 (N_37282,N_34195,N_34035);
nand U37283 (N_37283,N_34014,N_34456);
nand U37284 (N_37284,N_34850,N_34966);
and U37285 (N_37285,N_35926,N_34397);
nor U37286 (N_37286,N_34360,N_34335);
xor U37287 (N_37287,N_34686,N_34245);
or U37288 (N_37288,N_35381,N_34296);
or U37289 (N_37289,N_34505,N_34955);
nor U37290 (N_37290,N_35857,N_34411);
or U37291 (N_37291,N_34410,N_35695);
or U37292 (N_37292,N_35142,N_34519);
and U37293 (N_37293,N_35557,N_34773);
nand U37294 (N_37294,N_35679,N_34337);
nand U37295 (N_37295,N_34458,N_35839);
xor U37296 (N_37296,N_35115,N_34154);
or U37297 (N_37297,N_35969,N_35368);
nand U37298 (N_37298,N_35353,N_34293);
nand U37299 (N_37299,N_34750,N_34645);
nand U37300 (N_37300,N_35833,N_34745);
xnor U37301 (N_37301,N_34727,N_35711);
xor U37302 (N_37302,N_34223,N_35620);
or U37303 (N_37303,N_35715,N_34963);
and U37304 (N_37304,N_34042,N_35999);
xnor U37305 (N_37305,N_34218,N_34360);
or U37306 (N_37306,N_35354,N_34034);
and U37307 (N_37307,N_34325,N_35891);
xor U37308 (N_37308,N_35538,N_34754);
and U37309 (N_37309,N_34554,N_35356);
or U37310 (N_37310,N_34790,N_35139);
or U37311 (N_37311,N_34459,N_34932);
nor U37312 (N_37312,N_35605,N_35529);
or U37313 (N_37313,N_34161,N_35289);
xor U37314 (N_37314,N_35431,N_34890);
xor U37315 (N_37315,N_34255,N_34595);
xor U37316 (N_37316,N_35587,N_35898);
nand U37317 (N_37317,N_35889,N_34240);
nand U37318 (N_37318,N_35376,N_34666);
nand U37319 (N_37319,N_35128,N_35774);
or U37320 (N_37320,N_34842,N_34470);
xnor U37321 (N_37321,N_35760,N_35771);
nand U37322 (N_37322,N_34783,N_34537);
or U37323 (N_37323,N_35740,N_35224);
or U37324 (N_37324,N_35539,N_35859);
nor U37325 (N_37325,N_35236,N_35538);
xnor U37326 (N_37326,N_34761,N_34674);
or U37327 (N_37327,N_35597,N_35097);
nand U37328 (N_37328,N_34803,N_35242);
or U37329 (N_37329,N_34955,N_34057);
xnor U37330 (N_37330,N_34566,N_34987);
nor U37331 (N_37331,N_35706,N_34527);
xor U37332 (N_37332,N_34025,N_34819);
or U37333 (N_37333,N_35495,N_34449);
nand U37334 (N_37334,N_34816,N_34750);
or U37335 (N_37335,N_34060,N_35587);
xnor U37336 (N_37336,N_35727,N_35828);
nor U37337 (N_37337,N_34061,N_35899);
xor U37338 (N_37338,N_34998,N_34869);
or U37339 (N_37339,N_35042,N_35613);
or U37340 (N_37340,N_35492,N_35425);
nand U37341 (N_37341,N_35245,N_34179);
and U37342 (N_37342,N_35138,N_34408);
or U37343 (N_37343,N_34096,N_35798);
nand U37344 (N_37344,N_34181,N_34625);
and U37345 (N_37345,N_35708,N_34584);
xor U37346 (N_37346,N_34055,N_35876);
nor U37347 (N_37347,N_34662,N_34807);
nor U37348 (N_37348,N_34072,N_34901);
nand U37349 (N_37349,N_35914,N_35114);
nand U37350 (N_37350,N_35530,N_34235);
xor U37351 (N_37351,N_34729,N_34736);
nand U37352 (N_37352,N_35512,N_35586);
nor U37353 (N_37353,N_34826,N_35547);
nor U37354 (N_37354,N_35951,N_34003);
or U37355 (N_37355,N_35784,N_35769);
nand U37356 (N_37356,N_34582,N_35049);
or U37357 (N_37357,N_34438,N_34330);
and U37358 (N_37358,N_35621,N_35168);
nand U37359 (N_37359,N_35815,N_35549);
nor U37360 (N_37360,N_34815,N_34626);
and U37361 (N_37361,N_35863,N_34927);
and U37362 (N_37362,N_34558,N_34563);
or U37363 (N_37363,N_35859,N_34243);
xor U37364 (N_37364,N_35898,N_35369);
or U37365 (N_37365,N_34892,N_34775);
and U37366 (N_37366,N_34990,N_34788);
and U37367 (N_37367,N_35349,N_34432);
and U37368 (N_37368,N_35491,N_35760);
and U37369 (N_37369,N_34119,N_35464);
xor U37370 (N_37370,N_34072,N_34733);
xnor U37371 (N_37371,N_35713,N_35983);
nor U37372 (N_37372,N_35783,N_34734);
nand U37373 (N_37373,N_35021,N_34618);
nor U37374 (N_37374,N_34177,N_35598);
or U37375 (N_37375,N_34858,N_35811);
nand U37376 (N_37376,N_35523,N_35406);
xnor U37377 (N_37377,N_34974,N_35512);
nor U37378 (N_37378,N_34498,N_35460);
nor U37379 (N_37379,N_34274,N_34211);
nor U37380 (N_37380,N_35946,N_34909);
xnor U37381 (N_37381,N_34028,N_34090);
and U37382 (N_37382,N_35369,N_35873);
or U37383 (N_37383,N_34856,N_34391);
nand U37384 (N_37384,N_34231,N_34268);
nand U37385 (N_37385,N_35932,N_34742);
nand U37386 (N_37386,N_35514,N_35603);
nand U37387 (N_37387,N_34977,N_34919);
nor U37388 (N_37388,N_35707,N_35416);
and U37389 (N_37389,N_34333,N_35555);
and U37390 (N_37390,N_34168,N_35234);
nor U37391 (N_37391,N_34325,N_35080);
and U37392 (N_37392,N_34397,N_34201);
xnor U37393 (N_37393,N_34481,N_34062);
xnor U37394 (N_37394,N_34958,N_34439);
and U37395 (N_37395,N_35086,N_34385);
xnor U37396 (N_37396,N_34276,N_34157);
nand U37397 (N_37397,N_35558,N_35949);
xnor U37398 (N_37398,N_34828,N_35174);
and U37399 (N_37399,N_34588,N_35131);
or U37400 (N_37400,N_35504,N_35888);
and U37401 (N_37401,N_35884,N_34912);
nand U37402 (N_37402,N_35107,N_34722);
and U37403 (N_37403,N_35841,N_35166);
xnor U37404 (N_37404,N_35794,N_34130);
nor U37405 (N_37405,N_35312,N_35018);
xnor U37406 (N_37406,N_34123,N_35686);
nand U37407 (N_37407,N_35581,N_35823);
and U37408 (N_37408,N_35870,N_34041);
xor U37409 (N_37409,N_35395,N_34532);
and U37410 (N_37410,N_35930,N_34410);
nand U37411 (N_37411,N_34494,N_34620);
nor U37412 (N_37412,N_35173,N_34428);
nand U37413 (N_37413,N_34972,N_35527);
nor U37414 (N_37414,N_35953,N_35770);
nand U37415 (N_37415,N_35097,N_35894);
and U37416 (N_37416,N_35555,N_34121);
xor U37417 (N_37417,N_35843,N_35524);
nor U37418 (N_37418,N_34381,N_35088);
nand U37419 (N_37419,N_35119,N_35810);
or U37420 (N_37420,N_34339,N_34179);
nor U37421 (N_37421,N_35102,N_35314);
or U37422 (N_37422,N_35578,N_34050);
or U37423 (N_37423,N_35475,N_35811);
and U37424 (N_37424,N_34604,N_35417);
xnor U37425 (N_37425,N_34280,N_34254);
xor U37426 (N_37426,N_35165,N_34420);
xnor U37427 (N_37427,N_35590,N_34460);
nand U37428 (N_37428,N_35699,N_35052);
nor U37429 (N_37429,N_35145,N_35904);
nor U37430 (N_37430,N_35530,N_34479);
and U37431 (N_37431,N_34858,N_34885);
nor U37432 (N_37432,N_35627,N_34592);
or U37433 (N_37433,N_35091,N_34377);
nand U37434 (N_37434,N_35170,N_34146);
nand U37435 (N_37435,N_34940,N_34502);
or U37436 (N_37436,N_34143,N_35296);
nand U37437 (N_37437,N_34508,N_35793);
and U37438 (N_37438,N_34866,N_35561);
xor U37439 (N_37439,N_34415,N_34300);
xor U37440 (N_37440,N_35673,N_34777);
xor U37441 (N_37441,N_35238,N_35196);
or U37442 (N_37442,N_35387,N_34961);
xnor U37443 (N_37443,N_34645,N_34673);
nor U37444 (N_37444,N_34044,N_34393);
nor U37445 (N_37445,N_34667,N_35629);
nor U37446 (N_37446,N_34401,N_35326);
nand U37447 (N_37447,N_34356,N_35317);
nor U37448 (N_37448,N_35810,N_34332);
or U37449 (N_37449,N_35359,N_34580);
nand U37450 (N_37450,N_35185,N_34007);
and U37451 (N_37451,N_35869,N_34050);
or U37452 (N_37452,N_35233,N_34558);
xnor U37453 (N_37453,N_34568,N_35911);
xor U37454 (N_37454,N_34596,N_35265);
xor U37455 (N_37455,N_35161,N_34792);
nor U37456 (N_37456,N_35306,N_35623);
xor U37457 (N_37457,N_35759,N_35555);
xnor U37458 (N_37458,N_34949,N_34105);
nor U37459 (N_37459,N_35855,N_34464);
nand U37460 (N_37460,N_35731,N_35077);
xor U37461 (N_37461,N_35104,N_34097);
or U37462 (N_37462,N_34058,N_35330);
nor U37463 (N_37463,N_34999,N_34069);
or U37464 (N_37464,N_35854,N_34364);
xnor U37465 (N_37465,N_34187,N_35486);
or U37466 (N_37466,N_34177,N_35619);
nor U37467 (N_37467,N_35506,N_35980);
and U37468 (N_37468,N_34487,N_34474);
and U37469 (N_37469,N_34040,N_34866);
nand U37470 (N_37470,N_34950,N_34298);
and U37471 (N_37471,N_35773,N_35626);
or U37472 (N_37472,N_35038,N_34744);
and U37473 (N_37473,N_35839,N_35210);
xor U37474 (N_37474,N_35599,N_35138);
and U37475 (N_37475,N_35421,N_34662);
nor U37476 (N_37476,N_35026,N_35318);
and U37477 (N_37477,N_35132,N_35032);
and U37478 (N_37478,N_34189,N_34436);
or U37479 (N_37479,N_35419,N_34037);
nor U37480 (N_37480,N_35976,N_34347);
and U37481 (N_37481,N_35205,N_34308);
nor U37482 (N_37482,N_34765,N_34629);
or U37483 (N_37483,N_34587,N_35124);
nor U37484 (N_37484,N_35692,N_34921);
and U37485 (N_37485,N_35193,N_34299);
nor U37486 (N_37486,N_35045,N_35841);
nor U37487 (N_37487,N_35585,N_34069);
xor U37488 (N_37488,N_35543,N_35570);
or U37489 (N_37489,N_34067,N_34823);
nand U37490 (N_37490,N_35343,N_35918);
or U37491 (N_37491,N_34944,N_34233);
xnor U37492 (N_37492,N_34865,N_34964);
xnor U37493 (N_37493,N_34988,N_34878);
nor U37494 (N_37494,N_34750,N_34082);
xor U37495 (N_37495,N_35437,N_34167);
nand U37496 (N_37496,N_35166,N_34891);
and U37497 (N_37497,N_34490,N_35879);
and U37498 (N_37498,N_34284,N_34136);
nand U37499 (N_37499,N_35097,N_35859);
nor U37500 (N_37500,N_34258,N_34075);
and U37501 (N_37501,N_35909,N_34505);
and U37502 (N_37502,N_35608,N_35890);
xnor U37503 (N_37503,N_35367,N_35424);
and U37504 (N_37504,N_34576,N_35669);
nand U37505 (N_37505,N_35868,N_35507);
nor U37506 (N_37506,N_34828,N_34354);
or U37507 (N_37507,N_34999,N_34122);
xnor U37508 (N_37508,N_34763,N_34017);
or U37509 (N_37509,N_35381,N_35542);
and U37510 (N_37510,N_35865,N_35881);
nand U37511 (N_37511,N_34704,N_35329);
nor U37512 (N_37512,N_34728,N_35744);
nor U37513 (N_37513,N_34375,N_35307);
nor U37514 (N_37514,N_35288,N_35652);
nor U37515 (N_37515,N_34425,N_35368);
and U37516 (N_37516,N_35428,N_34700);
nor U37517 (N_37517,N_35336,N_34557);
and U37518 (N_37518,N_35231,N_34472);
or U37519 (N_37519,N_34412,N_35985);
xnor U37520 (N_37520,N_34044,N_34928);
nor U37521 (N_37521,N_35207,N_35427);
nand U37522 (N_37522,N_34337,N_34208);
nor U37523 (N_37523,N_34038,N_34303);
or U37524 (N_37524,N_34949,N_35249);
nor U37525 (N_37525,N_35361,N_34295);
nand U37526 (N_37526,N_35588,N_35292);
xnor U37527 (N_37527,N_35261,N_35035);
xnor U37528 (N_37528,N_34284,N_35674);
and U37529 (N_37529,N_34514,N_35387);
xnor U37530 (N_37530,N_34518,N_34861);
or U37531 (N_37531,N_34993,N_34907);
xnor U37532 (N_37532,N_35405,N_35846);
or U37533 (N_37533,N_34265,N_34767);
or U37534 (N_37534,N_34503,N_35552);
or U37535 (N_37535,N_34036,N_35195);
and U37536 (N_37536,N_35940,N_34007);
or U37537 (N_37537,N_34577,N_34203);
nand U37538 (N_37538,N_35891,N_35650);
xor U37539 (N_37539,N_35322,N_35692);
xor U37540 (N_37540,N_35428,N_34192);
nand U37541 (N_37541,N_35381,N_34705);
nor U37542 (N_37542,N_35789,N_34643);
and U37543 (N_37543,N_35860,N_34730);
nand U37544 (N_37544,N_34627,N_34578);
or U37545 (N_37545,N_35985,N_34001);
or U37546 (N_37546,N_34032,N_34518);
nor U37547 (N_37547,N_35832,N_34347);
or U37548 (N_37548,N_34158,N_34619);
and U37549 (N_37549,N_35949,N_35276);
and U37550 (N_37550,N_35667,N_35771);
nor U37551 (N_37551,N_34459,N_34519);
xnor U37552 (N_37552,N_35498,N_34289);
nor U37553 (N_37553,N_35907,N_35023);
or U37554 (N_37554,N_34943,N_35454);
xnor U37555 (N_37555,N_35320,N_34905);
nand U37556 (N_37556,N_35759,N_35901);
nor U37557 (N_37557,N_35052,N_35105);
nor U37558 (N_37558,N_34899,N_34560);
xnor U37559 (N_37559,N_34961,N_34397);
and U37560 (N_37560,N_34010,N_35776);
nand U37561 (N_37561,N_35302,N_35855);
xnor U37562 (N_37562,N_34132,N_34533);
and U37563 (N_37563,N_34708,N_34521);
xnor U37564 (N_37564,N_35930,N_34917);
or U37565 (N_37565,N_35648,N_35884);
nor U37566 (N_37566,N_35909,N_35361);
nor U37567 (N_37567,N_34545,N_35856);
and U37568 (N_37568,N_35868,N_35125);
or U37569 (N_37569,N_34290,N_35724);
nand U37570 (N_37570,N_35648,N_34752);
nor U37571 (N_37571,N_34764,N_35800);
or U37572 (N_37572,N_34209,N_34754);
and U37573 (N_37573,N_35848,N_34402);
and U37574 (N_37574,N_35412,N_35687);
and U37575 (N_37575,N_34809,N_34228);
or U37576 (N_37576,N_35174,N_34911);
or U37577 (N_37577,N_35230,N_34494);
or U37578 (N_37578,N_35276,N_35340);
nor U37579 (N_37579,N_35176,N_34112);
and U37580 (N_37580,N_35078,N_34642);
nand U37581 (N_37581,N_35473,N_34885);
or U37582 (N_37582,N_35617,N_34937);
or U37583 (N_37583,N_34758,N_34870);
or U37584 (N_37584,N_34730,N_35630);
xnor U37585 (N_37585,N_35602,N_34287);
and U37586 (N_37586,N_35663,N_34325);
nor U37587 (N_37587,N_34352,N_35176);
nand U37588 (N_37588,N_34812,N_35275);
nor U37589 (N_37589,N_35786,N_35524);
nand U37590 (N_37590,N_35500,N_35012);
and U37591 (N_37591,N_34171,N_34507);
nor U37592 (N_37592,N_35332,N_34232);
and U37593 (N_37593,N_34721,N_34801);
nand U37594 (N_37594,N_35898,N_34931);
and U37595 (N_37595,N_35105,N_34438);
or U37596 (N_37596,N_35926,N_35305);
nor U37597 (N_37597,N_35007,N_34402);
nor U37598 (N_37598,N_35460,N_35359);
or U37599 (N_37599,N_34340,N_34034);
xnor U37600 (N_37600,N_35143,N_34802);
xnor U37601 (N_37601,N_35212,N_35266);
nand U37602 (N_37602,N_34183,N_34597);
xor U37603 (N_37603,N_34096,N_34674);
nand U37604 (N_37604,N_34273,N_35088);
or U37605 (N_37605,N_35056,N_35695);
xnor U37606 (N_37606,N_35354,N_35088);
xor U37607 (N_37607,N_34703,N_35574);
xnor U37608 (N_37608,N_35253,N_34850);
xor U37609 (N_37609,N_34035,N_34613);
xnor U37610 (N_37610,N_35887,N_34241);
nor U37611 (N_37611,N_35015,N_35551);
xor U37612 (N_37612,N_34218,N_34404);
xnor U37613 (N_37613,N_34774,N_34376);
and U37614 (N_37614,N_34464,N_35666);
xor U37615 (N_37615,N_34746,N_35534);
and U37616 (N_37616,N_34733,N_35015);
nor U37617 (N_37617,N_34252,N_34145);
and U37618 (N_37618,N_35542,N_35938);
and U37619 (N_37619,N_34321,N_35454);
or U37620 (N_37620,N_35797,N_34665);
and U37621 (N_37621,N_34160,N_34845);
xnor U37622 (N_37622,N_34870,N_35775);
nor U37623 (N_37623,N_34019,N_34040);
or U37624 (N_37624,N_34337,N_34853);
nand U37625 (N_37625,N_34498,N_35263);
xor U37626 (N_37626,N_34971,N_35170);
nand U37627 (N_37627,N_35924,N_35796);
nand U37628 (N_37628,N_34558,N_35429);
and U37629 (N_37629,N_34819,N_34285);
or U37630 (N_37630,N_34720,N_34300);
nand U37631 (N_37631,N_35814,N_34044);
or U37632 (N_37632,N_34665,N_35653);
nand U37633 (N_37633,N_35810,N_34783);
or U37634 (N_37634,N_35238,N_35083);
and U37635 (N_37635,N_34200,N_34689);
or U37636 (N_37636,N_34909,N_35488);
and U37637 (N_37637,N_34097,N_34969);
xor U37638 (N_37638,N_35109,N_34117);
xor U37639 (N_37639,N_34172,N_34803);
nor U37640 (N_37640,N_34607,N_34135);
nor U37641 (N_37641,N_35081,N_34423);
xnor U37642 (N_37642,N_34797,N_35108);
and U37643 (N_37643,N_34462,N_34899);
or U37644 (N_37644,N_34474,N_35970);
and U37645 (N_37645,N_35674,N_35488);
nand U37646 (N_37646,N_35257,N_34290);
nor U37647 (N_37647,N_35598,N_34607);
nand U37648 (N_37648,N_34847,N_34977);
or U37649 (N_37649,N_34768,N_34631);
nand U37650 (N_37650,N_34210,N_35280);
nor U37651 (N_37651,N_34216,N_34432);
or U37652 (N_37652,N_34594,N_35373);
and U37653 (N_37653,N_35746,N_35305);
xnor U37654 (N_37654,N_34303,N_35466);
and U37655 (N_37655,N_35289,N_35139);
or U37656 (N_37656,N_35995,N_34289);
and U37657 (N_37657,N_35811,N_34279);
xor U37658 (N_37658,N_34715,N_34564);
nand U37659 (N_37659,N_35631,N_34159);
xor U37660 (N_37660,N_35256,N_35439);
or U37661 (N_37661,N_35581,N_35451);
nand U37662 (N_37662,N_34478,N_35856);
nand U37663 (N_37663,N_35127,N_34281);
xnor U37664 (N_37664,N_35580,N_34698);
and U37665 (N_37665,N_35730,N_34362);
and U37666 (N_37666,N_35317,N_34842);
or U37667 (N_37667,N_34892,N_34667);
nor U37668 (N_37668,N_34204,N_34392);
xnor U37669 (N_37669,N_34002,N_34020);
or U37670 (N_37670,N_34221,N_35088);
nor U37671 (N_37671,N_35181,N_35401);
nor U37672 (N_37672,N_34276,N_34269);
nand U37673 (N_37673,N_35979,N_35257);
or U37674 (N_37674,N_34268,N_34925);
xor U37675 (N_37675,N_35711,N_35117);
and U37676 (N_37676,N_34263,N_34223);
nor U37677 (N_37677,N_35335,N_34585);
xnor U37678 (N_37678,N_34583,N_34431);
or U37679 (N_37679,N_35500,N_35862);
nor U37680 (N_37680,N_35951,N_35966);
xor U37681 (N_37681,N_35418,N_34278);
nor U37682 (N_37682,N_34117,N_34752);
and U37683 (N_37683,N_35748,N_35685);
xnor U37684 (N_37684,N_35593,N_35072);
nor U37685 (N_37685,N_34525,N_35159);
xor U37686 (N_37686,N_34647,N_35842);
and U37687 (N_37687,N_34111,N_34911);
nor U37688 (N_37688,N_35267,N_35247);
nor U37689 (N_37689,N_34554,N_34917);
and U37690 (N_37690,N_34178,N_35944);
nand U37691 (N_37691,N_35781,N_35772);
and U37692 (N_37692,N_34029,N_34096);
xor U37693 (N_37693,N_34761,N_35414);
or U37694 (N_37694,N_34985,N_34675);
or U37695 (N_37695,N_35763,N_35902);
or U37696 (N_37696,N_35714,N_34703);
and U37697 (N_37697,N_34898,N_35894);
nor U37698 (N_37698,N_35317,N_35058);
and U37699 (N_37699,N_35849,N_34612);
nor U37700 (N_37700,N_34093,N_34948);
xor U37701 (N_37701,N_35502,N_35674);
and U37702 (N_37702,N_34715,N_35681);
or U37703 (N_37703,N_35229,N_35621);
or U37704 (N_37704,N_34548,N_34048);
or U37705 (N_37705,N_34770,N_35251);
or U37706 (N_37706,N_35618,N_34761);
xnor U37707 (N_37707,N_34263,N_34783);
and U37708 (N_37708,N_34863,N_34946);
and U37709 (N_37709,N_35728,N_34852);
or U37710 (N_37710,N_34786,N_34899);
and U37711 (N_37711,N_34665,N_34830);
xnor U37712 (N_37712,N_35845,N_35170);
xnor U37713 (N_37713,N_34858,N_34412);
or U37714 (N_37714,N_34036,N_35621);
nand U37715 (N_37715,N_35514,N_35664);
and U37716 (N_37716,N_34483,N_34114);
nand U37717 (N_37717,N_35900,N_34160);
or U37718 (N_37718,N_34304,N_34111);
xor U37719 (N_37719,N_35687,N_34742);
or U37720 (N_37720,N_34224,N_35504);
or U37721 (N_37721,N_34718,N_35173);
and U37722 (N_37722,N_34410,N_34898);
nand U37723 (N_37723,N_34332,N_35672);
or U37724 (N_37724,N_34094,N_34570);
xor U37725 (N_37725,N_35028,N_34830);
nor U37726 (N_37726,N_35187,N_35679);
nand U37727 (N_37727,N_35253,N_34158);
nand U37728 (N_37728,N_34005,N_35919);
xor U37729 (N_37729,N_34872,N_35173);
nand U37730 (N_37730,N_35266,N_35836);
nor U37731 (N_37731,N_35194,N_35107);
and U37732 (N_37732,N_34837,N_35668);
nand U37733 (N_37733,N_35679,N_35400);
nor U37734 (N_37734,N_34450,N_34201);
nand U37735 (N_37735,N_34674,N_35878);
xor U37736 (N_37736,N_35793,N_34145);
nor U37737 (N_37737,N_34564,N_35206);
nand U37738 (N_37738,N_34674,N_35884);
nor U37739 (N_37739,N_35473,N_34095);
and U37740 (N_37740,N_35237,N_34760);
xor U37741 (N_37741,N_35025,N_34015);
and U37742 (N_37742,N_34524,N_34239);
xor U37743 (N_37743,N_35156,N_34183);
nand U37744 (N_37744,N_34066,N_35584);
xnor U37745 (N_37745,N_35755,N_35476);
or U37746 (N_37746,N_34864,N_34165);
and U37747 (N_37747,N_35131,N_34194);
or U37748 (N_37748,N_34425,N_34621);
or U37749 (N_37749,N_35667,N_35576);
nand U37750 (N_37750,N_35633,N_34211);
or U37751 (N_37751,N_34703,N_34212);
or U37752 (N_37752,N_35839,N_35149);
nand U37753 (N_37753,N_35588,N_35394);
or U37754 (N_37754,N_34851,N_35203);
and U37755 (N_37755,N_35000,N_35491);
or U37756 (N_37756,N_35459,N_34686);
or U37757 (N_37757,N_34093,N_35065);
and U37758 (N_37758,N_35815,N_35399);
nand U37759 (N_37759,N_35649,N_34177);
or U37760 (N_37760,N_35518,N_34582);
or U37761 (N_37761,N_34954,N_34894);
and U37762 (N_37762,N_35970,N_34327);
nand U37763 (N_37763,N_34567,N_35322);
xnor U37764 (N_37764,N_35251,N_35618);
and U37765 (N_37765,N_34530,N_35745);
xor U37766 (N_37766,N_35486,N_34293);
or U37767 (N_37767,N_34518,N_34189);
xor U37768 (N_37768,N_34237,N_34727);
xor U37769 (N_37769,N_34293,N_34905);
and U37770 (N_37770,N_34926,N_34240);
nor U37771 (N_37771,N_35853,N_34724);
nand U37772 (N_37772,N_35665,N_35662);
and U37773 (N_37773,N_35856,N_35771);
and U37774 (N_37774,N_34429,N_35213);
nand U37775 (N_37775,N_35195,N_35135);
nand U37776 (N_37776,N_34856,N_34641);
and U37777 (N_37777,N_34488,N_35387);
nand U37778 (N_37778,N_35103,N_35360);
nand U37779 (N_37779,N_35984,N_35380);
nand U37780 (N_37780,N_35631,N_34493);
nor U37781 (N_37781,N_35749,N_35511);
or U37782 (N_37782,N_35106,N_34059);
xor U37783 (N_37783,N_35498,N_35863);
nor U37784 (N_37784,N_34684,N_34286);
or U37785 (N_37785,N_35985,N_35478);
nor U37786 (N_37786,N_35689,N_35626);
and U37787 (N_37787,N_34408,N_34959);
nand U37788 (N_37788,N_35267,N_34976);
xnor U37789 (N_37789,N_34042,N_35233);
nor U37790 (N_37790,N_35319,N_35185);
and U37791 (N_37791,N_34826,N_35140);
and U37792 (N_37792,N_34970,N_35818);
or U37793 (N_37793,N_34724,N_34057);
and U37794 (N_37794,N_35000,N_35186);
nor U37795 (N_37795,N_35410,N_35647);
or U37796 (N_37796,N_34570,N_35794);
xor U37797 (N_37797,N_34717,N_35350);
and U37798 (N_37798,N_34003,N_34598);
and U37799 (N_37799,N_35453,N_35165);
xor U37800 (N_37800,N_35035,N_35198);
and U37801 (N_37801,N_35686,N_34925);
nor U37802 (N_37802,N_35261,N_34850);
and U37803 (N_37803,N_35012,N_34547);
nand U37804 (N_37804,N_34321,N_35675);
or U37805 (N_37805,N_35806,N_34668);
nand U37806 (N_37806,N_34707,N_35644);
and U37807 (N_37807,N_35125,N_35701);
and U37808 (N_37808,N_35836,N_35314);
nor U37809 (N_37809,N_35472,N_35353);
xnor U37810 (N_37810,N_34874,N_34415);
nor U37811 (N_37811,N_34220,N_35919);
xor U37812 (N_37812,N_34377,N_34406);
and U37813 (N_37813,N_34999,N_35458);
and U37814 (N_37814,N_35029,N_34475);
nand U37815 (N_37815,N_34180,N_34910);
and U37816 (N_37816,N_34744,N_34284);
or U37817 (N_37817,N_35398,N_34036);
nor U37818 (N_37818,N_34673,N_35297);
or U37819 (N_37819,N_34852,N_34306);
nand U37820 (N_37820,N_35671,N_34699);
nand U37821 (N_37821,N_34250,N_34954);
nand U37822 (N_37822,N_34519,N_35873);
nor U37823 (N_37823,N_35672,N_34979);
xor U37824 (N_37824,N_35827,N_35673);
or U37825 (N_37825,N_34686,N_34579);
or U37826 (N_37826,N_34491,N_34196);
and U37827 (N_37827,N_34330,N_34941);
and U37828 (N_37828,N_35772,N_35245);
and U37829 (N_37829,N_35369,N_34935);
xor U37830 (N_37830,N_35849,N_34232);
and U37831 (N_37831,N_34319,N_34734);
or U37832 (N_37832,N_34893,N_35188);
nand U37833 (N_37833,N_34306,N_35364);
or U37834 (N_37834,N_35462,N_35844);
nor U37835 (N_37835,N_35182,N_34156);
xnor U37836 (N_37836,N_34122,N_34550);
nor U37837 (N_37837,N_34844,N_35969);
or U37838 (N_37838,N_35794,N_35387);
nor U37839 (N_37839,N_34922,N_35568);
nor U37840 (N_37840,N_34830,N_34863);
xor U37841 (N_37841,N_34499,N_35408);
and U37842 (N_37842,N_34976,N_34568);
nand U37843 (N_37843,N_34577,N_34913);
nand U37844 (N_37844,N_35056,N_35059);
or U37845 (N_37845,N_35073,N_35324);
nand U37846 (N_37846,N_34832,N_35280);
or U37847 (N_37847,N_35177,N_34763);
nand U37848 (N_37848,N_34609,N_35561);
and U37849 (N_37849,N_34060,N_34776);
xor U37850 (N_37850,N_35916,N_35731);
nor U37851 (N_37851,N_34624,N_34675);
nand U37852 (N_37852,N_34512,N_34636);
xor U37853 (N_37853,N_35993,N_35930);
and U37854 (N_37854,N_35921,N_35561);
xnor U37855 (N_37855,N_34159,N_35055);
xor U37856 (N_37856,N_35558,N_34456);
and U37857 (N_37857,N_35917,N_35093);
xnor U37858 (N_37858,N_34075,N_35629);
xnor U37859 (N_37859,N_34648,N_35938);
nand U37860 (N_37860,N_34440,N_34210);
nor U37861 (N_37861,N_34512,N_35931);
xnor U37862 (N_37862,N_34748,N_34642);
and U37863 (N_37863,N_34314,N_34207);
and U37864 (N_37864,N_34165,N_34485);
xnor U37865 (N_37865,N_34100,N_34150);
or U37866 (N_37866,N_34701,N_34765);
nor U37867 (N_37867,N_34523,N_35046);
nor U37868 (N_37868,N_34793,N_35550);
or U37869 (N_37869,N_35967,N_35570);
nand U37870 (N_37870,N_34116,N_35006);
and U37871 (N_37871,N_35080,N_35078);
and U37872 (N_37872,N_34222,N_35990);
xnor U37873 (N_37873,N_34738,N_34551);
or U37874 (N_37874,N_35958,N_34473);
nor U37875 (N_37875,N_34619,N_34437);
nor U37876 (N_37876,N_35834,N_34644);
or U37877 (N_37877,N_34123,N_35644);
nand U37878 (N_37878,N_34162,N_35681);
nand U37879 (N_37879,N_35372,N_34012);
nand U37880 (N_37880,N_34836,N_35441);
and U37881 (N_37881,N_35549,N_34477);
nor U37882 (N_37882,N_35776,N_35127);
xnor U37883 (N_37883,N_34587,N_34022);
and U37884 (N_37884,N_35157,N_35952);
or U37885 (N_37885,N_34840,N_35235);
or U37886 (N_37886,N_34634,N_35172);
nor U37887 (N_37887,N_35142,N_34664);
and U37888 (N_37888,N_34809,N_34336);
and U37889 (N_37889,N_35409,N_34663);
xor U37890 (N_37890,N_35454,N_35675);
xnor U37891 (N_37891,N_35628,N_34567);
and U37892 (N_37892,N_35966,N_34225);
nand U37893 (N_37893,N_34120,N_34102);
and U37894 (N_37894,N_34325,N_34210);
and U37895 (N_37895,N_35458,N_35285);
xnor U37896 (N_37896,N_34027,N_35230);
nand U37897 (N_37897,N_35221,N_35299);
xnor U37898 (N_37898,N_34283,N_35525);
nor U37899 (N_37899,N_35534,N_34399);
xor U37900 (N_37900,N_34283,N_35313);
nand U37901 (N_37901,N_35601,N_35595);
or U37902 (N_37902,N_34416,N_35049);
xor U37903 (N_37903,N_34021,N_34673);
and U37904 (N_37904,N_34820,N_34439);
and U37905 (N_37905,N_34364,N_35226);
and U37906 (N_37906,N_35940,N_34457);
or U37907 (N_37907,N_35568,N_34464);
nor U37908 (N_37908,N_35316,N_35340);
and U37909 (N_37909,N_35119,N_35542);
and U37910 (N_37910,N_35744,N_35801);
xnor U37911 (N_37911,N_35866,N_35132);
xnor U37912 (N_37912,N_34098,N_35708);
or U37913 (N_37913,N_35111,N_34216);
xor U37914 (N_37914,N_34428,N_34111);
or U37915 (N_37915,N_35284,N_34270);
xnor U37916 (N_37916,N_35899,N_34759);
xnor U37917 (N_37917,N_34043,N_34087);
xnor U37918 (N_37918,N_34154,N_35501);
xnor U37919 (N_37919,N_34536,N_34815);
or U37920 (N_37920,N_35167,N_34013);
or U37921 (N_37921,N_34861,N_35437);
nor U37922 (N_37922,N_35592,N_35682);
nor U37923 (N_37923,N_34133,N_35644);
nand U37924 (N_37924,N_34940,N_34789);
xor U37925 (N_37925,N_34114,N_35043);
or U37926 (N_37926,N_34216,N_35328);
nand U37927 (N_37927,N_35968,N_35542);
and U37928 (N_37928,N_34704,N_34358);
xnor U37929 (N_37929,N_34483,N_35608);
or U37930 (N_37930,N_34895,N_34192);
or U37931 (N_37931,N_35361,N_35665);
and U37932 (N_37932,N_34641,N_34538);
nor U37933 (N_37933,N_35203,N_35202);
or U37934 (N_37934,N_35586,N_35912);
nand U37935 (N_37935,N_35067,N_34875);
and U37936 (N_37936,N_34659,N_35139);
nand U37937 (N_37937,N_34294,N_34164);
nand U37938 (N_37938,N_35292,N_34360);
and U37939 (N_37939,N_34514,N_35337);
and U37940 (N_37940,N_35221,N_34856);
nand U37941 (N_37941,N_35255,N_34335);
nor U37942 (N_37942,N_34661,N_35051);
and U37943 (N_37943,N_35361,N_35424);
nor U37944 (N_37944,N_34715,N_35241);
or U37945 (N_37945,N_35615,N_34594);
nor U37946 (N_37946,N_34105,N_34861);
xnor U37947 (N_37947,N_34765,N_35669);
or U37948 (N_37948,N_35144,N_34237);
nand U37949 (N_37949,N_34224,N_35487);
xnor U37950 (N_37950,N_35207,N_35247);
or U37951 (N_37951,N_35761,N_35682);
xor U37952 (N_37952,N_35057,N_35406);
or U37953 (N_37953,N_35207,N_35618);
or U37954 (N_37954,N_34177,N_34594);
xor U37955 (N_37955,N_35197,N_34605);
or U37956 (N_37956,N_34961,N_34005);
nand U37957 (N_37957,N_34461,N_35638);
xnor U37958 (N_37958,N_34667,N_34512);
and U37959 (N_37959,N_35216,N_35122);
and U37960 (N_37960,N_34838,N_35369);
nor U37961 (N_37961,N_35953,N_34437);
nand U37962 (N_37962,N_34097,N_34201);
or U37963 (N_37963,N_34398,N_34554);
xnor U37964 (N_37964,N_35250,N_34054);
nor U37965 (N_37965,N_34377,N_35718);
nand U37966 (N_37966,N_34307,N_34108);
or U37967 (N_37967,N_35460,N_35195);
nand U37968 (N_37968,N_35686,N_35595);
xnor U37969 (N_37969,N_34683,N_34762);
or U37970 (N_37970,N_35466,N_34396);
xnor U37971 (N_37971,N_35911,N_34484);
xnor U37972 (N_37972,N_34624,N_35858);
xnor U37973 (N_37973,N_35406,N_35226);
or U37974 (N_37974,N_35206,N_34147);
nor U37975 (N_37975,N_35514,N_35851);
xor U37976 (N_37976,N_34001,N_34542);
and U37977 (N_37977,N_34299,N_34747);
and U37978 (N_37978,N_35742,N_35279);
or U37979 (N_37979,N_34870,N_35051);
nand U37980 (N_37980,N_35714,N_35773);
nor U37981 (N_37981,N_35540,N_35613);
nor U37982 (N_37982,N_34133,N_35036);
and U37983 (N_37983,N_34603,N_35636);
xnor U37984 (N_37984,N_34975,N_34506);
nor U37985 (N_37985,N_34930,N_35699);
nand U37986 (N_37986,N_35398,N_35469);
xor U37987 (N_37987,N_34236,N_35327);
xor U37988 (N_37988,N_35536,N_34072);
and U37989 (N_37989,N_35853,N_35288);
and U37990 (N_37990,N_34971,N_34181);
xor U37991 (N_37991,N_34897,N_35576);
or U37992 (N_37992,N_35372,N_34005);
or U37993 (N_37993,N_34652,N_35357);
and U37994 (N_37994,N_35538,N_35026);
and U37995 (N_37995,N_34124,N_35759);
nor U37996 (N_37996,N_34183,N_35297);
nor U37997 (N_37997,N_35138,N_35224);
and U37998 (N_37998,N_34127,N_35532);
and U37999 (N_37999,N_34034,N_34554);
and U38000 (N_38000,N_37453,N_36550);
nand U38001 (N_38001,N_36686,N_36857);
and U38002 (N_38002,N_37665,N_37197);
xor U38003 (N_38003,N_36592,N_37915);
nor U38004 (N_38004,N_36246,N_37846);
or U38005 (N_38005,N_37299,N_36090);
and U38006 (N_38006,N_36134,N_36158);
nand U38007 (N_38007,N_36718,N_37536);
or U38008 (N_38008,N_36285,N_36093);
xor U38009 (N_38009,N_36363,N_36122);
xnor U38010 (N_38010,N_36851,N_37270);
nand U38011 (N_38011,N_37708,N_37007);
xor U38012 (N_38012,N_37698,N_37702);
or U38013 (N_38013,N_36775,N_36971);
nor U38014 (N_38014,N_37126,N_36199);
nand U38015 (N_38015,N_36482,N_37511);
nand U38016 (N_38016,N_36229,N_37857);
xnor U38017 (N_38017,N_37988,N_36140);
nand U38018 (N_38018,N_36888,N_36548);
xor U38019 (N_38019,N_36964,N_36803);
nor U38020 (N_38020,N_36405,N_37479);
xnor U38021 (N_38021,N_36388,N_36476);
nor U38022 (N_38022,N_36515,N_37165);
or U38023 (N_38023,N_36856,N_37827);
xor U38024 (N_38024,N_37447,N_37110);
xor U38025 (N_38025,N_37184,N_36316);
nand U38026 (N_38026,N_36027,N_36977);
or U38027 (N_38027,N_37381,N_36207);
nand U38028 (N_38028,N_36690,N_36738);
nand U38029 (N_38029,N_36596,N_37374);
nand U38030 (N_38030,N_36133,N_36214);
nand U38031 (N_38031,N_37085,N_36160);
and U38032 (N_38032,N_36120,N_37121);
nand U38033 (N_38033,N_37163,N_36716);
xnor U38034 (N_38034,N_37474,N_36731);
or U38035 (N_38035,N_36391,N_37866);
or U38036 (N_38036,N_36469,N_37319);
or U38037 (N_38037,N_37445,N_36322);
or U38038 (N_38038,N_37981,N_37002);
and U38039 (N_38039,N_36887,N_36142);
or U38040 (N_38040,N_37816,N_37397);
and U38041 (N_38041,N_37441,N_36944);
and U38042 (N_38042,N_36098,N_36565);
and U38043 (N_38043,N_36268,N_36830);
nand U38044 (N_38044,N_36138,N_37063);
or U38045 (N_38045,N_37781,N_37191);
and U38046 (N_38046,N_37854,N_36306);
or U38047 (N_38047,N_37567,N_36232);
and U38048 (N_38048,N_37412,N_36751);
xnor U38049 (N_38049,N_36466,N_37368);
xor U38050 (N_38050,N_37924,N_36886);
nor U38051 (N_38051,N_37001,N_37093);
xor U38052 (N_38052,N_37830,N_37545);
or U38053 (N_38053,N_36968,N_37304);
nor U38054 (N_38054,N_36769,N_36038);
or U38055 (N_38055,N_37497,N_36916);
nor U38056 (N_38056,N_37973,N_37751);
xnor U38057 (N_38057,N_36849,N_37463);
and U38058 (N_38058,N_36075,N_37181);
and U38059 (N_38059,N_37073,N_37354);
nand U38060 (N_38060,N_36054,N_36556);
and U38061 (N_38061,N_36959,N_37882);
nor U38062 (N_38062,N_36763,N_37573);
nor U38063 (N_38063,N_36957,N_37175);
and U38064 (N_38064,N_37097,N_37625);
or U38065 (N_38065,N_37145,N_36777);
xor U38066 (N_38066,N_36181,N_36765);
nand U38067 (N_38067,N_37266,N_36156);
nor U38068 (N_38068,N_37752,N_36371);
nand U38069 (N_38069,N_36096,N_37054);
xor U38070 (N_38070,N_37638,N_36904);
xor U38071 (N_38071,N_36774,N_37729);
nor U38072 (N_38072,N_37208,N_36755);
or U38073 (N_38073,N_37053,N_37860);
nor U38074 (N_38074,N_37903,N_37513);
and U38075 (N_38075,N_36875,N_37837);
nand U38076 (N_38076,N_37190,N_37488);
and U38077 (N_38077,N_37456,N_37839);
nor U38078 (N_38078,N_37321,N_37808);
nand U38079 (N_38079,N_37489,N_36077);
or U38080 (N_38080,N_37433,N_37177);
nand U38081 (N_38081,N_37146,N_36000);
or U38082 (N_38082,N_36015,N_37749);
or U38083 (N_38083,N_37164,N_37541);
or U38084 (N_38084,N_37448,N_37894);
xnor U38085 (N_38085,N_37438,N_36304);
xor U38086 (N_38086,N_36416,N_36983);
nand U38087 (N_38087,N_37595,N_36240);
nor U38088 (N_38088,N_37458,N_37239);
nor U38089 (N_38089,N_36114,N_36662);
and U38090 (N_38090,N_37080,N_36705);
or U38091 (N_38091,N_36128,N_37522);
xor U38092 (N_38092,N_37500,N_36118);
and U38093 (N_38093,N_36585,N_36664);
and U38094 (N_38094,N_37652,N_36242);
nor U38095 (N_38095,N_37057,N_37783);
nand U38096 (N_38096,N_36127,N_36056);
nand U38097 (N_38097,N_36935,N_37921);
and U38098 (N_38098,N_37566,N_37661);
nor U38099 (N_38099,N_37312,N_37284);
or U38100 (N_38100,N_36193,N_37858);
nor U38101 (N_38101,N_37020,N_37634);
and U38102 (N_38102,N_36897,N_37821);
nand U38103 (N_38103,N_37796,N_37482);
and U38104 (N_38104,N_36921,N_37991);
nor U38105 (N_38105,N_36280,N_37167);
xnor U38106 (N_38106,N_37280,N_37640);
nor U38107 (N_38107,N_36829,N_37809);
nor U38108 (N_38108,N_36922,N_36668);
nand U38109 (N_38109,N_36725,N_36636);
and U38110 (N_38110,N_36091,N_37913);
or U38111 (N_38111,N_37591,N_36761);
nand U38112 (N_38112,N_37834,N_37731);
nand U38113 (N_38113,N_36745,N_37738);
nand U38114 (N_38114,N_37597,N_36337);
xnor U38115 (N_38115,N_36454,N_36694);
nor U38116 (N_38116,N_37631,N_37250);
xor U38117 (N_38117,N_36043,N_36167);
xnor U38118 (N_38118,N_36575,N_36237);
nand U38119 (N_38119,N_36177,N_37570);
nand U38120 (N_38120,N_37347,N_37688);
nand U38121 (N_38121,N_36559,N_36828);
nor U38122 (N_38122,N_36419,N_36562);
or U38123 (N_38123,N_36825,N_36872);
nor U38124 (N_38124,N_37272,N_36221);
or U38125 (N_38125,N_36960,N_37606);
and U38126 (N_38126,N_37125,N_37389);
xnor U38127 (N_38127,N_36679,N_36894);
nor U38128 (N_38128,N_36182,N_37530);
or U38129 (N_38129,N_36506,N_36442);
nor U38130 (N_38130,N_36135,N_36014);
nand U38131 (N_38131,N_37695,N_36370);
or U38132 (N_38132,N_37826,N_37629);
or U38133 (N_38133,N_36447,N_36528);
nor U38134 (N_38134,N_36607,N_37247);
nor U38135 (N_38135,N_37955,N_36555);
and U38136 (N_38136,N_36748,N_36511);
nor U38137 (N_38137,N_36892,N_37743);
and U38138 (N_38138,N_37544,N_36995);
nor U38139 (N_38139,N_37758,N_37253);
xor U38140 (N_38140,N_36846,N_37432);
nor U38141 (N_38141,N_36800,N_37475);
nand U38142 (N_38142,N_36588,N_36009);
xnor U38143 (N_38143,N_36433,N_36319);
nand U38144 (N_38144,N_36527,N_37446);
xnor U38145 (N_38145,N_37295,N_37976);
xnor U38146 (N_38146,N_36450,N_36670);
and U38147 (N_38147,N_37936,N_36954);
and U38148 (N_38148,N_37192,N_37531);
nand U38149 (N_38149,N_36987,N_36005);
or U38150 (N_38150,N_36839,N_36247);
and U38151 (N_38151,N_37710,N_37185);
nand U38152 (N_38152,N_36196,N_37082);
xnor U38153 (N_38153,N_36248,N_37604);
and U38154 (N_38154,N_36730,N_36976);
nor U38155 (N_38155,N_37491,N_36378);
or U38156 (N_38156,N_36064,N_37733);
and U38157 (N_38157,N_37139,N_37662);
and U38158 (N_38158,N_36513,N_36833);
xnor U38159 (N_38159,N_37217,N_36552);
nand U38160 (N_38160,N_36991,N_37717);
nand U38161 (N_38161,N_36162,N_36947);
nor U38162 (N_38162,N_37271,N_36484);
xor U38163 (N_38163,N_36072,N_37296);
and U38164 (N_38164,N_36794,N_37352);
or U38165 (N_38165,N_37840,N_36564);
or U38166 (N_38166,N_36068,N_37943);
nor U38167 (N_38167,N_36898,N_36651);
nand U38168 (N_38168,N_36671,N_37766);
and U38169 (N_38169,N_37345,N_36786);
or U38170 (N_38170,N_36330,N_36583);
nand U38171 (N_38171,N_36202,N_36272);
xor U38172 (N_38172,N_36599,N_36545);
or U38173 (N_38173,N_37898,N_37200);
nand U38174 (N_38174,N_36423,N_37524);
nand U38175 (N_38175,N_37173,N_36571);
xnor U38176 (N_38176,N_37358,N_37170);
nand U38177 (N_38177,N_37876,N_37907);
or U38178 (N_38178,N_36974,N_37671);
and U38179 (N_38179,N_36462,N_36187);
nand U38180 (N_38180,N_37189,N_37293);
or U38181 (N_38181,N_37306,N_37770);
xnor U38182 (N_38182,N_36665,N_37257);
or U38183 (N_38183,N_36868,N_36346);
nor U38184 (N_38184,N_36847,N_37999);
xor U38185 (N_38185,N_36266,N_36656);
xnor U38186 (N_38186,N_36741,N_36325);
or U38187 (N_38187,N_36660,N_36270);
nand U38188 (N_38188,N_37212,N_37800);
nor U38189 (N_38189,N_36355,N_37643);
and U38190 (N_38190,N_37383,N_36963);
and U38191 (N_38191,N_36340,N_37158);
or U38192 (N_38192,N_37401,N_37194);
or U38193 (N_38193,N_37526,N_36809);
xnor U38194 (N_38194,N_36811,N_37867);
nor U38195 (N_38195,N_36498,N_37814);
nand U38196 (N_38196,N_37006,N_36648);
or U38197 (N_38197,N_37559,N_36175);
and U38198 (N_38198,N_37686,N_37685);
and U38199 (N_38199,N_36400,N_37843);
or U38200 (N_38200,N_36088,N_36468);
nand U38201 (N_38201,N_36842,N_36587);
nand U38202 (N_38202,N_37736,N_36866);
and U38203 (N_38203,N_37452,N_37405);
nand U38204 (N_38204,N_36130,N_36997);
nand U38205 (N_38205,N_36678,N_37162);
nand U38206 (N_38206,N_37238,N_36164);
xnor U38207 (N_38207,N_36576,N_37476);
xor U38208 (N_38208,N_37421,N_37654);
nor U38209 (N_38209,N_36453,N_37116);
nand U38210 (N_38210,N_37983,N_36905);
nor U38211 (N_38211,N_36750,N_36600);
and U38212 (N_38212,N_36899,N_37737);
or U38213 (N_38213,N_37734,N_36219);
nor U38214 (N_38214,N_37061,N_36037);
nand U38215 (N_38215,N_37375,N_36524);
and U38216 (N_38216,N_36464,N_37278);
xnor U38217 (N_38217,N_36696,N_36401);
or U38218 (N_38218,N_36951,N_36275);
xor U38219 (N_38219,N_36518,N_37336);
nand U38220 (N_38220,N_36802,N_36614);
xor U38221 (N_38221,N_37935,N_37307);
and U38222 (N_38222,N_37583,N_37017);
and U38223 (N_38223,N_36256,N_36883);
xor U38224 (N_38224,N_36840,N_36634);
or U38225 (N_38225,N_36402,N_37202);
or U38226 (N_38226,N_37885,N_37952);
xnor U38227 (N_38227,N_36150,N_37069);
and U38228 (N_38228,N_36929,N_36125);
or U38229 (N_38229,N_37546,N_36200);
and U38230 (N_38230,N_36906,N_37450);
nand U38231 (N_38231,N_36428,N_37269);
or U38232 (N_38232,N_36157,N_36999);
and U38233 (N_38233,N_36492,N_36055);
and U38234 (N_38234,N_36495,N_37178);
nand U38235 (N_38235,N_37392,N_36948);
nand U38236 (N_38236,N_37015,N_36299);
and U38237 (N_38237,N_36106,N_36642);
nor U38238 (N_38238,N_36172,N_37431);
xor U38239 (N_38239,N_37540,N_36822);
nand U38240 (N_38240,N_36826,N_37519);
or U38241 (N_38241,N_36624,N_36626);
xnor U38242 (N_38242,N_36305,N_36147);
xor U38243 (N_38243,N_37343,N_36420);
xnor U38244 (N_38244,N_36444,N_37118);
nand U38245 (N_38245,N_36016,N_36042);
nor U38246 (N_38246,N_37207,N_37950);
xor U38247 (N_38247,N_37424,N_37155);
or U38248 (N_38248,N_37213,N_37060);
nand U38249 (N_38249,N_36719,N_37908);
nand U38250 (N_38250,N_36525,N_37141);
nor U38251 (N_38251,N_36764,N_36163);
or U38252 (N_38252,N_36049,N_37616);
and U38253 (N_38253,N_37305,N_37615);
or U38254 (N_38254,N_37510,N_37772);
xnor U38255 (N_38255,N_36473,N_36680);
xnor U38256 (N_38256,N_37225,N_37620);
nand U38257 (N_38257,N_36967,N_36435);
nor U38258 (N_38258,N_36517,N_37941);
nand U38259 (N_38259,N_36688,N_37993);
nor U38260 (N_38260,N_36211,N_36558);
nand U38261 (N_38261,N_36001,N_37930);
and U38262 (N_38262,N_37459,N_37868);
nand U38263 (N_38263,N_37227,N_36647);
xnor U38264 (N_38264,N_37487,N_36782);
nor U38265 (N_38265,N_36982,N_37302);
nand U38266 (N_38266,N_37912,N_37386);
or U38267 (N_38267,N_36465,N_36943);
and U38268 (N_38268,N_37746,N_36279);
nand U38269 (N_38269,N_36500,N_37443);
nand U38270 (N_38270,N_36271,N_36394);
xnor U38271 (N_38271,N_36939,N_36235);
nand U38272 (N_38272,N_36815,N_36918);
nand U38273 (N_38273,N_36927,N_37696);
nand U38274 (N_38274,N_37504,N_36621);
or U38275 (N_38275,N_36308,N_37198);
nor U38276 (N_38276,N_37435,N_37948);
nor U38277 (N_38277,N_37251,N_37282);
and U38278 (N_38278,N_36836,N_37480);
nor U38279 (N_38279,N_37787,N_37290);
and U38280 (N_38280,N_36390,N_36737);
nand U38281 (N_38281,N_36099,N_36261);
nor U38282 (N_38282,N_36955,N_37967);
xnor U38283 (N_38283,N_36992,N_37856);
xnor U38284 (N_38284,N_37996,N_36611);
or U38285 (N_38285,N_37142,N_36180);
xor U38286 (N_38286,N_37939,N_37881);
nor U38287 (N_38287,N_37371,N_36165);
nor U38288 (N_38288,N_36823,N_36928);
nor U38289 (N_38289,N_36061,N_36641);
xnor U38290 (N_38290,N_36426,N_37823);
xor U38291 (N_38291,N_36084,N_37013);
nor U38292 (N_38292,N_36573,N_37979);
nor U38293 (N_38293,N_36205,N_36729);
or U38294 (N_38294,N_36734,N_36882);
xor U38295 (N_38295,N_36307,N_37848);
and U38296 (N_38296,N_37622,N_36744);
nand U38297 (N_38297,N_36885,N_37716);
nor U38298 (N_38298,N_36321,N_37958);
xnor U38299 (N_38299,N_37244,N_37434);
xor U38300 (N_38300,N_37810,N_37725);
and U38301 (N_38301,N_37376,N_36060);
xnor U38302 (N_38302,N_36488,N_37666);
nand U38303 (N_38303,N_37317,N_37019);
or U38304 (N_38304,N_36924,N_37949);
nand U38305 (N_38305,N_36097,N_37561);
nor U38306 (N_38306,N_37931,N_36501);
xnor U38307 (N_38307,N_37201,N_37148);
and U38308 (N_38308,N_36736,N_37124);
nor U38309 (N_38309,N_37310,N_36643);
and U38310 (N_38310,N_36313,N_37451);
or U38311 (N_38311,N_37515,N_36577);
xor U38312 (N_38312,N_37588,N_37070);
nor U38313 (N_38313,N_36377,N_36372);
xor U38314 (N_38314,N_36919,N_36101);
nand U38315 (N_38315,N_36123,N_37120);
or U38316 (N_38316,N_37131,N_36691);
nor U38317 (N_38317,N_36263,N_36108);
nand U38318 (N_38318,N_36233,N_36224);
nor U38319 (N_38319,N_37572,N_36612);
nor U38320 (N_38320,N_37436,N_37529);
nand U38321 (N_38321,N_36862,N_37641);
nor U38322 (N_38322,N_36066,N_37387);
and U38323 (N_38323,N_36590,N_36870);
and U38324 (N_38324,N_36732,N_36474);
xnor U38325 (N_38325,N_37799,N_36439);
nor U38326 (N_38326,N_36359,N_37829);
nand U38327 (N_38327,N_37267,N_37822);
and U38328 (N_38328,N_36215,N_36631);
nor U38329 (N_38329,N_37333,N_36243);
or U38330 (N_38330,N_37520,N_37393);
nor U38331 (N_38331,N_36386,N_37523);
nor U38332 (N_38332,N_37777,N_36654);
nor U38333 (N_38333,N_36630,N_36778);
nand U38334 (N_38334,N_37971,N_36923);
or U38335 (N_38335,N_36531,N_36148);
and U38336 (N_38336,N_37966,N_36768);
and U38337 (N_38337,N_36111,N_37713);
nor U38338 (N_38338,N_37340,N_37650);
and U38339 (N_38339,N_37875,N_36602);
or U38340 (N_38340,N_36458,N_37514);
nand U38341 (N_38341,N_36094,N_36645);
and U38342 (N_38342,N_37344,N_36812);
xor U38343 (N_38343,N_36519,N_37548);
nor U38344 (N_38344,N_37174,N_36936);
nor U38345 (N_38345,N_37797,N_37169);
or U38346 (N_38346,N_36153,N_37219);
nor U38347 (N_38347,N_37298,N_37975);
or U38348 (N_38348,N_36578,N_37832);
xnor U38349 (N_38349,N_37578,N_37029);
and U38350 (N_38350,N_37538,N_36877);
nand U38351 (N_38351,N_36429,N_37918);
or U38352 (N_38352,N_37419,N_37552);
nand U38353 (N_38353,N_36970,N_37329);
nor U38354 (N_38354,N_36735,N_37095);
nor U38355 (N_38355,N_37235,N_37537);
nor U38356 (N_38356,N_36855,N_37951);
nor U38357 (N_38357,N_36779,N_37547);
xnor U38358 (N_38358,N_36920,N_37642);
nand U38359 (N_38359,N_37571,N_37256);
nor U38360 (N_38360,N_36891,N_37838);
xor U38361 (N_38361,N_36278,N_36335);
and U38362 (N_38362,N_37301,N_36131);
and U38363 (N_38363,N_36483,N_36490);
or U38364 (N_38364,N_37929,N_36821);
nand U38365 (N_38365,N_37103,N_36950);
nor U38366 (N_38366,N_37653,N_37845);
or U38367 (N_38367,N_37074,N_37483);
nor U38368 (N_38368,N_36910,N_37982);
or U38369 (N_38369,N_37812,N_37264);
or U38370 (N_38370,N_37831,N_36740);
nor U38371 (N_38371,N_37824,N_37291);
xor U38372 (N_38372,N_36303,N_36282);
and U38373 (N_38373,N_37961,N_37044);
xnor U38374 (N_38374,N_37104,N_37068);
nand U38375 (N_38375,N_37075,N_36859);
nor U38376 (N_38376,N_37111,N_37933);
xnor U38377 (N_38377,N_36772,N_36436);
and U38378 (N_38378,N_37166,N_37932);
nor U38379 (N_38379,N_37090,N_37682);
or U38380 (N_38380,N_36551,N_36817);
nor U38381 (N_38381,N_37579,N_36301);
xor U38382 (N_38382,N_37330,N_36861);
or U38383 (N_38383,N_37292,N_36357);
nand U38384 (N_38384,N_36480,N_37630);
and U38385 (N_38385,N_36295,N_37584);
or U38386 (N_38386,N_37037,N_36913);
xor U38387 (N_38387,N_36220,N_36824);
xor U38388 (N_38388,N_37398,N_36186);
xnor U38389 (N_38389,N_37423,N_37112);
or U38390 (N_38390,N_36666,N_36685);
nor U38391 (N_38391,N_37954,N_36608);
and U38392 (N_38392,N_37362,N_36644);
and U38393 (N_38393,N_36721,N_37624);
and U38394 (N_38394,N_37214,N_37742);
or U38395 (N_38395,N_36789,N_37224);
nor U38396 (N_38396,N_36105,N_37621);
nand U38397 (N_38397,N_37956,N_36773);
or U38398 (N_38398,N_36461,N_36343);
xor U38399 (N_38399,N_36781,N_36339);
xor U38400 (N_38400,N_37473,N_36776);
nand U38401 (N_38401,N_37047,N_37804);
or U38402 (N_38402,N_37176,N_37687);
xor U38403 (N_38403,N_36813,N_37722);
nand U38404 (N_38404,N_36677,N_36598);
nand U38405 (N_38405,N_37833,N_37774);
nand U38406 (N_38406,N_37506,N_36427);
nor U38407 (N_38407,N_36451,N_36457);
or U38408 (N_38408,N_37626,N_37657);
nor U38409 (N_38409,N_36591,N_37396);
and U38410 (N_38410,N_37763,N_37632);
nor U38411 (N_38411,N_36616,N_37726);
nand U38412 (N_38412,N_37281,N_37350);
nand U38413 (N_38413,N_37516,N_36026);
and U38414 (N_38414,N_37805,N_36485);
or U38415 (N_38415,N_37633,N_36050);
and U38416 (N_38416,N_37689,N_36407);
or U38417 (N_38417,N_36456,N_36044);
nand U38418 (N_38418,N_37072,N_36692);
xor U38419 (N_38419,N_36998,N_37455);
nor U38420 (N_38420,N_37676,N_36129);
and U38421 (N_38421,N_36538,N_36979);
or U38422 (N_38422,N_36796,N_36874);
nand U38423 (N_38423,N_36076,N_36703);
nand U38424 (N_38424,N_37965,N_37254);
or U38425 (N_38425,N_36649,N_36623);
and U38426 (N_38426,N_37087,N_36362);
nand U38427 (N_38427,N_37471,N_36281);
or U38428 (N_38428,N_36900,N_36168);
nor U38429 (N_38429,N_36707,N_37378);
nor U38430 (N_38430,N_36854,N_37355);
nand U38431 (N_38431,N_36606,N_37346);
or U38432 (N_38432,N_36318,N_36414);
nor U38433 (N_38433,N_36958,N_36032);
xnor U38434 (N_38434,N_37549,N_37565);
xnor U38435 (N_38435,N_36880,N_37288);
nor U38436 (N_38436,N_37825,N_37106);
and U38437 (N_38437,N_36053,N_36714);
nor U38438 (N_38438,N_37113,N_37788);
and U38439 (N_38439,N_37819,N_36973);
xor U38440 (N_38440,N_37043,N_36361);
and U38441 (N_38441,N_36852,N_36526);
nand U38442 (N_38442,N_37998,N_37614);
and U38443 (N_38443,N_36294,N_37762);
nor U38444 (N_38444,N_37107,N_37079);
nand U38445 (N_38445,N_37563,N_36807);
nor U38446 (N_38446,N_37320,N_36546);
or U38447 (N_38447,N_36452,N_37357);
or U38448 (N_38448,N_37957,N_36568);
or U38449 (N_38449,N_37851,N_36615);
nand U38450 (N_38450,N_36700,N_36191);
or U38451 (N_38451,N_36569,N_36733);
nand U38452 (N_38452,N_37348,N_37795);
nand U38453 (N_38453,N_36675,N_36192);
or U38454 (N_38454,N_37580,N_37258);
or U38455 (N_38455,N_36188,N_37589);
or U38456 (N_38456,N_36702,N_36195);
and U38457 (N_38457,N_36865,N_36942);
nand U38458 (N_38458,N_36257,N_36204);
and U38459 (N_38459,N_37502,N_37384);
and U38460 (N_38460,N_37747,N_36421);
and U38461 (N_38461,N_36541,N_36806);
and U38462 (N_38462,N_36788,N_36659);
or U38463 (N_38463,N_36345,N_36292);
xor U38464 (N_38464,N_37741,N_36884);
nand U38465 (N_38465,N_36065,N_36350);
xor U38466 (N_38466,N_36635,N_37066);
nand U38467 (N_38467,N_37425,N_37995);
nand U38468 (N_38468,N_37909,N_37862);
nand U38469 (N_38469,N_36310,N_37042);
xnor U38470 (N_38470,N_36136,N_37969);
xnor U38471 (N_38471,N_37009,N_36259);
nor U38472 (N_38472,N_36946,N_37636);
or U38473 (N_38473,N_36236,N_36572);
or U38474 (N_38474,N_36446,N_36759);
or U38475 (N_38475,N_37052,N_37464);
nor U38476 (N_38476,N_37646,N_37062);
and U38477 (N_38477,N_37645,N_37880);
or U38478 (N_38478,N_37945,N_37243);
and U38479 (N_38479,N_36536,N_36810);
nor U38480 (N_38480,N_36673,N_37364);
nand U38481 (N_38481,N_36980,N_36742);
and U38482 (N_38482,N_37324,N_37428);
or U38483 (N_38483,N_37740,N_36493);
and U38484 (N_38484,N_36410,N_37422);
nand U38485 (N_38485,N_37779,N_36658);
and U38486 (N_38486,N_37323,N_37927);
or U38487 (N_38487,N_37366,N_36605);
nand U38488 (N_38488,N_36085,N_37083);
or U38489 (N_38489,N_36582,N_36080);
nand U38490 (N_38490,N_37236,N_36542);
nor U38491 (N_38491,N_37286,N_36352);
and U38492 (N_38492,N_37161,N_36708);
nor U38493 (N_38493,N_36757,N_37255);
xnor U38494 (N_38494,N_36198,N_37938);
nor U38495 (N_38495,N_36141,N_37245);
or U38496 (N_38496,N_36908,N_37922);
nor U38497 (N_38497,N_36639,N_36640);
or U38498 (N_38498,N_36253,N_36727);
or U38499 (N_38499,N_37096,N_36226);
or U38500 (N_38500,N_37730,N_37033);
or U38501 (N_38501,N_37149,N_37755);
nor U38502 (N_38502,N_37179,N_36393);
or U38503 (N_38503,N_36931,N_37115);
xor U38504 (N_38504,N_36687,N_36962);
or U38505 (N_38505,N_37134,N_36045);
nor U38506 (N_38506,N_37261,N_37992);
nand U38507 (N_38507,N_37801,N_36267);
nor U38508 (N_38508,N_37785,N_36539);
nand U38509 (N_38509,N_37486,N_37048);
nand U38510 (N_38510,N_36535,N_36154);
xor U38511 (N_38511,N_37128,N_37180);
nor U38512 (N_38512,N_36103,N_37539);
xnor U38513 (N_38513,N_37562,N_36503);
nand U38514 (N_38514,N_36273,N_36031);
or U38515 (N_38515,N_36533,N_36197);
and U38516 (N_38516,N_37656,N_36837);
or U38517 (N_38517,N_36379,N_37028);
nand U38518 (N_38518,N_37714,N_37897);
xor U38519 (N_38519,N_36553,N_36021);
or U38520 (N_38520,N_36601,N_36025);
nor U38521 (N_38521,N_37904,N_37887);
nand U38522 (N_38522,N_36933,N_37542);
or U38523 (N_38523,N_37429,N_36185);
nor U38524 (N_38524,N_37861,N_37046);
nand U38525 (N_38525,N_37495,N_36753);
xor U38526 (N_38526,N_37129,N_36367);
nor U38527 (N_38527,N_37325,N_37986);
or U38528 (N_38528,N_36724,N_36895);
or U38529 (N_38529,N_36034,N_36342);
and U38530 (N_38530,N_36547,N_36418);
nor U38531 (N_38531,N_36293,N_36260);
nor U38532 (N_38532,N_37454,N_37026);
nor U38533 (N_38533,N_36073,N_36383);
nand U38534 (N_38534,N_36432,N_37187);
nand U38535 (N_38535,N_36618,N_37870);
or U38536 (N_38536,N_36424,N_37910);
and U38537 (N_38537,N_36169,N_36107);
or U38538 (N_38538,N_36911,N_36440);
nand U38539 (N_38539,N_37263,N_36479);
nor U38540 (N_38540,N_37601,N_36477);
and U38541 (N_38541,N_37314,N_36889);
and U38542 (N_38542,N_36695,N_37803);
or U38543 (N_38543,N_36333,N_36230);
nand U38544 (N_38544,N_37792,N_36879);
or U38545 (N_38545,N_37667,N_37953);
and U38546 (N_38546,N_37311,N_37963);
or U38547 (N_38547,N_37417,N_36622);
nand U38548 (N_38548,N_36652,N_37039);
or U38549 (N_38549,N_37274,N_36041);
nor U38550 (N_38550,N_37771,N_36011);
and U38551 (N_38551,N_37649,N_36434);
and U38552 (N_38552,N_36509,N_37157);
nand U38553 (N_38553,N_36722,N_36693);
nor U38554 (N_38554,N_37186,N_37233);
xnor U38555 (N_38555,N_37203,N_37171);
nor U38556 (N_38556,N_37411,N_37813);
nor U38557 (N_38557,N_37415,N_37593);
nand U38558 (N_38558,N_37209,N_36184);
or U38559 (N_38559,N_37582,N_36269);
nand U38560 (N_38560,N_37050,N_37440);
or U38561 (N_38561,N_37603,N_36739);
or U38562 (N_38562,N_37210,N_37873);
nor U38563 (N_38563,N_36149,N_37294);
or U38564 (N_38564,N_36311,N_37490);
xor U38565 (N_38565,N_37853,N_36712);
xnor U38566 (N_38566,N_36331,N_37859);
nand U38567 (N_38567,N_37430,N_37928);
xnor U38568 (N_38568,N_36353,N_37234);
or U38569 (N_38569,N_37313,N_36063);
xnor U38570 (N_38570,N_36682,N_37521);
nor U38571 (N_38571,N_36790,N_37004);
or U38572 (N_38572,N_36586,N_37206);
nand U38573 (N_38573,N_36563,N_36317);
nand U38574 (N_38574,N_37628,N_36793);
or U38575 (N_38575,N_37156,N_36079);
and U38576 (N_38576,N_36089,N_37828);
xnor U38577 (N_38577,N_36805,N_37503);
and U38578 (N_38578,N_36554,N_36082);
and U38579 (N_38579,N_37872,N_36663);
or U38580 (N_38580,N_36067,N_36975);
and U38581 (N_38581,N_36143,N_37756);
xnor U38582 (N_38582,N_37679,N_36323);
nor U38583 (N_38583,N_37820,N_37659);
and U38584 (N_38584,N_37764,N_36579);
nand U38585 (N_38585,N_37444,N_36507);
or U38586 (N_38586,N_36276,N_36669);
and U38587 (N_38587,N_37493,N_36338);
nor U38588 (N_38588,N_36771,N_36347);
xor U38589 (N_38589,N_36985,N_37395);
nor U38590 (N_38590,N_37420,N_37150);
xnor U38591 (N_38591,N_36212,N_36241);
nand U38592 (N_38592,N_36010,N_37380);
nor U38593 (N_38593,N_36030,N_37049);
xnor U38594 (N_38594,N_37130,N_37154);
nor U38595 (N_38595,N_37022,N_37727);
and U38596 (N_38596,N_36754,N_36472);
xnor U38597 (N_38597,N_36382,N_36470);
or U38598 (N_38598,N_36858,N_37533);
nor U38599 (N_38599,N_37328,N_37407);
or U38600 (N_38600,N_37852,N_37663);
and U38601 (N_38601,N_37361,N_37609);
nand U38602 (N_38602,N_36574,N_37403);
xnor U38603 (N_38603,N_37308,N_37152);
nand U38604 (N_38604,N_37065,N_36239);
and U38605 (N_38605,N_36194,N_37027);
nor U38606 (N_38606,N_37944,N_36019);
and U38607 (N_38607,N_36024,N_36326);
nand U38608 (N_38608,N_36058,N_36201);
or U38609 (N_38609,N_36159,N_37576);
xnor U38610 (N_38610,N_36785,N_36092);
or U38611 (N_38611,N_36190,N_37466);
or U38612 (N_38612,N_36609,N_37410);
or U38613 (N_38613,N_36746,N_37794);
xor U38614 (N_38614,N_36981,N_37064);
nand U38615 (N_38615,N_36613,N_37211);
or U38616 (N_38616,N_36399,N_37560);
xor U38617 (N_38617,N_37372,N_37911);
and U38618 (N_38618,N_37008,N_36560);
nor U38619 (N_38619,N_37058,N_37172);
nor U38620 (N_38620,N_36006,N_37612);
xnor U38621 (N_38621,N_36039,N_37501);
or U38622 (N_38622,N_37081,N_36018);
nand U38623 (N_38623,N_36332,N_36767);
xor U38624 (N_38624,N_37119,N_37221);
xor U38625 (N_38625,N_37677,N_37757);
nand U38626 (N_38626,N_37744,N_37365);
nor U38627 (N_38627,N_36183,N_36445);
xor U38628 (N_38628,N_37359,N_36300);
xnor U38629 (N_38629,N_36597,N_37599);
and U38630 (N_38630,N_37318,N_37902);
nor U38631 (N_38631,N_36376,N_36711);
nand U38632 (N_38632,N_37160,N_36146);
nor U38633 (N_38633,N_37241,N_37003);
xor U38634 (N_38634,N_37874,N_36161);
or U38635 (N_38635,N_36499,N_36901);
or U38636 (N_38636,N_37086,N_37399);
nand U38637 (N_38637,N_37137,N_36683);
and U38638 (N_38638,N_37369,N_36814);
xor U38639 (N_38639,N_37195,N_37780);
nand U38640 (N_38640,N_37750,N_37332);
xnor U38641 (N_38641,N_36062,N_37449);
xnor U38642 (N_38642,N_37276,N_36628);
xnor U38643 (N_38643,N_37334,N_37715);
or U38644 (N_38644,N_37498,N_36593);
xor U38645 (N_38645,N_36994,N_36798);
nor U38646 (N_38646,N_36356,N_37926);
or U38647 (N_38647,N_37946,N_37220);
nor U38648 (N_38648,N_37525,N_36173);
and U38649 (N_38649,N_36956,N_36937);
xnor U38650 (N_38650,N_37285,N_37427);
nand U38651 (N_38651,N_36411,N_36348);
xor U38652 (N_38652,N_37228,N_37341);
nor U38653 (N_38653,N_37528,N_37618);
or U38654 (N_38654,N_37644,N_36132);
nor U38655 (N_38655,N_36448,N_37732);
and U38656 (N_38656,N_36437,N_37940);
and U38657 (N_38657,N_36832,N_36584);
or U38658 (N_38658,N_37639,N_37014);
nand U38659 (N_38659,N_36358,N_37590);
nand U38660 (N_38660,N_37602,N_36706);
xor U38661 (N_38661,N_37222,N_37051);
nand U38662 (N_38662,N_37249,N_37712);
nand U38663 (N_38663,N_37990,N_37720);
or U38664 (N_38664,N_36425,N_37024);
nand U38665 (N_38665,N_36869,N_37140);
nor U38666 (N_38666,N_36561,N_36835);
nor U38667 (N_38667,N_37159,N_37691);
or U38668 (N_38668,N_36972,N_37467);
nand U38669 (N_38669,N_36523,N_36381);
xor U38670 (N_38670,N_36965,N_37985);
or U38671 (N_38671,N_36699,N_36250);
xor U38672 (N_38672,N_36007,N_36478);
or U38673 (N_38673,N_37034,N_37262);
and U38674 (N_38674,N_37699,N_37554);
or U38675 (N_38675,N_36422,N_36397);
and U38676 (N_38676,N_37914,N_37509);
xor U38677 (N_38677,N_37108,N_37091);
nand U38678 (N_38678,N_37989,N_37575);
nand U38679 (N_38679,N_37855,N_37505);
nor U38680 (N_38680,N_36844,N_36415);
and U38681 (N_38681,N_36036,N_36231);
xnor U38682 (N_38682,N_37768,N_37032);
nor U38683 (N_38683,N_36521,N_37151);
nor U38684 (N_38684,N_36713,N_37775);
and U38685 (N_38685,N_37232,N_36344);
nor U38686 (N_38686,N_37252,N_36653);
and U38687 (N_38687,N_36915,N_36549);
nor U38688 (N_38688,N_37071,N_36657);
and U38689 (N_38689,N_37338,N_36848);
nand U38690 (N_38690,N_37697,N_36831);
xor U38691 (N_38691,N_36375,N_36406);
xnor U38692 (N_38692,N_37704,N_36341);
nand U38693 (N_38693,N_36655,N_37012);
and U38694 (N_38694,N_36459,N_37647);
or U38695 (N_38695,N_37786,N_37363);
xor U38696 (N_38696,N_36354,N_36417);
nand U38697 (N_38697,N_37793,N_37077);
nand U38698 (N_38698,N_36522,N_37481);
nand U38699 (N_38699,N_37373,N_37893);
and U38700 (N_38700,N_37105,N_37099);
xor U38701 (N_38701,N_36028,N_37404);
xnor U38702 (N_38702,N_36069,N_36620);
nand U38703 (N_38703,N_36244,N_36672);
nand U38704 (N_38704,N_36932,N_36510);
nor U38705 (N_38705,N_37675,N_37753);
and U38706 (N_38706,N_37895,N_36404);
nand U38707 (N_38707,N_36544,N_37216);
nor U38708 (N_38708,N_37367,N_36121);
and U38709 (N_38709,N_37277,N_37778);
or U38710 (N_38710,N_37970,N_36907);
and U38711 (N_38711,N_36217,N_36176);
and U38712 (N_38712,N_37442,N_36496);
nand U38713 (N_38713,N_36853,N_37863);
nor U38714 (N_38714,N_37672,N_36467);
nor U38715 (N_38715,N_37512,N_36179);
xor U38716 (N_38716,N_37402,N_37122);
or U38717 (N_38717,N_36726,N_36312);
nand U38718 (N_38718,N_36059,N_36819);
nand U38719 (N_38719,N_36115,N_36784);
xnor U38720 (N_38720,N_37462,N_36780);
nand U38721 (N_38721,N_36520,N_37568);
nand U38722 (N_38722,N_36283,N_36966);
nor U38723 (N_38723,N_37030,N_36697);
nor U38724 (N_38724,N_37135,N_36984);
or U38725 (N_38725,N_36941,N_36797);
and U38726 (N_38726,N_36431,N_37016);
and U38727 (N_38727,N_36917,N_36704);
or U38728 (N_38728,N_36139,N_36366);
xnor U38729 (N_38729,N_36249,N_36297);
or U38730 (N_38730,N_36403,N_37275);
nor U38731 (N_38731,N_36938,N_37553);
and U38732 (N_38732,N_37748,N_37229);
nand U38733 (N_38733,N_36914,N_37723);
nor U38734 (N_38734,N_36286,N_36667);
or U38735 (N_38735,N_37706,N_37098);
nand U38736 (N_38736,N_36514,N_37600);
and U38737 (N_38737,N_37842,N_36902);
and U38738 (N_38738,N_36717,N_36646);
nor U38739 (N_38739,N_36008,N_36385);
nor U38740 (N_38740,N_37413,N_36989);
xnor U38741 (N_38741,N_37133,N_36289);
xnor U38742 (N_38742,N_36570,N_36033);
and U38743 (N_38743,N_36698,N_37718);
nand U38744 (N_38744,N_36990,N_36566);
xor U38745 (N_38745,N_37492,N_37707);
xor U38746 (N_38746,N_36387,N_36530);
and U38747 (N_38747,N_37680,N_37906);
nand U38748 (N_38748,N_36953,N_37089);
and U38749 (N_38749,N_36209,N_37871);
xor U38750 (N_38750,N_36969,N_36783);
nand U38751 (N_38751,N_36013,N_37460);
xor U38752 (N_38752,N_37889,N_37608);
nand U38753 (N_38753,N_37204,N_36234);
nor U38754 (N_38754,N_37917,N_36816);
nand U38755 (N_38755,N_37789,N_37005);
xnor U38756 (N_38756,N_37188,N_37619);
nand U38757 (N_38757,N_37469,N_37683);
nand U38758 (N_38758,N_37240,N_37901);
or U38759 (N_38759,N_36747,N_36603);
xor U38760 (N_38760,N_37987,N_36792);
nor U38761 (N_38761,N_37218,N_36309);
or U38762 (N_38762,N_36291,N_37351);
nand U38763 (N_38763,N_37508,N_36684);
or U38764 (N_38764,N_37617,N_36003);
or U38765 (N_38765,N_37327,N_37193);
nor U38766 (N_38766,N_37920,N_37478);
xor U38767 (N_38767,N_36170,N_37205);
nand U38768 (N_38768,N_37183,N_37036);
xor U38769 (N_38769,N_36109,N_37899);
nor U38770 (N_38770,N_37864,N_36720);
xor U38771 (N_38771,N_36126,N_37038);
xor U38772 (N_38772,N_36252,N_36020);
nand U38773 (N_38773,N_37596,N_37892);
xor U38774 (N_38774,N_37242,N_37335);
and U38775 (N_38775,N_36328,N_36223);
and U38776 (N_38776,N_36993,N_36380);
nor U38777 (N_38777,N_36369,N_37470);
and U38778 (N_38778,N_37598,N_37959);
or U38779 (N_38779,N_36580,N_37353);
or U38780 (N_38780,N_36302,N_37611);
nor U38781 (N_38781,N_37692,N_36225);
nor U38782 (N_38782,N_36532,N_36890);
and U38783 (N_38783,N_36449,N_37811);
nand U38784 (N_38784,N_37592,N_36255);
nand U38785 (N_38785,N_37784,N_37147);
nand U38786 (N_38786,N_37472,N_37076);
or U38787 (N_38787,N_36327,N_36749);
or U38788 (N_38788,N_37673,N_36808);
or U38789 (N_38789,N_37199,N_36818);
nor U38790 (N_38790,N_37370,N_36681);
or U38791 (N_38791,N_36455,N_36743);
or U38792 (N_38792,N_37613,N_36930);
xnor U38793 (N_38793,N_36113,N_36296);
or U38794 (N_38794,N_37709,N_36873);
nor U38795 (N_38795,N_36638,N_37703);
nand U38796 (N_38796,N_37968,N_36756);
nand U38797 (N_38797,N_37627,N_36863);
xor U38798 (N_38798,N_36504,N_36505);
nand U38799 (N_38799,N_37694,N_37010);
nor U38800 (N_38800,N_36443,N_37287);
or U38801 (N_38801,N_36274,N_37078);
and U38802 (N_38802,N_36820,N_36137);
nor U38803 (N_38803,N_37056,N_37997);
xnor U38804 (N_38804,N_37669,N_36838);
xnor U38805 (N_38805,N_37972,N_36878);
nand U38806 (N_38806,N_36860,N_36537);
nor U38807 (N_38807,N_37919,N_36766);
or U38808 (N_38808,N_36413,N_37377);
and U38809 (N_38809,N_37331,N_36320);
and U38810 (N_38810,N_36368,N_37891);
and U38811 (N_38811,N_37791,N_36206);
nand U38812 (N_38812,N_36035,N_37088);
xor U38813 (N_38813,N_37835,N_37760);
or U38814 (N_38814,N_37196,N_37836);
nor U38815 (N_38815,N_36762,N_36218);
xnor U38816 (N_38816,N_36051,N_36804);
xnor U38817 (N_38817,N_37623,N_37040);
xnor U38818 (N_38818,N_36398,N_36491);
and U38819 (N_38819,N_37268,N_37847);
or U38820 (N_38820,N_37585,N_36112);
xor U38821 (N_38821,N_37259,N_37153);
and U38822 (N_38822,N_36567,N_36227);
xor U38823 (N_38823,N_36314,N_37655);
and U38824 (N_38824,N_37532,N_37942);
nor U38825 (N_38825,N_36512,N_37994);
and U38826 (N_38826,N_36222,N_37517);
nor U38827 (N_38827,N_37230,N_37316);
and U38828 (N_38828,N_36277,N_36119);
nor U38829 (N_38829,N_36408,N_36627);
nand U38830 (N_38830,N_37283,N_37705);
or U38831 (N_38831,N_37138,N_37144);
xor U38832 (N_38832,N_36945,N_37494);
nand U38833 (N_38833,N_36144,N_36728);
xnor U38834 (N_38834,N_36040,N_37577);
nand U38835 (N_38835,N_37558,N_36083);
nor U38836 (N_38836,N_37728,N_37815);
or U38837 (N_38837,N_36074,N_37759);
or U38838 (N_38838,N_36475,N_37721);
xor U38839 (N_38839,N_37117,N_36834);
nor U38840 (N_38840,N_37569,N_37123);
and U38841 (N_38841,N_37900,N_36174);
and U38842 (N_38842,N_36373,N_37527);
and U38843 (N_38843,N_36795,N_36110);
or U38844 (N_38844,N_36710,N_36254);
xor U38845 (N_38845,N_36048,N_37248);
or U38846 (N_38846,N_37635,N_37587);
and U38847 (N_38847,N_37101,N_36799);
nand U38848 (N_38848,N_36117,N_37182);
nand U38849 (N_38849,N_37841,N_37406);
nor U38850 (N_38850,N_37023,N_36071);
and U38851 (N_38851,N_36723,N_36046);
or U38852 (N_38852,N_37877,N_36002);
and U38853 (N_38853,N_37408,N_37962);
xnor U38854 (N_38854,N_36460,N_36298);
nor U38855 (N_38855,N_36324,N_36463);
and U38856 (N_38856,N_36934,N_36095);
xor U38857 (N_38857,N_36017,N_37000);
nand U38858 (N_38858,N_37782,N_37391);
and U38859 (N_38859,N_36412,N_36497);
nand U38860 (N_38860,N_36487,N_37886);
and U38861 (N_38861,N_37610,N_37094);
nor U38862 (N_38862,N_37418,N_36543);
or U38863 (N_38863,N_37260,N_37092);
or U38864 (N_38864,N_37461,N_37309);
or U38865 (N_38865,N_36637,N_37790);
nand U38866 (N_38866,N_36489,N_37700);
nor U38867 (N_38867,N_36349,N_37574);
nor U38868 (N_38868,N_36104,N_36988);
or U38869 (N_38869,N_37400,N_36978);
xnor U38870 (N_38870,N_37297,N_36471);
nor U38871 (N_38871,N_37660,N_36329);
nor U38872 (N_38872,N_37231,N_36392);
xnor U38873 (N_38873,N_37802,N_37658);
nand U38874 (N_38874,N_36086,N_37670);
nor U38875 (N_38875,N_36100,N_37439);
nor U38876 (N_38876,N_37681,N_37765);
xnor U38877 (N_38877,N_37315,N_37581);
xnor U38878 (N_38878,N_37817,N_37360);
and U38879 (N_38879,N_36395,N_36481);
and U38880 (N_38880,N_37416,N_37977);
and U38881 (N_38881,N_37067,N_36912);
nand U38882 (N_38882,N_37890,N_36715);
or U38883 (N_38883,N_37798,N_37925);
nand U38884 (N_38884,N_36078,N_36258);
nor U38885 (N_38885,N_36430,N_37322);
xnor U38886 (N_38886,N_37974,N_36508);
nor U38887 (N_38887,N_36265,N_36604);
nor U38888 (N_38888,N_37409,N_36760);
xnor U38889 (N_38889,N_36166,N_37109);
xnor U38890 (N_38890,N_37980,N_37143);
or U38891 (N_38891,N_37849,N_36617);
nor U38892 (N_38892,N_36087,N_37934);
xnor U38893 (N_38893,N_37923,N_37916);
or U38894 (N_38894,N_36189,N_37879);
nor U38895 (N_38895,N_37850,N_37607);
nor U38896 (N_38896,N_36029,N_37168);
nor U38897 (N_38897,N_37739,N_36843);
nand U38898 (N_38898,N_37648,N_36441);
xnor U38899 (N_38899,N_37059,N_36409);
and U38900 (N_38900,N_36925,N_37550);
nor U38901 (N_38901,N_36384,N_36208);
and U38902 (N_38902,N_36004,N_37507);
nor U38903 (N_38903,N_37484,N_37237);
and U38904 (N_38904,N_36502,N_37651);
and U38905 (N_38905,N_36057,N_37884);
xor U38906 (N_38906,N_37883,N_36023);
nand U38907 (N_38907,N_37300,N_36876);
nand U38908 (N_38908,N_36047,N_36801);
nand U38909 (N_38909,N_36288,N_37535);
nand U38910 (N_38910,N_37136,N_36290);
nand U38911 (N_38911,N_36633,N_37382);
nor U38912 (N_38912,N_36787,N_37114);
or U38913 (N_38913,N_36486,N_37865);
nor U38914 (N_38914,N_36893,N_37468);
nand U38915 (N_38915,N_37534,N_36940);
xnor U38916 (N_38916,N_37388,N_37984);
nand U38917 (N_38917,N_37674,N_37035);
and U38918 (N_38918,N_36336,N_36557);
nand U38919 (N_38919,N_36245,N_36070);
nor U38920 (N_38920,N_37693,N_36909);
nand U38921 (N_38921,N_36360,N_37226);
nor U38922 (N_38922,N_37102,N_36374);
xnor U38923 (N_38923,N_37084,N_37543);
xnor U38924 (N_38924,N_37807,N_37339);
nand U38925 (N_38925,N_36213,N_37477);
and U38926 (N_38926,N_36203,N_37031);
or U38927 (N_38927,N_37342,N_37385);
and U38928 (N_38928,N_37279,N_37937);
nor U38929 (N_38929,N_36178,N_37132);
nor U38930 (N_38930,N_36145,N_37964);
and U38931 (N_38931,N_36758,N_36516);
nand U38932 (N_38932,N_37761,N_37905);
or U38933 (N_38933,N_37045,N_36155);
and U38934 (N_38934,N_37457,N_37394);
nor U38935 (N_38935,N_36674,N_36871);
and U38936 (N_38936,N_36676,N_36124);
nand U38937 (N_38937,N_36845,N_37678);
and U38938 (N_38938,N_36529,N_37499);
or U38939 (N_38939,N_37564,N_37557);
or U38940 (N_38940,N_37303,N_36632);
or U38941 (N_38941,N_37711,N_37246);
xnor U38942 (N_38942,N_36287,N_37337);
or U38943 (N_38943,N_37767,N_37011);
or U38944 (N_38944,N_36494,N_36171);
nand U38945 (N_38945,N_36864,N_36365);
or U38946 (N_38946,N_36589,N_36228);
nor U38947 (N_38947,N_36364,N_36903);
or U38948 (N_38948,N_37684,N_36629);
and U38949 (N_38949,N_37586,N_36841);
xor U38950 (N_38950,N_36081,N_36625);
nor U38951 (N_38951,N_37127,N_36540);
nand U38952 (N_38952,N_37349,N_36251);
and U38953 (N_38953,N_37818,N_36770);
nand U38954 (N_38954,N_37806,N_37379);
and U38955 (N_38955,N_36594,N_37888);
nand U38956 (N_38956,N_36216,N_36850);
or U38957 (N_38957,N_37637,N_36238);
nand U38958 (N_38958,N_36610,N_37869);
and U38959 (N_38959,N_37556,N_36262);
xor U38960 (N_38960,N_37426,N_36661);
xor U38961 (N_38961,N_37223,N_37960);
nand U38962 (N_38962,N_36102,N_36791);
nand U38963 (N_38963,N_36284,N_37041);
xnor U38964 (N_38964,N_37668,N_36650);
or U38965 (N_38965,N_37414,N_36827);
or U38966 (N_38966,N_36709,N_36052);
or U38967 (N_38967,N_37555,N_37055);
nand U38968 (N_38968,N_37551,N_37485);
or U38969 (N_38969,N_36867,N_37724);
and U38970 (N_38970,N_37947,N_36881);
nor U38971 (N_38971,N_37496,N_36389);
nand U38972 (N_38972,N_37465,N_36926);
nor U38973 (N_38973,N_37978,N_37754);
xnor U38974 (N_38974,N_36595,N_37776);
and U38975 (N_38975,N_37896,N_37437);
xnor U38976 (N_38976,N_36022,N_36351);
and U38977 (N_38977,N_37265,N_37025);
or U38978 (N_38978,N_37878,N_36949);
or U38979 (N_38979,N_37701,N_36116);
or U38980 (N_38980,N_36619,N_37356);
and U38981 (N_38981,N_36152,N_36996);
nand U38982 (N_38982,N_36210,N_36752);
nand U38983 (N_38983,N_37605,N_37273);
or U38984 (N_38984,N_36334,N_37021);
nor U38985 (N_38985,N_37719,N_36534);
nor U38986 (N_38986,N_36689,N_37594);
nor U38987 (N_38987,N_37735,N_36896);
nor U38988 (N_38988,N_37390,N_36012);
nor U38989 (N_38989,N_37326,N_37215);
or U38990 (N_38990,N_37664,N_36701);
and U38991 (N_38991,N_37690,N_36581);
or U38992 (N_38992,N_37289,N_37100);
nand U38993 (N_38993,N_36986,N_37769);
xnor U38994 (N_38994,N_37844,N_37518);
xor U38995 (N_38995,N_37018,N_37773);
xnor U38996 (N_38996,N_37745,N_36961);
nand U38997 (N_38997,N_36396,N_36151);
or U38998 (N_38998,N_36315,N_36952);
or U38999 (N_38999,N_36438,N_36264);
and U39000 (N_39000,N_36888,N_37610);
xor U39001 (N_39001,N_37446,N_36967);
nor U39002 (N_39002,N_36805,N_36052);
nand U39003 (N_39003,N_37471,N_37668);
or U39004 (N_39004,N_36560,N_37499);
or U39005 (N_39005,N_36976,N_37836);
nand U39006 (N_39006,N_36367,N_37768);
nand U39007 (N_39007,N_36683,N_37795);
nor U39008 (N_39008,N_36199,N_37848);
and U39009 (N_39009,N_37265,N_37196);
xnor U39010 (N_39010,N_36930,N_37835);
nand U39011 (N_39011,N_36069,N_36172);
or U39012 (N_39012,N_37713,N_36872);
xor U39013 (N_39013,N_36323,N_36868);
or U39014 (N_39014,N_37072,N_36351);
xor U39015 (N_39015,N_36502,N_36765);
nand U39016 (N_39016,N_37912,N_37806);
nand U39017 (N_39017,N_37286,N_36962);
nand U39018 (N_39018,N_36398,N_36981);
xnor U39019 (N_39019,N_36883,N_36207);
or U39020 (N_39020,N_36775,N_36928);
or U39021 (N_39021,N_37282,N_36434);
or U39022 (N_39022,N_36992,N_37770);
nor U39023 (N_39023,N_37364,N_37442);
and U39024 (N_39024,N_36193,N_37740);
and U39025 (N_39025,N_37651,N_36692);
nor U39026 (N_39026,N_37059,N_37584);
and U39027 (N_39027,N_37611,N_37001);
xor U39028 (N_39028,N_37292,N_36553);
xnor U39029 (N_39029,N_37635,N_36405);
and U39030 (N_39030,N_36031,N_36091);
nor U39031 (N_39031,N_37157,N_37324);
nand U39032 (N_39032,N_37025,N_36763);
and U39033 (N_39033,N_37110,N_37403);
xor U39034 (N_39034,N_36450,N_37544);
and U39035 (N_39035,N_36628,N_37891);
nor U39036 (N_39036,N_36128,N_36919);
and U39037 (N_39037,N_36519,N_36993);
and U39038 (N_39038,N_36115,N_37147);
xor U39039 (N_39039,N_37999,N_37360);
nor U39040 (N_39040,N_36530,N_37990);
nor U39041 (N_39041,N_36928,N_37074);
or U39042 (N_39042,N_36912,N_37119);
nor U39043 (N_39043,N_37614,N_36047);
xor U39044 (N_39044,N_37915,N_37693);
xor U39045 (N_39045,N_37758,N_37779);
nand U39046 (N_39046,N_36419,N_36616);
nor U39047 (N_39047,N_37379,N_37996);
nand U39048 (N_39048,N_36916,N_37395);
and U39049 (N_39049,N_36169,N_37593);
nand U39050 (N_39050,N_36108,N_36333);
and U39051 (N_39051,N_37616,N_36085);
nand U39052 (N_39052,N_37837,N_37957);
nor U39053 (N_39053,N_37115,N_37979);
nor U39054 (N_39054,N_36212,N_37662);
nand U39055 (N_39055,N_36841,N_36048);
and U39056 (N_39056,N_37870,N_37902);
and U39057 (N_39057,N_37100,N_36814);
nand U39058 (N_39058,N_36329,N_37754);
nor U39059 (N_39059,N_37077,N_36480);
or U39060 (N_39060,N_37885,N_37351);
nor U39061 (N_39061,N_36356,N_37612);
xor U39062 (N_39062,N_36381,N_36468);
xor U39063 (N_39063,N_36215,N_37489);
nor U39064 (N_39064,N_37394,N_37038);
and U39065 (N_39065,N_36774,N_37903);
or U39066 (N_39066,N_37968,N_36793);
nand U39067 (N_39067,N_36550,N_37415);
xnor U39068 (N_39068,N_37118,N_36753);
nor U39069 (N_39069,N_37591,N_36359);
or U39070 (N_39070,N_37057,N_37153);
xor U39071 (N_39071,N_36984,N_37337);
nand U39072 (N_39072,N_37350,N_37292);
xnor U39073 (N_39073,N_36781,N_36861);
and U39074 (N_39074,N_37037,N_36266);
or U39075 (N_39075,N_36762,N_36130);
nor U39076 (N_39076,N_37721,N_36080);
nand U39077 (N_39077,N_36493,N_36022);
xor U39078 (N_39078,N_36860,N_36043);
nand U39079 (N_39079,N_36645,N_36625);
nor U39080 (N_39080,N_36937,N_36731);
nor U39081 (N_39081,N_37771,N_37992);
xnor U39082 (N_39082,N_37752,N_37494);
or U39083 (N_39083,N_36722,N_37713);
or U39084 (N_39084,N_37631,N_37902);
nor U39085 (N_39085,N_36170,N_37162);
and U39086 (N_39086,N_37893,N_37302);
nand U39087 (N_39087,N_37183,N_37204);
nor U39088 (N_39088,N_36677,N_36470);
or U39089 (N_39089,N_36063,N_37175);
or U39090 (N_39090,N_36550,N_37950);
or U39091 (N_39091,N_36218,N_36058);
and U39092 (N_39092,N_37462,N_37410);
nand U39093 (N_39093,N_36135,N_37893);
xor U39094 (N_39094,N_36891,N_36375);
or U39095 (N_39095,N_36277,N_37671);
nand U39096 (N_39096,N_36231,N_36772);
nand U39097 (N_39097,N_36768,N_37791);
or U39098 (N_39098,N_36729,N_36711);
or U39099 (N_39099,N_37734,N_37313);
nor U39100 (N_39100,N_36834,N_36381);
nand U39101 (N_39101,N_36917,N_37288);
or U39102 (N_39102,N_36954,N_36044);
nand U39103 (N_39103,N_36346,N_37533);
xor U39104 (N_39104,N_36189,N_36128);
nand U39105 (N_39105,N_37939,N_36953);
nor U39106 (N_39106,N_36084,N_37960);
and U39107 (N_39107,N_36115,N_36683);
xor U39108 (N_39108,N_37151,N_36996);
xor U39109 (N_39109,N_36727,N_37708);
nand U39110 (N_39110,N_37099,N_37818);
nand U39111 (N_39111,N_36827,N_37276);
and U39112 (N_39112,N_37196,N_37964);
nand U39113 (N_39113,N_37589,N_36850);
and U39114 (N_39114,N_36469,N_36223);
xnor U39115 (N_39115,N_37628,N_36652);
xor U39116 (N_39116,N_36839,N_36629);
or U39117 (N_39117,N_37622,N_37573);
and U39118 (N_39118,N_37336,N_37124);
nor U39119 (N_39119,N_36817,N_36344);
and U39120 (N_39120,N_36543,N_37784);
xnor U39121 (N_39121,N_37511,N_37897);
or U39122 (N_39122,N_36972,N_36244);
nor U39123 (N_39123,N_37443,N_37359);
xor U39124 (N_39124,N_36620,N_36677);
xnor U39125 (N_39125,N_37541,N_37131);
or U39126 (N_39126,N_37936,N_37429);
nand U39127 (N_39127,N_37932,N_37323);
nand U39128 (N_39128,N_37080,N_36207);
nand U39129 (N_39129,N_37486,N_36490);
nand U39130 (N_39130,N_36697,N_36558);
or U39131 (N_39131,N_36757,N_36292);
or U39132 (N_39132,N_37429,N_36764);
xor U39133 (N_39133,N_37955,N_36159);
xnor U39134 (N_39134,N_36316,N_37196);
nand U39135 (N_39135,N_37456,N_37036);
and U39136 (N_39136,N_37076,N_36641);
xnor U39137 (N_39137,N_36440,N_36834);
nand U39138 (N_39138,N_36833,N_36503);
or U39139 (N_39139,N_36192,N_36475);
and U39140 (N_39140,N_37792,N_36394);
nor U39141 (N_39141,N_37453,N_36587);
xor U39142 (N_39142,N_36440,N_36410);
xnor U39143 (N_39143,N_36274,N_36433);
nand U39144 (N_39144,N_36164,N_37471);
nand U39145 (N_39145,N_36659,N_36957);
nor U39146 (N_39146,N_37198,N_37819);
and U39147 (N_39147,N_36933,N_36281);
nor U39148 (N_39148,N_36459,N_36385);
nand U39149 (N_39149,N_36406,N_37488);
xnor U39150 (N_39150,N_36067,N_37163);
xnor U39151 (N_39151,N_37232,N_36148);
xor U39152 (N_39152,N_37349,N_37886);
nor U39153 (N_39153,N_37209,N_37132);
nor U39154 (N_39154,N_36000,N_36530);
nor U39155 (N_39155,N_37079,N_37698);
nor U39156 (N_39156,N_36461,N_37229);
xnor U39157 (N_39157,N_37941,N_37543);
nand U39158 (N_39158,N_37241,N_36483);
and U39159 (N_39159,N_36722,N_36680);
nor U39160 (N_39160,N_37268,N_37149);
nor U39161 (N_39161,N_36651,N_37702);
nor U39162 (N_39162,N_36761,N_37788);
or U39163 (N_39163,N_37634,N_36316);
xnor U39164 (N_39164,N_36378,N_37229);
and U39165 (N_39165,N_36017,N_36867);
or U39166 (N_39166,N_37903,N_36476);
nand U39167 (N_39167,N_36490,N_36107);
nand U39168 (N_39168,N_37878,N_37592);
nand U39169 (N_39169,N_37674,N_36033);
xor U39170 (N_39170,N_36132,N_36435);
or U39171 (N_39171,N_37881,N_37427);
or U39172 (N_39172,N_37654,N_36891);
or U39173 (N_39173,N_37242,N_36679);
or U39174 (N_39174,N_36588,N_36879);
and U39175 (N_39175,N_36936,N_36984);
nor U39176 (N_39176,N_36603,N_37984);
or U39177 (N_39177,N_36653,N_37284);
nand U39178 (N_39178,N_36414,N_37705);
and U39179 (N_39179,N_37093,N_37213);
and U39180 (N_39180,N_36911,N_37044);
and U39181 (N_39181,N_37267,N_37633);
nor U39182 (N_39182,N_36071,N_36515);
nor U39183 (N_39183,N_37043,N_37192);
or U39184 (N_39184,N_36672,N_36771);
xnor U39185 (N_39185,N_36263,N_37486);
nand U39186 (N_39186,N_37669,N_36341);
nor U39187 (N_39187,N_36439,N_37215);
xor U39188 (N_39188,N_37181,N_37152);
or U39189 (N_39189,N_37313,N_37823);
nor U39190 (N_39190,N_37223,N_36248);
or U39191 (N_39191,N_37335,N_37954);
or U39192 (N_39192,N_37395,N_36396);
nor U39193 (N_39193,N_37249,N_36180);
and U39194 (N_39194,N_36563,N_36732);
nand U39195 (N_39195,N_36085,N_37127);
nor U39196 (N_39196,N_36384,N_37656);
xor U39197 (N_39197,N_36087,N_37810);
nand U39198 (N_39198,N_36818,N_36125);
xnor U39199 (N_39199,N_37624,N_36778);
and U39200 (N_39200,N_36699,N_37175);
nor U39201 (N_39201,N_36419,N_36997);
and U39202 (N_39202,N_36182,N_36366);
nor U39203 (N_39203,N_37967,N_36493);
nor U39204 (N_39204,N_37111,N_36251);
nand U39205 (N_39205,N_37382,N_36421);
nand U39206 (N_39206,N_36920,N_36750);
and U39207 (N_39207,N_37799,N_37117);
or U39208 (N_39208,N_37131,N_37905);
xor U39209 (N_39209,N_36266,N_37307);
nand U39210 (N_39210,N_37985,N_36334);
or U39211 (N_39211,N_37548,N_36349);
nor U39212 (N_39212,N_37813,N_37817);
xor U39213 (N_39213,N_37334,N_37455);
nand U39214 (N_39214,N_36783,N_36815);
or U39215 (N_39215,N_37440,N_37696);
nor U39216 (N_39216,N_37295,N_36743);
xnor U39217 (N_39217,N_36421,N_37933);
xnor U39218 (N_39218,N_37295,N_36430);
nor U39219 (N_39219,N_36540,N_36341);
nor U39220 (N_39220,N_36832,N_37299);
nand U39221 (N_39221,N_36563,N_37781);
nand U39222 (N_39222,N_37943,N_36254);
and U39223 (N_39223,N_36770,N_36167);
nor U39224 (N_39224,N_36843,N_36081);
and U39225 (N_39225,N_36509,N_36264);
and U39226 (N_39226,N_36738,N_37659);
or U39227 (N_39227,N_37001,N_36768);
nor U39228 (N_39228,N_37840,N_36148);
nor U39229 (N_39229,N_37526,N_36843);
nand U39230 (N_39230,N_36666,N_37865);
nand U39231 (N_39231,N_37753,N_36187);
or U39232 (N_39232,N_36715,N_37934);
xor U39233 (N_39233,N_37256,N_36799);
nand U39234 (N_39234,N_36299,N_37229);
nand U39235 (N_39235,N_37196,N_36842);
or U39236 (N_39236,N_37812,N_36818);
and U39237 (N_39237,N_36331,N_36492);
nor U39238 (N_39238,N_37827,N_36569);
nor U39239 (N_39239,N_36055,N_37390);
and U39240 (N_39240,N_36302,N_36834);
xor U39241 (N_39241,N_37309,N_37733);
or U39242 (N_39242,N_37089,N_37876);
xor U39243 (N_39243,N_36632,N_37514);
nor U39244 (N_39244,N_36726,N_37039);
nor U39245 (N_39245,N_37810,N_37424);
nand U39246 (N_39246,N_37059,N_37224);
nor U39247 (N_39247,N_37782,N_37810);
and U39248 (N_39248,N_37133,N_36023);
or U39249 (N_39249,N_37702,N_36171);
xnor U39250 (N_39250,N_37018,N_36702);
and U39251 (N_39251,N_36985,N_37953);
or U39252 (N_39252,N_36213,N_37005);
nand U39253 (N_39253,N_37522,N_37054);
or U39254 (N_39254,N_37070,N_37028);
and U39255 (N_39255,N_36701,N_37338);
nand U39256 (N_39256,N_37104,N_37510);
nand U39257 (N_39257,N_36495,N_36554);
and U39258 (N_39258,N_37661,N_36246);
nand U39259 (N_39259,N_36018,N_36824);
and U39260 (N_39260,N_36767,N_37953);
xor U39261 (N_39261,N_37415,N_37755);
or U39262 (N_39262,N_37899,N_37370);
nor U39263 (N_39263,N_36027,N_36596);
nor U39264 (N_39264,N_36968,N_36567);
nand U39265 (N_39265,N_37365,N_36593);
and U39266 (N_39266,N_37157,N_36105);
and U39267 (N_39267,N_37667,N_37099);
xor U39268 (N_39268,N_37909,N_36852);
xor U39269 (N_39269,N_36389,N_37765);
nor U39270 (N_39270,N_36158,N_36233);
nor U39271 (N_39271,N_36493,N_37199);
nor U39272 (N_39272,N_36397,N_36076);
xnor U39273 (N_39273,N_36441,N_36287);
nand U39274 (N_39274,N_36820,N_36320);
xor U39275 (N_39275,N_36804,N_37846);
nor U39276 (N_39276,N_36839,N_37083);
nor U39277 (N_39277,N_37094,N_36771);
xor U39278 (N_39278,N_36680,N_37669);
nand U39279 (N_39279,N_36505,N_36620);
nand U39280 (N_39280,N_36247,N_36841);
or U39281 (N_39281,N_36936,N_37718);
and U39282 (N_39282,N_36278,N_37061);
and U39283 (N_39283,N_37061,N_37664);
xnor U39284 (N_39284,N_36200,N_37559);
nand U39285 (N_39285,N_37667,N_36346);
nand U39286 (N_39286,N_36550,N_36609);
or U39287 (N_39287,N_37969,N_36986);
and U39288 (N_39288,N_37795,N_36626);
and U39289 (N_39289,N_37616,N_36463);
or U39290 (N_39290,N_37051,N_37837);
nor U39291 (N_39291,N_37582,N_36504);
or U39292 (N_39292,N_36528,N_37368);
nand U39293 (N_39293,N_36591,N_37337);
nand U39294 (N_39294,N_36262,N_36945);
xnor U39295 (N_39295,N_37743,N_36178);
and U39296 (N_39296,N_36238,N_36236);
xor U39297 (N_39297,N_37718,N_36643);
nor U39298 (N_39298,N_36445,N_37148);
nor U39299 (N_39299,N_36516,N_36978);
xnor U39300 (N_39300,N_37662,N_36829);
and U39301 (N_39301,N_36272,N_37159);
xnor U39302 (N_39302,N_37625,N_37026);
nand U39303 (N_39303,N_37780,N_37061);
nand U39304 (N_39304,N_37836,N_37738);
or U39305 (N_39305,N_37511,N_36874);
nor U39306 (N_39306,N_36928,N_36701);
and U39307 (N_39307,N_37204,N_36260);
nor U39308 (N_39308,N_36200,N_36030);
and U39309 (N_39309,N_37545,N_36738);
nand U39310 (N_39310,N_36295,N_36682);
and U39311 (N_39311,N_36045,N_36976);
nor U39312 (N_39312,N_37127,N_37759);
and U39313 (N_39313,N_37902,N_36346);
xor U39314 (N_39314,N_37388,N_37793);
or U39315 (N_39315,N_37863,N_36246);
xnor U39316 (N_39316,N_37091,N_37788);
xor U39317 (N_39317,N_37036,N_36678);
or U39318 (N_39318,N_37460,N_37720);
or U39319 (N_39319,N_36592,N_37502);
nor U39320 (N_39320,N_37380,N_37797);
nand U39321 (N_39321,N_36464,N_37337);
or U39322 (N_39322,N_37597,N_36562);
nand U39323 (N_39323,N_36992,N_36117);
nor U39324 (N_39324,N_36559,N_37686);
or U39325 (N_39325,N_36887,N_37082);
xnor U39326 (N_39326,N_37590,N_36556);
nor U39327 (N_39327,N_36520,N_36669);
xnor U39328 (N_39328,N_37387,N_36885);
nand U39329 (N_39329,N_36372,N_36165);
and U39330 (N_39330,N_36289,N_36256);
xnor U39331 (N_39331,N_36737,N_36595);
nor U39332 (N_39332,N_37578,N_36753);
and U39333 (N_39333,N_37636,N_36381);
nand U39334 (N_39334,N_37541,N_37461);
or U39335 (N_39335,N_37031,N_37099);
nand U39336 (N_39336,N_37047,N_37947);
or U39337 (N_39337,N_36533,N_37787);
or U39338 (N_39338,N_37716,N_37618);
nand U39339 (N_39339,N_37145,N_37566);
nand U39340 (N_39340,N_37311,N_36797);
and U39341 (N_39341,N_36428,N_36071);
nand U39342 (N_39342,N_36347,N_37936);
xor U39343 (N_39343,N_36745,N_36817);
nor U39344 (N_39344,N_37762,N_37322);
nand U39345 (N_39345,N_37554,N_36357);
and U39346 (N_39346,N_37982,N_37742);
and U39347 (N_39347,N_36443,N_36216);
nand U39348 (N_39348,N_37588,N_37256);
and U39349 (N_39349,N_36485,N_36475);
xor U39350 (N_39350,N_37130,N_36046);
or U39351 (N_39351,N_36771,N_37918);
or U39352 (N_39352,N_37590,N_36922);
xnor U39353 (N_39353,N_36428,N_36176);
or U39354 (N_39354,N_37287,N_36307);
xor U39355 (N_39355,N_36387,N_37673);
nand U39356 (N_39356,N_36240,N_37904);
nor U39357 (N_39357,N_36537,N_37869);
or U39358 (N_39358,N_36920,N_36676);
nand U39359 (N_39359,N_36815,N_36729);
or U39360 (N_39360,N_36808,N_36985);
or U39361 (N_39361,N_37041,N_37630);
and U39362 (N_39362,N_36552,N_37346);
nand U39363 (N_39363,N_36972,N_37013);
xnor U39364 (N_39364,N_37742,N_36644);
or U39365 (N_39365,N_36389,N_37990);
xnor U39366 (N_39366,N_36215,N_36196);
nor U39367 (N_39367,N_37088,N_37678);
nand U39368 (N_39368,N_37260,N_36526);
and U39369 (N_39369,N_37027,N_36469);
nand U39370 (N_39370,N_37776,N_36245);
nor U39371 (N_39371,N_36023,N_36985);
and U39372 (N_39372,N_37890,N_36871);
xnor U39373 (N_39373,N_36325,N_36805);
nand U39374 (N_39374,N_37077,N_37371);
nand U39375 (N_39375,N_36411,N_36619);
nand U39376 (N_39376,N_36212,N_36548);
or U39377 (N_39377,N_37954,N_37497);
or U39378 (N_39378,N_37602,N_37252);
xor U39379 (N_39379,N_36674,N_37303);
nor U39380 (N_39380,N_36356,N_37942);
nor U39381 (N_39381,N_36063,N_37764);
xor U39382 (N_39382,N_37297,N_36101);
nor U39383 (N_39383,N_37726,N_36415);
nand U39384 (N_39384,N_37255,N_36262);
nand U39385 (N_39385,N_36765,N_36132);
or U39386 (N_39386,N_37420,N_37145);
or U39387 (N_39387,N_37229,N_36840);
xor U39388 (N_39388,N_36078,N_37176);
xor U39389 (N_39389,N_37602,N_36365);
nand U39390 (N_39390,N_36505,N_36219);
nor U39391 (N_39391,N_36078,N_36098);
xnor U39392 (N_39392,N_37049,N_37759);
xnor U39393 (N_39393,N_36784,N_37338);
and U39394 (N_39394,N_37304,N_36401);
and U39395 (N_39395,N_36598,N_36459);
and U39396 (N_39396,N_36739,N_37479);
nand U39397 (N_39397,N_37404,N_37834);
or U39398 (N_39398,N_37131,N_36617);
xnor U39399 (N_39399,N_37746,N_36044);
nand U39400 (N_39400,N_37681,N_36489);
nor U39401 (N_39401,N_37043,N_36408);
or U39402 (N_39402,N_37133,N_36055);
nor U39403 (N_39403,N_37707,N_37701);
and U39404 (N_39404,N_37931,N_37387);
and U39405 (N_39405,N_36737,N_36723);
or U39406 (N_39406,N_37896,N_36358);
xor U39407 (N_39407,N_36542,N_36772);
or U39408 (N_39408,N_36913,N_37625);
nand U39409 (N_39409,N_37971,N_36063);
or U39410 (N_39410,N_37036,N_37985);
xnor U39411 (N_39411,N_36074,N_37750);
nor U39412 (N_39412,N_36645,N_36165);
and U39413 (N_39413,N_36623,N_37682);
xor U39414 (N_39414,N_36599,N_37464);
or U39415 (N_39415,N_37386,N_36942);
nor U39416 (N_39416,N_36197,N_36754);
or U39417 (N_39417,N_37514,N_36297);
or U39418 (N_39418,N_37930,N_36680);
nor U39419 (N_39419,N_36911,N_37468);
xor U39420 (N_39420,N_36925,N_36944);
nor U39421 (N_39421,N_36653,N_36096);
xnor U39422 (N_39422,N_37686,N_37625);
nor U39423 (N_39423,N_36238,N_36312);
xnor U39424 (N_39424,N_37254,N_36573);
and U39425 (N_39425,N_37785,N_37767);
or U39426 (N_39426,N_36491,N_37594);
nor U39427 (N_39427,N_36627,N_37223);
nand U39428 (N_39428,N_37604,N_37166);
or U39429 (N_39429,N_36096,N_36804);
and U39430 (N_39430,N_37932,N_37361);
nand U39431 (N_39431,N_37068,N_37062);
and U39432 (N_39432,N_37439,N_36944);
and U39433 (N_39433,N_37814,N_36699);
nand U39434 (N_39434,N_36460,N_36626);
xnor U39435 (N_39435,N_37556,N_36558);
and U39436 (N_39436,N_37562,N_37199);
nand U39437 (N_39437,N_37116,N_36905);
xor U39438 (N_39438,N_36787,N_37160);
xor U39439 (N_39439,N_36092,N_37688);
nand U39440 (N_39440,N_37900,N_37883);
and U39441 (N_39441,N_36817,N_37527);
nor U39442 (N_39442,N_37310,N_37509);
and U39443 (N_39443,N_36099,N_36877);
nand U39444 (N_39444,N_36847,N_36862);
and U39445 (N_39445,N_36930,N_37140);
and U39446 (N_39446,N_36537,N_36909);
nor U39447 (N_39447,N_36573,N_36483);
nand U39448 (N_39448,N_37285,N_37367);
xnor U39449 (N_39449,N_37420,N_37667);
xnor U39450 (N_39450,N_36300,N_37588);
nor U39451 (N_39451,N_37481,N_37881);
nor U39452 (N_39452,N_36520,N_36838);
nand U39453 (N_39453,N_36971,N_36442);
xor U39454 (N_39454,N_37660,N_36864);
or U39455 (N_39455,N_36872,N_37217);
nand U39456 (N_39456,N_36488,N_36682);
and U39457 (N_39457,N_36557,N_37636);
xnor U39458 (N_39458,N_36813,N_37145);
nand U39459 (N_39459,N_37651,N_36639);
nand U39460 (N_39460,N_36710,N_37461);
xnor U39461 (N_39461,N_37520,N_36944);
xor U39462 (N_39462,N_36537,N_37855);
nand U39463 (N_39463,N_37756,N_37074);
and U39464 (N_39464,N_36101,N_36935);
and U39465 (N_39465,N_36668,N_36030);
and U39466 (N_39466,N_37557,N_36484);
nor U39467 (N_39467,N_37935,N_37571);
nand U39468 (N_39468,N_36912,N_37590);
nand U39469 (N_39469,N_36022,N_37647);
xor U39470 (N_39470,N_37758,N_36757);
or U39471 (N_39471,N_36564,N_37574);
or U39472 (N_39472,N_37577,N_37477);
nor U39473 (N_39473,N_37303,N_37952);
nand U39474 (N_39474,N_36251,N_36451);
nand U39475 (N_39475,N_36828,N_36835);
nand U39476 (N_39476,N_36076,N_37813);
nor U39477 (N_39477,N_37924,N_36903);
and U39478 (N_39478,N_36088,N_37611);
and U39479 (N_39479,N_36947,N_36748);
or U39480 (N_39480,N_36999,N_37700);
nor U39481 (N_39481,N_36469,N_36722);
nand U39482 (N_39482,N_36975,N_37289);
or U39483 (N_39483,N_37975,N_37540);
xor U39484 (N_39484,N_37121,N_37593);
xor U39485 (N_39485,N_36626,N_36116);
nand U39486 (N_39486,N_37570,N_37551);
or U39487 (N_39487,N_37658,N_36075);
xnor U39488 (N_39488,N_36298,N_36399);
nor U39489 (N_39489,N_37812,N_37216);
and U39490 (N_39490,N_37874,N_37513);
nand U39491 (N_39491,N_37433,N_36393);
xnor U39492 (N_39492,N_37077,N_36211);
xnor U39493 (N_39493,N_37524,N_36827);
nand U39494 (N_39494,N_36295,N_36836);
or U39495 (N_39495,N_37557,N_37952);
and U39496 (N_39496,N_36624,N_37331);
nand U39497 (N_39497,N_37841,N_37469);
nand U39498 (N_39498,N_37027,N_37473);
and U39499 (N_39499,N_36789,N_37749);
xnor U39500 (N_39500,N_37004,N_36384);
xor U39501 (N_39501,N_36406,N_36743);
nor U39502 (N_39502,N_37023,N_36403);
nor U39503 (N_39503,N_36172,N_37219);
or U39504 (N_39504,N_37326,N_37930);
xor U39505 (N_39505,N_37178,N_37730);
nand U39506 (N_39506,N_36262,N_37282);
or U39507 (N_39507,N_36596,N_36464);
or U39508 (N_39508,N_37478,N_36312);
nand U39509 (N_39509,N_37621,N_36258);
and U39510 (N_39510,N_36935,N_37124);
nor U39511 (N_39511,N_36514,N_37077);
or U39512 (N_39512,N_37164,N_36827);
and U39513 (N_39513,N_37379,N_37941);
and U39514 (N_39514,N_37030,N_37954);
and U39515 (N_39515,N_36867,N_37620);
xnor U39516 (N_39516,N_37230,N_37528);
and U39517 (N_39517,N_36843,N_36660);
xor U39518 (N_39518,N_36213,N_36304);
or U39519 (N_39519,N_36412,N_37656);
or U39520 (N_39520,N_37360,N_36096);
and U39521 (N_39521,N_36561,N_37334);
or U39522 (N_39522,N_37153,N_36238);
nand U39523 (N_39523,N_37270,N_36097);
nand U39524 (N_39524,N_36293,N_37820);
nand U39525 (N_39525,N_36886,N_37826);
nand U39526 (N_39526,N_37279,N_36461);
nand U39527 (N_39527,N_36340,N_37085);
nand U39528 (N_39528,N_36579,N_36072);
xor U39529 (N_39529,N_36761,N_37301);
or U39530 (N_39530,N_37087,N_37331);
xor U39531 (N_39531,N_36783,N_37297);
nand U39532 (N_39532,N_37689,N_37046);
and U39533 (N_39533,N_37057,N_37440);
nor U39534 (N_39534,N_36831,N_37363);
nor U39535 (N_39535,N_36982,N_36500);
nand U39536 (N_39536,N_36541,N_36539);
nand U39537 (N_39537,N_36773,N_37880);
and U39538 (N_39538,N_36112,N_36731);
nor U39539 (N_39539,N_37242,N_36523);
nor U39540 (N_39540,N_36984,N_37448);
xnor U39541 (N_39541,N_37946,N_36850);
xnor U39542 (N_39542,N_37862,N_37527);
nand U39543 (N_39543,N_36588,N_36698);
nand U39544 (N_39544,N_36490,N_36255);
xor U39545 (N_39545,N_37329,N_37507);
or U39546 (N_39546,N_36771,N_36860);
or U39547 (N_39547,N_36610,N_36325);
nand U39548 (N_39548,N_37959,N_37171);
nor U39549 (N_39549,N_36555,N_37195);
nor U39550 (N_39550,N_37978,N_37511);
nor U39551 (N_39551,N_36591,N_37683);
and U39552 (N_39552,N_37174,N_37331);
and U39553 (N_39553,N_36326,N_36913);
and U39554 (N_39554,N_36071,N_36821);
or U39555 (N_39555,N_37327,N_37795);
and U39556 (N_39556,N_36384,N_37580);
nand U39557 (N_39557,N_37868,N_36472);
nand U39558 (N_39558,N_37366,N_36504);
xor U39559 (N_39559,N_37630,N_37006);
and U39560 (N_39560,N_37074,N_37921);
xnor U39561 (N_39561,N_36466,N_37325);
nand U39562 (N_39562,N_36613,N_36253);
and U39563 (N_39563,N_37275,N_36647);
nand U39564 (N_39564,N_37944,N_36522);
nor U39565 (N_39565,N_37115,N_36635);
and U39566 (N_39566,N_37031,N_37507);
xor U39567 (N_39567,N_37797,N_36089);
and U39568 (N_39568,N_36446,N_37285);
nand U39569 (N_39569,N_36487,N_37944);
xnor U39570 (N_39570,N_36612,N_36680);
and U39571 (N_39571,N_36319,N_36321);
nand U39572 (N_39572,N_37945,N_36967);
nand U39573 (N_39573,N_36479,N_37329);
and U39574 (N_39574,N_37108,N_37989);
or U39575 (N_39575,N_37801,N_36545);
nand U39576 (N_39576,N_37451,N_36709);
nor U39577 (N_39577,N_37040,N_36138);
xnor U39578 (N_39578,N_37234,N_37583);
nand U39579 (N_39579,N_36243,N_37604);
xor U39580 (N_39580,N_37712,N_36967);
xor U39581 (N_39581,N_36137,N_36943);
or U39582 (N_39582,N_36554,N_37792);
or U39583 (N_39583,N_37759,N_37201);
nor U39584 (N_39584,N_37766,N_37730);
xnor U39585 (N_39585,N_36635,N_36699);
or U39586 (N_39586,N_36642,N_36485);
xor U39587 (N_39587,N_36164,N_36835);
and U39588 (N_39588,N_37272,N_36199);
nor U39589 (N_39589,N_36400,N_37585);
or U39590 (N_39590,N_37212,N_36089);
nand U39591 (N_39591,N_37468,N_36409);
xor U39592 (N_39592,N_36278,N_36463);
nor U39593 (N_39593,N_37730,N_37159);
nor U39594 (N_39594,N_36707,N_37328);
or U39595 (N_39595,N_37053,N_36602);
and U39596 (N_39596,N_36459,N_37909);
nor U39597 (N_39597,N_37739,N_37225);
nand U39598 (N_39598,N_37420,N_37140);
or U39599 (N_39599,N_36151,N_36208);
nor U39600 (N_39600,N_36456,N_36056);
and U39601 (N_39601,N_36291,N_37739);
and U39602 (N_39602,N_37534,N_37699);
and U39603 (N_39603,N_36066,N_36433);
nand U39604 (N_39604,N_37052,N_37810);
and U39605 (N_39605,N_37754,N_36019);
and U39606 (N_39606,N_37127,N_36589);
and U39607 (N_39607,N_37995,N_37072);
or U39608 (N_39608,N_37018,N_37443);
nor U39609 (N_39609,N_37462,N_36842);
and U39610 (N_39610,N_37234,N_37889);
xnor U39611 (N_39611,N_37563,N_36273);
nand U39612 (N_39612,N_37422,N_37463);
and U39613 (N_39613,N_37443,N_36879);
or U39614 (N_39614,N_36527,N_37868);
and U39615 (N_39615,N_37079,N_37142);
or U39616 (N_39616,N_36960,N_37560);
and U39617 (N_39617,N_37200,N_36444);
nor U39618 (N_39618,N_36699,N_36994);
or U39619 (N_39619,N_36433,N_36977);
nand U39620 (N_39620,N_36105,N_36248);
xor U39621 (N_39621,N_36595,N_36096);
xor U39622 (N_39622,N_37563,N_37472);
nand U39623 (N_39623,N_37311,N_36701);
nand U39624 (N_39624,N_36017,N_37869);
nand U39625 (N_39625,N_36655,N_37538);
and U39626 (N_39626,N_36433,N_36812);
nor U39627 (N_39627,N_37294,N_36924);
nand U39628 (N_39628,N_37589,N_37101);
nand U39629 (N_39629,N_36507,N_37546);
nand U39630 (N_39630,N_37865,N_36166);
or U39631 (N_39631,N_36137,N_36541);
nand U39632 (N_39632,N_37006,N_37749);
nand U39633 (N_39633,N_36380,N_36819);
nand U39634 (N_39634,N_37197,N_37176);
nand U39635 (N_39635,N_37883,N_36840);
nor U39636 (N_39636,N_37473,N_37204);
nand U39637 (N_39637,N_36617,N_36612);
and U39638 (N_39638,N_37572,N_37587);
xnor U39639 (N_39639,N_36128,N_37351);
or U39640 (N_39640,N_36632,N_37515);
or U39641 (N_39641,N_37475,N_36382);
xor U39642 (N_39642,N_36543,N_36160);
nand U39643 (N_39643,N_36008,N_37597);
nor U39644 (N_39644,N_36053,N_37414);
and U39645 (N_39645,N_36292,N_36569);
xnor U39646 (N_39646,N_36423,N_37131);
nand U39647 (N_39647,N_37590,N_37026);
nand U39648 (N_39648,N_36745,N_37049);
and U39649 (N_39649,N_36932,N_37647);
nand U39650 (N_39650,N_36366,N_36222);
and U39651 (N_39651,N_36037,N_36457);
nand U39652 (N_39652,N_36896,N_36480);
nand U39653 (N_39653,N_37476,N_36658);
and U39654 (N_39654,N_36405,N_36684);
nor U39655 (N_39655,N_37817,N_37434);
and U39656 (N_39656,N_37807,N_37038);
nor U39657 (N_39657,N_36264,N_37351);
xnor U39658 (N_39658,N_36818,N_36057);
and U39659 (N_39659,N_37933,N_37827);
and U39660 (N_39660,N_37652,N_36154);
and U39661 (N_39661,N_37149,N_37186);
nand U39662 (N_39662,N_37625,N_36459);
xor U39663 (N_39663,N_36374,N_37009);
and U39664 (N_39664,N_37228,N_37982);
nor U39665 (N_39665,N_37274,N_36342);
and U39666 (N_39666,N_36081,N_37435);
xor U39667 (N_39667,N_36205,N_36421);
or U39668 (N_39668,N_36133,N_37887);
or U39669 (N_39669,N_37358,N_36471);
or U39670 (N_39670,N_37562,N_37397);
xnor U39671 (N_39671,N_36733,N_37807);
nor U39672 (N_39672,N_37259,N_37681);
nand U39673 (N_39673,N_37163,N_36304);
nor U39674 (N_39674,N_37736,N_36112);
or U39675 (N_39675,N_36918,N_37043);
or U39676 (N_39676,N_36060,N_37670);
or U39677 (N_39677,N_37080,N_36769);
nor U39678 (N_39678,N_37411,N_37267);
nand U39679 (N_39679,N_36598,N_37849);
or U39680 (N_39680,N_37303,N_37947);
nor U39681 (N_39681,N_36181,N_37121);
and U39682 (N_39682,N_36707,N_36690);
nor U39683 (N_39683,N_37860,N_37619);
xor U39684 (N_39684,N_36842,N_37799);
nor U39685 (N_39685,N_36728,N_37678);
nand U39686 (N_39686,N_36663,N_36212);
nand U39687 (N_39687,N_36578,N_36149);
or U39688 (N_39688,N_37104,N_36579);
xnor U39689 (N_39689,N_36623,N_36941);
xor U39690 (N_39690,N_37434,N_36955);
nor U39691 (N_39691,N_36622,N_36877);
xnor U39692 (N_39692,N_36253,N_36688);
xor U39693 (N_39693,N_37880,N_37730);
nor U39694 (N_39694,N_37465,N_37210);
and U39695 (N_39695,N_37967,N_36048);
nor U39696 (N_39696,N_37043,N_37620);
or U39697 (N_39697,N_36523,N_36319);
or U39698 (N_39698,N_36152,N_37215);
nand U39699 (N_39699,N_36466,N_37870);
and U39700 (N_39700,N_36643,N_37385);
nor U39701 (N_39701,N_37809,N_36462);
xnor U39702 (N_39702,N_36319,N_37797);
or U39703 (N_39703,N_36480,N_37873);
nor U39704 (N_39704,N_37065,N_36073);
and U39705 (N_39705,N_36414,N_36673);
xor U39706 (N_39706,N_36178,N_36958);
nor U39707 (N_39707,N_36590,N_37525);
nor U39708 (N_39708,N_36073,N_36299);
xnor U39709 (N_39709,N_36745,N_36532);
nor U39710 (N_39710,N_37480,N_36655);
xnor U39711 (N_39711,N_37168,N_36342);
and U39712 (N_39712,N_36036,N_36030);
nor U39713 (N_39713,N_36840,N_37108);
nand U39714 (N_39714,N_37884,N_37500);
nor U39715 (N_39715,N_36065,N_36940);
and U39716 (N_39716,N_37295,N_37120);
or U39717 (N_39717,N_37680,N_37490);
xnor U39718 (N_39718,N_37173,N_37029);
nand U39719 (N_39719,N_37948,N_36155);
nand U39720 (N_39720,N_37755,N_37562);
and U39721 (N_39721,N_36183,N_37139);
nor U39722 (N_39722,N_37713,N_37763);
and U39723 (N_39723,N_37650,N_36758);
nand U39724 (N_39724,N_36457,N_36218);
nand U39725 (N_39725,N_36262,N_37434);
xnor U39726 (N_39726,N_37591,N_36686);
and U39727 (N_39727,N_37810,N_37206);
nor U39728 (N_39728,N_36194,N_37642);
nor U39729 (N_39729,N_36947,N_37185);
and U39730 (N_39730,N_36294,N_36192);
or U39731 (N_39731,N_37937,N_36277);
nand U39732 (N_39732,N_37403,N_37823);
and U39733 (N_39733,N_37696,N_36891);
xnor U39734 (N_39734,N_37876,N_36137);
nand U39735 (N_39735,N_36708,N_37236);
xnor U39736 (N_39736,N_36515,N_36463);
xnor U39737 (N_39737,N_36962,N_37816);
nor U39738 (N_39738,N_37488,N_36148);
nand U39739 (N_39739,N_36831,N_37388);
nor U39740 (N_39740,N_36418,N_36280);
and U39741 (N_39741,N_37173,N_36020);
and U39742 (N_39742,N_36397,N_37121);
nor U39743 (N_39743,N_37088,N_37560);
and U39744 (N_39744,N_37224,N_36166);
nand U39745 (N_39745,N_37569,N_37266);
and U39746 (N_39746,N_37405,N_36376);
or U39747 (N_39747,N_37219,N_37671);
nand U39748 (N_39748,N_36308,N_36516);
or U39749 (N_39749,N_36612,N_37522);
nor U39750 (N_39750,N_36117,N_37221);
xor U39751 (N_39751,N_36595,N_37235);
or U39752 (N_39752,N_37181,N_37773);
or U39753 (N_39753,N_37306,N_37457);
nor U39754 (N_39754,N_36243,N_36484);
nand U39755 (N_39755,N_37932,N_36238);
nand U39756 (N_39756,N_36877,N_37880);
nor U39757 (N_39757,N_36975,N_37473);
and U39758 (N_39758,N_37813,N_36526);
nand U39759 (N_39759,N_37490,N_37457);
nor U39760 (N_39760,N_36484,N_37745);
or U39761 (N_39761,N_36247,N_36902);
nor U39762 (N_39762,N_36956,N_36367);
nor U39763 (N_39763,N_36215,N_36120);
and U39764 (N_39764,N_37452,N_36793);
or U39765 (N_39765,N_37925,N_36983);
or U39766 (N_39766,N_37784,N_37881);
or U39767 (N_39767,N_37825,N_37121);
or U39768 (N_39768,N_36363,N_36772);
or U39769 (N_39769,N_36829,N_37520);
nand U39770 (N_39770,N_37483,N_37672);
xor U39771 (N_39771,N_37421,N_37916);
xor U39772 (N_39772,N_36054,N_36945);
xnor U39773 (N_39773,N_37409,N_36978);
nand U39774 (N_39774,N_37799,N_37464);
nand U39775 (N_39775,N_37876,N_37721);
or U39776 (N_39776,N_37270,N_37470);
xor U39777 (N_39777,N_37920,N_37100);
nand U39778 (N_39778,N_37046,N_36269);
and U39779 (N_39779,N_36326,N_36666);
nand U39780 (N_39780,N_36670,N_36714);
and U39781 (N_39781,N_37049,N_36318);
xor U39782 (N_39782,N_37643,N_36126);
or U39783 (N_39783,N_37345,N_37160);
xnor U39784 (N_39784,N_37000,N_36758);
nand U39785 (N_39785,N_37846,N_37064);
nor U39786 (N_39786,N_36747,N_37348);
and U39787 (N_39787,N_37249,N_36033);
xor U39788 (N_39788,N_37017,N_37727);
or U39789 (N_39789,N_37281,N_37315);
nor U39790 (N_39790,N_36090,N_36806);
xnor U39791 (N_39791,N_36209,N_36076);
and U39792 (N_39792,N_36857,N_37448);
nor U39793 (N_39793,N_36973,N_37118);
nand U39794 (N_39794,N_37996,N_36038);
xnor U39795 (N_39795,N_37115,N_37237);
or U39796 (N_39796,N_36714,N_36007);
xor U39797 (N_39797,N_37750,N_37086);
nand U39798 (N_39798,N_36907,N_36309);
or U39799 (N_39799,N_36732,N_36135);
or U39800 (N_39800,N_36836,N_37588);
nor U39801 (N_39801,N_36270,N_37753);
nor U39802 (N_39802,N_37753,N_36965);
and U39803 (N_39803,N_37017,N_37014);
and U39804 (N_39804,N_36548,N_37005);
nand U39805 (N_39805,N_37403,N_37429);
and U39806 (N_39806,N_36994,N_37057);
nand U39807 (N_39807,N_37318,N_37914);
xnor U39808 (N_39808,N_37750,N_36630);
and U39809 (N_39809,N_36960,N_36063);
or U39810 (N_39810,N_37511,N_37616);
xor U39811 (N_39811,N_36208,N_36137);
and U39812 (N_39812,N_37205,N_36862);
nand U39813 (N_39813,N_37246,N_37725);
and U39814 (N_39814,N_36122,N_37277);
or U39815 (N_39815,N_37285,N_36833);
nand U39816 (N_39816,N_36548,N_37475);
xnor U39817 (N_39817,N_36152,N_37031);
or U39818 (N_39818,N_37148,N_36929);
nand U39819 (N_39819,N_37397,N_37359);
or U39820 (N_39820,N_36473,N_36670);
xnor U39821 (N_39821,N_36096,N_37047);
or U39822 (N_39822,N_37309,N_36052);
or U39823 (N_39823,N_36131,N_36898);
nand U39824 (N_39824,N_36958,N_37357);
xnor U39825 (N_39825,N_36368,N_36904);
nor U39826 (N_39826,N_37369,N_37615);
and U39827 (N_39827,N_37938,N_37142);
nand U39828 (N_39828,N_36315,N_37581);
nor U39829 (N_39829,N_36382,N_36390);
or U39830 (N_39830,N_36419,N_36298);
and U39831 (N_39831,N_36232,N_37805);
nand U39832 (N_39832,N_36375,N_37845);
or U39833 (N_39833,N_36764,N_36691);
nor U39834 (N_39834,N_37659,N_37169);
nor U39835 (N_39835,N_36009,N_37151);
nor U39836 (N_39836,N_37806,N_37343);
nor U39837 (N_39837,N_36408,N_36690);
nand U39838 (N_39838,N_37814,N_36399);
xor U39839 (N_39839,N_36488,N_36776);
nand U39840 (N_39840,N_36559,N_36099);
nor U39841 (N_39841,N_37184,N_36973);
and U39842 (N_39842,N_37441,N_37290);
xnor U39843 (N_39843,N_37740,N_36922);
nand U39844 (N_39844,N_37361,N_36995);
and U39845 (N_39845,N_37923,N_36474);
or U39846 (N_39846,N_36010,N_37869);
or U39847 (N_39847,N_37083,N_37439);
or U39848 (N_39848,N_37316,N_36876);
nand U39849 (N_39849,N_36141,N_37345);
xnor U39850 (N_39850,N_37386,N_37602);
nand U39851 (N_39851,N_36885,N_36085);
nor U39852 (N_39852,N_37774,N_36660);
or U39853 (N_39853,N_36316,N_36877);
xor U39854 (N_39854,N_36358,N_37936);
xnor U39855 (N_39855,N_37049,N_37494);
and U39856 (N_39856,N_36520,N_37921);
and U39857 (N_39857,N_36088,N_37023);
nand U39858 (N_39858,N_37448,N_37410);
and U39859 (N_39859,N_37041,N_37206);
nand U39860 (N_39860,N_37384,N_37313);
xnor U39861 (N_39861,N_36523,N_37289);
and U39862 (N_39862,N_37224,N_37145);
or U39863 (N_39863,N_37524,N_37507);
or U39864 (N_39864,N_36725,N_36126);
nor U39865 (N_39865,N_36031,N_37387);
nand U39866 (N_39866,N_37838,N_37405);
nand U39867 (N_39867,N_36036,N_36691);
nor U39868 (N_39868,N_37791,N_37420);
nor U39869 (N_39869,N_36764,N_37098);
and U39870 (N_39870,N_37592,N_36248);
xor U39871 (N_39871,N_36426,N_37028);
nor U39872 (N_39872,N_37225,N_37622);
nor U39873 (N_39873,N_37389,N_37880);
or U39874 (N_39874,N_36530,N_36621);
xnor U39875 (N_39875,N_36190,N_37737);
and U39876 (N_39876,N_37466,N_37312);
xor U39877 (N_39877,N_37600,N_37045);
and U39878 (N_39878,N_36934,N_36688);
xor U39879 (N_39879,N_37369,N_36329);
nor U39880 (N_39880,N_36594,N_36832);
and U39881 (N_39881,N_37502,N_36141);
nor U39882 (N_39882,N_36494,N_36392);
and U39883 (N_39883,N_36664,N_36796);
xnor U39884 (N_39884,N_36864,N_37647);
or U39885 (N_39885,N_37680,N_37628);
or U39886 (N_39886,N_36345,N_36636);
or U39887 (N_39887,N_37274,N_36937);
or U39888 (N_39888,N_36313,N_36647);
nor U39889 (N_39889,N_36482,N_36702);
and U39890 (N_39890,N_37522,N_36543);
xnor U39891 (N_39891,N_37451,N_36635);
nand U39892 (N_39892,N_36850,N_36321);
nand U39893 (N_39893,N_36870,N_37448);
nor U39894 (N_39894,N_36403,N_37117);
nor U39895 (N_39895,N_36553,N_36063);
nor U39896 (N_39896,N_37899,N_37860);
xnor U39897 (N_39897,N_36440,N_37931);
or U39898 (N_39898,N_37763,N_37376);
or U39899 (N_39899,N_36807,N_36610);
nand U39900 (N_39900,N_37982,N_36354);
nand U39901 (N_39901,N_37223,N_37364);
and U39902 (N_39902,N_36277,N_37158);
or U39903 (N_39903,N_37710,N_37462);
xor U39904 (N_39904,N_36344,N_37075);
nor U39905 (N_39905,N_37477,N_37505);
nand U39906 (N_39906,N_37918,N_37875);
nand U39907 (N_39907,N_37903,N_37706);
and U39908 (N_39908,N_37505,N_36654);
or U39909 (N_39909,N_36412,N_36331);
nand U39910 (N_39910,N_37624,N_36952);
or U39911 (N_39911,N_36050,N_37960);
nor U39912 (N_39912,N_36296,N_36375);
or U39913 (N_39913,N_36701,N_37936);
nand U39914 (N_39914,N_36483,N_36794);
nand U39915 (N_39915,N_36704,N_37808);
or U39916 (N_39916,N_36377,N_36952);
nor U39917 (N_39917,N_37504,N_36336);
nand U39918 (N_39918,N_37378,N_36704);
or U39919 (N_39919,N_37358,N_36806);
and U39920 (N_39920,N_37132,N_36228);
or U39921 (N_39921,N_37218,N_36909);
and U39922 (N_39922,N_37228,N_36019);
and U39923 (N_39923,N_37506,N_36081);
and U39924 (N_39924,N_36548,N_37268);
or U39925 (N_39925,N_37141,N_37542);
xor U39926 (N_39926,N_36831,N_36083);
nand U39927 (N_39927,N_36991,N_37712);
and U39928 (N_39928,N_36346,N_36900);
xnor U39929 (N_39929,N_37950,N_37862);
xor U39930 (N_39930,N_37054,N_36153);
and U39931 (N_39931,N_36913,N_36518);
nand U39932 (N_39932,N_37242,N_37776);
or U39933 (N_39933,N_37274,N_37358);
nand U39934 (N_39934,N_37670,N_37336);
nor U39935 (N_39935,N_36254,N_37098);
and U39936 (N_39936,N_36404,N_37803);
xnor U39937 (N_39937,N_37278,N_37639);
and U39938 (N_39938,N_36081,N_36407);
and U39939 (N_39939,N_37075,N_37842);
and U39940 (N_39940,N_36921,N_37469);
or U39941 (N_39941,N_36866,N_37295);
or U39942 (N_39942,N_36141,N_37088);
nor U39943 (N_39943,N_37774,N_36649);
nand U39944 (N_39944,N_36074,N_36375);
nor U39945 (N_39945,N_36165,N_37684);
nor U39946 (N_39946,N_37757,N_36826);
xor U39947 (N_39947,N_37511,N_37782);
nor U39948 (N_39948,N_36394,N_36445);
and U39949 (N_39949,N_36381,N_36035);
xnor U39950 (N_39950,N_36523,N_37098);
or U39951 (N_39951,N_36079,N_36328);
xnor U39952 (N_39952,N_36325,N_36337);
nand U39953 (N_39953,N_36180,N_36518);
and U39954 (N_39954,N_37542,N_37227);
xor U39955 (N_39955,N_36069,N_37099);
or U39956 (N_39956,N_37745,N_37376);
or U39957 (N_39957,N_36426,N_36291);
xnor U39958 (N_39958,N_36034,N_37058);
nor U39959 (N_39959,N_36644,N_36026);
nor U39960 (N_39960,N_36981,N_36188);
nor U39961 (N_39961,N_37107,N_37186);
nand U39962 (N_39962,N_37689,N_37796);
nor U39963 (N_39963,N_37771,N_36382);
and U39964 (N_39964,N_36712,N_36156);
or U39965 (N_39965,N_36639,N_37913);
or U39966 (N_39966,N_37889,N_37634);
nor U39967 (N_39967,N_37641,N_36564);
xnor U39968 (N_39968,N_36725,N_36812);
and U39969 (N_39969,N_37240,N_36441);
xor U39970 (N_39970,N_37256,N_36743);
nand U39971 (N_39971,N_36067,N_37984);
xor U39972 (N_39972,N_37004,N_37367);
xnor U39973 (N_39973,N_37754,N_36399);
and U39974 (N_39974,N_37457,N_37381);
nand U39975 (N_39975,N_37751,N_36417);
nand U39976 (N_39976,N_37288,N_36403);
and U39977 (N_39977,N_37322,N_37017);
and U39978 (N_39978,N_36735,N_36296);
xnor U39979 (N_39979,N_37128,N_36901);
nand U39980 (N_39980,N_37779,N_37741);
or U39981 (N_39981,N_36514,N_36017);
and U39982 (N_39982,N_37134,N_37071);
nand U39983 (N_39983,N_36798,N_37481);
nor U39984 (N_39984,N_36969,N_37890);
nor U39985 (N_39985,N_36067,N_36076);
or U39986 (N_39986,N_36952,N_37712);
xnor U39987 (N_39987,N_36583,N_36900);
xor U39988 (N_39988,N_36771,N_37618);
or U39989 (N_39989,N_36760,N_37489);
or U39990 (N_39990,N_36806,N_37247);
xnor U39991 (N_39991,N_36384,N_36363);
and U39992 (N_39992,N_36226,N_37932);
and U39993 (N_39993,N_37613,N_36560);
nor U39994 (N_39994,N_36367,N_37716);
nand U39995 (N_39995,N_37225,N_36995);
xnor U39996 (N_39996,N_36052,N_37437);
nand U39997 (N_39997,N_36164,N_37041);
or U39998 (N_39998,N_37072,N_37467);
nor U39999 (N_39999,N_37144,N_36863);
and U40000 (N_40000,N_39544,N_38593);
nor U40001 (N_40001,N_38331,N_39465);
nand U40002 (N_40002,N_39485,N_38700);
and U40003 (N_40003,N_39385,N_39846);
xnor U40004 (N_40004,N_39219,N_38466);
nand U40005 (N_40005,N_38195,N_39608);
nor U40006 (N_40006,N_38302,N_38543);
or U40007 (N_40007,N_39508,N_38896);
nor U40008 (N_40008,N_39640,N_39678);
nand U40009 (N_40009,N_39979,N_39148);
or U40010 (N_40010,N_38962,N_39830);
nand U40011 (N_40011,N_39627,N_39383);
nand U40012 (N_40012,N_39428,N_38831);
or U40013 (N_40013,N_39228,N_38203);
and U40014 (N_40014,N_38645,N_39123);
or U40015 (N_40015,N_38018,N_38559);
nand U40016 (N_40016,N_39154,N_39657);
xnor U40017 (N_40017,N_38628,N_38855);
nand U40018 (N_40018,N_38416,N_39201);
and U40019 (N_40019,N_38879,N_39746);
or U40020 (N_40020,N_39269,N_38950);
or U40021 (N_40021,N_38997,N_38754);
or U40022 (N_40022,N_39563,N_38257);
xor U40023 (N_40023,N_38961,N_38605);
or U40024 (N_40024,N_39764,N_39570);
and U40025 (N_40025,N_39361,N_38650);
xnor U40026 (N_40026,N_38584,N_39708);
nor U40027 (N_40027,N_39929,N_38964);
or U40028 (N_40028,N_39005,N_39324);
xnor U40029 (N_40029,N_38782,N_38552);
or U40030 (N_40030,N_38542,N_38457);
nand U40031 (N_40031,N_38901,N_38238);
nand U40032 (N_40032,N_38285,N_38274);
or U40033 (N_40033,N_38536,N_39216);
and U40034 (N_40034,N_39258,N_39651);
or U40035 (N_40035,N_38159,N_38732);
xnor U40036 (N_40036,N_39558,N_38562);
and U40037 (N_40037,N_39514,N_38833);
or U40038 (N_40038,N_39593,N_39326);
and U40039 (N_40039,N_39480,N_39643);
nand U40040 (N_40040,N_38882,N_39795);
nand U40041 (N_40041,N_38972,N_38503);
and U40042 (N_40042,N_38734,N_39995);
or U40043 (N_40043,N_39623,N_39065);
and U40044 (N_40044,N_39461,N_39016);
nand U40045 (N_40045,N_38380,N_39373);
and U40046 (N_40046,N_38521,N_38321);
nand U40047 (N_40047,N_39853,N_39624);
xor U40048 (N_40048,N_39828,N_39701);
nor U40049 (N_40049,N_38277,N_39015);
nand U40050 (N_40050,N_38809,N_39868);
nor U40051 (N_40051,N_39445,N_39852);
or U40052 (N_40052,N_39063,N_39820);
nand U40053 (N_40053,N_38804,N_39547);
or U40054 (N_40054,N_38706,N_39191);
or U40055 (N_40055,N_38060,N_38468);
nand U40056 (N_40056,N_39441,N_39838);
xor U40057 (N_40057,N_39469,N_39859);
nor U40058 (N_40058,N_39376,N_38318);
and U40059 (N_40059,N_39943,N_38307);
xor U40060 (N_40060,N_39082,N_39215);
xnor U40061 (N_40061,N_39128,N_39030);
nand U40062 (N_40062,N_39458,N_38558);
nand U40063 (N_40063,N_39909,N_39032);
and U40064 (N_40064,N_39025,N_39143);
and U40065 (N_40065,N_39520,N_38270);
nand U40066 (N_40066,N_38723,N_39295);
or U40067 (N_40067,N_38191,N_38422);
nand U40068 (N_40068,N_38472,N_38927);
and U40069 (N_40069,N_39056,N_38080);
xor U40070 (N_40070,N_39773,N_39618);
nor U40071 (N_40071,N_38737,N_39038);
xor U40072 (N_40072,N_38414,N_38792);
and U40073 (N_40073,N_38642,N_38326);
nor U40074 (N_40074,N_39274,N_39387);
xor U40075 (N_40075,N_38504,N_39546);
nor U40076 (N_40076,N_39422,N_38739);
xor U40077 (N_40077,N_39724,N_39778);
or U40078 (N_40078,N_39367,N_38899);
nor U40079 (N_40079,N_38527,N_39506);
and U40080 (N_40080,N_39247,N_39450);
nand U40081 (N_40081,N_38058,N_38614);
nand U40082 (N_40082,N_39914,N_38954);
or U40083 (N_40083,N_38683,N_38785);
xor U40084 (N_40084,N_38462,N_39847);
xor U40085 (N_40085,N_38924,N_38673);
nand U40086 (N_40086,N_39007,N_39069);
or U40087 (N_40087,N_39446,N_39978);
nor U40088 (N_40088,N_38555,N_39283);
nor U40089 (N_40089,N_38115,N_38801);
nand U40090 (N_40090,N_38398,N_39109);
nor U40091 (N_40091,N_39139,N_38744);
xnor U40092 (N_40092,N_38769,N_39682);
and U40093 (N_40093,N_39741,N_39991);
xnor U40094 (N_40094,N_38889,N_38418);
or U40095 (N_40095,N_39865,N_39052);
nor U40096 (N_40096,N_39581,N_38288);
xor U40097 (N_40097,N_39960,N_38629);
xnor U40098 (N_40098,N_39060,N_39039);
xnor U40099 (N_40099,N_38498,N_38222);
and U40100 (N_40100,N_38588,N_38677);
or U40101 (N_40101,N_39931,N_39115);
nor U40102 (N_40102,N_39177,N_38531);
and U40103 (N_40103,N_38190,N_39070);
xor U40104 (N_40104,N_39455,N_38768);
nor U40105 (N_40105,N_39013,N_38862);
nor U40106 (N_40106,N_38158,N_39529);
or U40107 (N_40107,N_39769,N_38750);
nor U40108 (N_40108,N_39181,N_39055);
and U40109 (N_40109,N_38082,N_38685);
nand U40110 (N_40110,N_39475,N_39925);
nand U40111 (N_40111,N_39084,N_39057);
nand U40112 (N_40112,N_39111,N_39067);
nand U40113 (N_40113,N_38044,N_38957);
or U40114 (N_40114,N_38884,N_38229);
or U40115 (N_40115,N_39183,N_39474);
xnor U40116 (N_40116,N_39410,N_38424);
nand U40117 (N_40117,N_38956,N_39249);
or U40118 (N_40118,N_39604,N_39275);
and U40119 (N_40119,N_39281,N_39985);
and U40120 (N_40120,N_38161,N_38590);
or U40121 (N_40121,N_38039,N_39483);
xnor U40122 (N_40122,N_39142,N_38284);
xnor U40123 (N_40123,N_39615,N_38660);
xnor U40124 (N_40124,N_39347,N_39849);
and U40125 (N_40125,N_39531,N_39433);
or U40126 (N_40126,N_39008,N_39185);
or U40127 (N_40127,N_39806,N_38120);
or U40128 (N_40128,N_38054,N_39649);
and U40129 (N_40129,N_39759,N_39045);
and U40130 (N_40130,N_39158,N_39346);
nor U40131 (N_40131,N_39218,N_38143);
nor U40132 (N_40132,N_38554,N_39522);
nor U40133 (N_40133,N_38929,N_38985);
xnor U40134 (N_40134,N_38824,N_38902);
nand U40135 (N_40135,N_39756,N_39232);
and U40136 (N_40136,N_39194,N_39074);
nand U40137 (N_40137,N_38881,N_38266);
xor U40138 (N_40138,N_39681,N_38609);
or U40139 (N_40139,N_39356,N_39954);
xor U40140 (N_40140,N_39323,N_39389);
xnor U40141 (N_40141,N_38295,N_39984);
xor U40142 (N_40142,N_39031,N_38800);
nand U40143 (N_40143,N_39166,N_38421);
nor U40144 (N_40144,N_39730,N_38453);
xor U40145 (N_40145,N_38656,N_39377);
and U40146 (N_40146,N_38979,N_38539);
or U40147 (N_40147,N_38196,N_39368);
xnor U40148 (N_40148,N_38779,N_38217);
nor U40149 (N_40149,N_39336,N_38566);
or U40150 (N_40150,N_38933,N_39573);
xor U40151 (N_40151,N_38601,N_38168);
xor U40152 (N_40152,N_39340,N_38965);
or U40153 (N_40153,N_39878,N_38033);
nor U40154 (N_40154,N_38736,N_39692);
xnor U40155 (N_40155,N_38662,N_38727);
and U40156 (N_40156,N_38808,N_38514);
nor U40157 (N_40157,N_38942,N_38960);
nor U40158 (N_40158,N_39226,N_38124);
nor U40159 (N_40159,N_39941,N_39910);
or U40160 (N_40160,N_39350,N_38166);
xor U40161 (N_40161,N_38306,N_38897);
nor U40162 (N_40162,N_38205,N_38846);
and U40163 (N_40163,N_39983,N_38705);
and U40164 (N_40164,N_39528,N_39525);
nand U40165 (N_40165,N_39947,N_39816);
or U40166 (N_40166,N_38894,N_39685);
nand U40167 (N_40167,N_38001,N_39767);
or U40168 (N_40168,N_38218,N_39918);
nor U40169 (N_40169,N_39920,N_38572);
xnor U40170 (N_40170,N_38814,N_38339);
nor U40171 (N_40171,N_38608,N_39120);
or U40172 (N_40172,N_39845,N_38637);
or U40173 (N_40173,N_38821,N_39851);
or U40174 (N_40174,N_38878,N_38286);
xnor U40175 (N_40175,N_38387,N_39321);
xor U40176 (N_40176,N_38621,N_38141);
nor U40177 (N_40177,N_38915,N_39409);
xor U40178 (N_40178,N_39273,N_38099);
nor U40179 (N_40179,N_38016,N_39230);
nand U40180 (N_40180,N_38299,N_39584);
and U40181 (N_40181,N_38496,N_39899);
nor U40182 (N_40182,N_39707,N_38027);
xnor U40183 (N_40183,N_38223,N_38056);
and U40184 (N_40184,N_39398,N_38234);
or U40185 (N_40185,N_39279,N_39253);
nor U40186 (N_40186,N_38130,N_38678);
and U40187 (N_40187,N_39205,N_38428);
nand U40188 (N_40188,N_38771,N_38322);
or U40189 (N_40189,N_38759,N_39538);
nor U40190 (N_40190,N_39526,N_39020);
nand U40191 (N_40191,N_39975,N_38697);
nor U40192 (N_40192,N_38966,N_39319);
or U40193 (N_40193,N_39904,N_39535);
or U40194 (N_40194,N_39872,N_38912);
nand U40195 (N_40195,N_38169,N_38085);
nor U40196 (N_40196,N_38842,N_39486);
nand U40197 (N_40197,N_39196,N_38072);
and U40198 (N_40198,N_39251,N_39192);
or U40199 (N_40199,N_39690,N_39470);
and U40200 (N_40200,N_38999,N_39698);
and U40201 (N_40201,N_38361,N_39532);
nor U40202 (N_40202,N_39857,N_38308);
and U40203 (N_40203,N_38653,N_38461);
nand U40204 (N_40204,N_39245,N_39411);
and U40205 (N_40205,N_38061,N_39588);
and U40206 (N_40206,N_39293,N_39507);
nor U40207 (N_40207,N_39444,N_38908);
and U40208 (N_40208,N_38372,N_39309);
xnor U40209 (N_40209,N_38606,N_38078);
and U40210 (N_40210,N_39793,N_38256);
nand U40211 (N_40211,N_38490,N_38740);
and U40212 (N_40212,N_38332,N_38548);
nand U40213 (N_40213,N_39337,N_39949);
nor U40214 (N_40214,N_39802,N_38847);
and U40215 (N_40215,N_39772,N_39203);
nor U40216 (N_40216,N_38731,N_38093);
and U40217 (N_40217,N_39271,N_38793);
nor U40218 (N_40218,N_39568,N_39787);
and U40219 (N_40219,N_38427,N_38356);
nor U40220 (N_40220,N_39644,N_38029);
xor U40221 (N_40221,N_38176,N_38200);
nand U40222 (N_40222,N_38703,N_39944);
and U40223 (N_40223,N_39147,N_38350);
xor U40224 (N_40224,N_39647,N_38946);
xor U40225 (N_40225,N_39453,N_38360);
or U40226 (N_40226,N_38556,N_39727);
nor U40227 (N_40227,N_38474,N_39962);
nand U40228 (N_40228,N_39945,N_38377);
or U40229 (N_40229,N_38921,N_38487);
nand U40230 (N_40230,N_39482,N_38760);
nand U40231 (N_40231,N_38941,N_39355);
xnor U40232 (N_40232,N_39571,N_39360);
xnor U40233 (N_40233,N_39262,N_39138);
or U40234 (N_40234,N_38136,N_39722);
and U40235 (N_40235,N_38146,N_38342);
xor U40236 (N_40236,N_39322,N_38850);
xnor U40237 (N_40237,N_39823,N_39102);
or U40238 (N_40238,N_39992,N_38478);
nand U40239 (N_40239,N_39462,N_39108);
and U40240 (N_40240,N_38355,N_38042);
xor U40241 (N_40241,N_38005,N_39178);
nor U40242 (N_40242,N_39782,N_39189);
and U40243 (N_40243,N_39753,N_38682);
or U40244 (N_40244,N_39221,N_39856);
and U40245 (N_40245,N_39699,N_38989);
nor U40246 (N_40246,N_39748,N_39905);
xor U40247 (N_40247,N_38240,N_38892);
xor U40248 (N_40248,N_39210,N_39307);
nor U40249 (N_40249,N_39233,N_39654);
xor U40250 (N_40250,N_38173,N_39705);
nand U40251 (N_40251,N_38907,N_38669);
nor U40252 (N_40252,N_39098,N_38599);
or U40253 (N_40253,N_38518,N_38788);
nand U40254 (N_40254,N_39740,N_39035);
xnor U40255 (N_40255,N_38108,N_39897);
nor U40256 (N_40256,N_38224,N_38425);
xor U40257 (N_40257,N_39695,N_38188);
nor U40258 (N_40258,N_38951,N_39915);
or U40259 (N_40259,N_38932,N_39107);
xnor U40260 (N_40260,N_38171,N_39993);
xor U40261 (N_40261,N_38037,N_38362);
nand U40262 (N_40262,N_39449,N_38103);
xnor U40263 (N_40263,N_39917,N_38272);
nor U40264 (N_40264,N_39146,N_39404);
nor U40265 (N_40265,N_39501,N_39677);
and U40266 (N_40266,N_38340,N_38963);
or U40267 (N_40267,N_39997,N_39697);
or U40268 (N_40268,N_39184,N_38648);
xnor U40269 (N_40269,N_39548,N_39413);
xnor U40270 (N_40270,N_38297,N_39700);
and U40271 (N_40271,N_38649,N_38646);
and U40272 (N_40272,N_38106,N_38413);
xor U40273 (N_40273,N_39110,N_39155);
or U40274 (N_40274,N_38402,N_38347);
or U40275 (N_40275,N_38097,N_38305);
nand U40276 (N_40276,N_39238,N_39371);
or U40277 (N_40277,N_38442,N_39399);
nand U40278 (N_40278,N_39352,N_38119);
xor U40279 (N_40279,N_39041,N_39620);
nand U40280 (N_40280,N_38247,N_38470);
nand U40281 (N_40281,N_38412,N_39592);
and U40282 (N_40282,N_38829,N_38631);
and U40283 (N_40283,N_38110,N_39405);
nand U40284 (N_40284,N_39105,N_39390);
nand U40285 (N_40285,N_39605,N_39270);
xnor U40286 (N_40286,N_38845,N_39260);
xor U40287 (N_40287,N_39932,N_38351);
nor U40288 (N_40288,N_39840,N_38565);
or U40289 (N_40289,N_39048,N_38184);
and U40290 (N_40290,N_39564,N_38625);
or U40291 (N_40291,N_39792,N_39438);
xnor U40292 (N_40292,N_39781,N_38452);
and U40293 (N_40293,N_38762,N_38563);
and U40294 (N_40294,N_38681,N_38291);
xnor U40295 (N_40295,N_39254,N_38081);
nand U40296 (N_40296,N_39658,N_39095);
or U40297 (N_40297,N_38944,N_39952);
or U40298 (N_40298,N_38167,N_39933);
and U40299 (N_40299,N_38242,N_38324);
xnor U40300 (N_40300,N_39292,N_39642);
xnor U40301 (N_40301,N_39824,N_38877);
xor U40302 (N_40302,N_39188,N_39619);
and U40303 (N_40303,N_39159,N_38102);
xnor U40304 (N_40304,N_38992,N_38447);
and U40305 (N_40305,N_38463,N_38043);
xnor U40306 (N_40306,N_39661,N_39810);
xnor U40307 (N_40307,N_39716,N_39908);
nor U40308 (N_40308,N_38510,N_38499);
xnor U40309 (N_40309,N_39287,N_39901);
nand U40310 (N_40310,N_38764,N_38079);
or U40311 (N_40311,N_39611,N_39179);
nor U40312 (N_40312,N_38024,N_39870);
nand U40313 (N_40313,N_39328,N_38666);
or U40314 (N_40314,N_38450,N_39112);
or U40315 (N_40315,N_38014,N_38047);
xnor U40316 (N_40316,N_39671,N_38393);
nor U40317 (N_40317,N_38836,N_38987);
and U40318 (N_40318,N_39655,N_38485);
and U40319 (N_40319,N_38893,N_39091);
and U40320 (N_40320,N_39988,N_39382);
and U40321 (N_40321,N_38181,N_39092);
nand U40322 (N_40322,N_39848,N_38010);
and U40323 (N_40323,N_39022,N_38382);
nand U40324 (N_40324,N_38155,N_39175);
and U40325 (N_40325,N_39898,N_39459);
and U40326 (N_40326,N_38651,N_38525);
nor U40327 (N_40327,N_38512,N_39684);
nor U40328 (N_40328,N_38761,N_39841);
or U40329 (N_40329,N_38870,N_39771);
nand U40330 (N_40330,N_39893,N_39660);
or U40331 (N_40331,N_38226,N_38214);
nor U40332 (N_40332,N_38207,N_38886);
and U40333 (N_40333,N_39687,N_39970);
xnor U40334 (N_40334,N_38330,N_38919);
xor U40335 (N_40335,N_38585,N_38945);
nand U40336 (N_40336,N_38128,N_39986);
xnor U40337 (N_40337,N_38235,N_39980);
and U40338 (N_40338,N_38062,N_39419);
xor U40339 (N_40339,N_39311,N_38883);
or U40340 (N_40340,N_38509,N_38185);
xnor U40341 (N_40341,N_38445,N_38652);
or U40342 (N_40342,N_38564,N_38349);
nor U40343 (N_40343,N_38125,N_39044);
or U40344 (N_40344,N_38797,N_39776);
nor U40345 (N_40345,N_38333,N_38654);
xnor U40346 (N_40346,N_38664,N_39613);
nand U40347 (N_40347,N_39648,N_39752);
nand U40348 (N_40348,N_39565,N_38123);
and U40349 (N_40349,N_38852,N_38087);
or U40350 (N_40350,N_38610,N_38827);
nor U40351 (N_40351,N_38368,N_39645);
nor U40352 (N_40352,N_38454,N_38905);
and U40353 (N_40353,N_39327,N_39141);
and U40354 (N_40354,N_38311,N_38210);
and U40355 (N_40355,N_39930,N_39530);
or U40356 (N_40356,N_38507,N_38679);
nor U40357 (N_40357,N_38114,N_38034);
nand U40358 (N_40358,N_38243,N_39276);
nor U40359 (N_40359,N_38871,N_38738);
or U40360 (N_40360,N_38943,N_39585);
and U40361 (N_40361,N_38665,N_38613);
xnor U40362 (N_40362,N_39598,N_38315);
xor U40363 (N_40363,N_38083,N_39173);
or U40364 (N_40364,N_39693,N_38177);
xor U40365 (N_40365,N_39637,N_39521);
xor U40366 (N_40366,N_39042,N_39948);
nand U40367 (N_40367,N_39879,N_38245);
nand U40368 (N_40368,N_39436,N_38689);
nor U40369 (N_40369,N_39892,N_38742);
or U40370 (N_40370,N_39014,N_38157);
nand U40371 (N_40371,N_39332,N_38201);
and U40372 (N_40372,N_38269,N_39672);
nor U40373 (N_40373,N_39523,N_39843);
nor U40374 (N_40374,N_38670,N_39320);
or U40375 (N_40375,N_38611,N_39762);
or U40376 (N_40376,N_38859,N_38502);
xor U40377 (N_40377,N_38696,N_39447);
and U40378 (N_40378,N_38420,N_38598);
nor U40379 (N_40379,N_38948,N_39132);
and U40380 (N_40380,N_39610,N_38105);
and U40381 (N_40381,N_39799,N_38730);
nor U40382 (N_40382,N_39479,N_38122);
xnor U40383 (N_40383,N_38367,N_39935);
xor U40384 (N_40384,N_39452,N_38780);
nand U40385 (N_40385,N_38436,N_38261);
and U40386 (N_40386,N_39811,N_39277);
or U40387 (N_40387,N_39302,N_38456);
and U40388 (N_40388,N_38230,N_38888);
nand U40389 (N_40389,N_38404,N_39348);
nand U40390 (N_40390,N_39435,N_38832);
xnor U40391 (N_40391,N_38647,N_39813);
nor U40392 (N_40392,N_39683,N_39628);
nor U40393 (N_40393,N_38885,N_39875);
xor U40394 (N_40394,N_39308,N_38301);
or U40395 (N_40395,N_39854,N_39263);
nor U40396 (N_40396,N_38505,N_38440);
and U40397 (N_40397,N_38594,N_38383);
or U40398 (N_40398,N_38358,N_38341);
nor U40399 (N_40399,N_38688,N_38517);
and U40400 (N_40400,N_38237,N_38684);
and U40401 (N_40401,N_39464,N_39406);
nand U40402 (N_40402,N_38603,N_39599);
nand U40403 (N_40403,N_39891,N_38763);
and U40404 (N_40404,N_39537,N_38553);
and U40405 (N_40405,N_39488,N_39888);
nand U40406 (N_40406,N_38417,N_39424);
or U40407 (N_40407,N_39539,N_39556);
and U40408 (N_40408,N_39834,N_39403);
xor U40409 (N_40409,N_38091,N_39837);
nand U40410 (N_40410,N_38008,N_38174);
or U40411 (N_40411,N_38492,N_38074);
or U40412 (N_40412,N_39500,N_38506);
nand U40413 (N_40413,N_39807,N_38751);
xnor U40414 (N_40414,N_38092,N_38025);
and U40415 (N_40415,N_39825,N_38117);
xor U40416 (N_40416,N_38783,N_38303);
nor U40417 (N_40417,N_39629,N_38415);
xnor U40418 (N_40418,N_38596,N_38515);
nand U40419 (N_40419,N_38077,N_39751);
xnor U40420 (N_40420,N_39712,N_39476);
or U40421 (N_40421,N_39364,N_39632);
nand U40422 (N_40422,N_39567,N_39517);
or U40423 (N_40423,N_38296,N_38019);
xor U40424 (N_40424,N_38276,N_38426);
and U40425 (N_40425,N_39156,N_38577);
xnor U40426 (N_40426,N_38511,N_39803);
or U40427 (N_40427,N_38695,N_38244);
and U40428 (N_40428,N_38973,N_39938);
and U40429 (N_40429,N_38746,N_38917);
nand U40430 (N_40430,N_38920,N_39577);
nand U40431 (N_40431,N_38163,N_39527);
nor U40432 (N_40432,N_39096,N_38982);
nor U40433 (N_40433,N_38547,N_39460);
or U40434 (N_40434,N_38038,N_39118);
nor U40435 (N_40435,N_38644,N_38142);
or U40436 (N_40436,N_38709,N_39421);
or U40437 (N_40437,N_38071,N_39420);
nand U40438 (N_40438,N_38733,N_38756);
xor U40439 (N_40439,N_39334,N_38813);
xor U40440 (N_40440,N_39089,N_39395);
nand U40441 (N_40441,N_39036,N_38874);
nand U40442 (N_40442,N_39267,N_39939);
xor U40443 (N_40443,N_38796,N_39186);
xor U40444 (N_40444,N_39026,N_38459);
xor U40445 (N_40445,N_38051,N_39796);
nor U40446 (N_40446,N_39490,N_39440);
xor U40447 (N_40447,N_38263,N_39209);
or U40448 (N_40448,N_39703,N_39116);
or U40449 (N_40449,N_39516,N_39609);
nand U40450 (N_40450,N_39443,N_38467);
or U40451 (N_40451,N_39425,N_39075);
nand U40452 (N_40452,N_38994,N_38934);
xor U40453 (N_40453,N_39229,N_39922);
or U40454 (N_40454,N_39626,N_38258);
or U40455 (N_40455,N_39027,N_38493);
xnor U40456 (N_40456,N_38930,N_39207);
xor U40457 (N_40457,N_39250,N_38523);
xor U40458 (N_40458,N_38273,N_39600);
and U40459 (N_40459,N_39457,N_39714);
xnor U40460 (N_40460,N_38617,N_38743);
and U40461 (N_40461,N_39844,N_38403);
xnor U40462 (N_40462,N_38365,N_38620);
or U40463 (N_40463,N_38817,N_39497);
nand U40464 (N_40464,N_39393,N_38289);
or U40465 (N_40465,N_39818,N_38003);
or U40466 (N_40466,N_38784,N_38127);
or U40467 (N_40467,N_38635,N_39887);
xor U40468 (N_40468,N_39912,N_38250);
or U40469 (N_40469,N_39068,N_38352);
xor U40470 (N_40470,N_39085,N_39797);
nor U40471 (N_40471,N_38209,N_39294);
and U40472 (N_40472,N_39214,N_39162);
nor U40473 (N_40473,N_39630,N_39551);
or U40474 (N_40474,N_38795,N_38489);
or U40475 (N_40475,N_39131,N_39342);
xnor U40476 (N_40476,N_39919,N_39890);
nand U40477 (N_40477,N_39959,N_38765);
nor U40478 (N_40478,N_38755,N_38069);
or U40479 (N_40479,N_38345,N_38712);
nor U40480 (N_40480,N_39873,N_39037);
nand U40481 (N_40481,N_39220,N_39963);
nand U40482 (N_40482,N_39656,N_39282);
nand U40483 (N_40483,N_39001,N_39549);
nor U40484 (N_40484,N_39650,N_38002);
and U40485 (N_40485,N_39972,N_39002);
or U40486 (N_40486,N_39955,N_38320);
xor U40487 (N_40487,N_38535,N_38570);
xnor U40488 (N_40488,N_38052,N_39272);
nand U40489 (N_40489,N_39950,N_39053);
or U40490 (N_40490,N_38011,N_39786);
nand U40491 (N_40491,N_39987,N_38815);
and U40492 (N_40492,N_38589,N_38710);
xnor U40493 (N_40493,N_38676,N_39953);
or U40494 (N_40494,N_39686,N_38702);
and U40495 (N_40495,N_39338,N_38189);
nor U40496 (N_40496,N_39244,N_39161);
xor U40497 (N_40497,N_39726,N_39235);
nand U40498 (N_40498,N_39006,N_39241);
and U40499 (N_40499,N_39417,N_38373);
or U40500 (N_40500,N_39386,N_38501);
nor U40501 (N_40501,N_38843,N_39301);
xnor U40502 (N_40502,N_39582,N_38013);
xor U40503 (N_40503,N_38446,N_39896);
nand U40504 (N_40504,N_39004,N_39614);
nand U40505 (N_40505,N_38023,N_38578);
or U40506 (N_40506,N_38508,N_38206);
xor U40507 (N_40507,N_38538,N_39572);
and U40508 (N_40508,N_38281,N_38208);
nand U40509 (N_40509,N_38694,N_39809);
or U40510 (N_40510,N_39638,N_38477);
nor U40511 (N_40511,N_39858,N_38455);
or U40512 (N_40512,N_39426,N_39861);
xnor U40513 (N_40513,N_39193,N_38334);
nor U40514 (N_40514,N_39401,N_39822);
nand U40515 (N_40515,N_38410,N_39408);
nor U40516 (N_40516,N_39554,N_39578);
nand U40517 (N_40517,N_38323,N_39829);
xor U40518 (N_40518,N_39576,N_39903);
nor U40519 (N_40519,N_39296,N_39090);
and U40520 (N_40520,N_38947,N_38991);
nand U40521 (N_40521,N_39855,N_39864);
or U40522 (N_40522,N_38327,N_39553);
nand U40523 (N_40523,N_38668,N_39911);
nor U40524 (N_40524,N_39248,N_38290);
xor U40525 (N_40525,N_39087,N_39400);
and U40526 (N_40526,N_38798,N_39906);
xnor U40527 (N_40527,N_38822,N_39256);
nor U40528 (N_40528,N_38135,N_38781);
nor U40529 (N_40529,N_38838,N_39958);
or U40530 (N_40530,N_38265,N_38232);
xnor U40531 (N_40531,N_39021,N_38026);
nor U40532 (N_40532,N_38260,N_38627);
xor U40533 (N_40533,N_38312,N_39874);
nor U40534 (N_40534,N_38968,N_39761);
nand U40535 (N_40535,N_38519,N_38707);
or U40536 (N_40536,N_39288,N_38280);
nand U40537 (N_40537,N_38748,N_39495);
xor U40538 (N_40538,N_38031,N_39153);
or U40539 (N_40539,N_39560,N_39814);
or U40540 (N_40540,N_39145,N_38483);
or U40541 (N_40541,N_38111,N_39616);
nor U40542 (N_40542,N_38335,N_39804);
nand U40543 (N_40543,N_38622,N_38399);
nand U40544 (N_40544,N_39134,N_38619);
and U40545 (N_40545,N_39487,N_38568);
xnor U40546 (N_40546,N_38970,N_39237);
nor U40547 (N_40547,N_39715,N_39354);
nand U40548 (N_40548,N_39575,N_39040);
or U40549 (N_40549,N_39774,N_39489);
and U40550 (N_40550,N_38595,N_39639);
and U40551 (N_40551,N_39505,N_39492);
nand U40552 (N_40552,N_38179,N_38811);
nor U40553 (N_40553,N_39339,N_38213);
or U40554 (N_40554,N_39977,N_39545);
or U40555 (N_40555,N_39524,N_39885);
or U40556 (N_40556,N_38819,N_39496);
xor U40557 (N_40557,N_38549,N_39836);
or U40558 (N_40558,N_39174,N_39136);
and U40559 (N_40559,N_39504,N_39093);
and U40560 (N_40560,N_38252,N_39511);
xor U40561 (N_40561,N_38239,N_38435);
and U40562 (N_40562,N_38000,N_39329);
and U40563 (N_40563,N_38394,N_38586);
nor U40564 (N_40564,N_38392,N_38036);
nor U40565 (N_40565,N_39928,N_39330);
and U40566 (N_40566,N_39344,N_38346);
xnor U40567 (N_40567,N_38262,N_39003);
nor U40568 (N_40568,N_39827,N_39880);
nor U40569 (N_40569,N_38640,N_38292);
xnor U40570 (N_40570,N_38657,N_38253);
nand U40571 (N_40571,N_39202,N_38204);
or U40572 (N_40572,N_38065,N_39380);
nand U40573 (N_40573,N_38236,N_39043);
nand U40574 (N_40574,N_39937,N_39213);
nor U40575 (N_40575,N_38152,N_38408);
nand U40576 (N_40576,N_39552,N_38587);
and U40577 (N_40577,N_38098,N_39137);
and U40578 (N_40578,N_38820,N_39916);
nor U40579 (N_40579,N_39176,N_38906);
xnor U40580 (N_40580,N_39788,N_38571);
or U40581 (N_40581,N_39314,N_39595);
and U40582 (N_40582,N_38221,N_39491);
nand U40583 (N_40583,N_39135,N_39467);
xnor U40584 (N_40584,N_39631,N_39736);
nand U40585 (N_40585,N_39924,N_39305);
nor U40586 (N_40586,N_38495,N_38104);
nor U40587 (N_40587,N_39821,N_39583);
nand U40588 (N_40588,N_39934,N_39559);
xor U40589 (N_40589,N_39484,N_39757);
nor U40590 (N_40590,N_39499,N_39391);
nor U40591 (N_40591,N_38494,N_38357);
nand U40592 (N_40592,N_38363,N_39881);
or U40593 (N_40593,N_38914,N_38144);
xor U40594 (N_40594,N_38145,N_38041);
nand U40595 (N_40595,N_39086,N_38325);
xnor U40596 (N_40596,N_39513,N_38279);
or U40597 (N_40597,N_38776,N_38856);
xnor U40598 (N_40598,N_39080,N_38940);
or U40599 (N_40599,N_39180,N_38259);
and U40600 (N_40600,N_39167,N_39981);
xnor U40601 (N_40601,N_38766,N_39622);
xnor U40602 (N_40602,N_39009,N_38534);
xnor U40603 (N_40603,N_39882,N_38579);
nand U40604 (N_40604,N_39190,N_39735);
or U40605 (N_40605,N_38928,N_38423);
and U40606 (N_40606,N_38219,N_39812);
nand U40607 (N_40607,N_38215,N_38148);
nor U40608 (N_40608,N_38643,N_38012);
nand U40609 (N_40609,N_38865,N_39378);
nand U40610 (N_40610,N_39133,N_39125);
or U40611 (N_40611,N_39129,N_39617);
nor U40612 (N_40612,N_39612,N_39662);
nand U40613 (N_40613,N_38704,N_38583);
nor U40614 (N_40614,N_38624,N_39169);
and U40615 (N_40615,N_39602,N_38431);
or U40616 (N_40616,N_39783,N_39636);
or U40617 (N_40617,N_38314,N_38154);
or U40618 (N_40618,N_38406,N_38747);
nor U40619 (N_40619,N_39242,N_38317);
xor U40620 (N_40620,N_39240,N_38248);
nor U40621 (N_40621,N_39728,N_38530);
xnor U40622 (N_40622,N_39028,N_39555);
nor U40623 (N_40623,N_39171,N_38868);
or U40624 (N_40624,N_38532,N_38958);
and U40625 (N_40625,N_39097,N_38227);
nand U40626 (N_40626,N_38369,N_39494);
or U40627 (N_40627,N_38395,N_38728);
nor U40628 (N_40628,N_38988,N_38255);
nand U40629 (N_40629,N_38050,N_38658);
xnor U40630 (N_40630,N_39819,N_39099);
nor U40631 (N_40631,N_39366,N_38810);
xor U40632 (N_40632,N_38381,N_38895);
nor U40633 (N_40633,N_38197,N_39280);
and U40634 (N_40634,N_38283,N_38839);
nor U40635 (N_40635,N_38094,N_38116);
and U40636 (N_40636,N_38486,N_39396);
nor U40637 (N_40637,N_39737,N_38156);
and U40638 (N_40638,N_38006,N_39353);
nand U40639 (N_40639,N_39990,N_39734);
nor U40640 (N_40640,N_38867,N_38429);
xnor U40641 (N_40641,N_38767,N_39676);
xor U40642 (N_40642,N_39860,N_38557);
or U40643 (N_40643,N_39743,N_38939);
nand U40644 (N_40644,N_39742,N_38212);
xor U40645 (N_40645,N_39747,N_39266);
nand U40646 (N_40646,N_38186,N_39076);
xnor U40647 (N_40647,N_38790,N_39867);
nand U40648 (N_40648,N_39303,N_39473);
and U40649 (N_40649,N_38537,N_38473);
and U40650 (N_40650,N_39101,N_38089);
or U40651 (N_40651,N_39312,N_39763);
nor U40652 (N_40652,N_38545,N_38757);
and U40653 (N_40653,N_38147,N_39777);
nand U40654 (N_40654,N_39999,N_39286);
nor U40655 (N_40655,N_38913,N_39349);
nor U40656 (N_40656,N_38981,N_39946);
xnor U40657 (N_40657,N_38030,N_38898);
nand U40658 (N_40658,N_39392,N_39493);
or U40659 (N_40659,N_39711,N_39124);
nand U40660 (N_40660,N_39785,N_39359);
nor U40661 (N_40661,N_39510,N_39372);
nor U40662 (N_40662,N_39635,N_39335);
and U40663 (N_40663,N_39994,N_38004);
nand U40664 (N_40664,N_39369,N_39206);
or U40665 (N_40665,N_38246,N_39072);
or U40666 (N_40666,N_39688,N_38675);
nand U40667 (N_40667,N_38522,N_38995);
xnor U40668 (N_40668,N_38851,N_38983);
xnor U40669 (N_40669,N_39760,N_38419);
xor U40670 (N_40670,N_38112,N_38986);
or U40671 (N_40671,N_39083,N_39961);
nand U40672 (N_40672,N_39088,N_38132);
xnor U40673 (N_40673,N_39871,N_38708);
nor U40674 (N_40674,N_38095,N_38866);
xnor U40675 (N_40675,N_39427,N_39313);
nor U40676 (N_40676,N_38618,N_38343);
and U40677 (N_40677,N_39691,N_38837);
or U40678 (N_40678,N_39942,N_38729);
or U40679 (N_40679,N_38480,N_38691);
nor U40680 (N_40680,N_39050,N_39317);
and U40681 (N_40681,N_38687,N_38741);
nand U40682 (N_40682,N_39754,N_39877);
nor U40683 (N_40683,N_38672,N_38978);
nand U40684 (N_40684,N_38581,N_39432);
nand U40685 (N_40685,N_38816,N_38497);
or U40686 (N_40686,N_38546,N_38268);
and U40687 (N_40687,N_38969,N_38353);
or U40688 (N_40688,N_38967,N_38384);
or U40689 (N_40689,N_39884,N_38374);
xor U40690 (N_40690,N_39315,N_39866);
and U40691 (N_40691,N_38726,N_38984);
xnor U40692 (N_40692,N_38225,N_38149);
and U40693 (N_40693,N_38432,N_38922);
nor U40694 (N_40694,N_38977,N_38469);
nand U40695 (N_40695,N_38828,N_39217);
and U40696 (N_40696,N_39130,N_39729);
nand U40697 (N_40697,N_39478,N_38778);
xor U40698 (N_40698,N_39850,N_39379);
xnor U40699 (N_40699,N_38304,N_38890);
or U40700 (N_40700,N_39375,N_39160);
nand U40701 (N_40701,N_38375,N_38385);
or U40702 (N_40702,N_39374,N_38430);
xor U40703 (N_40703,N_38582,N_39394);
and U40704 (N_40704,N_39755,N_39832);
xor U40705 (N_40705,N_38164,N_38550);
nor U40706 (N_40706,N_38465,N_39264);
and U40707 (N_40707,N_39310,N_39255);
and U40708 (N_40708,N_39512,N_39017);
nand U40709 (N_40709,N_39029,N_39151);
nor U40710 (N_40710,N_39224,N_39587);
nand U40711 (N_40711,N_39114,N_39634);
nand U40712 (N_40712,N_39779,N_39739);
xor U40713 (N_40713,N_39826,N_39704);
and U40714 (N_40714,N_38998,N_38528);
or U40715 (N_40715,N_39252,N_38777);
nand U40716 (N_40716,N_38251,N_38389);
and U40717 (N_40717,N_39550,N_39749);
nor U40718 (N_40718,N_39212,N_38411);
nor U40719 (N_40719,N_38719,N_38386);
nor U40720 (N_40720,N_38575,N_39325);
or U40721 (N_40721,N_39557,N_39718);
nand U40722 (N_40722,N_39223,N_39594);
nor U40723 (N_40723,N_38923,N_39345);
and U40724 (N_40724,N_39341,N_39725);
nor U40725 (N_40725,N_38067,N_38137);
and U40726 (N_40726,N_39434,N_38667);
nor U40727 (N_40727,N_39049,N_38786);
or U40728 (N_40728,N_39291,N_39964);
nand U40729 (N_40729,N_38160,N_38220);
nor U40730 (N_40730,N_39717,N_39603);
nor U40731 (N_40731,N_38316,N_38900);
nand U40732 (N_40732,N_39936,N_38659);
or U40733 (N_40733,N_38597,N_39306);
and U40734 (N_40734,N_39236,N_38671);
nand U40735 (N_40735,N_38275,N_39163);
nor U40736 (N_40736,N_39702,N_39199);
xnor U40737 (N_40737,N_39641,N_39104);
and U40738 (N_40738,N_39831,N_38264);
nor U40739 (N_40739,N_39876,N_39668);
or U40740 (N_40740,N_39710,N_38359);
nand U40741 (N_40741,N_39680,N_39018);
and U40742 (N_40742,N_38633,N_38909);
and U40743 (N_40743,N_39384,N_38448);
nand U40744 (N_40744,N_39081,N_38231);
xor U40745 (N_40745,N_38853,N_39051);
or U40746 (N_40746,N_39569,N_38861);
nand U40747 (N_40747,N_38153,N_38444);
and U40748 (N_40748,N_39974,N_38513);
or U40749 (N_40749,N_39119,N_39808);
nand U40750 (N_40750,N_39590,N_38282);
and U40751 (N_40751,N_38714,N_38772);
xnor U40752 (N_40752,N_38192,N_39299);
or U40753 (N_40753,N_38309,N_38370);
and U40754 (N_40754,N_39407,N_38053);
nand U40755 (N_40755,N_39140,N_38980);
nand U40756 (N_40756,N_39957,N_39454);
nand U40757 (N_40757,N_38996,N_38602);
nor U40758 (N_40758,N_39062,N_38720);
or U40759 (N_40759,N_39973,N_39333);
nand U40760 (N_40760,N_38376,N_39534);
or U40761 (N_40761,N_39121,N_39996);
xnor U40762 (N_40762,N_39894,N_39046);
nor U40763 (N_40763,N_39418,N_39078);
nor U40764 (N_40764,N_39103,N_39106);
xnor U40765 (N_40765,N_38482,N_38133);
nor U40766 (N_40766,N_39515,N_39694);
and U40767 (N_40767,N_39768,N_38600);
and U40768 (N_40768,N_38287,N_39239);
nor U40769 (N_40769,N_39669,N_38770);
nor U40770 (N_40770,N_38835,N_38910);
nand U40771 (N_40771,N_39388,N_39540);
xnor U40772 (N_40772,N_38278,N_38107);
nand U40773 (N_40773,N_39331,N_39073);
nor U40774 (N_40774,N_39061,N_38066);
nand U40775 (N_40775,N_38749,N_38063);
nand U40776 (N_40776,N_39211,N_38544);
nor U40777 (N_40777,N_39471,N_39625);
or U40778 (N_40778,N_38955,N_39113);
nor U40779 (N_40779,N_38854,N_39149);
nand U40780 (N_40780,N_39466,N_38400);
or U40781 (N_40781,N_38366,N_38787);
or U40782 (N_40782,N_38388,N_39503);
nand U40783 (N_40783,N_39198,N_39227);
nand U40784 (N_40784,N_38860,N_38165);
or U40785 (N_40785,N_39775,N_38849);
xnor U40786 (N_40786,N_38604,N_39182);
and U40787 (N_40787,N_39208,N_38397);
nand U40788 (N_40788,N_39956,N_38294);
or U40789 (N_40789,N_39071,N_38918);
xnor U40790 (N_40790,N_38634,N_39863);
or U40791 (N_40791,N_39646,N_39397);
nand U40792 (N_40792,N_39365,N_39745);
nor U40793 (N_40793,N_38500,N_38131);
nand U40794 (N_40794,N_39607,N_38100);
nand U40795 (N_40795,N_39430,N_38698);
xor U40796 (N_40796,N_39351,N_39562);
nand U40797 (N_40797,N_38178,N_38310);
xnor U40798 (N_40798,N_38194,N_39566);
or U40799 (N_40799,N_39058,N_39463);
nand U40800 (N_40800,N_38717,N_38396);
or U40801 (N_40801,N_38344,N_38064);
or U40802 (N_40802,N_38086,N_39670);
nor U40803 (N_40803,N_39416,N_38150);
or U40804 (N_40804,N_38935,N_38328);
xor U40805 (N_40805,N_38925,N_39502);
xnor U40806 (N_40806,N_39415,N_39801);
nand U40807 (N_40807,N_39429,N_39165);
nor U40808 (N_40808,N_39451,N_39789);
nand U40809 (N_40809,N_38401,N_39732);
nand U40810 (N_40810,N_39719,N_38175);
nand U40811 (N_40811,N_38484,N_39204);
or U40812 (N_40812,N_38791,N_38015);
xor U40813 (N_40813,N_39243,N_38319);
xnor U40814 (N_40814,N_38560,N_38834);
or U40815 (N_40815,N_38725,N_39653);
nand U40816 (N_40816,N_39921,N_38735);
xnor U40817 (N_40817,N_38638,N_38615);
nand U40818 (N_40818,N_39839,N_38364);
nor U40819 (N_40819,N_39689,N_38775);
and U40820 (N_40820,N_38113,N_39731);
xor U40821 (N_40821,N_38663,N_38576);
nand U40822 (N_40822,N_39370,N_38211);
xor U40823 (N_40823,N_39157,N_38551);
nor U40824 (N_40824,N_39448,N_39989);
xnor U40825 (N_40825,N_38887,N_38391);
or U40826 (N_40826,N_38692,N_38976);
and U40827 (N_40827,N_38118,N_39363);
or U40828 (N_40828,N_38789,N_39168);
nor U40829 (N_40829,N_38533,N_38434);
xor U40830 (N_40830,N_39094,N_38409);
xor U40831 (N_40831,N_38390,N_39601);
or U40832 (N_40832,N_38674,N_39316);
and U40833 (N_40833,N_38630,N_39765);
xnor U40834 (N_40834,N_38254,N_39589);
or U40835 (N_40835,N_39414,N_38336);
or U40836 (N_40836,N_38880,N_39357);
nor U40837 (N_40837,N_39883,N_38524);
or U40838 (N_40838,N_39034,N_39509);
xnor U40839 (N_40839,N_39431,N_38713);
nor U40840 (N_40840,N_38774,N_39606);
and U40841 (N_40841,N_38873,N_38475);
nor U40842 (N_40842,N_38180,N_39923);
and U40843 (N_40843,N_39150,N_38520);
nand U40844 (N_40844,N_39481,N_39290);
or U40845 (N_40845,N_39126,N_39667);
nand U40846 (N_40846,N_39197,N_38338);
and U40847 (N_40847,N_38573,N_38249);
nor U40848 (N_40848,N_38471,N_38198);
nand U40849 (N_40849,N_38045,N_38830);
and U40850 (N_40850,N_39835,N_39951);
nor U40851 (N_40851,N_38329,N_38202);
nand U40852 (N_40852,N_39663,N_39561);
or U40853 (N_40853,N_38059,N_38271);
xnor U40854 (N_40854,N_39437,N_39721);
xnor U40855 (N_40855,N_38216,N_39172);
or U40856 (N_40856,N_38953,N_38858);
and U40857 (N_40857,N_39542,N_39579);
and U40858 (N_40858,N_39633,N_39596);
nand U40859 (N_40859,N_39127,N_38721);
nor U40860 (N_40860,N_39679,N_38017);
or U40861 (N_40861,N_38233,N_39222);
nor U40862 (N_40862,N_39900,N_39024);
xor U40863 (N_40863,N_38464,N_38172);
nor U40864 (N_40864,N_38076,N_38574);
and U40865 (N_40865,N_39902,N_38020);
xnor U40866 (N_40866,N_39468,N_38458);
nor U40867 (N_40867,N_39591,N_39187);
nand U40868 (N_40868,N_39318,N_39971);
nor U40869 (N_40869,N_39967,N_39927);
or U40870 (N_40870,N_39709,N_39477);
and U40871 (N_40871,N_38378,N_38170);
or U40872 (N_40872,N_38437,N_38869);
nor U40873 (N_40873,N_39278,N_39019);
or U40874 (N_40874,N_38806,N_39077);
nand U40875 (N_40875,N_39666,N_38569);
nor U40876 (N_40876,N_38903,N_39304);
nand U40877 (N_40877,N_38641,N_39621);
xnor U40878 (N_40878,N_38009,N_38049);
or U40879 (N_40879,N_38701,N_39144);
or U40880 (N_40880,N_39442,N_39010);
xnor U40881 (N_40881,N_38876,N_39784);
or U40882 (N_40882,N_39122,N_38623);
nand U40883 (N_40883,N_38516,N_39652);
and U40884 (N_40884,N_38129,N_38526);
and U40885 (N_40885,N_39965,N_38690);
and U40886 (N_40886,N_38844,N_39895);
or U40887 (N_40887,N_39472,N_38863);
nand U40888 (N_40888,N_38540,N_38057);
xnor U40889 (N_40889,N_39833,N_39289);
or U40890 (N_40890,N_38715,N_38443);
nand U40891 (N_40891,N_39012,N_39750);
xnor U40892 (N_40892,N_39064,N_39966);
nor U40893 (N_40893,N_39696,N_39800);
nor U40894 (N_40894,N_38773,N_38718);
nor U40895 (N_40895,N_38567,N_38088);
xnor U40896 (N_40896,N_39439,N_39541);
or U40897 (N_40897,N_38182,N_39225);
nand U40898 (N_40898,N_39152,N_38974);
or U40899 (N_40899,N_38680,N_38993);
xor U40900 (N_40900,N_38758,N_39381);
and U40901 (N_40901,N_38711,N_38857);
nor U40902 (N_40902,N_38101,N_38639);
xnor U40903 (N_40903,N_39574,N_38541);
and U40904 (N_40904,N_39659,N_39285);
and U40905 (N_40905,N_38807,N_38959);
or U40906 (N_40906,N_39794,N_39268);
xnor U40907 (N_40907,N_39968,N_38607);
nor U40908 (N_40908,N_38183,N_38841);
nor U40909 (N_40909,N_39791,N_38904);
xor U40910 (N_40910,N_38716,N_39976);
nand U40911 (N_40911,N_38937,N_39706);
and U40912 (N_40912,N_38438,N_39246);
or U40913 (N_40913,N_38975,N_39798);
or U40914 (N_40914,N_39597,N_39402);
or U40915 (N_40915,N_38745,N_38090);
or U40916 (N_40916,N_38805,N_39261);
and U40917 (N_40917,N_38949,N_39744);
and U40918 (N_40918,N_38476,N_39586);
nor U40919 (N_40919,N_38241,N_38655);
nor U40920 (N_40920,N_38794,N_39456);
and U40921 (N_40921,N_38228,N_39164);
xnor U40922 (N_40922,N_38068,N_38407);
or U40923 (N_40923,N_39284,N_38371);
nor U40924 (N_40924,N_39869,N_39862);
nand U40925 (N_40925,N_38405,N_38848);
nand U40926 (N_40926,N_38891,N_39519);
nor U40927 (N_40927,N_38990,N_38799);
xor U40928 (N_40928,N_39543,N_39675);
xnor U40929 (N_40929,N_39011,N_38451);
nor U40930 (N_40930,N_38722,N_39200);
nor U40931 (N_40931,N_39033,N_39231);
or U40932 (N_40932,N_39170,N_39100);
nand U40933 (N_40933,N_39733,N_38931);
nand U40934 (N_40934,N_38035,N_38046);
or U40935 (N_40935,N_39738,N_38661);
and U40936 (N_40936,N_38139,N_38592);
nor U40937 (N_40937,N_38040,N_39982);
nor U40938 (N_40938,N_38802,N_39913);
and U40939 (N_40939,N_38070,N_39665);
nand U40940 (N_40940,N_38803,N_38379);
xnor U40941 (N_40941,N_38752,N_39758);
nand U40942 (N_40942,N_39423,N_38055);
nand U40943 (N_40943,N_39362,N_39998);
xnor U40944 (N_40944,N_38354,N_38812);
xnor U40945 (N_40945,N_38926,N_38840);
and U40946 (N_40946,N_38561,N_38028);
nor U40947 (N_40947,N_39117,N_39298);
nor U40948 (N_40948,N_38875,N_38084);
xor U40949 (N_40949,N_39343,N_38616);
and U40950 (N_40950,N_39059,N_38313);
nand U40951 (N_40951,N_38439,N_39234);
nand U40952 (N_40952,N_39842,N_38096);
xnor U40953 (N_40953,N_38193,N_39047);
and U40954 (N_40954,N_39713,N_39498);
nand U40955 (N_40955,N_38591,N_39533);
nand U40956 (N_40956,N_38007,N_38048);
nor U40957 (N_40957,N_38936,N_39412);
and U40958 (N_40958,N_38626,N_39674);
nand U40959 (N_40959,N_38724,N_38872);
nor U40960 (N_40960,N_38032,N_38162);
nor U40961 (N_40961,N_38823,N_38636);
and U40962 (N_40962,N_38298,N_39723);
or U40963 (N_40963,N_38126,N_39889);
or U40964 (N_40964,N_38686,N_39969);
xor U40965 (N_40965,N_38938,N_39536);
or U40966 (N_40966,N_38449,N_38134);
or U40967 (N_40967,N_38479,N_39518);
and U40968 (N_40968,N_38021,N_38460);
xnor U40969 (N_40969,N_38971,N_38693);
nor U40970 (N_40970,N_39817,N_39926);
nand U40971 (N_40971,N_38073,N_38911);
or U40972 (N_40972,N_38952,N_38121);
or U40973 (N_40973,N_39940,N_39673);
xor U40974 (N_40974,N_38612,N_39054);
and U40975 (N_40975,N_38199,N_38140);
nand U40976 (N_40976,N_38488,N_39259);
nand U40977 (N_40977,N_39358,N_39079);
xnor U40978 (N_40978,N_38022,N_38481);
or U40979 (N_40979,N_39580,N_39766);
and U40980 (N_40980,N_38529,N_38580);
nor U40981 (N_40981,N_39907,N_38864);
or U40982 (N_40982,N_39780,N_39195);
and U40983 (N_40983,N_39805,N_38826);
and U40984 (N_40984,N_38916,N_39790);
nor U40985 (N_40985,N_38267,N_39815);
and U40986 (N_40986,N_38348,N_38187);
nor U40987 (N_40987,N_39720,N_38825);
nand U40988 (N_40988,N_38632,N_38138);
and U40989 (N_40989,N_39886,N_39300);
xor U40990 (N_40990,N_38753,N_39664);
or U40991 (N_40991,N_39297,N_39257);
or U40992 (N_40992,N_39770,N_38491);
xor U40993 (N_40993,N_38433,N_38441);
and U40994 (N_40994,N_38075,N_39265);
and U40995 (N_40995,N_38337,N_38293);
or U40996 (N_40996,N_38818,N_38300);
or U40997 (N_40997,N_38151,N_38699);
nor U40998 (N_40998,N_38109,N_39066);
or U40999 (N_40999,N_39000,N_39023);
xnor U41000 (N_41000,N_38902,N_39169);
or U41001 (N_41001,N_39068,N_39286);
and U41002 (N_41002,N_39448,N_38056);
and U41003 (N_41003,N_39085,N_38948);
nand U41004 (N_41004,N_38594,N_39879);
or U41005 (N_41005,N_38676,N_38643);
nand U41006 (N_41006,N_39658,N_38453);
and U41007 (N_41007,N_39800,N_39943);
xor U41008 (N_41008,N_38697,N_38527);
nor U41009 (N_41009,N_38694,N_38406);
xnor U41010 (N_41010,N_39885,N_38693);
xor U41011 (N_41011,N_39337,N_38131);
nor U41012 (N_41012,N_38968,N_39468);
nor U41013 (N_41013,N_38049,N_39684);
or U41014 (N_41014,N_39645,N_38354);
or U41015 (N_41015,N_39314,N_38457);
nor U41016 (N_41016,N_38274,N_39264);
nand U41017 (N_41017,N_39066,N_39184);
xor U41018 (N_41018,N_38976,N_38420);
and U41019 (N_41019,N_39609,N_39250);
nor U41020 (N_41020,N_38799,N_39870);
or U41021 (N_41021,N_38118,N_39985);
nand U41022 (N_41022,N_38815,N_39216);
nand U41023 (N_41023,N_38116,N_38923);
or U41024 (N_41024,N_38990,N_39307);
and U41025 (N_41025,N_39675,N_38754);
xor U41026 (N_41026,N_38952,N_39144);
nor U41027 (N_41027,N_38311,N_39755);
xor U41028 (N_41028,N_38179,N_39739);
nor U41029 (N_41029,N_38252,N_38248);
nand U41030 (N_41030,N_39141,N_39479);
and U41031 (N_41031,N_39522,N_39191);
and U41032 (N_41032,N_39491,N_38294);
nand U41033 (N_41033,N_39108,N_39623);
and U41034 (N_41034,N_38891,N_39382);
xnor U41035 (N_41035,N_38970,N_38003);
or U41036 (N_41036,N_39753,N_39994);
or U41037 (N_41037,N_39952,N_39673);
xnor U41038 (N_41038,N_39975,N_39370);
and U41039 (N_41039,N_38829,N_39181);
nor U41040 (N_41040,N_38526,N_39188);
nor U41041 (N_41041,N_38421,N_39342);
or U41042 (N_41042,N_38860,N_39471);
nand U41043 (N_41043,N_39532,N_38563);
and U41044 (N_41044,N_38161,N_39897);
nand U41045 (N_41045,N_38884,N_38428);
nand U41046 (N_41046,N_39740,N_39923);
and U41047 (N_41047,N_38206,N_39566);
xnor U41048 (N_41048,N_38278,N_39213);
nor U41049 (N_41049,N_38467,N_39194);
or U41050 (N_41050,N_39908,N_39369);
nor U41051 (N_41051,N_38114,N_39687);
xnor U41052 (N_41052,N_39271,N_38195);
or U41053 (N_41053,N_39637,N_39682);
and U41054 (N_41054,N_39191,N_39002);
and U41055 (N_41055,N_38410,N_39425);
nand U41056 (N_41056,N_38668,N_39151);
nand U41057 (N_41057,N_39706,N_39597);
or U41058 (N_41058,N_38734,N_39522);
nand U41059 (N_41059,N_39917,N_38255);
nor U41060 (N_41060,N_38002,N_39935);
and U41061 (N_41061,N_38082,N_39718);
and U41062 (N_41062,N_38984,N_38109);
nor U41063 (N_41063,N_39941,N_38169);
and U41064 (N_41064,N_39750,N_38599);
nor U41065 (N_41065,N_38670,N_38974);
nand U41066 (N_41066,N_38614,N_38126);
or U41067 (N_41067,N_39038,N_39362);
xor U41068 (N_41068,N_39772,N_39738);
or U41069 (N_41069,N_39803,N_39813);
xnor U41070 (N_41070,N_39544,N_38170);
xnor U41071 (N_41071,N_39534,N_39537);
xor U41072 (N_41072,N_39491,N_39393);
nor U41073 (N_41073,N_39542,N_39953);
nand U41074 (N_41074,N_38875,N_39733);
nand U41075 (N_41075,N_39487,N_39982);
nor U41076 (N_41076,N_38782,N_38300);
nand U41077 (N_41077,N_39039,N_38988);
xnor U41078 (N_41078,N_39582,N_39316);
or U41079 (N_41079,N_39517,N_38145);
xnor U41080 (N_41080,N_38171,N_38824);
nor U41081 (N_41081,N_39037,N_39507);
or U41082 (N_41082,N_38309,N_39825);
nand U41083 (N_41083,N_38548,N_39183);
and U41084 (N_41084,N_38806,N_39449);
xor U41085 (N_41085,N_38369,N_39949);
xor U41086 (N_41086,N_39051,N_38493);
nand U41087 (N_41087,N_38466,N_38997);
nor U41088 (N_41088,N_38103,N_38828);
xor U41089 (N_41089,N_39640,N_38644);
and U41090 (N_41090,N_38911,N_39435);
xor U41091 (N_41091,N_38775,N_38785);
nand U41092 (N_41092,N_38190,N_39427);
nand U41093 (N_41093,N_39122,N_39856);
nand U41094 (N_41094,N_38229,N_38799);
xnor U41095 (N_41095,N_38609,N_39445);
xor U41096 (N_41096,N_39226,N_39947);
nor U41097 (N_41097,N_39951,N_38319);
or U41098 (N_41098,N_38451,N_39473);
and U41099 (N_41099,N_38013,N_38599);
nand U41100 (N_41100,N_39966,N_39585);
xor U41101 (N_41101,N_39435,N_39603);
nor U41102 (N_41102,N_38121,N_39076);
nand U41103 (N_41103,N_38689,N_38688);
or U41104 (N_41104,N_39985,N_39988);
and U41105 (N_41105,N_39910,N_38587);
xor U41106 (N_41106,N_39491,N_39130);
xor U41107 (N_41107,N_38958,N_39142);
xor U41108 (N_41108,N_39161,N_39043);
nand U41109 (N_41109,N_38038,N_38814);
or U41110 (N_41110,N_39545,N_38013);
xor U41111 (N_41111,N_38365,N_39547);
nand U41112 (N_41112,N_38224,N_39321);
nor U41113 (N_41113,N_38570,N_39523);
or U41114 (N_41114,N_38549,N_39255);
and U41115 (N_41115,N_39534,N_39759);
xor U41116 (N_41116,N_39618,N_39477);
and U41117 (N_41117,N_39517,N_38060);
nor U41118 (N_41118,N_38828,N_39739);
and U41119 (N_41119,N_39457,N_38320);
or U41120 (N_41120,N_38797,N_39808);
or U41121 (N_41121,N_39746,N_38234);
xnor U41122 (N_41122,N_38904,N_38984);
or U41123 (N_41123,N_38022,N_39001);
nor U41124 (N_41124,N_39115,N_38455);
and U41125 (N_41125,N_39166,N_39204);
nand U41126 (N_41126,N_38599,N_38637);
xor U41127 (N_41127,N_39212,N_38152);
nor U41128 (N_41128,N_38110,N_38146);
and U41129 (N_41129,N_38422,N_38585);
nand U41130 (N_41130,N_38645,N_38989);
or U41131 (N_41131,N_39727,N_38067);
nor U41132 (N_41132,N_39210,N_38487);
xnor U41133 (N_41133,N_39454,N_38956);
nor U41134 (N_41134,N_39719,N_39357);
or U41135 (N_41135,N_39982,N_39541);
nor U41136 (N_41136,N_38951,N_38629);
or U41137 (N_41137,N_38225,N_38445);
nor U41138 (N_41138,N_39271,N_38194);
and U41139 (N_41139,N_38823,N_38708);
and U41140 (N_41140,N_38098,N_38368);
xor U41141 (N_41141,N_38121,N_39579);
or U41142 (N_41142,N_38125,N_38973);
and U41143 (N_41143,N_39114,N_38295);
and U41144 (N_41144,N_39480,N_38913);
and U41145 (N_41145,N_39539,N_39512);
xnor U41146 (N_41146,N_39580,N_39482);
nor U41147 (N_41147,N_39967,N_38219);
nor U41148 (N_41148,N_38097,N_39674);
xnor U41149 (N_41149,N_38137,N_38952);
or U41150 (N_41150,N_38169,N_38087);
or U41151 (N_41151,N_38560,N_38607);
nor U41152 (N_41152,N_39830,N_39150);
or U41153 (N_41153,N_39209,N_39487);
and U41154 (N_41154,N_39663,N_38806);
nand U41155 (N_41155,N_39672,N_38381);
nand U41156 (N_41156,N_38261,N_39919);
nor U41157 (N_41157,N_39525,N_38968);
nor U41158 (N_41158,N_38153,N_38030);
and U41159 (N_41159,N_38121,N_39685);
and U41160 (N_41160,N_38734,N_39762);
nor U41161 (N_41161,N_38242,N_39221);
and U41162 (N_41162,N_38077,N_39829);
or U41163 (N_41163,N_38266,N_38357);
nand U41164 (N_41164,N_38838,N_38222);
and U41165 (N_41165,N_39419,N_38570);
or U41166 (N_41166,N_39085,N_39069);
nand U41167 (N_41167,N_38277,N_39304);
nor U41168 (N_41168,N_38067,N_39437);
and U41169 (N_41169,N_38531,N_39412);
and U41170 (N_41170,N_39626,N_38559);
nand U41171 (N_41171,N_38571,N_38545);
xor U41172 (N_41172,N_39722,N_39292);
and U41173 (N_41173,N_39856,N_38689);
nand U41174 (N_41174,N_38027,N_39186);
or U41175 (N_41175,N_39088,N_38785);
nor U41176 (N_41176,N_39363,N_39302);
and U41177 (N_41177,N_38734,N_38785);
or U41178 (N_41178,N_39107,N_38796);
nand U41179 (N_41179,N_38363,N_39686);
nand U41180 (N_41180,N_38892,N_38599);
or U41181 (N_41181,N_39058,N_39122);
and U41182 (N_41182,N_39388,N_38690);
or U41183 (N_41183,N_39766,N_39880);
nand U41184 (N_41184,N_38106,N_38028);
and U41185 (N_41185,N_39222,N_39698);
nand U41186 (N_41186,N_39339,N_39954);
xor U41187 (N_41187,N_38606,N_38985);
nor U41188 (N_41188,N_38771,N_38818);
and U41189 (N_41189,N_38152,N_38962);
and U41190 (N_41190,N_38630,N_38796);
and U41191 (N_41191,N_38165,N_38962);
xor U41192 (N_41192,N_39117,N_38488);
nor U41193 (N_41193,N_38641,N_38107);
nand U41194 (N_41194,N_38786,N_39741);
or U41195 (N_41195,N_39991,N_38670);
nand U41196 (N_41196,N_39461,N_38426);
nor U41197 (N_41197,N_38754,N_38378);
and U41198 (N_41198,N_38564,N_38682);
nand U41199 (N_41199,N_39226,N_39089);
nand U41200 (N_41200,N_39008,N_39609);
xor U41201 (N_41201,N_38552,N_38851);
and U41202 (N_41202,N_39065,N_39155);
and U41203 (N_41203,N_39977,N_38006);
and U41204 (N_41204,N_39361,N_39647);
or U41205 (N_41205,N_38921,N_38834);
nor U41206 (N_41206,N_38630,N_39501);
nand U41207 (N_41207,N_39058,N_38224);
nor U41208 (N_41208,N_38250,N_38710);
nor U41209 (N_41209,N_38002,N_38752);
xor U41210 (N_41210,N_38819,N_39165);
xnor U41211 (N_41211,N_39287,N_38110);
xor U41212 (N_41212,N_39310,N_38133);
or U41213 (N_41213,N_38467,N_39187);
or U41214 (N_41214,N_38227,N_38553);
and U41215 (N_41215,N_39769,N_39170);
xnor U41216 (N_41216,N_38749,N_38754);
xor U41217 (N_41217,N_39140,N_39545);
xor U41218 (N_41218,N_39720,N_38082);
nor U41219 (N_41219,N_39528,N_38218);
nand U41220 (N_41220,N_39752,N_38812);
nand U41221 (N_41221,N_38025,N_39672);
or U41222 (N_41222,N_38713,N_38840);
nor U41223 (N_41223,N_38643,N_38016);
nand U41224 (N_41224,N_38767,N_39953);
and U41225 (N_41225,N_39019,N_38733);
and U41226 (N_41226,N_39440,N_38577);
and U41227 (N_41227,N_38944,N_39074);
and U41228 (N_41228,N_38474,N_39781);
nand U41229 (N_41229,N_38797,N_38331);
and U41230 (N_41230,N_38395,N_39881);
and U41231 (N_41231,N_38926,N_39705);
and U41232 (N_41232,N_39244,N_39641);
nand U41233 (N_41233,N_39844,N_39524);
xor U41234 (N_41234,N_39091,N_38558);
xor U41235 (N_41235,N_38203,N_39148);
or U41236 (N_41236,N_39954,N_38278);
and U41237 (N_41237,N_38435,N_39526);
and U41238 (N_41238,N_38844,N_39724);
nor U41239 (N_41239,N_39651,N_38699);
or U41240 (N_41240,N_38158,N_38053);
and U41241 (N_41241,N_39457,N_39072);
nor U41242 (N_41242,N_39055,N_38885);
nor U41243 (N_41243,N_38460,N_39836);
and U41244 (N_41244,N_39819,N_39889);
nand U41245 (N_41245,N_38085,N_39499);
or U41246 (N_41246,N_39208,N_38059);
nor U41247 (N_41247,N_39428,N_38857);
nand U41248 (N_41248,N_39028,N_38285);
and U41249 (N_41249,N_39406,N_38832);
nor U41250 (N_41250,N_38051,N_39921);
nor U41251 (N_41251,N_39191,N_39708);
nand U41252 (N_41252,N_38961,N_39924);
xor U41253 (N_41253,N_39311,N_39967);
xor U41254 (N_41254,N_39746,N_38827);
and U41255 (N_41255,N_38422,N_39297);
or U41256 (N_41256,N_38084,N_38235);
or U41257 (N_41257,N_38772,N_39599);
and U41258 (N_41258,N_38858,N_38794);
nand U41259 (N_41259,N_39913,N_39719);
nor U41260 (N_41260,N_38535,N_39240);
xnor U41261 (N_41261,N_38657,N_39491);
xnor U41262 (N_41262,N_38912,N_38957);
or U41263 (N_41263,N_39653,N_39598);
and U41264 (N_41264,N_38942,N_39531);
xnor U41265 (N_41265,N_39349,N_38228);
or U41266 (N_41266,N_39396,N_39080);
nor U41267 (N_41267,N_38079,N_38744);
xor U41268 (N_41268,N_39315,N_38702);
nand U41269 (N_41269,N_38910,N_39778);
xnor U41270 (N_41270,N_39939,N_39515);
nor U41271 (N_41271,N_39864,N_39743);
nand U41272 (N_41272,N_38906,N_39926);
nand U41273 (N_41273,N_38994,N_39235);
or U41274 (N_41274,N_38592,N_39620);
xor U41275 (N_41275,N_38360,N_39033);
nand U41276 (N_41276,N_39833,N_38726);
nor U41277 (N_41277,N_39232,N_38163);
nand U41278 (N_41278,N_39755,N_39566);
and U41279 (N_41279,N_38829,N_38710);
nand U41280 (N_41280,N_38726,N_39811);
nand U41281 (N_41281,N_39419,N_39628);
xnor U41282 (N_41282,N_38960,N_38531);
or U41283 (N_41283,N_38500,N_38186);
nand U41284 (N_41284,N_38272,N_39454);
or U41285 (N_41285,N_39671,N_39069);
and U41286 (N_41286,N_39257,N_39089);
or U41287 (N_41287,N_38762,N_38988);
xor U41288 (N_41288,N_39750,N_39627);
or U41289 (N_41289,N_39099,N_38917);
nor U41290 (N_41290,N_38695,N_39551);
nand U41291 (N_41291,N_38259,N_38233);
nand U41292 (N_41292,N_39695,N_38462);
and U41293 (N_41293,N_38888,N_38448);
and U41294 (N_41294,N_38901,N_38268);
nand U41295 (N_41295,N_38414,N_39628);
nand U41296 (N_41296,N_39874,N_39272);
nor U41297 (N_41297,N_38412,N_38227);
xor U41298 (N_41298,N_38919,N_39492);
and U41299 (N_41299,N_38602,N_38913);
nor U41300 (N_41300,N_38831,N_38287);
nand U41301 (N_41301,N_38835,N_39104);
xor U41302 (N_41302,N_39334,N_38647);
xnor U41303 (N_41303,N_39997,N_38689);
nand U41304 (N_41304,N_39585,N_39551);
nor U41305 (N_41305,N_39079,N_38876);
nor U41306 (N_41306,N_38954,N_39091);
nand U41307 (N_41307,N_39023,N_39176);
xor U41308 (N_41308,N_39051,N_38723);
nor U41309 (N_41309,N_38969,N_38190);
nor U41310 (N_41310,N_39606,N_39084);
nor U41311 (N_41311,N_38344,N_39363);
nand U41312 (N_41312,N_39927,N_38167);
xor U41313 (N_41313,N_39974,N_39184);
xnor U41314 (N_41314,N_38750,N_38590);
xnor U41315 (N_41315,N_38026,N_38517);
and U41316 (N_41316,N_39262,N_39648);
and U41317 (N_41317,N_38208,N_39643);
nor U41318 (N_41318,N_39298,N_39664);
or U41319 (N_41319,N_38609,N_38565);
xnor U41320 (N_41320,N_39566,N_38267);
xnor U41321 (N_41321,N_39262,N_38525);
nand U41322 (N_41322,N_39848,N_38189);
nor U41323 (N_41323,N_39443,N_38139);
nor U41324 (N_41324,N_38992,N_38147);
nand U41325 (N_41325,N_38704,N_39910);
or U41326 (N_41326,N_39234,N_38781);
xnor U41327 (N_41327,N_39713,N_38370);
nor U41328 (N_41328,N_38665,N_38195);
and U41329 (N_41329,N_38265,N_38742);
or U41330 (N_41330,N_38702,N_38296);
nand U41331 (N_41331,N_39423,N_39875);
nand U41332 (N_41332,N_38505,N_39958);
and U41333 (N_41333,N_38941,N_38913);
nand U41334 (N_41334,N_39926,N_39551);
nor U41335 (N_41335,N_39508,N_38461);
nand U41336 (N_41336,N_38824,N_38357);
nand U41337 (N_41337,N_39943,N_38489);
or U41338 (N_41338,N_38723,N_38476);
nor U41339 (N_41339,N_39449,N_38969);
and U41340 (N_41340,N_39334,N_38076);
nand U41341 (N_41341,N_38916,N_39670);
or U41342 (N_41342,N_38741,N_39121);
xor U41343 (N_41343,N_38607,N_38719);
nand U41344 (N_41344,N_38772,N_39194);
or U41345 (N_41345,N_38653,N_39397);
and U41346 (N_41346,N_38916,N_38422);
or U41347 (N_41347,N_39969,N_39064);
and U41348 (N_41348,N_38245,N_39975);
or U41349 (N_41349,N_38994,N_39186);
nor U41350 (N_41350,N_38107,N_39323);
xnor U41351 (N_41351,N_39340,N_39212);
nand U41352 (N_41352,N_38289,N_38183);
and U41353 (N_41353,N_39295,N_38216);
or U41354 (N_41354,N_38274,N_39646);
xor U41355 (N_41355,N_38993,N_39359);
xor U41356 (N_41356,N_39686,N_38341);
xnor U41357 (N_41357,N_38974,N_39257);
xor U41358 (N_41358,N_38428,N_38405);
or U41359 (N_41359,N_39472,N_38091);
nor U41360 (N_41360,N_38100,N_39168);
or U41361 (N_41361,N_38390,N_39200);
or U41362 (N_41362,N_38112,N_38770);
and U41363 (N_41363,N_39517,N_39608);
or U41364 (N_41364,N_39064,N_38358);
nor U41365 (N_41365,N_38330,N_38960);
or U41366 (N_41366,N_38279,N_39865);
or U41367 (N_41367,N_39240,N_38918);
nand U41368 (N_41368,N_39191,N_39084);
or U41369 (N_41369,N_39212,N_39299);
nor U41370 (N_41370,N_38005,N_39553);
and U41371 (N_41371,N_39485,N_38842);
and U41372 (N_41372,N_38680,N_39495);
xnor U41373 (N_41373,N_38919,N_38413);
nand U41374 (N_41374,N_39461,N_38896);
or U41375 (N_41375,N_39510,N_38962);
nand U41376 (N_41376,N_38180,N_39442);
xor U41377 (N_41377,N_38793,N_38210);
nor U41378 (N_41378,N_38640,N_39829);
and U41379 (N_41379,N_39289,N_39705);
nor U41380 (N_41380,N_38336,N_38171);
xnor U41381 (N_41381,N_39970,N_39980);
xnor U41382 (N_41382,N_39635,N_39486);
or U41383 (N_41383,N_38231,N_38822);
nor U41384 (N_41384,N_39575,N_38229);
xnor U41385 (N_41385,N_38857,N_39100);
nor U41386 (N_41386,N_39376,N_38072);
and U41387 (N_41387,N_38367,N_39466);
or U41388 (N_41388,N_38421,N_38468);
nor U41389 (N_41389,N_38994,N_39196);
nand U41390 (N_41390,N_39476,N_39797);
or U41391 (N_41391,N_39470,N_39168);
xor U41392 (N_41392,N_39419,N_39034);
and U41393 (N_41393,N_39461,N_39475);
nand U41394 (N_41394,N_39518,N_39849);
or U41395 (N_41395,N_38628,N_39378);
or U41396 (N_41396,N_39133,N_38827);
xnor U41397 (N_41397,N_39096,N_38456);
xnor U41398 (N_41398,N_38972,N_39819);
and U41399 (N_41399,N_38891,N_39007);
or U41400 (N_41400,N_39551,N_39165);
nand U41401 (N_41401,N_38657,N_38116);
and U41402 (N_41402,N_38225,N_39946);
xor U41403 (N_41403,N_38330,N_38206);
and U41404 (N_41404,N_39977,N_38831);
and U41405 (N_41405,N_38962,N_38312);
or U41406 (N_41406,N_38312,N_38168);
xnor U41407 (N_41407,N_38892,N_39249);
nand U41408 (N_41408,N_38362,N_38912);
and U41409 (N_41409,N_38484,N_38958);
nand U41410 (N_41410,N_38344,N_38967);
and U41411 (N_41411,N_38165,N_39413);
nand U41412 (N_41412,N_38505,N_39781);
and U41413 (N_41413,N_38647,N_39511);
nand U41414 (N_41414,N_38302,N_38328);
and U41415 (N_41415,N_38314,N_38088);
and U41416 (N_41416,N_39984,N_38334);
xnor U41417 (N_41417,N_38939,N_39945);
nand U41418 (N_41418,N_39418,N_39817);
xor U41419 (N_41419,N_39398,N_38601);
or U41420 (N_41420,N_39860,N_38876);
or U41421 (N_41421,N_39180,N_39154);
nor U41422 (N_41422,N_38454,N_38139);
nor U41423 (N_41423,N_38377,N_39061);
nand U41424 (N_41424,N_38147,N_39611);
and U41425 (N_41425,N_38208,N_38435);
or U41426 (N_41426,N_39875,N_39299);
nand U41427 (N_41427,N_39651,N_38748);
nand U41428 (N_41428,N_38750,N_38308);
xnor U41429 (N_41429,N_38721,N_38282);
or U41430 (N_41430,N_38495,N_39750);
nor U41431 (N_41431,N_39858,N_39456);
nor U41432 (N_41432,N_38593,N_38772);
and U41433 (N_41433,N_39493,N_38752);
nor U41434 (N_41434,N_39577,N_39878);
xnor U41435 (N_41435,N_39287,N_39369);
xnor U41436 (N_41436,N_38704,N_38939);
and U41437 (N_41437,N_38958,N_38292);
xor U41438 (N_41438,N_39393,N_38899);
xnor U41439 (N_41439,N_38100,N_38202);
and U41440 (N_41440,N_39540,N_38427);
nor U41441 (N_41441,N_38912,N_38737);
and U41442 (N_41442,N_39439,N_39531);
nand U41443 (N_41443,N_39839,N_39937);
or U41444 (N_41444,N_39272,N_39374);
nand U41445 (N_41445,N_39054,N_38646);
xnor U41446 (N_41446,N_38607,N_38022);
or U41447 (N_41447,N_39753,N_39513);
and U41448 (N_41448,N_38348,N_39633);
or U41449 (N_41449,N_38845,N_39846);
and U41450 (N_41450,N_39223,N_39172);
nand U41451 (N_41451,N_39215,N_39033);
and U41452 (N_41452,N_39381,N_39109);
or U41453 (N_41453,N_38685,N_38255);
nor U41454 (N_41454,N_39939,N_38809);
xnor U41455 (N_41455,N_39850,N_39433);
xnor U41456 (N_41456,N_38098,N_38760);
nor U41457 (N_41457,N_38136,N_39596);
nand U41458 (N_41458,N_38327,N_39324);
and U41459 (N_41459,N_39868,N_38651);
xnor U41460 (N_41460,N_39490,N_39472);
or U41461 (N_41461,N_38931,N_39087);
xor U41462 (N_41462,N_39627,N_38238);
and U41463 (N_41463,N_39363,N_38215);
xor U41464 (N_41464,N_39717,N_39739);
xnor U41465 (N_41465,N_38173,N_38640);
or U41466 (N_41466,N_38021,N_39993);
xnor U41467 (N_41467,N_39497,N_39944);
nand U41468 (N_41468,N_39540,N_39155);
nor U41469 (N_41469,N_39227,N_39275);
xor U41470 (N_41470,N_38056,N_39527);
nand U41471 (N_41471,N_38446,N_38859);
nor U41472 (N_41472,N_38594,N_38157);
and U41473 (N_41473,N_39984,N_39442);
or U41474 (N_41474,N_38945,N_39174);
and U41475 (N_41475,N_38456,N_39091);
nor U41476 (N_41476,N_39095,N_39565);
or U41477 (N_41477,N_39632,N_39616);
and U41478 (N_41478,N_38411,N_39643);
nor U41479 (N_41479,N_38755,N_38878);
and U41480 (N_41480,N_38197,N_38690);
or U41481 (N_41481,N_38945,N_38152);
xnor U41482 (N_41482,N_38569,N_38326);
nor U41483 (N_41483,N_38943,N_38215);
or U41484 (N_41484,N_38545,N_39918);
and U41485 (N_41485,N_38857,N_38127);
xnor U41486 (N_41486,N_38011,N_38207);
or U41487 (N_41487,N_39175,N_39340);
and U41488 (N_41488,N_39782,N_39459);
or U41489 (N_41489,N_38178,N_38870);
nand U41490 (N_41490,N_39511,N_38048);
nand U41491 (N_41491,N_38764,N_38215);
xor U41492 (N_41492,N_39491,N_38982);
and U41493 (N_41493,N_38277,N_39144);
xor U41494 (N_41494,N_38443,N_38065);
nor U41495 (N_41495,N_38151,N_39925);
and U41496 (N_41496,N_39635,N_39614);
nor U41497 (N_41497,N_38777,N_38181);
or U41498 (N_41498,N_39558,N_39260);
and U41499 (N_41499,N_38258,N_38874);
and U41500 (N_41500,N_38336,N_38562);
nand U41501 (N_41501,N_39638,N_38036);
nand U41502 (N_41502,N_39470,N_39997);
xor U41503 (N_41503,N_39145,N_38823);
nor U41504 (N_41504,N_39250,N_39562);
or U41505 (N_41505,N_38578,N_38523);
xor U41506 (N_41506,N_39616,N_38106);
nor U41507 (N_41507,N_39226,N_39280);
and U41508 (N_41508,N_39106,N_39516);
and U41509 (N_41509,N_39477,N_39162);
nor U41510 (N_41510,N_38914,N_38566);
nor U41511 (N_41511,N_38636,N_39892);
and U41512 (N_41512,N_38732,N_39542);
nor U41513 (N_41513,N_39093,N_38338);
nand U41514 (N_41514,N_39107,N_39272);
xor U41515 (N_41515,N_39269,N_39604);
or U41516 (N_41516,N_39858,N_39006);
or U41517 (N_41517,N_39128,N_38269);
xor U41518 (N_41518,N_38782,N_38407);
or U41519 (N_41519,N_38383,N_39626);
nor U41520 (N_41520,N_38888,N_39195);
xnor U41521 (N_41521,N_38018,N_39491);
or U41522 (N_41522,N_39892,N_39028);
or U41523 (N_41523,N_38983,N_38763);
xor U41524 (N_41524,N_39094,N_39545);
nand U41525 (N_41525,N_38466,N_38991);
nor U41526 (N_41526,N_39489,N_38993);
or U41527 (N_41527,N_39428,N_38169);
and U41528 (N_41528,N_39667,N_38981);
nand U41529 (N_41529,N_38342,N_39166);
or U41530 (N_41530,N_39270,N_38844);
nor U41531 (N_41531,N_38032,N_38503);
nand U41532 (N_41532,N_39388,N_38158);
or U41533 (N_41533,N_38588,N_38481);
xor U41534 (N_41534,N_38895,N_39367);
nand U41535 (N_41535,N_39714,N_39343);
xor U41536 (N_41536,N_39633,N_38915);
nor U41537 (N_41537,N_39163,N_39446);
or U41538 (N_41538,N_39745,N_39712);
xnor U41539 (N_41539,N_38846,N_39768);
nor U41540 (N_41540,N_39699,N_38624);
and U41541 (N_41541,N_38540,N_38438);
or U41542 (N_41542,N_39741,N_38148);
nand U41543 (N_41543,N_38343,N_39034);
nand U41544 (N_41544,N_38813,N_39322);
and U41545 (N_41545,N_38450,N_39636);
nand U41546 (N_41546,N_38085,N_38141);
nand U41547 (N_41547,N_38806,N_39007);
xor U41548 (N_41548,N_38938,N_39056);
nor U41549 (N_41549,N_38248,N_39650);
and U41550 (N_41550,N_38009,N_39780);
and U41551 (N_41551,N_39012,N_39062);
xor U41552 (N_41552,N_38328,N_39087);
and U41553 (N_41553,N_39754,N_39557);
nand U41554 (N_41554,N_38847,N_38723);
and U41555 (N_41555,N_39049,N_38466);
xor U41556 (N_41556,N_38201,N_38648);
or U41557 (N_41557,N_38665,N_39182);
or U41558 (N_41558,N_38732,N_38510);
or U41559 (N_41559,N_38516,N_39798);
nand U41560 (N_41560,N_39778,N_39156);
or U41561 (N_41561,N_39087,N_39914);
or U41562 (N_41562,N_38478,N_39395);
xor U41563 (N_41563,N_38851,N_39611);
xnor U41564 (N_41564,N_39417,N_39215);
and U41565 (N_41565,N_38441,N_38388);
nand U41566 (N_41566,N_39009,N_39827);
nand U41567 (N_41567,N_38141,N_38973);
nor U41568 (N_41568,N_38984,N_39939);
nand U41569 (N_41569,N_39332,N_39785);
xor U41570 (N_41570,N_38091,N_38923);
and U41571 (N_41571,N_39793,N_38069);
nor U41572 (N_41572,N_38398,N_39483);
or U41573 (N_41573,N_38219,N_38028);
or U41574 (N_41574,N_39682,N_38307);
nor U41575 (N_41575,N_38260,N_38340);
nand U41576 (N_41576,N_38391,N_38302);
and U41577 (N_41577,N_39928,N_38953);
and U41578 (N_41578,N_39416,N_39970);
xnor U41579 (N_41579,N_39524,N_39268);
nor U41580 (N_41580,N_39216,N_38526);
xor U41581 (N_41581,N_38829,N_39003);
or U41582 (N_41582,N_39687,N_38357);
xor U41583 (N_41583,N_39965,N_38818);
nor U41584 (N_41584,N_39783,N_39442);
or U41585 (N_41585,N_38120,N_39372);
xnor U41586 (N_41586,N_39594,N_38508);
or U41587 (N_41587,N_39800,N_38018);
xnor U41588 (N_41588,N_39429,N_38155);
and U41589 (N_41589,N_38042,N_38791);
and U41590 (N_41590,N_38578,N_39074);
nand U41591 (N_41591,N_38084,N_39404);
or U41592 (N_41592,N_38362,N_38463);
and U41593 (N_41593,N_39287,N_38229);
or U41594 (N_41594,N_38257,N_39430);
nand U41595 (N_41595,N_39339,N_39723);
nor U41596 (N_41596,N_38887,N_39570);
nor U41597 (N_41597,N_39581,N_38562);
or U41598 (N_41598,N_39419,N_38401);
or U41599 (N_41599,N_39100,N_39888);
nor U41600 (N_41600,N_39454,N_38527);
xor U41601 (N_41601,N_39155,N_38365);
nand U41602 (N_41602,N_38021,N_38246);
and U41603 (N_41603,N_38317,N_39802);
and U41604 (N_41604,N_38210,N_38540);
or U41605 (N_41605,N_38988,N_39963);
nor U41606 (N_41606,N_39390,N_39339);
xor U41607 (N_41607,N_38360,N_38607);
and U41608 (N_41608,N_38398,N_39376);
nor U41609 (N_41609,N_38546,N_38626);
nor U41610 (N_41610,N_39386,N_39066);
nand U41611 (N_41611,N_38746,N_38367);
nand U41612 (N_41612,N_38883,N_38751);
or U41613 (N_41613,N_38220,N_39867);
xor U41614 (N_41614,N_38721,N_39273);
nor U41615 (N_41615,N_38223,N_38501);
nand U41616 (N_41616,N_39441,N_38040);
or U41617 (N_41617,N_39492,N_38686);
xnor U41618 (N_41618,N_39732,N_38865);
and U41619 (N_41619,N_39367,N_38567);
xor U41620 (N_41620,N_38764,N_39885);
or U41621 (N_41621,N_39837,N_39174);
or U41622 (N_41622,N_38487,N_38521);
or U41623 (N_41623,N_39926,N_38792);
nand U41624 (N_41624,N_39288,N_38969);
xnor U41625 (N_41625,N_39302,N_39887);
nand U41626 (N_41626,N_38415,N_39735);
xnor U41627 (N_41627,N_39054,N_38688);
xnor U41628 (N_41628,N_39035,N_39962);
nand U41629 (N_41629,N_39030,N_39612);
or U41630 (N_41630,N_38713,N_38410);
or U41631 (N_41631,N_39418,N_38101);
or U41632 (N_41632,N_38857,N_38853);
nor U41633 (N_41633,N_38387,N_38616);
and U41634 (N_41634,N_39710,N_38554);
or U41635 (N_41635,N_38020,N_39654);
or U41636 (N_41636,N_39588,N_39061);
nor U41637 (N_41637,N_39580,N_38894);
or U41638 (N_41638,N_38312,N_39203);
and U41639 (N_41639,N_39434,N_39881);
xnor U41640 (N_41640,N_38914,N_38948);
and U41641 (N_41641,N_38095,N_39519);
and U41642 (N_41642,N_39073,N_39543);
xor U41643 (N_41643,N_39756,N_38660);
xnor U41644 (N_41644,N_39593,N_39735);
or U41645 (N_41645,N_39961,N_39115);
nor U41646 (N_41646,N_38353,N_39108);
nand U41647 (N_41647,N_38503,N_39922);
nor U41648 (N_41648,N_39063,N_38426);
or U41649 (N_41649,N_39084,N_38907);
and U41650 (N_41650,N_38350,N_39117);
nand U41651 (N_41651,N_39969,N_38703);
xnor U41652 (N_41652,N_39580,N_38202);
nor U41653 (N_41653,N_39052,N_38072);
or U41654 (N_41654,N_38334,N_39954);
nand U41655 (N_41655,N_38125,N_38476);
and U41656 (N_41656,N_39186,N_39257);
xnor U41657 (N_41657,N_39258,N_38755);
and U41658 (N_41658,N_38933,N_38617);
nand U41659 (N_41659,N_39140,N_39315);
xor U41660 (N_41660,N_38087,N_39601);
or U41661 (N_41661,N_38218,N_38331);
xnor U41662 (N_41662,N_38754,N_38438);
or U41663 (N_41663,N_38827,N_38192);
nand U41664 (N_41664,N_38731,N_39211);
nand U41665 (N_41665,N_39145,N_38751);
nor U41666 (N_41666,N_38744,N_39186);
nor U41667 (N_41667,N_39647,N_39178);
nand U41668 (N_41668,N_38393,N_38140);
and U41669 (N_41669,N_39143,N_39398);
xnor U41670 (N_41670,N_39936,N_39606);
nor U41671 (N_41671,N_39328,N_39164);
nand U41672 (N_41672,N_39359,N_38930);
nand U41673 (N_41673,N_39705,N_39382);
or U41674 (N_41674,N_38449,N_38071);
nor U41675 (N_41675,N_38989,N_38849);
nor U41676 (N_41676,N_39479,N_38543);
nor U41677 (N_41677,N_39540,N_38595);
or U41678 (N_41678,N_39032,N_38468);
nor U41679 (N_41679,N_39652,N_39098);
nand U41680 (N_41680,N_38299,N_39544);
nor U41681 (N_41681,N_39008,N_38425);
nor U41682 (N_41682,N_39535,N_39986);
nand U41683 (N_41683,N_39881,N_38839);
xor U41684 (N_41684,N_39284,N_38457);
xnor U41685 (N_41685,N_38855,N_38596);
nand U41686 (N_41686,N_39403,N_38568);
or U41687 (N_41687,N_38100,N_39256);
and U41688 (N_41688,N_39504,N_39532);
nor U41689 (N_41689,N_38515,N_38465);
or U41690 (N_41690,N_38102,N_38083);
and U41691 (N_41691,N_38240,N_38915);
nand U41692 (N_41692,N_39812,N_39686);
nand U41693 (N_41693,N_39400,N_38347);
xnor U41694 (N_41694,N_38226,N_38296);
and U41695 (N_41695,N_39621,N_38212);
or U41696 (N_41696,N_39284,N_38546);
or U41697 (N_41697,N_38060,N_38284);
or U41698 (N_41698,N_38061,N_38769);
or U41699 (N_41699,N_39682,N_38830);
and U41700 (N_41700,N_39972,N_39981);
nor U41701 (N_41701,N_38218,N_39414);
and U41702 (N_41702,N_38457,N_38097);
and U41703 (N_41703,N_38780,N_38797);
and U41704 (N_41704,N_38574,N_38619);
xnor U41705 (N_41705,N_38674,N_38521);
nand U41706 (N_41706,N_38993,N_38669);
nor U41707 (N_41707,N_38749,N_39462);
nor U41708 (N_41708,N_39342,N_39022);
xnor U41709 (N_41709,N_38685,N_39689);
nor U41710 (N_41710,N_38117,N_39418);
nand U41711 (N_41711,N_38227,N_39774);
and U41712 (N_41712,N_39611,N_39806);
or U41713 (N_41713,N_38811,N_39456);
nand U41714 (N_41714,N_38742,N_39310);
xnor U41715 (N_41715,N_38694,N_38303);
and U41716 (N_41716,N_38801,N_38503);
nand U41717 (N_41717,N_38114,N_38157);
or U41718 (N_41718,N_38025,N_39852);
nand U41719 (N_41719,N_38383,N_39189);
nand U41720 (N_41720,N_39985,N_38049);
xor U41721 (N_41721,N_39078,N_39623);
nand U41722 (N_41722,N_39117,N_39732);
or U41723 (N_41723,N_38884,N_38421);
nand U41724 (N_41724,N_39016,N_39319);
nor U41725 (N_41725,N_39715,N_39797);
nand U41726 (N_41726,N_38438,N_39146);
nand U41727 (N_41727,N_38007,N_39522);
nor U41728 (N_41728,N_39942,N_38170);
nand U41729 (N_41729,N_38183,N_38144);
nand U41730 (N_41730,N_38150,N_38123);
or U41731 (N_41731,N_38854,N_39837);
or U41732 (N_41732,N_39613,N_38572);
nor U41733 (N_41733,N_38646,N_38011);
xor U41734 (N_41734,N_39725,N_39936);
or U41735 (N_41735,N_38593,N_39558);
and U41736 (N_41736,N_38649,N_39666);
nand U41737 (N_41737,N_39393,N_39315);
xnor U41738 (N_41738,N_39176,N_38448);
or U41739 (N_41739,N_38552,N_38578);
nand U41740 (N_41740,N_39715,N_38960);
nor U41741 (N_41741,N_39502,N_39468);
or U41742 (N_41742,N_39833,N_39196);
nor U41743 (N_41743,N_39744,N_39677);
xor U41744 (N_41744,N_38184,N_39826);
or U41745 (N_41745,N_39048,N_39484);
nand U41746 (N_41746,N_38884,N_39909);
nand U41747 (N_41747,N_39760,N_39045);
nand U41748 (N_41748,N_39446,N_39115);
xnor U41749 (N_41749,N_39373,N_39501);
or U41750 (N_41750,N_39373,N_39176);
or U41751 (N_41751,N_39707,N_39850);
nor U41752 (N_41752,N_38695,N_39264);
xnor U41753 (N_41753,N_39716,N_38297);
xnor U41754 (N_41754,N_39872,N_39366);
nand U41755 (N_41755,N_39280,N_38104);
nor U41756 (N_41756,N_39624,N_38878);
xor U41757 (N_41757,N_39141,N_39952);
nor U41758 (N_41758,N_38662,N_38954);
or U41759 (N_41759,N_38654,N_39699);
or U41760 (N_41760,N_38689,N_39964);
nor U41761 (N_41761,N_39446,N_39518);
nand U41762 (N_41762,N_38138,N_38636);
nor U41763 (N_41763,N_38156,N_39291);
xor U41764 (N_41764,N_38979,N_38203);
and U41765 (N_41765,N_38050,N_39709);
xnor U41766 (N_41766,N_38812,N_38662);
or U41767 (N_41767,N_38735,N_39762);
nand U41768 (N_41768,N_39685,N_38337);
nor U41769 (N_41769,N_38553,N_38447);
xor U41770 (N_41770,N_39295,N_39665);
nand U41771 (N_41771,N_38488,N_38990);
nor U41772 (N_41772,N_39622,N_39743);
nand U41773 (N_41773,N_39001,N_38369);
xor U41774 (N_41774,N_38114,N_39955);
or U41775 (N_41775,N_39241,N_39757);
nand U41776 (N_41776,N_39601,N_38899);
and U41777 (N_41777,N_39085,N_39282);
nand U41778 (N_41778,N_38650,N_39180);
or U41779 (N_41779,N_38500,N_38400);
and U41780 (N_41780,N_39658,N_38728);
xnor U41781 (N_41781,N_39384,N_38460);
and U41782 (N_41782,N_38958,N_39747);
and U41783 (N_41783,N_39339,N_39422);
and U41784 (N_41784,N_39281,N_38622);
nand U41785 (N_41785,N_38041,N_39139);
or U41786 (N_41786,N_39299,N_38629);
nor U41787 (N_41787,N_39551,N_39015);
nor U41788 (N_41788,N_38300,N_38784);
nor U41789 (N_41789,N_38838,N_38301);
and U41790 (N_41790,N_39799,N_39035);
nor U41791 (N_41791,N_38908,N_38204);
nand U41792 (N_41792,N_39283,N_39038);
or U41793 (N_41793,N_39659,N_38183);
nand U41794 (N_41794,N_38640,N_38224);
xnor U41795 (N_41795,N_39693,N_39173);
and U41796 (N_41796,N_39803,N_39633);
and U41797 (N_41797,N_39938,N_39251);
or U41798 (N_41798,N_38143,N_38088);
nand U41799 (N_41799,N_38772,N_38483);
and U41800 (N_41800,N_39287,N_39626);
nor U41801 (N_41801,N_39793,N_38929);
and U41802 (N_41802,N_38375,N_39766);
xnor U41803 (N_41803,N_38556,N_38734);
nand U41804 (N_41804,N_39634,N_39232);
nand U41805 (N_41805,N_39865,N_39478);
nor U41806 (N_41806,N_39480,N_39619);
and U41807 (N_41807,N_39032,N_39292);
and U41808 (N_41808,N_39673,N_38425);
or U41809 (N_41809,N_38918,N_38031);
nor U41810 (N_41810,N_38969,N_38776);
or U41811 (N_41811,N_38280,N_38716);
xnor U41812 (N_41812,N_38039,N_38035);
xnor U41813 (N_41813,N_39689,N_38503);
nand U41814 (N_41814,N_39359,N_38336);
and U41815 (N_41815,N_38967,N_38728);
or U41816 (N_41816,N_38769,N_38981);
nor U41817 (N_41817,N_39038,N_38844);
nor U41818 (N_41818,N_38827,N_39227);
or U41819 (N_41819,N_39010,N_39260);
xor U41820 (N_41820,N_39820,N_38732);
xor U41821 (N_41821,N_38751,N_38813);
and U41822 (N_41822,N_38279,N_39832);
or U41823 (N_41823,N_39641,N_38549);
and U41824 (N_41824,N_39054,N_38593);
or U41825 (N_41825,N_39734,N_39366);
and U41826 (N_41826,N_39145,N_38025);
nand U41827 (N_41827,N_38118,N_38563);
nand U41828 (N_41828,N_39678,N_39628);
or U41829 (N_41829,N_38949,N_38043);
nand U41830 (N_41830,N_38949,N_38703);
nand U41831 (N_41831,N_38413,N_39626);
nor U41832 (N_41832,N_39576,N_38793);
nand U41833 (N_41833,N_38919,N_38366);
or U41834 (N_41834,N_39504,N_38063);
nand U41835 (N_41835,N_38639,N_39557);
nor U41836 (N_41836,N_38769,N_38483);
or U41837 (N_41837,N_38509,N_39800);
or U41838 (N_41838,N_38021,N_39002);
and U41839 (N_41839,N_39535,N_38971);
nand U41840 (N_41840,N_39235,N_39245);
nor U41841 (N_41841,N_39481,N_39648);
xnor U41842 (N_41842,N_38176,N_39856);
xnor U41843 (N_41843,N_39794,N_39003);
nand U41844 (N_41844,N_38918,N_39338);
and U41845 (N_41845,N_38030,N_38363);
nand U41846 (N_41846,N_39481,N_39974);
and U41847 (N_41847,N_39942,N_38698);
nor U41848 (N_41848,N_38977,N_38487);
and U41849 (N_41849,N_39385,N_39111);
and U41850 (N_41850,N_38488,N_39700);
nand U41851 (N_41851,N_39793,N_39043);
and U41852 (N_41852,N_38998,N_38624);
and U41853 (N_41853,N_39106,N_38828);
and U41854 (N_41854,N_38331,N_38537);
and U41855 (N_41855,N_38029,N_38187);
nand U41856 (N_41856,N_38770,N_38668);
nand U41857 (N_41857,N_38671,N_38557);
or U41858 (N_41858,N_39941,N_39998);
and U41859 (N_41859,N_38809,N_39509);
nor U41860 (N_41860,N_38661,N_38697);
nand U41861 (N_41861,N_39068,N_38965);
nand U41862 (N_41862,N_38664,N_38085);
xnor U41863 (N_41863,N_39401,N_38354);
or U41864 (N_41864,N_39259,N_39401);
nand U41865 (N_41865,N_39676,N_39121);
nand U41866 (N_41866,N_38062,N_39591);
nor U41867 (N_41867,N_39820,N_38990);
nor U41868 (N_41868,N_38545,N_38217);
nand U41869 (N_41869,N_39607,N_38392);
nand U41870 (N_41870,N_39852,N_39957);
nor U41871 (N_41871,N_39309,N_38390);
and U41872 (N_41872,N_38587,N_39828);
nand U41873 (N_41873,N_38457,N_39398);
nor U41874 (N_41874,N_38858,N_39886);
xor U41875 (N_41875,N_39242,N_39981);
xor U41876 (N_41876,N_38802,N_38105);
or U41877 (N_41877,N_39653,N_39054);
xnor U41878 (N_41878,N_38228,N_39036);
and U41879 (N_41879,N_39386,N_38119);
or U41880 (N_41880,N_39179,N_38731);
and U41881 (N_41881,N_39704,N_39827);
xnor U41882 (N_41882,N_38329,N_39999);
and U41883 (N_41883,N_38777,N_39624);
xor U41884 (N_41884,N_38000,N_38265);
or U41885 (N_41885,N_39855,N_38795);
or U41886 (N_41886,N_39901,N_39849);
xor U41887 (N_41887,N_38045,N_39205);
or U41888 (N_41888,N_39948,N_39945);
or U41889 (N_41889,N_38955,N_39039);
nand U41890 (N_41890,N_39781,N_39189);
nor U41891 (N_41891,N_39003,N_39082);
nand U41892 (N_41892,N_38236,N_39083);
or U41893 (N_41893,N_39000,N_39994);
nor U41894 (N_41894,N_38224,N_38366);
nand U41895 (N_41895,N_39046,N_39249);
and U41896 (N_41896,N_38243,N_38418);
nand U41897 (N_41897,N_38806,N_38310);
nor U41898 (N_41898,N_38072,N_38625);
xor U41899 (N_41899,N_38139,N_39517);
xnor U41900 (N_41900,N_39920,N_39308);
xor U41901 (N_41901,N_39347,N_38750);
and U41902 (N_41902,N_39341,N_39784);
nor U41903 (N_41903,N_39191,N_38449);
and U41904 (N_41904,N_38608,N_38287);
nand U41905 (N_41905,N_38781,N_38097);
nor U41906 (N_41906,N_39836,N_38497);
and U41907 (N_41907,N_39258,N_38597);
and U41908 (N_41908,N_38863,N_39293);
or U41909 (N_41909,N_38480,N_39457);
or U41910 (N_41910,N_38776,N_38071);
and U41911 (N_41911,N_38022,N_39531);
or U41912 (N_41912,N_38992,N_38686);
nand U41913 (N_41913,N_39516,N_39211);
xnor U41914 (N_41914,N_38608,N_38206);
nor U41915 (N_41915,N_39795,N_38005);
and U41916 (N_41916,N_39015,N_39484);
nor U41917 (N_41917,N_38755,N_39597);
and U41918 (N_41918,N_38475,N_39427);
xnor U41919 (N_41919,N_39096,N_38656);
and U41920 (N_41920,N_38466,N_39038);
and U41921 (N_41921,N_39193,N_39156);
nor U41922 (N_41922,N_39946,N_39326);
and U41923 (N_41923,N_39202,N_39292);
or U41924 (N_41924,N_39542,N_39350);
nand U41925 (N_41925,N_39455,N_38337);
nor U41926 (N_41926,N_39797,N_39575);
nor U41927 (N_41927,N_39959,N_38291);
and U41928 (N_41928,N_39068,N_38065);
nand U41929 (N_41929,N_38705,N_39059);
nand U41930 (N_41930,N_38678,N_39175);
xnor U41931 (N_41931,N_38485,N_38636);
or U41932 (N_41932,N_39420,N_38581);
or U41933 (N_41933,N_38719,N_38122);
xnor U41934 (N_41934,N_38855,N_39846);
or U41935 (N_41935,N_39876,N_38519);
nor U41936 (N_41936,N_38766,N_38874);
nor U41937 (N_41937,N_39023,N_39405);
and U41938 (N_41938,N_38717,N_38895);
or U41939 (N_41939,N_39623,N_38786);
and U41940 (N_41940,N_38010,N_39227);
and U41941 (N_41941,N_38006,N_39432);
or U41942 (N_41942,N_39233,N_39740);
nor U41943 (N_41943,N_38603,N_38795);
xor U41944 (N_41944,N_38346,N_39123);
and U41945 (N_41945,N_38601,N_38190);
nor U41946 (N_41946,N_38242,N_39816);
nand U41947 (N_41947,N_38269,N_38081);
xor U41948 (N_41948,N_38507,N_39422);
xor U41949 (N_41949,N_39178,N_38418);
and U41950 (N_41950,N_38013,N_39414);
or U41951 (N_41951,N_39642,N_39720);
or U41952 (N_41952,N_39742,N_39514);
nand U41953 (N_41953,N_39855,N_39452);
xnor U41954 (N_41954,N_38901,N_38794);
and U41955 (N_41955,N_39831,N_38490);
nor U41956 (N_41956,N_38239,N_39172);
nor U41957 (N_41957,N_39278,N_38136);
and U41958 (N_41958,N_38553,N_38875);
and U41959 (N_41959,N_38833,N_39072);
xor U41960 (N_41960,N_38055,N_38209);
and U41961 (N_41961,N_39617,N_38758);
nor U41962 (N_41962,N_38797,N_39757);
xnor U41963 (N_41963,N_39149,N_39473);
xor U41964 (N_41964,N_38425,N_38381);
or U41965 (N_41965,N_39562,N_39083);
or U41966 (N_41966,N_39292,N_38579);
nand U41967 (N_41967,N_39185,N_38270);
xor U41968 (N_41968,N_39533,N_38992);
or U41969 (N_41969,N_38909,N_39229);
and U41970 (N_41970,N_39686,N_39681);
and U41971 (N_41971,N_38729,N_38172);
nor U41972 (N_41972,N_39736,N_39505);
or U41973 (N_41973,N_38778,N_38887);
nor U41974 (N_41974,N_39455,N_38566);
xor U41975 (N_41975,N_39063,N_39257);
or U41976 (N_41976,N_39670,N_38515);
nand U41977 (N_41977,N_39875,N_38822);
nor U41978 (N_41978,N_39241,N_38230);
and U41979 (N_41979,N_39309,N_38136);
nor U41980 (N_41980,N_39242,N_39119);
and U41981 (N_41981,N_39778,N_39269);
nor U41982 (N_41982,N_38404,N_38555);
nand U41983 (N_41983,N_39443,N_39263);
or U41984 (N_41984,N_39706,N_39713);
xnor U41985 (N_41985,N_38376,N_39894);
and U41986 (N_41986,N_39283,N_38518);
and U41987 (N_41987,N_38550,N_38759);
nor U41988 (N_41988,N_39222,N_39814);
nor U41989 (N_41989,N_38894,N_39043);
nor U41990 (N_41990,N_38248,N_39177);
nor U41991 (N_41991,N_39799,N_38795);
xor U41992 (N_41992,N_38225,N_39685);
and U41993 (N_41993,N_39462,N_38767);
nand U41994 (N_41994,N_38019,N_39910);
and U41995 (N_41995,N_39407,N_39773);
nand U41996 (N_41996,N_38101,N_38331);
and U41997 (N_41997,N_39896,N_38458);
and U41998 (N_41998,N_38857,N_38256);
xnor U41999 (N_41999,N_39103,N_38623);
nor U42000 (N_42000,N_40239,N_40537);
and U42001 (N_42001,N_41202,N_40842);
nor U42002 (N_42002,N_41816,N_41193);
nor U42003 (N_42003,N_41228,N_40492);
nand U42004 (N_42004,N_40070,N_41917);
nand U42005 (N_42005,N_40730,N_40408);
nor U42006 (N_42006,N_41119,N_40467);
or U42007 (N_42007,N_41968,N_40757);
nor U42008 (N_42008,N_40963,N_41627);
and U42009 (N_42009,N_41155,N_41858);
or U42010 (N_42010,N_41961,N_41292);
nor U42011 (N_42011,N_40728,N_40485);
xnor U42012 (N_42012,N_41597,N_41371);
nand U42013 (N_42013,N_40732,N_41906);
or U42014 (N_42014,N_40826,N_41183);
nand U42015 (N_42015,N_41636,N_40369);
nand U42016 (N_42016,N_41601,N_40954);
xor U42017 (N_42017,N_41680,N_40869);
nand U42018 (N_42018,N_41755,N_41459);
xnor U42019 (N_42019,N_40406,N_41139);
xnor U42020 (N_42020,N_40082,N_40405);
nor U42021 (N_42021,N_40221,N_41199);
and U42022 (N_42022,N_40603,N_40468);
nand U42023 (N_42023,N_41167,N_40303);
nand U42024 (N_42024,N_40004,N_40225);
or U42025 (N_42025,N_40392,N_40249);
or U42026 (N_42026,N_40165,N_40804);
nor U42027 (N_42027,N_41837,N_41914);
or U42028 (N_42028,N_40762,N_40719);
nand U42029 (N_42029,N_40543,N_41232);
nor U42030 (N_42030,N_40563,N_41399);
nand U42031 (N_42031,N_40731,N_41084);
or U42032 (N_42032,N_40117,N_40981);
xnor U42033 (N_42033,N_40651,N_40993);
nand U42034 (N_42034,N_40726,N_41972);
and U42035 (N_42035,N_40496,N_41019);
nand U42036 (N_42036,N_40042,N_40850);
or U42037 (N_42037,N_40803,N_41197);
xor U42038 (N_42038,N_40794,N_40860);
nor U42039 (N_42039,N_40815,N_40489);
or U42040 (N_42040,N_41231,N_41840);
or U42041 (N_42041,N_40520,N_41358);
xnor U42042 (N_42042,N_40367,N_41066);
xnor U42043 (N_42043,N_41951,N_41591);
or U42044 (N_42044,N_40959,N_40856);
xor U42045 (N_42045,N_40930,N_41419);
and U42046 (N_42046,N_40798,N_40894);
and U42047 (N_42047,N_41373,N_40770);
nand U42048 (N_42048,N_41915,N_40482);
and U42049 (N_42049,N_40896,N_41469);
xor U42050 (N_42050,N_40355,N_40351);
and U42051 (N_42051,N_40232,N_40991);
nor U42052 (N_42052,N_40189,N_41833);
or U42053 (N_42053,N_41261,N_41963);
nor U42054 (N_42054,N_41815,N_40703);
nor U42055 (N_42055,N_40578,N_41409);
xnor U42056 (N_42056,N_41608,N_41493);
xnor U42057 (N_42057,N_41630,N_40783);
nand U42058 (N_42058,N_41294,N_40641);
and U42059 (N_42059,N_40559,N_40386);
nand U42060 (N_42060,N_41556,N_40618);
nor U42061 (N_42061,N_40668,N_41763);
xor U42062 (N_42062,N_41614,N_41310);
nand U42063 (N_42063,N_40420,N_40634);
nand U42064 (N_42064,N_41845,N_41401);
and U42065 (N_42065,N_40056,N_41296);
nand U42066 (N_42066,N_41235,N_41234);
and U42067 (N_42067,N_40148,N_40756);
xnor U42068 (N_42068,N_41902,N_41892);
nand U42069 (N_42069,N_40902,N_40847);
and U42070 (N_42070,N_41583,N_41730);
xor U42071 (N_42071,N_41617,N_40390);
and U42072 (N_42072,N_41854,N_40407);
nand U42073 (N_42073,N_40067,N_41782);
and U42074 (N_42074,N_40129,N_40216);
nor U42075 (N_42075,N_40150,N_40704);
nand U42076 (N_42076,N_41668,N_41021);
or U42077 (N_42077,N_41561,N_40648);
xor U42078 (N_42078,N_40718,N_41092);
nor U42079 (N_42079,N_40280,N_40617);
xor U42080 (N_42080,N_41780,N_41102);
or U42081 (N_42081,N_40060,N_41637);
or U42082 (N_42082,N_40620,N_41670);
nand U42083 (N_42083,N_40435,N_41513);
nand U42084 (N_42084,N_40671,N_40933);
nand U42085 (N_42085,N_41027,N_41030);
and U42086 (N_42086,N_41884,N_40733);
xor U42087 (N_42087,N_41623,N_40034);
and U42088 (N_42088,N_41101,N_40130);
and U42089 (N_42089,N_41303,N_41511);
nor U42090 (N_42090,N_40147,N_40895);
nand U42091 (N_42091,N_40062,N_41694);
and U42092 (N_42092,N_41501,N_40104);
and U42093 (N_42093,N_40497,N_40336);
xor U42094 (N_42094,N_41908,N_41153);
nor U42095 (N_42095,N_41457,N_41652);
nor U42096 (N_42096,N_41465,N_40453);
and U42097 (N_42097,N_40928,N_41046);
and U42098 (N_42098,N_41146,N_40059);
xnor U42099 (N_42099,N_41315,N_40400);
and U42100 (N_42100,N_40315,N_40901);
nand U42101 (N_42101,N_40200,N_41650);
or U42102 (N_42102,N_40025,N_41689);
xnor U42103 (N_42103,N_41322,N_41307);
nand U42104 (N_42104,N_41135,N_41477);
and U42105 (N_42105,N_40831,N_41244);
or U42106 (N_42106,N_41194,N_41372);
and U42107 (N_42107,N_40352,N_40793);
or U42108 (N_42108,N_41787,N_40058);
xnor U42109 (N_42109,N_41069,N_41293);
or U42110 (N_42110,N_41796,N_40590);
nand U42111 (N_42111,N_40428,N_41860);
nand U42112 (N_42112,N_41034,N_41390);
nor U42113 (N_42113,N_40698,N_40570);
nor U42114 (N_42114,N_41640,N_41662);
and U42115 (N_42115,N_40548,N_41000);
xnor U42116 (N_42116,N_40643,N_41578);
or U42117 (N_42117,N_41215,N_41661);
nand U42118 (N_42118,N_40961,N_40994);
xor U42119 (N_42119,N_41281,N_40207);
and U42120 (N_42120,N_41181,N_40153);
nand U42121 (N_42121,N_41891,N_41605);
xnor U42122 (N_42122,N_41642,N_41012);
and U42123 (N_42123,N_40596,N_41022);
or U42124 (N_42124,N_41909,N_41391);
and U42125 (N_42125,N_41814,N_40413);
or U42126 (N_42126,N_40396,N_40914);
and U42127 (N_42127,N_40103,N_41276);
nand U42128 (N_42128,N_41570,N_41471);
nand U42129 (N_42129,N_41881,N_41064);
nor U42130 (N_42130,N_40461,N_40627);
nand U42131 (N_42131,N_40734,N_41347);
xor U42132 (N_42132,N_40683,N_41203);
xor U42133 (N_42133,N_40136,N_40658);
nand U42134 (N_42134,N_41912,N_41430);
and U42135 (N_42135,N_40133,N_41517);
or U42136 (N_42136,N_41077,N_40608);
nand U42137 (N_42137,N_40688,N_41674);
or U42138 (N_42138,N_40795,N_40848);
xnor U42139 (N_42139,N_40662,N_40913);
nand U42140 (N_42140,N_41045,N_40823);
nand U42141 (N_42141,N_41052,N_41999);
or U42142 (N_42142,N_41790,N_41638);
xor U42143 (N_42143,N_40329,N_41005);
xnor U42144 (N_42144,N_41132,N_40217);
or U42145 (N_42145,N_41934,N_40260);
nor U42146 (N_42146,N_40927,N_41770);
and U42147 (N_42147,N_41725,N_40265);
xor U42148 (N_42148,N_40247,N_40046);
or U42149 (N_42149,N_40785,N_40455);
or U42150 (N_42150,N_40594,N_40495);
xor U42151 (N_42151,N_41384,N_41624);
xor U42152 (N_42152,N_41693,N_40715);
and U42153 (N_42153,N_41211,N_41622);
or U42154 (N_42154,N_40121,N_41079);
xnor U42155 (N_42155,N_41828,N_40502);
nand U42156 (N_42156,N_41427,N_41568);
and U42157 (N_42157,N_40910,N_40882);
or U42158 (N_42158,N_40615,N_40614);
or U42159 (N_42159,N_41849,N_41415);
xor U42160 (N_42160,N_41946,N_40131);
and U42161 (N_42161,N_40965,N_41380);
or U42162 (N_42162,N_41646,N_41086);
or U42163 (N_42163,N_40021,N_41160);
nor U42164 (N_42164,N_41374,N_41318);
xor U42165 (N_42165,N_40972,N_41644);
or U42166 (N_42166,N_40909,N_41308);
nand U42167 (N_42167,N_41118,N_40955);
or U42168 (N_42168,N_40100,N_40986);
nand U42169 (N_42169,N_40096,N_40393);
xor U42170 (N_42170,N_41502,N_40676);
nand U42171 (N_42171,N_40223,N_41089);
nand U42172 (N_42172,N_41708,N_40547);
or U42173 (N_42173,N_41474,N_40305);
xor U42174 (N_42174,N_41533,N_40654);
or U42175 (N_42175,N_41351,N_40743);
nand U42176 (N_42176,N_40213,N_41547);
or U42177 (N_42177,N_40904,N_40899);
xor U42178 (N_42178,N_41074,N_40094);
and U42179 (N_42179,N_41768,N_41248);
or U42180 (N_42180,N_40645,N_40487);
nand U42181 (N_42181,N_40636,N_40619);
nand U42182 (N_42182,N_41346,N_41579);
nor U42183 (N_42183,N_40198,N_40979);
nor U42184 (N_42184,N_40344,N_40810);
nand U42185 (N_42185,N_40112,N_40178);
nand U42186 (N_42186,N_41700,N_40414);
and U42187 (N_42187,N_40720,N_40323);
xor U42188 (N_42188,N_41889,N_41168);
nand U42189 (N_42189,N_41800,N_40817);
nor U42190 (N_42190,N_40918,N_41539);
and U42191 (N_42191,N_41606,N_41076);
nor U42192 (N_42192,N_41788,N_41421);
nor U42193 (N_42193,N_40253,N_41242);
and U42194 (N_42194,N_41841,N_40182);
xnor U42195 (N_42195,N_41407,N_41300);
and U42196 (N_42196,N_40786,N_40050);
or U42197 (N_42197,N_40833,N_41658);
nand U42198 (N_42198,N_41195,N_40318);
and U42199 (N_42199,N_41263,N_41222);
nor U42200 (N_42200,N_41776,N_40481);
or U42201 (N_42201,N_41134,N_40019);
nor U42202 (N_42202,N_40188,N_41037);
xor U42203 (N_42203,N_41072,N_41099);
nand U42204 (N_42204,N_41872,N_41857);
nor U42205 (N_42205,N_40208,N_40088);
xnor U42206 (N_42206,N_40048,N_41070);
and U42207 (N_42207,N_41486,N_41697);
and U42208 (N_42208,N_40983,N_41283);
xor U42209 (N_42209,N_41594,N_40637);
or U42210 (N_42210,N_40790,N_40859);
nand U42211 (N_42211,N_40383,N_41530);
or U42212 (N_42212,N_40639,N_41733);
nand U42213 (N_42213,N_40426,N_40095);
or U42214 (N_42214,N_41799,N_40119);
xnor U42215 (N_42215,N_41621,N_40261);
xnor U42216 (N_42216,N_41309,N_40337);
xnor U42217 (N_42217,N_40539,N_41769);
nand U42218 (N_42218,N_40602,N_40195);
or U42219 (N_42219,N_40843,N_41746);
xor U42220 (N_42220,N_41278,N_40205);
or U42221 (N_42221,N_40814,N_40358);
and U42222 (N_42222,N_41317,N_40294);
and U42223 (N_42223,N_40713,N_40974);
or U42224 (N_42224,N_41789,N_41795);
and U42225 (N_42225,N_40777,N_41552);
nand U42226 (N_42226,N_41122,N_40488);
xnor U42227 (N_42227,N_40171,N_40997);
xnor U42228 (N_42228,N_40044,N_40716);
or U42229 (N_42229,N_41903,N_40015);
or U42230 (N_42230,N_41060,N_40419);
and U42231 (N_42231,N_40958,N_41894);
nor U42232 (N_42232,N_40439,N_40572);
nand U42233 (N_42233,N_41206,N_41343);
nor U42234 (N_42234,N_40109,N_40739);
or U42235 (N_42235,N_40682,N_40236);
and U42236 (N_42236,N_40533,N_40747);
nand U42237 (N_42237,N_40063,N_41435);
nor U42238 (N_42238,N_41357,N_40191);
nand U42239 (N_42239,N_40475,N_40222);
nand U42240 (N_42240,N_40126,N_40154);
xor U42241 (N_42241,N_41613,N_41957);
and U42242 (N_42242,N_40346,N_40258);
xnor U42243 (N_42243,N_41143,N_41080);
nor U42244 (N_42244,N_41747,N_40268);
and U42245 (N_42245,N_41103,N_41006);
or U42246 (N_42246,N_41492,N_41632);
nand U42247 (N_42247,N_40008,N_41824);
and U42248 (N_42248,N_41128,N_40052);
and U42249 (N_42249,N_40569,N_40255);
nand U42250 (N_42250,N_40600,N_40145);
xnor U42251 (N_42251,N_41057,N_40418);
nand U42252 (N_42252,N_40544,N_41679);
nor U42253 (N_42253,N_41282,N_41114);
nor U42254 (N_42254,N_41531,N_40558);
xor U42255 (N_42255,N_40234,N_40861);
or U42256 (N_42256,N_40621,N_40160);
nand U42257 (N_42257,N_41068,N_40343);
nor U42258 (N_42258,N_40445,N_41440);
nor U42259 (N_42259,N_40291,N_41479);
or U42260 (N_42260,N_40878,N_41573);
or U42261 (N_42261,N_40851,N_40169);
nor U42262 (N_42262,N_41284,N_41130);
and U42263 (N_42263,N_41847,N_40252);
or U42264 (N_42264,N_41596,N_41190);
nor U42265 (N_42265,N_41345,N_40277);
or U42266 (N_42266,N_41853,N_40923);
xnor U42267 (N_42267,N_41496,N_40956);
or U42268 (N_42268,N_40526,N_41745);
xnor U42269 (N_42269,N_40484,N_41748);
xor U42270 (N_42270,N_40708,N_41911);
or U42271 (N_42271,N_41370,N_40338);
or U42272 (N_42272,N_41353,N_40146);
nand U42273 (N_42273,N_41138,N_41805);
xor U42274 (N_42274,N_40259,N_40555);
xor U42275 (N_42275,N_41255,N_40384);
nand U42276 (N_42276,N_40561,N_41223);
nand U42277 (N_42277,N_41285,N_41984);
xnor U42278 (N_42278,N_41483,N_41204);
or U42279 (N_42279,N_40211,N_40349);
nand U42280 (N_42280,N_40672,N_40283);
nand U42281 (N_42281,N_40068,N_41110);
and U42282 (N_42282,N_40812,N_41274);
and U42283 (N_42283,N_41151,N_40309);
nand U42284 (N_42284,N_40663,N_40964);
or U42285 (N_42285,N_40542,N_41529);
and U42286 (N_42286,N_41259,N_41843);
xnor U42287 (N_42287,N_40952,N_41402);
xnor U42288 (N_42288,N_40506,N_41324);
or U42289 (N_42289,N_41991,N_41250);
and U42290 (N_42290,N_41610,N_41018);
or U42291 (N_42291,N_41224,N_40254);
and U42292 (N_42292,N_41166,N_41855);
nand U42293 (N_42293,N_40201,N_40697);
or U42294 (N_42294,N_40078,N_41707);
or U42295 (N_42295,N_41731,N_40028);
or U42296 (N_42296,N_41470,N_40272);
and U42297 (N_42297,N_40741,N_41761);
or U42298 (N_42298,N_40264,N_40545);
xnor U42299 (N_42299,N_40281,N_41813);
and U42300 (N_42300,N_41218,N_41869);
xor U42301 (N_42301,N_41628,N_41995);
or U42302 (N_42302,N_40238,N_40335);
nand U42303 (N_42303,N_41559,N_40771);
and U42304 (N_42304,N_40298,N_40745);
nand U42305 (N_42305,N_40348,N_41097);
and U42306 (N_42306,N_40016,N_41988);
xor U42307 (N_42307,N_41834,N_41412);
and U42308 (N_42308,N_40900,N_40565);
nand U42309 (N_42309,N_41649,N_40871);
xor U42310 (N_42310,N_41467,N_41749);
and U42311 (N_42311,N_41260,N_41550);
nor U42312 (N_42312,N_41701,N_40120);
nand U42313 (N_42313,N_41408,N_41953);
xor U42314 (N_42314,N_40554,N_41221);
nand U42315 (N_42315,N_40454,N_41480);
nor U42316 (N_42316,N_40992,N_41767);
and U42317 (N_42317,N_41049,N_40655);
xnor U42318 (N_42318,N_40401,N_41544);
and U42319 (N_42319,N_40159,N_40480);
nand U42320 (N_42320,N_41716,N_40702);
or U42321 (N_42321,N_40051,N_40834);
or U42322 (N_42322,N_40185,N_41335);
nor U42323 (N_42323,N_41952,N_41548);
nor U42324 (N_42324,N_40076,N_41148);
nand U42325 (N_42325,N_40006,N_41955);
and U42326 (N_42326,N_40791,N_41907);
nor U42327 (N_42327,N_41212,N_40322);
and U42328 (N_42328,N_41537,N_41269);
nor U42329 (N_42329,N_40152,N_41161);
or U42330 (N_42330,N_41712,N_41239);
xor U42331 (N_42331,N_40907,N_41312);
xnor U42332 (N_42332,N_41004,N_40778);
nand U42333 (N_42333,N_40632,N_40789);
or U42334 (N_42334,N_41979,N_40376);
nor U42335 (N_42335,N_41014,N_41386);
or U42336 (N_42336,N_40389,N_41806);
xor U42337 (N_42337,N_40940,N_41081);
or U42338 (N_42338,N_41750,N_41519);
nand U42339 (N_42339,N_41185,N_41987);
xnor U42340 (N_42340,N_41172,N_40334);
nand U42341 (N_42341,N_41523,N_41265);
xor U42342 (N_42342,N_41448,N_41311);
xnor U42343 (N_42343,N_41923,N_41425);
nor U42344 (N_42344,N_40278,N_41029);
nand U42345 (N_42345,N_41209,N_41829);
nor U42346 (N_42346,N_41672,N_40233);
and U42347 (N_42347,N_41862,N_41607);
xnor U42348 (N_42348,N_40362,N_40302);
nor U42349 (N_42349,N_41938,N_40161);
nor U42350 (N_42350,N_40379,N_40382);
nor U42351 (N_42351,N_40622,N_41641);
nand U42352 (N_42352,N_40018,N_41048);
xor U42353 (N_42353,N_40518,N_40598);
xnor U42354 (N_42354,N_40538,N_41367);
nor U42355 (N_42355,N_40522,N_41592);
xnor U42356 (N_42356,N_40748,N_41098);
nor U42357 (N_42357,N_40949,N_41595);
nor U42358 (N_42358,N_41482,N_40628);
nor U42359 (N_42359,N_40670,N_40700);
and U42360 (N_42360,N_41512,N_41618);
or U42361 (N_42361,N_40585,N_41365);
nand U42362 (N_42362,N_41176,N_40677);
nand U42363 (N_42363,N_40297,N_40167);
or U42364 (N_42364,N_41330,N_40839);
and U42365 (N_42365,N_40361,N_40532);
nor U42366 (N_42366,N_40027,N_41772);
xor U42367 (N_42367,N_41002,N_40037);
or U42368 (N_42368,N_40231,N_40415);
and U42369 (N_42369,N_41313,N_41779);
nor U42370 (N_42370,N_41025,N_40101);
and U42371 (N_42371,N_40511,N_40380);
and U42372 (N_42372,N_40988,N_40135);
xor U42373 (N_42373,N_40498,N_41563);
and U42374 (N_42374,N_40727,N_41422);
xor U42375 (N_42375,N_40036,N_40581);
and U42376 (N_42376,N_40549,N_40875);
xor U42377 (N_42377,N_40512,N_40141);
nand U42378 (N_42378,N_40080,N_41704);
or U42379 (N_42379,N_40827,N_40127);
and U42380 (N_42380,N_40661,N_41339);
and U42381 (N_42381,N_40157,N_41673);
xnor U42382 (N_42382,N_40033,N_40057);
xnor U42383 (N_42383,N_41085,N_40073);
or U42384 (N_42384,N_41352,N_41585);
or U42385 (N_42385,N_40517,N_40444);
or U42386 (N_42386,N_40434,N_40087);
and U42387 (N_42387,N_40002,N_40462);
nor U42388 (N_42388,N_40235,N_41379);
or U42389 (N_42389,N_40043,N_40079);
and U42390 (N_42390,N_41572,N_41921);
xnor U42391 (N_42391,N_40776,N_40045);
nand U42392 (N_42392,N_40686,N_40364);
nand U42393 (N_42393,N_40653,N_41503);
xnor U42394 (N_42394,N_40611,N_40372);
or U42395 (N_42395,N_41893,N_41126);
xnor U42396 (N_42396,N_41580,N_41931);
or U42397 (N_42397,N_40772,N_40394);
or U42398 (N_42398,N_41207,N_40915);
nor U42399 (N_42399,N_41942,N_40177);
nand U42400 (N_42400,N_41088,N_41851);
nor U42401 (N_42401,N_41065,N_41551);
and U42402 (N_42402,N_40229,N_41803);
xor U42403 (N_42403,N_41577,N_40363);
and U42404 (N_42404,N_40665,N_41297);
or U42405 (N_42405,N_41035,N_41288);
and U42406 (N_42406,N_41735,N_41818);
and U42407 (N_42407,N_41944,N_41522);
xnor U42408 (N_42408,N_41526,N_40753);
and U42409 (N_42409,N_40942,N_41127);
and U42410 (N_42410,N_41378,N_41238);
and U42411 (N_42411,N_40164,N_41514);
nand U42412 (N_42412,N_40519,N_40138);
nand U42413 (N_42413,N_40465,N_41809);
nor U42414 (N_42414,N_40365,N_41041);
nand U42415 (N_42415,N_41376,N_40564);
and U42416 (N_42416,N_40787,N_41775);
xnor U42417 (N_42417,N_41090,N_40000);
nor U42418 (N_42418,N_41055,N_41387);
and U42419 (N_42419,N_40287,N_40054);
xor U42420 (N_42420,N_40921,N_40174);
and U42421 (N_42421,N_40314,N_40903);
xnor U42422 (N_42422,N_41885,N_41091);
or U42423 (N_42423,N_40353,N_40797);
or U42424 (N_42424,N_41233,N_40411);
nor U42425 (N_42425,N_41710,N_41040);
and U42426 (N_42426,N_41877,N_41977);
nand U42427 (N_42427,N_40646,N_41444);
nand U42428 (N_42428,N_41994,N_40685);
nand U42429 (N_42429,N_40736,N_41752);
xnor U42430 (N_42430,N_41949,N_40106);
and U42431 (N_42431,N_41028,N_40024);
and U42432 (N_42432,N_40179,N_41383);
or U42433 (N_42433,N_41129,N_40083);
and U42434 (N_42434,N_41369,N_40881);
nand U42435 (N_42435,N_40477,N_41781);
nor U42436 (N_42436,N_41534,N_40071);
or U42437 (N_42437,N_41158,N_40540);
xor U42438 (N_42438,N_41655,N_41901);
xor U42439 (N_42439,N_41913,N_41890);
and U42440 (N_42440,N_40011,N_41846);
xor U42441 (N_42441,N_40948,N_41823);
nor U42442 (N_42442,N_40982,N_40694);
and U42443 (N_42443,N_41536,N_41200);
xor U42444 (N_42444,N_40505,N_40391);
or U42445 (N_42445,N_41688,N_40709);
nor U42446 (N_42446,N_40317,N_40706);
xor U42447 (N_42447,N_41325,N_41436);
or U42448 (N_42448,N_41588,N_40387);
nor U42449 (N_42449,N_40802,N_40830);
nand U42450 (N_42450,N_40328,N_41878);
nand U42451 (N_42451,N_41115,N_41927);
nand U42452 (N_42452,N_40966,N_40950);
nor U42453 (N_42453,N_40858,N_41007);
nor U42454 (N_42454,N_41498,N_41342);
nand U42455 (N_42455,N_41416,N_41744);
nand U42456 (N_42456,N_41241,N_41565);
and U42457 (N_42457,N_41447,N_41867);
nor U42458 (N_42458,N_40752,N_40852);
nor U42459 (N_42459,N_40500,N_40717);
or U42460 (N_42460,N_40203,N_41187);
xnor U42461 (N_42461,N_41797,N_40557);
nand U42462 (N_42462,N_40113,N_41609);
xor U42463 (N_42463,N_41026,N_40529);
xnor U42464 (N_42464,N_40404,N_41031);
xnor U42465 (N_42465,N_40257,N_41320);
nor U42466 (N_42466,N_41567,N_41414);
nand U42467 (N_42467,N_40324,N_41462);
nor U42468 (N_42468,N_40746,N_41625);
and U42469 (N_42469,N_40656,N_41192);
and U42470 (N_42470,N_40735,N_41898);
and U42471 (N_42471,N_41997,N_41714);
or U42472 (N_42472,N_41692,N_40629);
xor U42473 (N_42473,N_40166,N_40199);
xnor U42474 (N_42474,N_41822,N_40173);
xor U42475 (N_42475,N_40560,N_40673);
nand U42476 (N_42476,N_40995,N_41032);
and U42477 (N_42477,N_40398,N_40635);
xor U42478 (N_42478,N_40749,N_41237);
nand U42479 (N_42479,N_41487,N_40829);
xnor U42480 (N_42480,N_41771,N_41327);
nand U42481 (N_42481,N_40168,N_41417);
nor U42482 (N_42482,N_41112,N_41978);
or U42483 (N_42483,N_40290,N_41574);
and U42484 (N_42484,N_40644,N_41439);
or U42485 (N_42485,N_41724,N_40210);
and U42486 (N_42486,N_40669,N_41581);
nand U42487 (N_42487,N_41827,N_40657);
and U42488 (N_42488,N_41291,N_41665);
xnor U42489 (N_42489,N_41943,N_40226);
nand U42490 (N_42490,N_41686,N_40381);
nor U42491 (N_42491,N_40722,N_40605);
and U42492 (N_42492,N_41058,N_41945);
xor U42493 (N_42493,N_40111,N_40055);
or U42494 (N_42494,N_40009,N_41794);
or U42495 (N_42495,N_40911,N_40808);
or U42496 (N_42496,N_40868,N_41476);
xnor U42497 (N_42497,N_40237,N_41586);
xor U42498 (N_42498,N_40796,N_40587);
xnor U42499 (N_42499,N_41366,N_40642);
and U42500 (N_42500,N_41381,N_40760);
nand U42501 (N_42501,N_41441,N_40282);
or U42502 (N_42502,N_40470,N_40666);
nor U42503 (N_42503,N_40388,N_41804);
or U42504 (N_42504,N_40340,N_41087);
or U42505 (N_42505,N_40696,N_41545);
xnor U42506 (N_42506,N_40820,N_41169);
nor U42507 (N_42507,N_41420,N_40219);
nor U42508 (N_42508,N_41321,N_40224);
and U42509 (N_42509,N_40494,N_40443);
nand U42510 (N_42510,N_40197,N_41899);
nand U42511 (N_42511,N_40593,N_41866);
nor U42512 (N_42512,N_40417,N_40325);
and U42513 (N_42513,N_41410,N_41532);
nand U42514 (N_42514,N_41718,N_41590);
nand U42515 (N_42515,N_40887,N_41125);
nand U42516 (N_42516,N_41765,N_40840);
nand U42517 (N_42517,N_40674,N_40086);
and U42518 (N_42518,N_41450,N_40528);
or U42519 (N_42519,N_41524,N_41377);
and U42520 (N_42520,N_41024,N_41880);
or U42521 (N_42521,N_41554,N_40667);
nand U42522 (N_42522,N_41445,N_41717);
nand U42523 (N_42523,N_40473,N_41976);
and U42524 (N_42524,N_41758,N_41230);
nand U42525 (N_42525,N_40562,N_41267);
or U42526 (N_42526,N_40595,N_40692);
xnor U42527 (N_42527,N_41705,N_41198);
or U42528 (N_42528,N_40262,N_40535);
nor U42529 (N_42529,N_40091,N_41729);
nand U42530 (N_42530,N_40320,N_41930);
nand U42531 (N_42531,N_40759,N_41393);
nor U42532 (N_42532,N_40501,N_40333);
and U42533 (N_42533,N_41684,N_40610);
and U42534 (N_42534,N_40660,N_40906);
nor U42535 (N_42535,N_41405,N_40275);
and U42536 (N_42536,N_41253,N_40107);
nor U42537 (N_42537,N_40531,N_41344);
and U42538 (N_42538,N_41817,N_41145);
and U42539 (N_42539,N_41919,N_41734);
or U42540 (N_42540,N_40271,N_41737);
xor U42541 (N_42541,N_41836,N_40809);
nor U42542 (N_42542,N_41905,N_41452);
and U42543 (N_42543,N_41631,N_40514);
nand U42544 (N_42544,N_40705,N_40510);
nor U42545 (N_42545,N_41826,N_41461);
xnor U42546 (N_42546,N_40601,N_41182);
nor U42547 (N_42547,N_41406,N_41271);
and U42548 (N_42548,N_40568,N_41879);
nand U42549 (N_42549,N_40920,N_40516);
and U42550 (N_42550,N_40929,N_40821);
nor U42551 (N_42551,N_40084,N_41396);
and U42552 (N_42552,N_40493,N_40678);
and U42553 (N_42553,N_40339,N_41071);
nand U42554 (N_42554,N_41990,N_41015);
nand U42555 (N_42555,N_40064,N_41142);
and U42556 (N_42556,N_41727,N_41683);
xor U42557 (N_42557,N_40170,N_40527);
and U42558 (N_42558,N_41722,N_40447);
nor U42559 (N_42559,N_40969,N_40960);
or U42560 (N_42560,N_41852,N_40984);
nand U42561 (N_42561,N_41695,N_40354);
xnor U42562 (N_42562,N_41777,N_41773);
or U42563 (N_42563,N_40108,N_41456);
xor U42564 (N_42564,N_41810,N_41404);
or U42565 (N_42565,N_40689,N_41666);
nand U42566 (N_42566,N_40250,N_40451);
or U42567 (N_42567,N_41210,N_41998);
nor U42568 (N_42568,N_41188,N_41008);
xnor U42569 (N_42569,N_41864,N_41654);
or U42570 (N_42570,N_41121,N_40591);
or U42571 (N_42571,N_41338,N_41540);
and U42572 (N_42572,N_41918,N_41152);
nand U42573 (N_42573,N_41760,N_41616);
and U42574 (N_42574,N_40864,N_41549);
or U42575 (N_42575,N_41243,N_41056);
nor U42576 (N_42576,N_40761,N_41333);
nor U42577 (N_42577,N_41350,N_40312);
and U42578 (N_42578,N_41812,N_41516);
nor U42579 (N_42579,N_41216,N_40245);
xnor U42580 (N_42580,N_40240,N_40575);
nand U42581 (N_42581,N_41392,N_41117);
and U42582 (N_42582,N_41489,N_40140);
and U42583 (N_42583,N_40970,N_41349);
nor U42584 (N_42584,N_41664,N_41510);
nand U42585 (N_42585,N_40853,N_40742);
nor U42586 (N_42586,N_41506,N_40385);
xor U42587 (N_42587,N_41560,N_40592);
xor U42588 (N_42588,N_40040,N_40597);
and U42589 (N_42589,N_40898,N_40711);
xor U42590 (N_42590,N_40123,N_41653);
nand U42591 (N_42591,N_41699,N_40293);
nand U42592 (N_42592,N_41116,N_40241);
nor U42593 (N_42593,N_41301,N_40458);
xnor U42594 (N_42594,N_41154,N_41690);
or U42595 (N_42595,N_41054,N_41562);
or U42596 (N_42596,N_40460,N_40576);
nand U42597 (N_42597,N_41720,N_40457);
and U42598 (N_42598,N_40023,N_40825);
xor U42599 (N_42599,N_41001,N_40566);
nor U42600 (N_42600,N_41394,N_40128);
xor U42601 (N_42601,N_40202,N_41948);
nand U42602 (N_42602,N_41289,N_41302);
and U42603 (N_42603,N_41442,N_40919);
nor U42604 (N_42604,N_40172,N_41842);
and U42605 (N_42605,N_41047,N_40890);
or U42606 (N_42606,N_40775,N_41227);
or U42607 (N_42607,N_41400,N_40144);
xnor U42608 (N_42608,N_40124,N_41706);
xnor U42609 (N_42609,N_41633,N_40659);
and U42610 (N_42610,N_41784,N_41106);
xnor U42611 (N_42611,N_41713,N_41982);
xnor U42612 (N_42612,N_40640,N_40935);
or U42613 (N_42613,N_40436,N_40985);
and U42614 (N_42614,N_40813,N_40922);
xnor U42615 (N_42615,N_41821,N_41895);
nor U42616 (N_42616,N_40630,N_41888);
and U42617 (N_42617,N_41558,N_40679);
and U42618 (N_42618,N_40577,N_40183);
and U42619 (N_42619,N_40701,N_40824);
nor U42620 (N_42620,N_40212,N_41290);
xor U42621 (N_42621,N_41326,N_41454);
or U42622 (N_42622,N_40699,N_41793);
nand U42623 (N_42623,N_41865,N_41108);
nor U42624 (N_42624,N_40276,N_41507);
and U42625 (N_42625,N_40712,N_41839);
nor U42626 (N_42626,N_40951,N_41508);
nor U42627 (N_42627,N_41933,N_40299);
and U42628 (N_42628,N_40370,N_40838);
or U42629 (N_42629,N_40765,N_40541);
nor U42630 (N_42630,N_40944,N_40574);
or U42631 (N_42631,N_40474,N_41715);
xor U42632 (N_42632,N_40256,N_40625);
xnor U42633 (N_42633,N_40521,N_41604);
nor U42634 (N_42634,N_41709,N_41651);
or U42635 (N_42635,N_40884,N_40421);
or U42636 (N_42636,N_41783,N_40916);
xnor U42637 (N_42637,N_40181,N_40962);
nand U42638 (N_42638,N_41095,N_41397);
or U42639 (N_42639,N_41437,N_41696);
or U42640 (N_42640,N_41602,N_41543);
nand U42641 (N_42641,N_41993,N_40041);
and U42642 (N_42642,N_40880,N_40805);
and U42643 (N_42643,N_41647,N_40924);
and U42644 (N_42644,N_40857,N_40891);
or U42645 (N_42645,N_41856,N_40779);
or U42646 (N_42646,N_41093,N_40680);
nor U42647 (N_42647,N_41932,N_41557);
xor U42648 (N_42648,N_41036,N_41165);
xnor U42649 (N_42649,N_40865,N_41225);
nand U42650 (N_42650,N_40990,N_41756);
xnor U42651 (N_42651,N_40464,N_41615);
and U42652 (N_42652,N_41546,N_40266);
nand U42653 (N_42653,N_40204,N_40729);
nor U42654 (N_42654,N_40368,N_41340);
xor U42655 (N_42655,N_40626,N_41463);
or U42656 (N_42656,N_41011,N_41922);
or U42657 (N_42657,N_40737,N_41323);
nand U42658 (N_42658,N_40513,N_41786);
and U42659 (N_42659,N_41220,N_40801);
nor U42660 (N_42660,N_41355,N_41460);
or U42661 (N_42661,N_40912,N_41759);
and U42662 (N_42662,N_41778,N_41164);
nand U42663 (N_42663,N_41171,N_40975);
nor U42664 (N_42664,N_40652,N_40438);
and U42665 (N_42665,N_40767,N_41105);
or U42666 (N_42666,N_41656,N_40483);
or U42667 (N_42667,N_41109,N_40893);
nand U42668 (N_42668,N_41639,N_40781);
or U42669 (N_42669,N_40883,N_40799);
or U42670 (N_42670,N_41598,N_40606);
nand U42671 (N_42671,N_41337,N_40691);
and U42672 (N_42672,N_41149,N_40486);
nor U42673 (N_42673,N_40751,N_40410);
or U42674 (N_42674,N_41832,N_41509);
xnor U42675 (N_42675,N_41051,N_41438);
xor U42676 (N_42676,N_40244,N_40936);
nand U42677 (N_42677,N_41053,N_41268);
and U42678 (N_42678,N_41256,N_40684);
or U42679 (N_42679,N_41835,N_41140);
xor U42680 (N_42680,N_40026,N_40289);
or U42681 (N_42681,N_40307,N_41676);
nor U42682 (N_42682,N_40459,N_41120);
nor U42683 (N_42683,N_40430,N_40295);
nor U42684 (N_42684,N_40149,N_41886);
nor U42685 (N_42685,N_40163,N_40509);
nor U42686 (N_42686,N_41348,N_41900);
nor U42687 (N_42687,N_41468,N_41726);
or U42688 (N_42688,N_40837,N_40114);
nor U42689 (N_42689,N_41719,N_40105);
nor U42690 (N_42690,N_41434,N_41453);
nand U42691 (N_42691,N_41868,N_40755);
nor U42692 (N_42692,N_40609,N_41481);
and U42693 (N_42693,N_40675,N_40681);
and U42694 (N_42694,N_40134,N_40081);
nand U42695 (N_42695,N_40553,N_41657);
and U42696 (N_42696,N_41941,N_41451);
nor U42697 (N_42697,N_41073,N_40116);
or U42698 (N_42698,N_41078,N_41251);
nand U42699 (N_42699,N_40375,N_41003);
or U42700 (N_42700,N_41947,N_40012);
nor U42701 (N_42701,N_40695,N_41663);
and U42702 (N_42702,N_41426,N_40807);
nor U42703 (N_42703,N_40999,N_41691);
nand U42704 (N_42704,N_40623,N_41920);
xnor U42705 (N_42705,N_40740,N_40077);
nor U42706 (N_42706,N_40267,N_40099);
or U42707 (N_42707,N_40350,N_41314);
and U42708 (N_42708,N_40889,N_40209);
nor U42709 (N_42709,N_41488,N_40586);
or U42710 (N_42710,N_40074,N_41926);
nand U42711 (N_42711,N_41964,N_40550);
and U42712 (N_42712,N_41721,N_41831);
nand U42713 (N_42713,N_41575,N_40347);
or U42714 (N_42714,N_40769,N_41163);
nor U42715 (N_42715,N_41175,N_41356);
or U42716 (N_42716,N_41629,N_41044);
or U42717 (N_42717,N_40186,N_41473);
and U42718 (N_42718,N_40849,N_41364);
nor U42719 (N_42719,N_40633,N_41279);
xor U42720 (N_42720,N_41542,N_41671);
and U42721 (N_42721,N_40613,N_41754);
nand U42722 (N_42722,N_40466,N_40841);
xor U42723 (N_42723,N_41939,N_41494);
or U42724 (N_42724,N_41863,N_40269);
nor U42725 (N_42725,N_40013,N_41050);
xnor U42726 (N_42726,N_41280,N_41429);
or U42727 (N_42727,N_41023,N_40589);
nand U42728 (N_42728,N_40788,N_40332);
nor U42729 (N_42729,N_41217,N_41133);
xor U42730 (N_42730,N_41500,N_40925);
or U42731 (N_42731,N_40007,N_40863);
or U42732 (N_42732,N_41587,N_40968);
or U42733 (N_42733,N_40507,N_40053);
or U42734 (N_42734,N_40321,N_40429);
or U42735 (N_42735,N_40230,N_41424);
nand U42736 (N_42736,N_41490,N_41753);
and U42737 (N_42737,N_40061,N_40132);
nand U42738 (N_42738,N_41388,N_41687);
or U42739 (N_42739,N_41458,N_41910);
nand U42740 (N_42740,N_40151,N_40845);
nor U42741 (N_42741,N_40780,N_41141);
and U42742 (N_42742,N_40987,N_40359);
nand U42743 (N_42743,N_40284,N_40403);
nand U42744 (N_42744,N_40273,N_41527);
nand U42745 (N_42745,N_40980,N_40504);
or U42746 (N_42746,N_41186,N_40412);
nor U42747 (N_42747,N_40158,N_40176);
and U42748 (N_42748,N_40828,N_40003);
or U42749 (N_42749,N_41094,N_41236);
or U42750 (N_42750,N_41681,N_40877);
or U42751 (N_42751,N_40989,N_40996);
nor U42752 (N_42752,N_41385,N_40366);
and U42753 (N_42753,N_41535,N_40313);
xnor U42754 (N_42754,N_41566,N_41331);
and U42755 (N_42755,N_41648,N_41966);
and U42756 (N_42756,N_40854,N_40017);
or U42757 (N_42757,N_41830,N_40624);
nand U42758 (N_42758,N_40750,N_41971);
xor U42759 (N_42759,N_40946,N_41272);
or U42760 (N_42760,N_40175,N_40908);
nor U42761 (N_42761,N_40649,N_41981);
nor U42762 (N_42762,N_40248,N_40867);
xor U42763 (N_42763,N_40873,N_41593);
nand U42764 (N_42764,N_41266,N_40816);
xnor U42765 (N_42765,N_40075,N_41887);
or U42766 (N_42766,N_40441,N_41792);
nor U42767 (N_42767,N_41589,N_40327);
xnor U42768 (N_42768,N_41033,N_41973);
or U42769 (N_42769,N_41111,N_40341);
and U42770 (N_42770,N_41063,N_41825);
xor U42771 (N_42771,N_41196,N_41062);
and U42772 (N_42772,N_40888,N_41455);
or U42773 (N_42773,N_40612,N_40976);
or U42774 (N_42774,N_40784,N_41685);
and U42775 (N_42775,N_40345,N_40886);
nor U42776 (N_42776,N_41428,N_41738);
or U42777 (N_42777,N_41929,N_41728);
nand U42778 (N_42778,N_40744,N_41801);
or U42779 (N_42779,N_40723,N_41924);
nor U42780 (N_42780,N_41928,N_41478);
xnor U42781 (N_42781,N_40218,N_40693);
nor U42782 (N_42782,N_41262,N_41361);
nor U42783 (N_42783,N_41774,N_40286);
and U42784 (N_42784,N_40471,N_41403);
xnor U42785 (N_42785,N_40472,N_41965);
nor U42786 (N_42786,N_40499,N_41131);
nor U42787 (N_42787,N_41850,N_40356);
xnor U42788 (N_42788,N_41328,N_41739);
nor U42789 (N_42789,N_41896,N_41732);
nor U42790 (N_42790,N_40524,N_41107);
xnor U42791 (N_42791,N_40448,N_41277);
xor U42792 (N_42792,N_40102,N_40288);
nor U42793 (N_42793,N_41059,N_40162);
nand U42794 (N_42794,N_40098,N_40431);
nand U42795 (N_42795,N_41144,N_40072);
and U42796 (N_42796,N_41247,N_40125);
nand U42797 (N_42797,N_40917,N_40931);
and U42798 (N_42798,N_40819,N_40001);
xnor U42799 (N_42799,N_41555,N_41245);
or U42800 (N_42800,N_41213,N_41083);
or U42801 (N_42801,N_41541,N_41316);
nand U42802 (N_42802,N_40432,N_40090);
nand U42803 (N_42803,N_40331,N_40523);
nand U42804 (N_42804,N_40876,N_40582);
xor U42805 (N_42805,N_41411,N_40242);
nand U42806 (N_42806,N_40616,N_40093);
and U42807 (N_42807,N_40947,N_41295);
xor U42808 (N_42808,N_41711,N_41208);
or U42809 (N_42809,N_40556,N_41897);
nand U42810 (N_42810,N_40433,N_41677);
nand U42811 (N_42811,N_41702,N_40939);
and U42812 (N_42812,N_40270,N_41354);
xor U42813 (N_42813,N_40758,N_41205);
and U42814 (N_42814,N_40664,N_40069);
nor U42815 (N_42815,N_41682,N_40953);
or U42816 (N_42816,N_40773,N_41940);
nand U42817 (N_42817,N_40416,N_41201);
nor U42818 (N_42818,N_41418,N_41871);
and U42819 (N_42819,N_40806,N_41246);
nand U42820 (N_42820,N_40479,N_41975);
nor U42821 (N_42821,N_41061,N_41582);
xnor U42822 (N_42822,N_41431,N_41703);
and U42823 (N_42823,N_40038,N_40967);
or U42824 (N_42824,N_40243,N_40115);
nor U42825 (N_42825,N_41937,N_40978);
nand U42826 (N_42826,N_41762,N_41904);
xor U42827 (N_42827,N_41848,N_41360);
and U42828 (N_42828,N_40422,N_40377);
and U42829 (N_42829,N_40724,N_40525);
xnor U42830 (N_42830,N_40316,N_41009);
nand U42831 (N_42831,N_41433,N_41743);
nand U42832 (N_42832,N_40721,N_41667);
nand U42833 (N_42833,N_40194,N_41273);
nand U42834 (N_42834,N_40862,N_41954);
or U42835 (N_42835,N_41757,N_40879);
xor U42836 (N_42836,N_41620,N_40552);
and U42837 (N_42837,N_41958,N_40192);
xnor U42838 (N_42838,N_41569,N_41270);
nand U42839 (N_42839,N_40926,N_41472);
or U42840 (N_42840,N_41043,N_40206);
nand U42841 (N_42841,N_41495,N_40110);
xor U42842 (N_42842,N_40279,N_41226);
or U42843 (N_42843,N_40934,N_41382);
and U42844 (N_42844,N_41980,N_40811);
and U42845 (N_42845,N_41785,N_41252);
and U42846 (N_42846,N_41039,N_41861);
and U42847 (N_42847,N_40546,N_41191);
nor U42848 (N_42848,N_41599,N_41016);
nor U42849 (N_42849,N_40423,N_40022);
nand U42850 (N_42850,N_40047,N_41791);
nand U42851 (N_42851,N_41660,N_40832);
and U42852 (N_42852,N_40897,N_40285);
xor U42853 (N_42853,N_40571,N_41807);
or U42854 (N_42854,N_40768,N_40326);
and U42855 (N_42855,N_41515,N_41017);
or U42856 (N_42856,N_41764,N_40725);
nor U42857 (N_42857,N_41104,N_40446);
and U42858 (N_42858,N_41485,N_41184);
or U42859 (N_42859,N_40836,N_41304);
or U42860 (N_42860,N_41038,N_41874);
nand U42861 (N_42861,N_41611,N_41214);
nand U42862 (N_42862,N_41375,N_41013);
nor U42863 (N_42863,N_40469,N_40190);
and U42864 (N_42864,N_41258,N_40650);
nand U42865 (N_42865,N_41299,N_40020);
or U42866 (N_42866,N_41876,N_40306);
xnor U42867 (N_42867,N_40998,N_41571);
xnor U42868 (N_42868,N_40330,N_41249);
xor U42869 (N_42869,N_41179,N_41859);
or U42870 (N_42870,N_41020,N_41766);
or U42871 (N_42871,N_41612,N_40714);
nand U42872 (N_42872,N_40957,N_40800);
or U42873 (N_42873,N_41150,N_41819);
nor U42874 (N_42874,N_41413,N_41986);
or U42875 (N_42875,N_40973,N_41974);
nand U42876 (N_42876,N_41286,N_40822);
or U42877 (N_42877,N_40515,N_40450);
xor U42878 (N_42878,N_40754,N_41723);
nor U42879 (N_42879,N_41042,N_40607);
nor U42880 (N_42880,N_41600,N_40905);
and U42881 (N_42881,N_40228,N_41564);
and U42882 (N_42882,N_41096,N_40409);
nor U42883 (N_42883,N_40456,N_41925);
or U42884 (N_42884,N_40227,N_41798);
and U42885 (N_42885,N_41177,N_40085);
and U42886 (N_42886,N_40274,N_40764);
xnor U42887 (N_42887,N_40156,N_41883);
or U42888 (N_42888,N_40792,N_41808);
and U42889 (N_42889,N_40573,N_40308);
nor U42890 (N_42890,N_40010,N_41100);
or U42891 (N_42891,N_41983,N_41742);
xor U42892 (N_42892,N_41219,N_41170);
xor U42893 (N_42893,N_41254,N_40246);
nor U42894 (N_42894,N_40452,N_41520);
nor U42895 (N_42895,N_41137,N_40463);
xor U42896 (N_42896,N_40030,N_41870);
nor U42897 (N_42897,N_40360,N_41464);
and U42898 (N_42898,N_41698,N_41950);
or U42899 (N_42899,N_40122,N_41619);
nand U42900 (N_42900,N_41174,N_40604);
or U42901 (N_42901,N_40184,N_40301);
or U42902 (N_42902,N_41882,N_41178);
xor U42903 (N_42903,N_40143,N_40971);
nand U42904 (N_42904,N_41264,N_41363);
and U42905 (N_42905,N_40476,N_40296);
nand U42906 (N_42906,N_41669,N_40937);
or U42907 (N_42907,N_41635,N_41319);
xnor U42908 (N_42908,N_40738,N_41173);
nand U42909 (N_42909,N_40932,N_40357);
and U42910 (N_42910,N_40599,N_41626);
nand U42911 (N_42911,N_41082,N_40065);
nor U42912 (N_42912,N_40092,N_41521);
nand U42913 (N_42913,N_41985,N_41802);
nor U42914 (N_42914,N_41553,N_40139);
xor U42915 (N_42915,N_41741,N_41935);
and U42916 (N_42916,N_40311,N_40142);
xor U42917 (N_42917,N_40491,N_41010);
and U42918 (N_42918,N_40647,N_40399);
nand U42919 (N_42919,N_41157,N_41067);
xnor U42920 (N_42920,N_41491,N_40977);
and U42921 (N_42921,N_40892,N_40872);
xnor U42922 (N_42922,N_40220,N_40005);
xnor U42923 (N_42923,N_40371,N_41475);
xor U42924 (N_42924,N_41359,N_40029);
nand U42925 (N_42925,N_40378,N_41659);
nor U42926 (N_42926,N_40196,N_41518);
and U42927 (N_42927,N_41341,N_41525);
or U42928 (N_42928,N_41956,N_40251);
and U42929 (N_42929,N_41189,N_41287);
xnor U42930 (N_42930,N_41395,N_41740);
or U42931 (N_42931,N_41423,N_40846);
or U42932 (N_42932,N_40534,N_41838);
xor U42933 (N_42933,N_41751,N_40032);
nand U42934 (N_42934,N_40031,N_41446);
xnor U42935 (N_42935,N_41499,N_40943);
nor U42936 (N_42936,N_41811,N_40580);
xnor U42937 (N_42937,N_41329,N_40766);
xnor U42938 (N_42938,N_41992,N_40567);
or U42939 (N_42939,N_40193,N_40442);
nor U42940 (N_42940,N_41113,N_41432);
xor U42941 (N_42941,N_40342,N_40874);
xnor U42942 (N_42942,N_41240,N_40774);
nand U42943 (N_42943,N_40039,N_40304);
nand U42944 (N_42944,N_40402,N_40397);
or U42945 (N_42945,N_41960,N_41820);
or U42946 (N_42946,N_40374,N_41497);
xnor U42947 (N_42947,N_41229,N_41916);
and U42948 (N_42948,N_41967,N_41959);
nand U42949 (N_42949,N_41368,N_40710);
nor U42950 (N_42950,N_40536,N_41576);
or U42951 (N_42951,N_40215,N_40588);
and U42952 (N_42952,N_40631,N_40449);
xor U42953 (N_42953,N_40292,N_40763);
xnor U42954 (N_42954,N_41678,N_40263);
and U42955 (N_42955,N_40551,N_41398);
nor U42956 (N_42956,N_40490,N_40584);
nor U42957 (N_42957,N_41298,N_41736);
nor U42958 (N_42958,N_40300,N_40214);
and U42959 (N_42959,N_41643,N_40319);
xnor U42960 (N_42960,N_41538,N_40310);
nor U42961 (N_42961,N_41466,N_40707);
and U42962 (N_42962,N_40844,N_41334);
xnor U42963 (N_42963,N_41389,N_41962);
or U42964 (N_42964,N_41634,N_41306);
or U42965 (N_42965,N_41504,N_40373);
xor U42966 (N_42966,N_41075,N_41124);
nand U42967 (N_42967,N_40687,N_41159);
nand U42968 (N_42968,N_40440,N_40137);
xnor U42969 (N_42969,N_40155,N_40478);
and U42970 (N_42970,N_41257,N_40424);
and U42971 (N_42971,N_40118,N_41332);
xor U42972 (N_42972,N_40885,N_41180);
and U42973 (N_42973,N_40066,N_41844);
and U42974 (N_42974,N_40690,N_40945);
or U42975 (N_42975,N_40180,N_40395);
and U42976 (N_42976,N_41123,N_40049);
or U42977 (N_42977,N_41603,N_40855);
xnor U42978 (N_42978,N_41362,N_40035);
xor U42979 (N_42979,N_41528,N_40782);
or U42980 (N_42980,N_40425,N_40014);
nor U42981 (N_42981,N_41275,N_41970);
nand U42982 (N_42982,N_40503,N_41449);
nor U42983 (N_42983,N_40427,N_40941);
xor U42984 (N_42984,N_41996,N_41336);
nand U42985 (N_42985,N_40579,N_41484);
or U42986 (N_42986,N_40870,N_41136);
xor U42987 (N_42987,N_40097,N_41675);
or U42988 (N_42988,N_41162,N_41443);
or U42989 (N_42989,N_40638,N_41645);
or U42990 (N_42990,N_40866,N_41936);
nand U42991 (N_42991,N_41875,N_40818);
nor U42992 (N_42992,N_40437,N_40187);
xor U42993 (N_42993,N_40835,N_40530);
nor U42994 (N_42994,N_41989,N_41584);
xnor U42995 (N_42995,N_41156,N_40583);
and U42996 (N_42996,N_41147,N_40089);
nor U42997 (N_42997,N_41873,N_40508);
nand U42998 (N_42998,N_40938,N_41969);
nor U42999 (N_42999,N_41505,N_41305);
or U43000 (N_43000,N_40634,N_40877);
or U43001 (N_43001,N_41322,N_41721);
xor U43002 (N_43002,N_41619,N_41923);
nand U43003 (N_43003,N_40879,N_41906);
xor U43004 (N_43004,N_40023,N_40916);
xor U43005 (N_43005,N_41983,N_40721);
or U43006 (N_43006,N_40826,N_40334);
and U43007 (N_43007,N_40449,N_40958);
and U43008 (N_43008,N_41990,N_40683);
xnor U43009 (N_43009,N_40020,N_41074);
xor U43010 (N_43010,N_41383,N_41995);
or U43011 (N_43011,N_41952,N_41138);
or U43012 (N_43012,N_40653,N_40039);
or U43013 (N_43013,N_41805,N_41986);
xnor U43014 (N_43014,N_41839,N_40402);
xnor U43015 (N_43015,N_40221,N_40587);
nand U43016 (N_43016,N_41414,N_41866);
and U43017 (N_43017,N_41397,N_41958);
xor U43018 (N_43018,N_41874,N_40667);
nand U43019 (N_43019,N_40629,N_40980);
nand U43020 (N_43020,N_40787,N_40658);
nor U43021 (N_43021,N_40762,N_40150);
and U43022 (N_43022,N_41268,N_41673);
nand U43023 (N_43023,N_41378,N_40000);
nor U43024 (N_43024,N_41553,N_41367);
nor U43025 (N_43025,N_41229,N_41627);
xor U43026 (N_43026,N_40840,N_41741);
and U43027 (N_43027,N_41241,N_41586);
and U43028 (N_43028,N_40367,N_40474);
and U43029 (N_43029,N_41174,N_40358);
or U43030 (N_43030,N_41636,N_40622);
xnor U43031 (N_43031,N_40142,N_40937);
and U43032 (N_43032,N_41867,N_40475);
and U43033 (N_43033,N_41314,N_40474);
xor U43034 (N_43034,N_40539,N_41130);
and U43035 (N_43035,N_41024,N_41409);
xnor U43036 (N_43036,N_40713,N_41867);
and U43037 (N_43037,N_40529,N_40716);
and U43038 (N_43038,N_40428,N_40002);
nand U43039 (N_43039,N_41549,N_40696);
and U43040 (N_43040,N_41382,N_41080);
nand U43041 (N_43041,N_41882,N_40367);
nand U43042 (N_43042,N_40330,N_40164);
nor U43043 (N_43043,N_41209,N_41138);
or U43044 (N_43044,N_41377,N_41072);
or U43045 (N_43045,N_40640,N_41482);
xnor U43046 (N_43046,N_41785,N_41839);
nand U43047 (N_43047,N_40867,N_41418);
or U43048 (N_43048,N_40530,N_40754);
nand U43049 (N_43049,N_40996,N_40776);
and U43050 (N_43050,N_41377,N_40884);
and U43051 (N_43051,N_40595,N_40362);
xnor U43052 (N_43052,N_40135,N_40442);
nor U43053 (N_43053,N_41023,N_40544);
and U43054 (N_43054,N_40335,N_40480);
nor U43055 (N_43055,N_41069,N_40619);
or U43056 (N_43056,N_40646,N_40109);
or U43057 (N_43057,N_40034,N_40004);
or U43058 (N_43058,N_40360,N_41166);
or U43059 (N_43059,N_41447,N_41666);
nor U43060 (N_43060,N_41522,N_41981);
or U43061 (N_43061,N_40617,N_40152);
or U43062 (N_43062,N_40606,N_41579);
or U43063 (N_43063,N_40069,N_40445);
xor U43064 (N_43064,N_40873,N_40503);
and U43065 (N_43065,N_41205,N_40865);
or U43066 (N_43066,N_41513,N_41926);
and U43067 (N_43067,N_40303,N_41020);
nor U43068 (N_43068,N_41598,N_41364);
nor U43069 (N_43069,N_40034,N_41580);
xor U43070 (N_43070,N_41146,N_41235);
nand U43071 (N_43071,N_41293,N_40857);
xnor U43072 (N_43072,N_41992,N_41742);
and U43073 (N_43073,N_41130,N_40109);
and U43074 (N_43074,N_41055,N_41974);
or U43075 (N_43075,N_40735,N_40543);
nand U43076 (N_43076,N_41017,N_40366);
xnor U43077 (N_43077,N_41191,N_41531);
xor U43078 (N_43078,N_40646,N_41472);
nor U43079 (N_43079,N_41400,N_41132);
nor U43080 (N_43080,N_40913,N_41179);
or U43081 (N_43081,N_41605,N_41640);
nor U43082 (N_43082,N_41817,N_40965);
or U43083 (N_43083,N_41968,N_41847);
or U43084 (N_43084,N_40500,N_41732);
xor U43085 (N_43085,N_40909,N_40663);
nor U43086 (N_43086,N_40491,N_40514);
nor U43087 (N_43087,N_41762,N_41058);
nor U43088 (N_43088,N_41134,N_40830);
xor U43089 (N_43089,N_40593,N_41231);
xnor U43090 (N_43090,N_41313,N_41660);
and U43091 (N_43091,N_40125,N_41529);
nand U43092 (N_43092,N_40317,N_41357);
nand U43093 (N_43093,N_40630,N_41647);
or U43094 (N_43094,N_41639,N_41809);
and U43095 (N_43095,N_41465,N_40258);
and U43096 (N_43096,N_40851,N_41368);
or U43097 (N_43097,N_41113,N_41191);
xnor U43098 (N_43098,N_41885,N_41781);
or U43099 (N_43099,N_41338,N_40840);
nor U43100 (N_43100,N_40022,N_41400);
nor U43101 (N_43101,N_41899,N_40746);
xnor U43102 (N_43102,N_41018,N_41453);
or U43103 (N_43103,N_40842,N_40945);
or U43104 (N_43104,N_41669,N_40827);
nand U43105 (N_43105,N_41926,N_40667);
or U43106 (N_43106,N_40702,N_40712);
or U43107 (N_43107,N_40961,N_40134);
nand U43108 (N_43108,N_41899,N_41353);
and U43109 (N_43109,N_41111,N_40535);
nand U43110 (N_43110,N_41478,N_40539);
xnor U43111 (N_43111,N_41802,N_40398);
nor U43112 (N_43112,N_41623,N_40893);
xor U43113 (N_43113,N_41733,N_41825);
xor U43114 (N_43114,N_41245,N_40837);
xor U43115 (N_43115,N_41923,N_40765);
xnor U43116 (N_43116,N_40237,N_40507);
xor U43117 (N_43117,N_41159,N_40107);
nand U43118 (N_43118,N_41043,N_40986);
nand U43119 (N_43119,N_41897,N_40150);
or U43120 (N_43120,N_40239,N_40977);
xor U43121 (N_43121,N_41301,N_41762);
nand U43122 (N_43122,N_40175,N_40419);
nor U43123 (N_43123,N_40030,N_40766);
xnor U43124 (N_43124,N_41139,N_40219);
nor U43125 (N_43125,N_40139,N_40961);
nand U43126 (N_43126,N_41802,N_41674);
and U43127 (N_43127,N_40426,N_41135);
nand U43128 (N_43128,N_41019,N_41931);
nand U43129 (N_43129,N_40978,N_41018);
or U43130 (N_43130,N_41635,N_40458);
nor U43131 (N_43131,N_40234,N_41343);
nor U43132 (N_43132,N_40742,N_40774);
nor U43133 (N_43133,N_41291,N_41950);
nand U43134 (N_43134,N_41661,N_40306);
nor U43135 (N_43135,N_41611,N_41341);
nand U43136 (N_43136,N_41004,N_40687);
nand U43137 (N_43137,N_41506,N_41112);
nand U43138 (N_43138,N_40925,N_40516);
nor U43139 (N_43139,N_40657,N_41243);
xor U43140 (N_43140,N_40905,N_41804);
and U43141 (N_43141,N_41408,N_40864);
nor U43142 (N_43142,N_40083,N_41052);
xnor U43143 (N_43143,N_41065,N_40187);
nor U43144 (N_43144,N_40334,N_40261);
nor U43145 (N_43145,N_41229,N_40071);
or U43146 (N_43146,N_41820,N_40177);
nor U43147 (N_43147,N_40946,N_40629);
nor U43148 (N_43148,N_40119,N_40706);
nand U43149 (N_43149,N_41069,N_41173);
and U43150 (N_43150,N_41598,N_41662);
xnor U43151 (N_43151,N_41412,N_41219);
nand U43152 (N_43152,N_40559,N_41014);
nand U43153 (N_43153,N_40069,N_41511);
xnor U43154 (N_43154,N_40038,N_41335);
xnor U43155 (N_43155,N_41493,N_41278);
nand U43156 (N_43156,N_41144,N_41551);
or U43157 (N_43157,N_41452,N_40654);
xnor U43158 (N_43158,N_41614,N_40874);
nor U43159 (N_43159,N_40815,N_40293);
nor U43160 (N_43160,N_40570,N_41275);
xor U43161 (N_43161,N_40711,N_40817);
nor U43162 (N_43162,N_41989,N_41036);
or U43163 (N_43163,N_40609,N_41522);
or U43164 (N_43164,N_40221,N_41285);
nor U43165 (N_43165,N_41904,N_40903);
xor U43166 (N_43166,N_41159,N_40772);
nand U43167 (N_43167,N_41346,N_41072);
nand U43168 (N_43168,N_41653,N_40208);
or U43169 (N_43169,N_40267,N_40123);
or U43170 (N_43170,N_41522,N_41537);
and U43171 (N_43171,N_41005,N_40793);
or U43172 (N_43172,N_40709,N_41178);
xor U43173 (N_43173,N_41779,N_40529);
and U43174 (N_43174,N_40994,N_40910);
nor U43175 (N_43175,N_41592,N_41833);
xor U43176 (N_43176,N_40900,N_41179);
nand U43177 (N_43177,N_41050,N_40481);
nand U43178 (N_43178,N_41618,N_41655);
and U43179 (N_43179,N_41199,N_40773);
nand U43180 (N_43180,N_41807,N_40750);
or U43181 (N_43181,N_41609,N_41455);
nand U43182 (N_43182,N_41184,N_41905);
and U43183 (N_43183,N_40178,N_41220);
or U43184 (N_43184,N_41318,N_41037);
or U43185 (N_43185,N_41613,N_41263);
xnor U43186 (N_43186,N_40473,N_40265);
or U43187 (N_43187,N_41771,N_40060);
xnor U43188 (N_43188,N_41742,N_40484);
or U43189 (N_43189,N_41573,N_41653);
nor U43190 (N_43190,N_41732,N_40668);
xnor U43191 (N_43191,N_40330,N_41911);
or U43192 (N_43192,N_41366,N_41076);
nand U43193 (N_43193,N_40560,N_41155);
xor U43194 (N_43194,N_40656,N_40787);
or U43195 (N_43195,N_41258,N_40153);
and U43196 (N_43196,N_41553,N_40674);
and U43197 (N_43197,N_40985,N_40963);
xor U43198 (N_43198,N_40462,N_40814);
and U43199 (N_43199,N_41351,N_41628);
and U43200 (N_43200,N_40715,N_41022);
and U43201 (N_43201,N_40342,N_41165);
nand U43202 (N_43202,N_40464,N_40784);
nand U43203 (N_43203,N_40339,N_40856);
or U43204 (N_43204,N_40606,N_41622);
or U43205 (N_43205,N_41391,N_40185);
nand U43206 (N_43206,N_41179,N_41519);
and U43207 (N_43207,N_41884,N_41270);
nand U43208 (N_43208,N_40554,N_40785);
nor U43209 (N_43209,N_40921,N_40560);
and U43210 (N_43210,N_41031,N_41403);
nand U43211 (N_43211,N_41335,N_40975);
nor U43212 (N_43212,N_41122,N_40232);
and U43213 (N_43213,N_41394,N_41162);
or U43214 (N_43214,N_41869,N_41412);
or U43215 (N_43215,N_41885,N_41759);
or U43216 (N_43216,N_40173,N_40049);
or U43217 (N_43217,N_41338,N_41554);
xor U43218 (N_43218,N_40216,N_40418);
or U43219 (N_43219,N_41062,N_40079);
nor U43220 (N_43220,N_41023,N_41539);
nor U43221 (N_43221,N_41319,N_40566);
or U43222 (N_43222,N_40343,N_40328);
xnor U43223 (N_43223,N_40456,N_41179);
xor U43224 (N_43224,N_40986,N_41415);
or U43225 (N_43225,N_40822,N_41484);
and U43226 (N_43226,N_41841,N_40250);
nor U43227 (N_43227,N_41002,N_41135);
and U43228 (N_43228,N_41324,N_41736);
nor U43229 (N_43229,N_41714,N_40341);
or U43230 (N_43230,N_40886,N_40781);
or U43231 (N_43231,N_40794,N_41810);
and U43232 (N_43232,N_41213,N_40226);
xor U43233 (N_43233,N_40493,N_41441);
or U43234 (N_43234,N_41725,N_41198);
or U43235 (N_43235,N_41808,N_40015);
or U43236 (N_43236,N_41209,N_40941);
nand U43237 (N_43237,N_40004,N_41308);
or U43238 (N_43238,N_41605,N_41956);
and U43239 (N_43239,N_40844,N_41552);
or U43240 (N_43240,N_40700,N_41535);
and U43241 (N_43241,N_41535,N_40556);
and U43242 (N_43242,N_41392,N_40789);
nand U43243 (N_43243,N_40972,N_41936);
nand U43244 (N_43244,N_40515,N_41687);
xnor U43245 (N_43245,N_40416,N_40400);
xor U43246 (N_43246,N_40570,N_40722);
xor U43247 (N_43247,N_40281,N_41926);
nor U43248 (N_43248,N_40132,N_41218);
and U43249 (N_43249,N_41625,N_41032);
nor U43250 (N_43250,N_41166,N_40127);
or U43251 (N_43251,N_40890,N_40449);
xor U43252 (N_43252,N_41572,N_40960);
xor U43253 (N_43253,N_41601,N_41051);
nor U43254 (N_43254,N_41675,N_40871);
nor U43255 (N_43255,N_40676,N_41905);
or U43256 (N_43256,N_41537,N_41371);
xor U43257 (N_43257,N_40404,N_40678);
nand U43258 (N_43258,N_40026,N_40588);
and U43259 (N_43259,N_40107,N_40020);
nor U43260 (N_43260,N_40525,N_40720);
xor U43261 (N_43261,N_40602,N_40923);
and U43262 (N_43262,N_40583,N_40079);
xor U43263 (N_43263,N_40230,N_41067);
xor U43264 (N_43264,N_40042,N_41655);
nor U43265 (N_43265,N_40919,N_41729);
nor U43266 (N_43266,N_41006,N_41685);
and U43267 (N_43267,N_41085,N_40849);
nand U43268 (N_43268,N_40507,N_41829);
nand U43269 (N_43269,N_40127,N_41075);
or U43270 (N_43270,N_40497,N_40592);
and U43271 (N_43271,N_41798,N_41055);
xnor U43272 (N_43272,N_40549,N_40692);
xor U43273 (N_43273,N_40226,N_40611);
or U43274 (N_43274,N_41090,N_40165);
and U43275 (N_43275,N_41996,N_41494);
or U43276 (N_43276,N_40882,N_40101);
and U43277 (N_43277,N_40055,N_41996);
nor U43278 (N_43278,N_40047,N_41554);
nor U43279 (N_43279,N_41475,N_41667);
nand U43280 (N_43280,N_40830,N_41986);
and U43281 (N_43281,N_40258,N_41516);
or U43282 (N_43282,N_41191,N_40845);
nand U43283 (N_43283,N_41829,N_40370);
or U43284 (N_43284,N_41477,N_41252);
and U43285 (N_43285,N_41097,N_40113);
or U43286 (N_43286,N_41927,N_40929);
and U43287 (N_43287,N_40925,N_41195);
nand U43288 (N_43288,N_41324,N_41509);
or U43289 (N_43289,N_40688,N_40810);
xor U43290 (N_43290,N_40242,N_40649);
and U43291 (N_43291,N_40308,N_41995);
nand U43292 (N_43292,N_40857,N_41092);
and U43293 (N_43293,N_40358,N_40720);
nor U43294 (N_43294,N_40522,N_41176);
and U43295 (N_43295,N_41171,N_41440);
and U43296 (N_43296,N_40779,N_41574);
and U43297 (N_43297,N_41597,N_41041);
nand U43298 (N_43298,N_41819,N_40060);
nand U43299 (N_43299,N_40002,N_40700);
xnor U43300 (N_43300,N_41475,N_40746);
xor U43301 (N_43301,N_40200,N_40474);
and U43302 (N_43302,N_40006,N_40881);
xor U43303 (N_43303,N_41421,N_41767);
and U43304 (N_43304,N_40833,N_40282);
xor U43305 (N_43305,N_40054,N_40478);
nor U43306 (N_43306,N_40126,N_40709);
nor U43307 (N_43307,N_41671,N_40172);
xor U43308 (N_43308,N_40247,N_41310);
and U43309 (N_43309,N_40942,N_41731);
nor U43310 (N_43310,N_41252,N_40844);
xor U43311 (N_43311,N_40468,N_41401);
xnor U43312 (N_43312,N_41968,N_41585);
nor U43313 (N_43313,N_41174,N_40730);
xnor U43314 (N_43314,N_40336,N_40253);
nor U43315 (N_43315,N_41471,N_40978);
nand U43316 (N_43316,N_41253,N_40383);
and U43317 (N_43317,N_41816,N_41732);
xnor U43318 (N_43318,N_41556,N_40147);
nor U43319 (N_43319,N_41684,N_40393);
nand U43320 (N_43320,N_41199,N_41614);
or U43321 (N_43321,N_41127,N_40615);
xnor U43322 (N_43322,N_40736,N_40925);
or U43323 (N_43323,N_41695,N_41567);
or U43324 (N_43324,N_40097,N_40320);
and U43325 (N_43325,N_40755,N_40503);
and U43326 (N_43326,N_40054,N_40189);
nand U43327 (N_43327,N_40828,N_41298);
and U43328 (N_43328,N_41332,N_41042);
or U43329 (N_43329,N_41893,N_41217);
nand U43330 (N_43330,N_41261,N_41748);
xor U43331 (N_43331,N_40517,N_40503);
and U43332 (N_43332,N_41253,N_40378);
and U43333 (N_43333,N_40994,N_40198);
and U43334 (N_43334,N_41042,N_41830);
and U43335 (N_43335,N_40138,N_41701);
or U43336 (N_43336,N_40400,N_41046);
or U43337 (N_43337,N_40426,N_40839);
and U43338 (N_43338,N_41745,N_40035);
nor U43339 (N_43339,N_40279,N_40941);
or U43340 (N_43340,N_40528,N_41408);
or U43341 (N_43341,N_40897,N_41843);
nand U43342 (N_43342,N_41785,N_40066);
xor U43343 (N_43343,N_41621,N_41389);
nor U43344 (N_43344,N_40895,N_40112);
xor U43345 (N_43345,N_41621,N_41705);
and U43346 (N_43346,N_41113,N_40110);
nand U43347 (N_43347,N_40223,N_41291);
nor U43348 (N_43348,N_41516,N_40268);
nor U43349 (N_43349,N_40081,N_40096);
xor U43350 (N_43350,N_41339,N_40840);
or U43351 (N_43351,N_41560,N_40334);
or U43352 (N_43352,N_40924,N_41889);
nand U43353 (N_43353,N_41007,N_41806);
xnor U43354 (N_43354,N_41377,N_40903);
nor U43355 (N_43355,N_40446,N_41385);
nor U43356 (N_43356,N_40162,N_40960);
and U43357 (N_43357,N_41194,N_41653);
xnor U43358 (N_43358,N_41195,N_40874);
xor U43359 (N_43359,N_40293,N_41862);
xnor U43360 (N_43360,N_40199,N_41097);
xor U43361 (N_43361,N_41508,N_40308);
nand U43362 (N_43362,N_40474,N_40416);
nand U43363 (N_43363,N_40684,N_40117);
xnor U43364 (N_43364,N_41382,N_41009);
nand U43365 (N_43365,N_40077,N_40598);
xnor U43366 (N_43366,N_41635,N_40526);
xnor U43367 (N_43367,N_40165,N_41970);
and U43368 (N_43368,N_40477,N_40799);
and U43369 (N_43369,N_41302,N_41654);
or U43370 (N_43370,N_41914,N_40869);
nor U43371 (N_43371,N_41456,N_40425);
and U43372 (N_43372,N_41675,N_41823);
and U43373 (N_43373,N_40559,N_40487);
xnor U43374 (N_43374,N_41397,N_40502);
nor U43375 (N_43375,N_40987,N_41798);
or U43376 (N_43376,N_41509,N_40630);
nand U43377 (N_43377,N_41198,N_41184);
xnor U43378 (N_43378,N_40202,N_41299);
nor U43379 (N_43379,N_40082,N_40858);
nor U43380 (N_43380,N_41789,N_41657);
or U43381 (N_43381,N_40373,N_40360);
or U43382 (N_43382,N_40014,N_41094);
nor U43383 (N_43383,N_40836,N_41434);
nand U43384 (N_43384,N_41132,N_41803);
and U43385 (N_43385,N_40491,N_40487);
xnor U43386 (N_43386,N_41755,N_40971);
nor U43387 (N_43387,N_40404,N_40640);
nor U43388 (N_43388,N_40241,N_40295);
xor U43389 (N_43389,N_40246,N_41808);
xor U43390 (N_43390,N_41346,N_41321);
and U43391 (N_43391,N_41313,N_41733);
or U43392 (N_43392,N_40632,N_40450);
and U43393 (N_43393,N_41309,N_41837);
or U43394 (N_43394,N_40300,N_40571);
or U43395 (N_43395,N_40109,N_41703);
nand U43396 (N_43396,N_40434,N_40740);
nand U43397 (N_43397,N_41313,N_40670);
or U43398 (N_43398,N_41432,N_41349);
xnor U43399 (N_43399,N_40558,N_41048);
and U43400 (N_43400,N_41711,N_41057);
and U43401 (N_43401,N_40646,N_41531);
xnor U43402 (N_43402,N_40863,N_40481);
and U43403 (N_43403,N_41385,N_41430);
or U43404 (N_43404,N_41742,N_40603);
xor U43405 (N_43405,N_41872,N_40024);
nor U43406 (N_43406,N_41527,N_40806);
nor U43407 (N_43407,N_41874,N_40647);
nand U43408 (N_43408,N_40829,N_40242);
nand U43409 (N_43409,N_40328,N_40999);
nand U43410 (N_43410,N_41583,N_40938);
or U43411 (N_43411,N_41421,N_41248);
and U43412 (N_43412,N_40785,N_41795);
and U43413 (N_43413,N_41822,N_41082);
or U43414 (N_43414,N_40565,N_40916);
nor U43415 (N_43415,N_40539,N_41001);
xor U43416 (N_43416,N_40300,N_40491);
xor U43417 (N_43417,N_40081,N_40780);
nor U43418 (N_43418,N_41737,N_40241);
and U43419 (N_43419,N_40578,N_41449);
xor U43420 (N_43420,N_41839,N_40262);
nor U43421 (N_43421,N_41119,N_40953);
or U43422 (N_43422,N_41889,N_40229);
xnor U43423 (N_43423,N_41412,N_40097);
nor U43424 (N_43424,N_40339,N_40912);
or U43425 (N_43425,N_41576,N_40953);
or U43426 (N_43426,N_41400,N_41730);
xor U43427 (N_43427,N_41994,N_40877);
xnor U43428 (N_43428,N_41759,N_41429);
or U43429 (N_43429,N_40305,N_40390);
or U43430 (N_43430,N_41612,N_40380);
nand U43431 (N_43431,N_41538,N_40293);
and U43432 (N_43432,N_40221,N_41746);
and U43433 (N_43433,N_40646,N_40898);
and U43434 (N_43434,N_41237,N_40342);
nand U43435 (N_43435,N_41854,N_41351);
nor U43436 (N_43436,N_41177,N_41937);
nor U43437 (N_43437,N_40673,N_41126);
or U43438 (N_43438,N_41399,N_40781);
or U43439 (N_43439,N_40220,N_40495);
xor U43440 (N_43440,N_41874,N_41948);
nor U43441 (N_43441,N_41369,N_41335);
nor U43442 (N_43442,N_41787,N_41918);
nor U43443 (N_43443,N_41833,N_41710);
xnor U43444 (N_43444,N_40099,N_41903);
nand U43445 (N_43445,N_41885,N_41458);
or U43446 (N_43446,N_40964,N_41760);
or U43447 (N_43447,N_41457,N_41192);
nor U43448 (N_43448,N_41356,N_40593);
nand U43449 (N_43449,N_41591,N_41278);
nor U43450 (N_43450,N_40697,N_41848);
and U43451 (N_43451,N_40669,N_40942);
nor U43452 (N_43452,N_40742,N_40320);
nor U43453 (N_43453,N_41809,N_40524);
or U43454 (N_43454,N_40927,N_40528);
nand U43455 (N_43455,N_40580,N_41136);
or U43456 (N_43456,N_41587,N_40441);
nand U43457 (N_43457,N_41313,N_41413);
or U43458 (N_43458,N_41124,N_40385);
nor U43459 (N_43459,N_40678,N_40324);
nand U43460 (N_43460,N_41511,N_41660);
and U43461 (N_43461,N_40004,N_40345);
or U43462 (N_43462,N_41219,N_41111);
xor U43463 (N_43463,N_41352,N_40368);
nand U43464 (N_43464,N_40287,N_41214);
and U43465 (N_43465,N_40560,N_41315);
and U43466 (N_43466,N_41725,N_41396);
xnor U43467 (N_43467,N_41788,N_40291);
nand U43468 (N_43468,N_41589,N_41976);
nor U43469 (N_43469,N_41374,N_40088);
nor U43470 (N_43470,N_41482,N_41191);
or U43471 (N_43471,N_40367,N_41164);
nand U43472 (N_43472,N_40279,N_41698);
nor U43473 (N_43473,N_40968,N_41641);
or U43474 (N_43474,N_41654,N_41214);
and U43475 (N_43475,N_41890,N_41166);
and U43476 (N_43476,N_40424,N_40198);
or U43477 (N_43477,N_40459,N_40900);
or U43478 (N_43478,N_41176,N_40507);
and U43479 (N_43479,N_41580,N_41315);
and U43480 (N_43480,N_41496,N_40847);
xor U43481 (N_43481,N_41258,N_41459);
nor U43482 (N_43482,N_41170,N_41241);
and U43483 (N_43483,N_40442,N_41280);
xor U43484 (N_43484,N_41461,N_41096);
nand U43485 (N_43485,N_40284,N_40737);
and U43486 (N_43486,N_41127,N_40859);
nand U43487 (N_43487,N_41932,N_41873);
or U43488 (N_43488,N_40503,N_41683);
or U43489 (N_43489,N_40821,N_41184);
nand U43490 (N_43490,N_40719,N_41029);
nand U43491 (N_43491,N_40364,N_40254);
and U43492 (N_43492,N_41660,N_41361);
and U43493 (N_43493,N_41648,N_41390);
xnor U43494 (N_43494,N_41297,N_41951);
xnor U43495 (N_43495,N_40580,N_40072);
nor U43496 (N_43496,N_41082,N_41239);
xor U43497 (N_43497,N_41512,N_40064);
xnor U43498 (N_43498,N_40035,N_41889);
xor U43499 (N_43499,N_41959,N_41356);
nand U43500 (N_43500,N_40466,N_41542);
nand U43501 (N_43501,N_40369,N_40402);
nand U43502 (N_43502,N_40284,N_40524);
and U43503 (N_43503,N_41011,N_41817);
nor U43504 (N_43504,N_41163,N_41342);
xor U43505 (N_43505,N_41202,N_41109);
or U43506 (N_43506,N_40244,N_41460);
xor U43507 (N_43507,N_40661,N_41218);
or U43508 (N_43508,N_40761,N_40115);
xor U43509 (N_43509,N_40042,N_41605);
or U43510 (N_43510,N_40922,N_41134);
or U43511 (N_43511,N_40084,N_41380);
and U43512 (N_43512,N_40553,N_40951);
nand U43513 (N_43513,N_40551,N_41564);
and U43514 (N_43514,N_41427,N_41132);
or U43515 (N_43515,N_40624,N_40736);
xnor U43516 (N_43516,N_41065,N_40719);
nor U43517 (N_43517,N_41107,N_41664);
and U43518 (N_43518,N_41473,N_40545);
xnor U43519 (N_43519,N_40495,N_40093);
and U43520 (N_43520,N_41331,N_40092);
or U43521 (N_43521,N_41257,N_41081);
xnor U43522 (N_43522,N_41934,N_41663);
and U43523 (N_43523,N_40123,N_40868);
nand U43524 (N_43524,N_40493,N_41477);
or U43525 (N_43525,N_40769,N_41225);
or U43526 (N_43526,N_41220,N_40066);
nand U43527 (N_43527,N_41309,N_40878);
xor U43528 (N_43528,N_41802,N_40998);
nor U43529 (N_43529,N_40110,N_40507);
or U43530 (N_43530,N_40960,N_40872);
nor U43531 (N_43531,N_40874,N_40665);
or U43532 (N_43532,N_41584,N_41003);
xnor U43533 (N_43533,N_40028,N_41887);
or U43534 (N_43534,N_41962,N_41406);
and U43535 (N_43535,N_40213,N_40850);
or U43536 (N_43536,N_40623,N_41825);
xor U43537 (N_43537,N_41507,N_40215);
nand U43538 (N_43538,N_40023,N_40621);
xnor U43539 (N_43539,N_40956,N_40701);
nor U43540 (N_43540,N_40055,N_41967);
and U43541 (N_43541,N_40150,N_40411);
nand U43542 (N_43542,N_40258,N_41060);
xnor U43543 (N_43543,N_40799,N_40440);
xor U43544 (N_43544,N_41486,N_40664);
and U43545 (N_43545,N_40828,N_41350);
or U43546 (N_43546,N_41383,N_40025);
nor U43547 (N_43547,N_40487,N_40576);
nand U43548 (N_43548,N_41895,N_41258);
xnor U43549 (N_43549,N_41023,N_41842);
or U43550 (N_43550,N_41250,N_41525);
and U43551 (N_43551,N_40904,N_41882);
nor U43552 (N_43552,N_41884,N_40533);
nand U43553 (N_43553,N_41841,N_40585);
or U43554 (N_43554,N_41163,N_40082);
xnor U43555 (N_43555,N_40806,N_41291);
nor U43556 (N_43556,N_41283,N_40375);
xnor U43557 (N_43557,N_40272,N_40872);
or U43558 (N_43558,N_41001,N_40862);
nand U43559 (N_43559,N_40849,N_41371);
and U43560 (N_43560,N_40540,N_41677);
xor U43561 (N_43561,N_40138,N_40756);
or U43562 (N_43562,N_40315,N_41709);
or U43563 (N_43563,N_41428,N_41218);
nor U43564 (N_43564,N_40805,N_40151);
nand U43565 (N_43565,N_40801,N_41379);
xnor U43566 (N_43566,N_40382,N_41639);
nor U43567 (N_43567,N_41359,N_40300);
and U43568 (N_43568,N_41051,N_41826);
xnor U43569 (N_43569,N_40983,N_40013);
and U43570 (N_43570,N_41814,N_41986);
nor U43571 (N_43571,N_41327,N_41151);
and U43572 (N_43572,N_41799,N_40331);
nand U43573 (N_43573,N_40728,N_40218);
and U43574 (N_43574,N_40207,N_40364);
xnor U43575 (N_43575,N_40657,N_40363);
nor U43576 (N_43576,N_41861,N_41422);
nand U43577 (N_43577,N_41551,N_41945);
or U43578 (N_43578,N_41911,N_40185);
nor U43579 (N_43579,N_40283,N_40622);
and U43580 (N_43580,N_40957,N_41575);
and U43581 (N_43581,N_40238,N_40746);
nor U43582 (N_43582,N_40783,N_41647);
or U43583 (N_43583,N_41063,N_41656);
and U43584 (N_43584,N_40973,N_40797);
or U43585 (N_43585,N_41367,N_41461);
and U43586 (N_43586,N_41250,N_41911);
or U43587 (N_43587,N_41033,N_41126);
nor U43588 (N_43588,N_41267,N_41239);
nand U43589 (N_43589,N_40280,N_40211);
and U43590 (N_43590,N_41211,N_40500);
or U43591 (N_43591,N_40728,N_41748);
nor U43592 (N_43592,N_40604,N_41088);
nor U43593 (N_43593,N_41912,N_41019);
nand U43594 (N_43594,N_41978,N_40408);
or U43595 (N_43595,N_41654,N_41568);
xor U43596 (N_43596,N_40875,N_41677);
and U43597 (N_43597,N_40900,N_40765);
or U43598 (N_43598,N_41590,N_41760);
or U43599 (N_43599,N_41032,N_40664);
nor U43600 (N_43600,N_40537,N_40416);
or U43601 (N_43601,N_40200,N_41134);
xor U43602 (N_43602,N_41379,N_40088);
xor U43603 (N_43603,N_41336,N_41549);
and U43604 (N_43604,N_40134,N_41092);
nor U43605 (N_43605,N_41772,N_41490);
xor U43606 (N_43606,N_40493,N_41853);
nor U43607 (N_43607,N_41138,N_41863);
xnor U43608 (N_43608,N_40957,N_41771);
xnor U43609 (N_43609,N_40062,N_41695);
or U43610 (N_43610,N_41974,N_40192);
nor U43611 (N_43611,N_41590,N_41422);
and U43612 (N_43612,N_40912,N_41878);
and U43613 (N_43613,N_40393,N_40475);
nand U43614 (N_43614,N_40468,N_41182);
xnor U43615 (N_43615,N_40711,N_41137);
and U43616 (N_43616,N_41292,N_41663);
and U43617 (N_43617,N_40906,N_41306);
and U43618 (N_43618,N_40314,N_40898);
and U43619 (N_43619,N_41154,N_41632);
and U43620 (N_43620,N_41977,N_41911);
or U43621 (N_43621,N_41064,N_40711);
nor U43622 (N_43622,N_41479,N_41250);
or U43623 (N_43623,N_40775,N_41557);
nor U43624 (N_43624,N_41747,N_41408);
or U43625 (N_43625,N_41671,N_40027);
and U43626 (N_43626,N_41156,N_41100);
nor U43627 (N_43627,N_41651,N_41706);
nor U43628 (N_43628,N_41059,N_40916);
xnor U43629 (N_43629,N_40368,N_41811);
and U43630 (N_43630,N_41011,N_40410);
xnor U43631 (N_43631,N_40827,N_40525);
and U43632 (N_43632,N_40334,N_41307);
xor U43633 (N_43633,N_40765,N_41325);
nor U43634 (N_43634,N_41532,N_41224);
nor U43635 (N_43635,N_40172,N_40808);
or U43636 (N_43636,N_40380,N_40266);
or U43637 (N_43637,N_40565,N_40332);
and U43638 (N_43638,N_40136,N_41740);
nor U43639 (N_43639,N_40103,N_40783);
nand U43640 (N_43640,N_41186,N_41426);
xor U43641 (N_43641,N_40635,N_41821);
nor U43642 (N_43642,N_40904,N_40956);
nand U43643 (N_43643,N_40997,N_41693);
or U43644 (N_43644,N_41625,N_40577);
xnor U43645 (N_43645,N_41515,N_41676);
or U43646 (N_43646,N_40323,N_41166);
nor U43647 (N_43647,N_41575,N_41549);
nor U43648 (N_43648,N_41119,N_40745);
nand U43649 (N_43649,N_40399,N_40280);
nand U43650 (N_43650,N_41858,N_40986);
nor U43651 (N_43651,N_41374,N_40154);
and U43652 (N_43652,N_40896,N_40964);
xor U43653 (N_43653,N_40885,N_40445);
and U43654 (N_43654,N_41871,N_41553);
nor U43655 (N_43655,N_40389,N_41349);
xor U43656 (N_43656,N_41128,N_40033);
nand U43657 (N_43657,N_40582,N_41747);
or U43658 (N_43658,N_40011,N_40098);
nand U43659 (N_43659,N_40900,N_40367);
nor U43660 (N_43660,N_41952,N_41976);
nand U43661 (N_43661,N_41555,N_41061);
or U43662 (N_43662,N_41543,N_41135);
xnor U43663 (N_43663,N_41094,N_41083);
xor U43664 (N_43664,N_41228,N_40475);
xnor U43665 (N_43665,N_41421,N_40095);
xnor U43666 (N_43666,N_40087,N_41460);
nor U43667 (N_43667,N_41761,N_40989);
and U43668 (N_43668,N_40265,N_40414);
and U43669 (N_43669,N_41832,N_41450);
and U43670 (N_43670,N_41422,N_41753);
nand U43671 (N_43671,N_41939,N_40904);
and U43672 (N_43672,N_41242,N_41570);
xor U43673 (N_43673,N_40552,N_40754);
and U43674 (N_43674,N_40341,N_40513);
xnor U43675 (N_43675,N_40071,N_41464);
nor U43676 (N_43676,N_41676,N_41946);
and U43677 (N_43677,N_40854,N_40907);
nor U43678 (N_43678,N_41076,N_41697);
nand U43679 (N_43679,N_41868,N_40248);
nand U43680 (N_43680,N_41398,N_40618);
xnor U43681 (N_43681,N_40464,N_40305);
nand U43682 (N_43682,N_41230,N_40691);
nand U43683 (N_43683,N_41343,N_40120);
nand U43684 (N_43684,N_41713,N_40367);
nor U43685 (N_43685,N_40499,N_41206);
nor U43686 (N_43686,N_40732,N_40752);
or U43687 (N_43687,N_40638,N_40440);
xnor U43688 (N_43688,N_40995,N_40370);
nand U43689 (N_43689,N_41357,N_40819);
nand U43690 (N_43690,N_40133,N_40958);
xor U43691 (N_43691,N_40086,N_40705);
and U43692 (N_43692,N_41475,N_41293);
or U43693 (N_43693,N_41643,N_41400);
or U43694 (N_43694,N_41077,N_41080);
or U43695 (N_43695,N_41673,N_41197);
nand U43696 (N_43696,N_41815,N_41266);
and U43697 (N_43697,N_40666,N_40931);
xor U43698 (N_43698,N_41257,N_41105);
and U43699 (N_43699,N_41580,N_40605);
xnor U43700 (N_43700,N_40420,N_41890);
nor U43701 (N_43701,N_41686,N_41795);
and U43702 (N_43702,N_41531,N_40713);
nand U43703 (N_43703,N_41064,N_41307);
nand U43704 (N_43704,N_40367,N_40982);
xnor U43705 (N_43705,N_40816,N_41863);
nand U43706 (N_43706,N_40641,N_41104);
xor U43707 (N_43707,N_40383,N_40394);
nand U43708 (N_43708,N_41905,N_40466);
nor U43709 (N_43709,N_40429,N_40092);
or U43710 (N_43710,N_40266,N_41264);
or U43711 (N_43711,N_41196,N_41049);
nand U43712 (N_43712,N_41345,N_40195);
and U43713 (N_43713,N_40745,N_40648);
and U43714 (N_43714,N_41170,N_41884);
nor U43715 (N_43715,N_40854,N_41418);
or U43716 (N_43716,N_40000,N_41379);
nand U43717 (N_43717,N_41901,N_40351);
nor U43718 (N_43718,N_41244,N_40782);
nand U43719 (N_43719,N_41310,N_40381);
and U43720 (N_43720,N_41563,N_40706);
xor U43721 (N_43721,N_41777,N_41296);
xor U43722 (N_43722,N_41884,N_41885);
and U43723 (N_43723,N_41555,N_40084);
nor U43724 (N_43724,N_40612,N_40584);
nor U43725 (N_43725,N_40963,N_41124);
or U43726 (N_43726,N_40194,N_41041);
and U43727 (N_43727,N_41701,N_40974);
or U43728 (N_43728,N_40125,N_40362);
or U43729 (N_43729,N_41981,N_41866);
xnor U43730 (N_43730,N_40004,N_40703);
xor U43731 (N_43731,N_40330,N_41217);
or U43732 (N_43732,N_41528,N_40593);
or U43733 (N_43733,N_40661,N_40528);
nand U43734 (N_43734,N_40703,N_41226);
and U43735 (N_43735,N_41736,N_40475);
nor U43736 (N_43736,N_41442,N_41905);
nor U43737 (N_43737,N_41015,N_40360);
nand U43738 (N_43738,N_40740,N_41299);
or U43739 (N_43739,N_41189,N_41567);
nor U43740 (N_43740,N_40248,N_41811);
and U43741 (N_43741,N_41850,N_41302);
xor U43742 (N_43742,N_41808,N_41797);
xnor U43743 (N_43743,N_41876,N_40654);
xnor U43744 (N_43744,N_41028,N_40847);
nand U43745 (N_43745,N_40644,N_40491);
xnor U43746 (N_43746,N_40698,N_40056);
and U43747 (N_43747,N_40964,N_40471);
nand U43748 (N_43748,N_40581,N_41913);
xnor U43749 (N_43749,N_40573,N_40075);
and U43750 (N_43750,N_41520,N_41803);
nor U43751 (N_43751,N_40315,N_41283);
nand U43752 (N_43752,N_41907,N_40361);
nor U43753 (N_43753,N_40837,N_40471);
nor U43754 (N_43754,N_41834,N_41099);
xor U43755 (N_43755,N_40182,N_41215);
xnor U43756 (N_43756,N_40525,N_40505);
or U43757 (N_43757,N_41095,N_41592);
nand U43758 (N_43758,N_41085,N_40084);
and U43759 (N_43759,N_40342,N_40285);
and U43760 (N_43760,N_40095,N_40770);
nand U43761 (N_43761,N_41140,N_41650);
and U43762 (N_43762,N_41868,N_41254);
or U43763 (N_43763,N_40238,N_40970);
xor U43764 (N_43764,N_41718,N_41168);
and U43765 (N_43765,N_40452,N_41846);
xnor U43766 (N_43766,N_40379,N_41386);
xor U43767 (N_43767,N_40886,N_41543);
and U43768 (N_43768,N_40819,N_41355);
and U43769 (N_43769,N_41103,N_40730);
nor U43770 (N_43770,N_41060,N_40706);
nor U43771 (N_43771,N_40620,N_40836);
or U43772 (N_43772,N_41946,N_40125);
xnor U43773 (N_43773,N_40028,N_40648);
xnor U43774 (N_43774,N_40426,N_40646);
xor U43775 (N_43775,N_41815,N_41549);
nor U43776 (N_43776,N_41321,N_41549);
xor U43777 (N_43777,N_41025,N_41865);
nor U43778 (N_43778,N_41597,N_40378);
nor U43779 (N_43779,N_40564,N_40243);
and U43780 (N_43780,N_40233,N_41641);
or U43781 (N_43781,N_40750,N_40571);
nor U43782 (N_43782,N_41989,N_41762);
or U43783 (N_43783,N_40481,N_41211);
and U43784 (N_43784,N_41924,N_40837);
nand U43785 (N_43785,N_41378,N_40517);
and U43786 (N_43786,N_41364,N_41518);
and U43787 (N_43787,N_40312,N_41739);
or U43788 (N_43788,N_41278,N_40103);
nor U43789 (N_43789,N_40106,N_40325);
xor U43790 (N_43790,N_40500,N_41343);
xor U43791 (N_43791,N_40713,N_40258);
or U43792 (N_43792,N_40668,N_40162);
xor U43793 (N_43793,N_41194,N_40140);
and U43794 (N_43794,N_41469,N_40599);
and U43795 (N_43795,N_40667,N_41002);
and U43796 (N_43796,N_40051,N_40836);
nor U43797 (N_43797,N_41476,N_41473);
and U43798 (N_43798,N_40567,N_41437);
or U43799 (N_43799,N_41549,N_40917);
or U43800 (N_43800,N_40673,N_40182);
nand U43801 (N_43801,N_40253,N_41968);
nor U43802 (N_43802,N_41760,N_41882);
nor U43803 (N_43803,N_40976,N_41356);
or U43804 (N_43804,N_40672,N_40121);
and U43805 (N_43805,N_40360,N_40515);
or U43806 (N_43806,N_41944,N_41566);
or U43807 (N_43807,N_41979,N_40513);
nor U43808 (N_43808,N_41192,N_40966);
xnor U43809 (N_43809,N_41532,N_40911);
and U43810 (N_43810,N_41170,N_40867);
and U43811 (N_43811,N_40181,N_41663);
and U43812 (N_43812,N_41443,N_41655);
nand U43813 (N_43813,N_41582,N_40381);
and U43814 (N_43814,N_41167,N_40804);
xnor U43815 (N_43815,N_40780,N_40518);
xor U43816 (N_43816,N_40829,N_41577);
and U43817 (N_43817,N_40782,N_41072);
or U43818 (N_43818,N_40703,N_41431);
nor U43819 (N_43819,N_41180,N_41434);
and U43820 (N_43820,N_40816,N_41798);
xnor U43821 (N_43821,N_41577,N_41969);
nand U43822 (N_43822,N_41213,N_40440);
and U43823 (N_43823,N_41285,N_40037);
nor U43824 (N_43824,N_41416,N_40622);
xor U43825 (N_43825,N_41811,N_41399);
nand U43826 (N_43826,N_41861,N_41814);
nand U43827 (N_43827,N_41595,N_40159);
and U43828 (N_43828,N_40597,N_41507);
and U43829 (N_43829,N_41364,N_40532);
or U43830 (N_43830,N_40907,N_41578);
and U43831 (N_43831,N_40693,N_40361);
nand U43832 (N_43832,N_40617,N_40361);
nand U43833 (N_43833,N_41224,N_40872);
nand U43834 (N_43834,N_40947,N_41095);
and U43835 (N_43835,N_41911,N_40686);
nand U43836 (N_43836,N_41419,N_40746);
and U43837 (N_43837,N_41991,N_40880);
nor U43838 (N_43838,N_40493,N_40119);
or U43839 (N_43839,N_40671,N_41284);
xnor U43840 (N_43840,N_41330,N_41572);
and U43841 (N_43841,N_41449,N_41252);
nor U43842 (N_43842,N_41028,N_40573);
nor U43843 (N_43843,N_41006,N_41297);
nor U43844 (N_43844,N_41915,N_41760);
nor U43845 (N_43845,N_41570,N_40409);
nand U43846 (N_43846,N_41987,N_41849);
nor U43847 (N_43847,N_40060,N_40440);
and U43848 (N_43848,N_41814,N_40803);
and U43849 (N_43849,N_40521,N_40088);
nand U43850 (N_43850,N_40622,N_41802);
and U43851 (N_43851,N_41250,N_41795);
xor U43852 (N_43852,N_40559,N_40724);
nand U43853 (N_43853,N_40928,N_41353);
or U43854 (N_43854,N_41274,N_41501);
nor U43855 (N_43855,N_40729,N_40086);
xnor U43856 (N_43856,N_41847,N_41275);
nor U43857 (N_43857,N_41684,N_40733);
and U43858 (N_43858,N_41071,N_40981);
nor U43859 (N_43859,N_41289,N_41332);
nor U43860 (N_43860,N_40895,N_41933);
xor U43861 (N_43861,N_41303,N_40625);
xor U43862 (N_43862,N_41239,N_40569);
nand U43863 (N_43863,N_40026,N_41963);
nor U43864 (N_43864,N_41622,N_40503);
or U43865 (N_43865,N_41386,N_41905);
xor U43866 (N_43866,N_40012,N_41573);
nand U43867 (N_43867,N_40379,N_41374);
or U43868 (N_43868,N_41534,N_40150);
nor U43869 (N_43869,N_40737,N_40223);
or U43870 (N_43870,N_40630,N_40466);
nand U43871 (N_43871,N_41500,N_41621);
or U43872 (N_43872,N_41322,N_40813);
and U43873 (N_43873,N_41372,N_40563);
and U43874 (N_43874,N_40458,N_41822);
or U43875 (N_43875,N_41068,N_40512);
and U43876 (N_43876,N_41381,N_41312);
or U43877 (N_43877,N_40004,N_41089);
xor U43878 (N_43878,N_41234,N_41991);
and U43879 (N_43879,N_40651,N_41610);
xnor U43880 (N_43880,N_41802,N_41378);
nand U43881 (N_43881,N_40702,N_40039);
nand U43882 (N_43882,N_41560,N_40852);
nor U43883 (N_43883,N_40137,N_40927);
xor U43884 (N_43884,N_41542,N_41736);
nor U43885 (N_43885,N_41949,N_40856);
or U43886 (N_43886,N_40204,N_40689);
nor U43887 (N_43887,N_41328,N_41322);
nand U43888 (N_43888,N_40120,N_41582);
nand U43889 (N_43889,N_40423,N_41855);
or U43890 (N_43890,N_40061,N_40208);
and U43891 (N_43891,N_41819,N_40439);
or U43892 (N_43892,N_41300,N_40230);
nor U43893 (N_43893,N_40303,N_41395);
nor U43894 (N_43894,N_41079,N_40954);
xnor U43895 (N_43895,N_40276,N_41476);
and U43896 (N_43896,N_40646,N_41705);
or U43897 (N_43897,N_40194,N_40299);
and U43898 (N_43898,N_41267,N_41053);
nand U43899 (N_43899,N_40920,N_40440);
or U43900 (N_43900,N_41407,N_41581);
or U43901 (N_43901,N_41831,N_41710);
nor U43902 (N_43902,N_40473,N_41009);
xnor U43903 (N_43903,N_41590,N_41767);
nand U43904 (N_43904,N_41346,N_40074);
nor U43905 (N_43905,N_40006,N_40870);
xnor U43906 (N_43906,N_41784,N_40087);
and U43907 (N_43907,N_40424,N_40776);
or U43908 (N_43908,N_40767,N_41025);
xnor U43909 (N_43909,N_41347,N_41381);
and U43910 (N_43910,N_40226,N_41188);
or U43911 (N_43911,N_40271,N_41357);
nor U43912 (N_43912,N_41228,N_41909);
or U43913 (N_43913,N_40269,N_40338);
or U43914 (N_43914,N_40010,N_40621);
or U43915 (N_43915,N_41988,N_41661);
and U43916 (N_43916,N_40910,N_40440);
nand U43917 (N_43917,N_40761,N_41237);
or U43918 (N_43918,N_40004,N_40562);
nor U43919 (N_43919,N_41217,N_41518);
or U43920 (N_43920,N_40181,N_40512);
nor U43921 (N_43921,N_41892,N_41720);
or U43922 (N_43922,N_41552,N_41545);
or U43923 (N_43923,N_40760,N_41710);
xor U43924 (N_43924,N_40542,N_40343);
nor U43925 (N_43925,N_40412,N_40388);
nor U43926 (N_43926,N_41689,N_41228);
nor U43927 (N_43927,N_40903,N_40744);
xnor U43928 (N_43928,N_41036,N_40458);
nor U43929 (N_43929,N_41871,N_40738);
xnor U43930 (N_43930,N_40841,N_41693);
nor U43931 (N_43931,N_41374,N_41744);
and U43932 (N_43932,N_40482,N_41092);
nor U43933 (N_43933,N_41814,N_40189);
nand U43934 (N_43934,N_40958,N_41815);
nand U43935 (N_43935,N_41555,N_41744);
nand U43936 (N_43936,N_41671,N_40907);
xor U43937 (N_43937,N_41290,N_40567);
nand U43938 (N_43938,N_41770,N_41005);
nor U43939 (N_43939,N_41812,N_40321);
and U43940 (N_43940,N_41141,N_41117);
or U43941 (N_43941,N_41964,N_41307);
and U43942 (N_43942,N_40937,N_40529);
or U43943 (N_43943,N_41191,N_41921);
nor U43944 (N_43944,N_40366,N_40008);
and U43945 (N_43945,N_40465,N_40138);
and U43946 (N_43946,N_41780,N_40543);
or U43947 (N_43947,N_41385,N_40519);
or U43948 (N_43948,N_40508,N_41828);
and U43949 (N_43949,N_41576,N_41470);
and U43950 (N_43950,N_40815,N_40129);
and U43951 (N_43951,N_41850,N_40679);
and U43952 (N_43952,N_40996,N_41739);
xor U43953 (N_43953,N_41682,N_41101);
and U43954 (N_43954,N_40375,N_41581);
xnor U43955 (N_43955,N_40407,N_41537);
and U43956 (N_43956,N_41774,N_41408);
nor U43957 (N_43957,N_40414,N_40666);
nand U43958 (N_43958,N_40211,N_41979);
nor U43959 (N_43959,N_41227,N_40920);
and U43960 (N_43960,N_40052,N_40834);
xnor U43961 (N_43961,N_40446,N_41202);
nor U43962 (N_43962,N_40376,N_41240);
xor U43963 (N_43963,N_40019,N_41100);
and U43964 (N_43964,N_41426,N_41556);
or U43965 (N_43965,N_41586,N_41062);
nand U43966 (N_43966,N_40872,N_41341);
and U43967 (N_43967,N_41907,N_40523);
xnor U43968 (N_43968,N_41312,N_41610);
nand U43969 (N_43969,N_41033,N_40608);
nand U43970 (N_43970,N_41358,N_41419);
or U43971 (N_43971,N_41510,N_40968);
nand U43972 (N_43972,N_40662,N_41317);
and U43973 (N_43973,N_40372,N_41225);
or U43974 (N_43974,N_41370,N_40820);
nand U43975 (N_43975,N_40453,N_40449);
nor U43976 (N_43976,N_40001,N_40568);
nor U43977 (N_43977,N_40973,N_41246);
nor U43978 (N_43978,N_40259,N_40235);
nor U43979 (N_43979,N_41630,N_40530);
nor U43980 (N_43980,N_40176,N_40776);
nand U43981 (N_43981,N_40840,N_41845);
or U43982 (N_43982,N_41646,N_41892);
xnor U43983 (N_43983,N_41135,N_40221);
nand U43984 (N_43984,N_40754,N_40194);
or U43985 (N_43985,N_40020,N_41588);
xnor U43986 (N_43986,N_40292,N_41385);
nand U43987 (N_43987,N_40721,N_40040);
xnor U43988 (N_43988,N_40363,N_41502);
nand U43989 (N_43989,N_40449,N_41961);
or U43990 (N_43990,N_40221,N_41514);
nand U43991 (N_43991,N_41092,N_40150);
or U43992 (N_43992,N_41008,N_41518);
xnor U43993 (N_43993,N_41777,N_41459);
xor U43994 (N_43994,N_40710,N_41986);
and U43995 (N_43995,N_41775,N_40070);
nor U43996 (N_43996,N_40941,N_40662);
xor U43997 (N_43997,N_41895,N_40034);
and U43998 (N_43998,N_41450,N_40122);
xnor U43999 (N_43999,N_40584,N_41163);
nand U44000 (N_44000,N_42621,N_42131);
nand U44001 (N_44001,N_42062,N_42307);
or U44002 (N_44002,N_43846,N_43956);
or U44003 (N_44003,N_43175,N_42392);
nand U44004 (N_44004,N_42344,N_42419);
xnor U44005 (N_44005,N_42961,N_43081);
xor U44006 (N_44006,N_43067,N_43545);
and U44007 (N_44007,N_43436,N_43162);
nand U44008 (N_44008,N_42539,N_43360);
nor U44009 (N_44009,N_43496,N_42266);
or U44010 (N_44010,N_43110,N_42100);
nand U44011 (N_44011,N_43996,N_43872);
nor U44012 (N_44012,N_43206,N_43517);
nand U44013 (N_44013,N_43873,N_43782);
nand U44014 (N_44014,N_42979,N_42046);
or U44015 (N_44015,N_42987,N_42689);
and U44016 (N_44016,N_42450,N_42826);
or U44017 (N_44017,N_43438,N_43239);
or U44018 (N_44018,N_42608,N_43124);
or U44019 (N_44019,N_42995,N_42099);
nor U44020 (N_44020,N_43020,N_42340);
nand U44021 (N_44021,N_42270,N_43988);
xnor U44022 (N_44022,N_42933,N_43421);
xor U44023 (N_44023,N_42636,N_42323);
nand U44024 (N_44024,N_43544,N_42895);
xor U44025 (N_44025,N_42187,N_42399);
and U44026 (N_44026,N_42715,N_43531);
and U44027 (N_44027,N_43828,N_43981);
and U44028 (N_44028,N_43464,N_42604);
or U44029 (N_44029,N_42506,N_42679);
nor U44030 (N_44030,N_43924,N_42626);
and U44031 (N_44031,N_43332,N_43039);
or U44032 (N_44032,N_43601,N_42547);
or U44033 (N_44033,N_42290,N_43387);
or U44034 (N_44034,N_42023,N_42338);
nand U44035 (N_44035,N_43346,N_43324);
or U44036 (N_44036,N_42137,N_42686);
or U44037 (N_44037,N_43082,N_42842);
nor U44038 (N_44038,N_42162,N_43701);
xnor U44039 (N_44039,N_42410,N_42512);
and U44040 (N_44040,N_43837,N_42646);
or U44041 (N_44041,N_43733,N_43275);
or U44042 (N_44042,N_43207,N_43942);
nand U44043 (N_44043,N_43220,N_43543);
nand U44044 (N_44044,N_42708,N_42225);
and U44045 (N_44045,N_42250,N_43695);
or U44046 (N_44046,N_42366,N_42537);
nand U44047 (N_44047,N_43718,N_42128);
nor U44048 (N_44048,N_43042,N_42601);
and U44049 (N_44049,N_42533,N_42739);
xor U44050 (N_44050,N_43209,N_42781);
and U44051 (N_44051,N_43224,N_42892);
nand U44052 (N_44052,N_43673,N_43474);
nand U44053 (N_44053,N_42520,N_42416);
or U44054 (N_44054,N_42513,N_43471);
or U44055 (N_44055,N_43547,N_43455);
nand U44056 (N_44056,N_42383,N_43613);
xor U44057 (N_44057,N_43909,N_43262);
xnor U44058 (N_44058,N_43505,N_42134);
nor U44059 (N_44059,N_43820,N_43740);
nor U44060 (N_44060,N_43252,N_43867);
xnor U44061 (N_44061,N_43378,N_42274);
and U44062 (N_44062,N_43064,N_43228);
xor U44063 (N_44063,N_43495,N_42069);
xnor U44064 (N_44064,N_43994,N_42996);
or U44065 (N_44065,N_42801,N_42784);
and U44066 (N_44066,N_42991,N_42582);
and U44067 (N_44067,N_43766,N_42977);
nor U44068 (N_44068,N_42171,N_42717);
or U44069 (N_44069,N_42075,N_43699);
nor U44070 (N_44070,N_43221,N_43935);
and U44071 (N_44071,N_43053,N_43112);
nor U44072 (N_44072,N_42551,N_42365);
and U44073 (N_44073,N_42030,N_42893);
or U44074 (N_44074,N_42792,N_43371);
xor U44075 (N_44075,N_42460,N_42321);
or U44076 (N_44076,N_43961,N_43071);
xor U44077 (N_44077,N_42106,N_43411);
nor U44078 (N_44078,N_43073,N_42959);
or U44079 (N_44079,N_43612,N_42249);
and U44080 (N_44080,N_42662,N_43927);
nor U44081 (N_44081,N_42643,N_43891);
xor U44082 (N_44082,N_42670,N_43434);
or U44083 (N_44083,N_43282,N_43598);
xor U44084 (N_44084,N_43018,N_43550);
nor U44085 (N_44085,N_42142,N_43466);
xnor U44086 (N_44086,N_43095,N_43085);
and U44087 (N_44087,N_42884,N_42754);
or U44088 (N_44088,N_42727,N_43204);
nor U44089 (N_44089,N_42605,N_42087);
and U44090 (N_44090,N_43687,N_43266);
or U44091 (N_44091,N_43934,N_42310);
nor U44092 (N_44092,N_42751,N_43458);
and U44093 (N_44093,N_42701,N_43803);
and U44094 (N_44094,N_42864,N_42793);
nand U44095 (N_44095,N_42967,N_43952);
nor U44096 (N_44096,N_42151,N_43274);
and U44097 (N_44097,N_42871,N_42259);
and U44098 (N_44098,N_43745,N_42090);
or U44099 (N_44099,N_42824,N_43088);
xnor U44100 (N_44100,N_43995,N_43549);
xnor U44101 (N_44101,N_43032,N_43164);
nand U44102 (N_44102,N_43717,N_43034);
and U44103 (N_44103,N_43509,N_43723);
nor U44104 (N_44104,N_43379,N_42080);
nand U44105 (N_44105,N_43280,N_43128);
and U44106 (N_44106,N_43140,N_42291);
nand U44107 (N_44107,N_42854,N_42822);
nor U44108 (N_44108,N_43491,N_43838);
nand U44109 (N_44109,N_42070,N_43972);
xnor U44110 (N_44110,N_43035,N_42029);
xnor U44111 (N_44111,N_42578,N_43494);
xor U44112 (N_44112,N_42200,N_43893);
nor U44113 (N_44113,N_43527,N_43542);
nor U44114 (N_44114,N_43991,N_43094);
nand U44115 (N_44115,N_42909,N_43932);
nand U44116 (N_44116,N_42060,N_42233);
nand U44117 (N_44117,N_43538,N_43072);
or U44118 (N_44118,N_42504,N_42101);
nor U44119 (N_44119,N_42294,N_43056);
nor U44120 (N_44120,N_42583,N_42944);
nand U44121 (N_44121,N_42089,N_42467);
nor U44122 (N_44122,N_42082,N_42839);
nor U44123 (N_44123,N_43815,N_42810);
or U44124 (N_44124,N_43345,N_43062);
nand U44125 (N_44125,N_43040,N_42345);
nand U44126 (N_44126,N_42865,N_43487);
or U44127 (N_44127,N_42245,N_42503);
and U44128 (N_44128,N_43394,N_42305);
nor U44129 (N_44129,N_42614,N_42063);
and U44130 (N_44130,N_43182,N_42386);
xor U44131 (N_44131,N_43727,N_42502);
nand U44132 (N_44132,N_42456,N_42086);
and U44133 (N_44133,N_43340,N_43615);
or U44134 (N_44134,N_43810,N_43233);
xnor U44135 (N_44135,N_43578,N_42960);
nor U44136 (N_44136,N_42038,N_42427);
xor U44137 (N_44137,N_43045,N_42789);
and U44138 (N_44138,N_43059,N_43962);
nand U44139 (N_44139,N_42630,N_43882);
nand U44140 (N_44140,N_43530,N_43851);
nand U44141 (N_44141,N_42451,N_43364);
xnor U44142 (N_44142,N_43533,N_43572);
or U44143 (N_44143,N_42804,N_42667);
nor U44144 (N_44144,N_42130,N_42753);
or U44145 (N_44145,N_43857,N_42415);
or U44146 (N_44146,N_43116,N_42546);
nor U44147 (N_44147,N_43048,N_42591);
nand U44148 (N_44148,N_43150,N_42396);
xor U44149 (N_44149,N_43693,N_43917);
xnor U44150 (N_44150,N_42420,N_43284);
or U44151 (N_44151,N_42828,N_42855);
and U44152 (N_44152,N_43675,N_42264);
xnor U44153 (N_44153,N_42102,N_42095);
and U44154 (N_44154,N_42375,N_42287);
nand U44155 (N_44155,N_43806,N_43084);
and U44156 (N_44156,N_43573,N_42774);
xor U44157 (N_44157,N_42722,N_42153);
nand U44158 (N_44158,N_42242,N_43419);
nand U44159 (N_44159,N_42756,N_42606);
nand U44160 (N_44160,N_42536,N_43512);
or U44161 (N_44161,N_42105,N_42692);
or U44162 (N_44162,N_43694,N_42508);
nand U44163 (N_44163,N_42769,N_43367);
nor U44164 (N_44164,N_42350,N_43377);
nor U44165 (N_44165,N_42501,N_42559);
or U44166 (N_44166,N_42829,N_42883);
and U44167 (N_44167,N_43422,N_42455);
nor U44168 (N_44168,N_42252,N_43634);
nand U44169 (N_44169,N_42992,N_43807);
xor U44170 (N_44170,N_43076,N_43606);
nand U44171 (N_44171,N_42542,N_43448);
or U44172 (N_44172,N_42093,N_42956);
xor U44173 (N_44173,N_43513,N_42555);
nor U44174 (N_44174,N_42232,N_42285);
nor U44175 (N_44175,N_43643,N_42115);
nor U44176 (N_44176,N_42619,N_42488);
or U44177 (N_44177,N_42726,N_43490);
xor U44178 (N_44178,N_43117,N_42586);
nor U44179 (N_44179,N_42429,N_43030);
and U44180 (N_44180,N_43715,N_42009);
nand U44181 (N_44181,N_43290,N_42728);
nor U44182 (N_44182,N_43516,N_43788);
nand U44183 (N_44183,N_42024,N_43721);
nand U44184 (N_44184,N_42900,N_43099);
nor U44185 (N_44185,N_43015,N_43257);
xnor U44186 (N_44186,N_42948,N_43485);
nand U44187 (N_44187,N_42048,N_43218);
or U44188 (N_44188,N_42665,N_42529);
and U44189 (N_44189,N_42697,N_43966);
xnor U44190 (N_44190,N_43472,N_42022);
nand U44191 (N_44191,N_43250,N_43482);
xnor U44192 (N_44192,N_42886,N_42440);
or U44193 (N_44193,N_42898,N_43534);
nand U44194 (N_44194,N_43597,N_43238);
and U44195 (N_44195,N_42858,N_42571);
or U44196 (N_44196,N_42940,N_42906);
or U44197 (N_44197,N_42120,N_43139);
or U44198 (N_44198,N_42421,N_42660);
and U44199 (N_44199,N_43920,N_42182);
nor U44200 (N_44200,N_43147,N_42470);
nor U44201 (N_44201,N_42866,N_42067);
or U44202 (N_44202,N_42928,N_42808);
xnor U44203 (N_44203,N_43347,N_43342);
and U44204 (N_44204,N_43753,N_42281);
xnor U44205 (N_44205,N_42704,N_42851);
and U44206 (N_44206,N_43603,N_43309);
xnor U44207 (N_44207,N_42320,N_43338);
and U44208 (N_44208,N_42339,N_43968);
nand U44209 (N_44209,N_43412,N_42318);
and U44210 (N_44210,N_42618,N_42723);
nor U44211 (N_44211,N_43594,N_42229);
nand U44212 (N_44212,N_43819,N_43213);
or U44213 (N_44213,N_43922,N_42325);
and U44214 (N_44214,N_43096,N_43013);
and U44215 (N_44215,N_42393,N_43362);
and U44216 (N_44216,N_42935,N_43826);
nand U44217 (N_44217,N_43781,N_43146);
xor U44218 (N_44218,N_43584,N_43017);
nor U44219 (N_44219,N_42327,N_42800);
xnor U44220 (N_44220,N_43575,N_43236);
or U44221 (N_44221,N_42872,N_43925);
xor U44222 (N_44222,N_43814,N_42224);
or U44223 (N_44223,N_42317,N_42355);
or U44224 (N_44224,N_42146,N_43794);
or U44225 (N_44225,N_43936,N_42141);
or U44226 (N_44226,N_42389,N_42004);
nand U44227 (N_44227,N_42112,N_43289);
or U44228 (N_44228,N_43525,N_43460);
or U44229 (N_44229,N_42277,N_43254);
or U44230 (N_44230,N_43319,N_43590);
and U44231 (N_44231,N_43748,N_43883);
or U44232 (N_44232,N_43208,N_43155);
nor U44233 (N_44233,N_43610,N_42199);
nand U44234 (N_44234,N_43977,N_42209);
nor U44235 (N_44235,N_42139,N_43058);
and U44236 (N_44236,N_42494,N_42525);
or U44237 (N_44237,N_43611,N_42005);
and U44238 (N_44238,N_43149,N_42113);
or U44239 (N_44239,N_42442,N_42714);
nand U44240 (N_44240,N_42170,N_42486);
nor U44241 (N_44241,N_42816,N_43514);
and U44242 (N_44242,N_43439,N_42477);
or U44243 (N_44243,N_43044,N_43014);
or U44244 (N_44244,N_42337,N_42836);
or U44245 (N_44245,N_42600,N_42984);
and U44246 (N_44246,N_42700,N_43344);
xor U44247 (N_44247,N_42603,N_42762);
nor U44248 (N_44248,N_43442,N_43716);
or U44249 (N_44249,N_42741,N_42351);
or U44250 (N_44250,N_43009,N_42179);
xor U44251 (N_44251,N_42878,N_42772);
nor U44252 (N_44252,N_42947,N_43349);
nand U44253 (N_44253,N_42138,N_42358);
or U44254 (N_44254,N_42193,N_43536);
xor U44255 (N_44255,N_43363,N_42805);
nor U44256 (N_44256,N_43944,N_42843);
nand U44257 (N_44257,N_43609,N_43772);
nor U44258 (N_44258,N_43417,N_43292);
nand U44259 (N_44259,N_43583,N_42856);
or U44260 (N_44260,N_42719,N_43993);
xnor U44261 (N_44261,N_42236,N_42584);
xnor U44262 (N_44262,N_43410,N_42292);
nand U44263 (N_44263,N_43736,N_42384);
or U44264 (N_44264,N_43260,N_43126);
or U44265 (N_44265,N_42914,N_42922);
or U44266 (N_44266,N_42219,N_43335);
nor U44267 (N_44267,N_43777,N_43385);
nand U44268 (N_44268,N_42234,N_43551);
nor U44269 (N_44269,N_43728,N_43582);
nor U44270 (N_44270,N_43180,N_42011);
or U44271 (N_44271,N_43690,N_42682);
or U44272 (N_44272,N_43350,N_43998);
nor U44273 (N_44273,N_43565,N_42316);
nand U44274 (N_44274,N_42255,N_43322);
nand U44275 (N_44275,N_42220,N_42484);
and U44276 (N_44276,N_43369,N_42212);
nor U44277 (N_44277,N_43051,N_42709);
xnor U44278 (N_44278,N_43423,N_42616);
or U44279 (N_44279,N_43674,N_42077);
xor U44280 (N_44280,N_42847,N_43918);
or U44281 (N_44281,N_42574,N_43089);
or U44282 (N_44282,N_43510,N_43231);
nand U44283 (N_44283,N_42196,N_42857);
xnor U44284 (N_44284,N_42482,N_43714);
nand U44285 (N_44285,N_42109,N_42370);
and U44286 (N_44286,N_42698,N_43878);
xnor U44287 (N_44287,N_42541,N_42336);
and U44288 (N_44288,N_43811,N_43554);
nand U44289 (N_44289,N_43604,N_42163);
nor U44290 (N_44290,N_42730,N_43227);
xnor U44291 (N_44291,N_43672,N_42204);
xnor U44292 (N_44292,N_43524,N_42406);
and U44293 (N_44293,N_42126,N_43800);
or U44294 (N_44294,N_42642,N_42713);
xor U44295 (N_44295,N_43910,N_42631);
nor U44296 (N_44296,N_43946,N_42381);
nor U44297 (N_44297,N_42990,N_42729);
nand U44298 (N_44298,N_43109,N_43237);
or U44299 (N_44299,N_42639,N_43090);
nor U44300 (N_44300,N_42590,N_42711);
or U44301 (N_44301,N_42088,N_43001);
nand U44302 (N_44302,N_42882,N_43852);
and U44303 (N_44303,N_42195,N_43200);
nor U44304 (N_44304,N_43398,N_42217);
or U44305 (N_44305,N_42716,N_43376);
xnor U44306 (N_44306,N_42577,N_43667);
or U44307 (N_44307,N_43930,N_42260);
xnor U44308 (N_44308,N_42066,N_42835);
nand U44309 (N_44309,N_43905,N_42083);
nor U44310 (N_44310,N_43468,N_42201);
nand U44311 (N_44311,N_42795,N_42210);
xnor U44312 (N_44312,N_43470,N_42638);
nor U44313 (N_44313,N_43562,N_42481);
nand U44314 (N_44314,N_42309,N_42184);
xor U44315 (N_44315,N_43348,N_43989);
nor U44316 (N_44316,N_43193,N_43300);
nand U44317 (N_44317,N_43560,N_43440);
xor U44318 (N_44318,N_42955,N_42827);
or U44319 (N_44319,N_43526,N_42174);
nand U44320 (N_44320,N_43003,N_43396);
xnor U44321 (N_44321,N_43884,N_42458);
nand U44322 (N_44322,N_43179,N_43092);
nand U44323 (N_44323,N_42438,N_42025);
or U44324 (N_44324,N_42013,N_42020);
and U44325 (N_44325,N_43774,N_43520);
and U44326 (N_44326,N_42957,N_42966);
xor U44327 (N_44327,N_43600,N_43523);
nor U44328 (N_44328,N_42687,N_43244);
xor U44329 (N_44329,N_43038,N_42258);
and U44330 (N_44330,N_43158,N_42760);
nor U44331 (N_44331,N_43314,N_43638);
nand U44332 (N_44332,N_43521,N_43426);
nand U44333 (N_44333,N_42441,N_43165);
nor U44334 (N_44334,N_42403,N_42937);
nand U44335 (N_44335,N_43689,N_43783);
xnor U44336 (N_44336,N_42941,N_43382);
and U44337 (N_44337,N_42357,N_42268);
or U44338 (N_44338,N_42054,N_42362);
and U44339 (N_44339,N_43005,N_42635);
nand U44340 (N_44340,N_43025,N_43087);
and U44341 (N_44341,N_43368,N_43401);
and U44342 (N_44342,N_42495,N_42404);
xnor U44343 (N_44343,N_43268,N_42908);
xnor U44344 (N_44344,N_42669,N_42263);
nor U44345 (N_44345,N_43686,N_43093);
xnor U44346 (N_44346,N_43418,N_43974);
and U44347 (N_44347,N_43668,N_43446);
xnor U44348 (N_44348,N_43608,N_42324);
and U44349 (N_44349,N_43651,N_42989);
xor U44350 (N_44350,N_42845,N_43476);
nor U44351 (N_44351,N_42019,N_42045);
nand U44352 (N_44352,N_43215,N_42167);
xor U44353 (N_44353,N_42887,N_42863);
nor U44354 (N_44354,N_42183,N_43901);
nand U44355 (N_44355,N_42850,N_43399);
nor U44356 (N_44356,N_43896,N_43160);
or U44357 (N_44357,N_43291,N_43450);
or U44358 (N_44358,N_42777,N_43163);
nor U44359 (N_44359,N_42147,N_42748);
xor U44360 (N_44360,N_42918,N_43190);
nor U44361 (N_44361,N_42581,N_43641);
or U44362 (N_44362,N_42830,N_42683);
nand U44363 (N_44363,N_42852,N_43692);
and U44364 (N_44364,N_42027,N_42594);
nor U44365 (N_44365,N_43189,N_42511);
and U44366 (N_44366,N_42738,N_42272);
nand U44367 (N_44367,N_43980,N_42040);
nor U44368 (N_44368,N_43768,N_42602);
nand U44369 (N_44369,N_42230,N_43311);
or U44370 (N_44370,N_42223,N_42471);
or U44371 (N_44371,N_42794,N_43123);
and U44372 (N_44372,N_42819,N_42433);
xnor U44373 (N_44373,N_43169,N_43395);
or U44374 (N_44374,N_43241,N_43636);
xnor U44375 (N_44375,N_43779,N_42862);
xnor U44376 (N_44376,N_43897,N_43965);
nand U44377 (N_44377,N_43743,N_43817);
xnor U44378 (N_44378,N_42731,N_42764);
nor U44379 (N_44379,N_43908,N_43862);
nand U44380 (N_44380,N_43913,N_42676);
or U44381 (N_44381,N_42859,N_43711);
xnor U44382 (N_44382,N_42962,N_43279);
nand U44383 (N_44383,N_43767,N_43240);
nor U44384 (N_44384,N_43397,N_43881);
nor U44385 (N_44385,N_42919,N_42622);
or U44386 (N_44386,N_42519,N_43469);
xor U44387 (N_44387,N_43522,N_43402);
or U44388 (N_44388,N_43447,N_42288);
and U44389 (N_44389,N_43122,N_42304);
nand U44390 (N_44390,N_43336,N_42592);
xor U44391 (N_44391,N_42656,N_42369);
and U44392 (N_44392,N_43131,N_43963);
nor U44393 (N_44393,N_43742,N_43478);
or U44394 (N_44394,N_42673,N_43958);
and U44395 (N_44395,N_42628,N_43619);
and U44396 (N_44396,N_43571,N_42097);
nand U44397 (N_44397,N_43329,N_42275);
or U44398 (N_44398,N_42319,N_43177);
and U44399 (N_44399,N_43443,N_42579);
xnor U44400 (N_44400,N_43926,N_42043);
and U44401 (N_44401,N_42205,N_42213);
and U44402 (N_44402,N_43272,N_42780);
and U44403 (N_44403,N_43790,N_42376);
or U44404 (N_44404,N_43245,N_42939);
or U44405 (N_44405,N_43276,N_43670);
nand U44406 (N_44406,N_43498,N_42159);
nor U44407 (N_44407,N_42874,N_43143);
or U44408 (N_44408,N_42480,N_43635);
nor U44409 (N_44409,N_42189,N_42071);
xnor U44410 (N_44410,N_42123,N_42752);
or U44411 (N_44411,N_43381,N_43293);
and U44412 (N_44412,N_42640,N_43201);
or U44413 (N_44413,N_42545,N_42968);
or U44414 (N_44414,N_43054,N_43984);
and U44415 (N_44415,N_42166,N_42761);
or U44416 (N_44416,N_42814,N_43312);
xor U44417 (N_44417,N_43049,N_42215);
or U44418 (N_44418,N_42790,N_42037);
xnor U44419 (N_44419,N_42889,N_43326);
nor U44420 (N_44420,N_43100,N_43586);
xnor U44421 (N_44421,N_42988,N_42273);
nor U44422 (N_44422,N_43372,N_43931);
xor U44423 (N_44423,N_42976,N_43880);
xor U44424 (N_44424,N_43771,N_42952);
and U44425 (N_44425,N_42791,N_43305);
and U44426 (N_44426,N_43626,N_43754);
and U44427 (N_44427,N_43113,N_43654);
nand U44428 (N_44428,N_43484,N_42148);
nor U44429 (N_44429,N_43392,N_43919);
nor U44430 (N_44430,N_42012,N_42565);
or U44431 (N_44431,N_42911,N_43557);
and U44432 (N_44432,N_43106,N_42500);
nand U44433 (N_44433,N_43269,N_43210);
xor U44434 (N_44434,N_42910,N_43202);
xor U44435 (N_44435,N_42931,N_42747);
nand U44436 (N_44436,N_42671,N_43313);
or U44437 (N_44437,N_42688,N_43429);
and U44438 (N_44438,N_43083,N_43595);
xnor U44439 (N_44439,N_43960,N_43135);
nor U44440 (N_44440,N_42107,N_43877);
nand U44441 (N_44441,N_42478,N_42188);
or U44442 (N_44442,N_42629,N_43341);
nor U44443 (N_44443,N_42133,N_43415);
xor U44444 (N_44444,N_43957,N_43178);
xor U44445 (N_44445,N_42749,N_43853);
xor U44446 (N_44446,N_42017,N_42524);
nor U44447 (N_44447,N_43849,N_43888);
and U44448 (N_44448,N_42462,N_43055);
and U44449 (N_44449,N_43142,N_43101);
and U44450 (N_44450,N_43663,N_42932);
xnor U44451 (N_44451,N_43389,N_43223);
nand U44452 (N_44452,N_43581,N_42228);
nand U44453 (N_44453,N_42057,N_42896);
or U44454 (N_44454,N_43705,N_43752);
or U44455 (N_44455,N_42509,N_43625);
xnor U44456 (N_44456,N_42981,N_42257);
nor U44457 (N_44457,N_42117,N_42530);
nor U44458 (N_44458,N_43688,N_42475);
nor U44459 (N_44459,N_42185,N_42768);
nand U44460 (N_44460,N_43869,N_42818);
nand U44461 (N_44461,N_43899,N_43004);
or U44462 (N_44462,N_43120,N_42554);
xnor U44463 (N_44463,N_42876,N_42437);
or U44464 (N_44464,N_43703,N_43744);
nor U44465 (N_44465,N_42568,N_42993);
and U44466 (N_44466,N_43229,N_42535);
and U44467 (N_44467,N_42468,N_42091);
or U44468 (N_44468,N_42103,N_43875);
nand U44469 (N_44469,N_43835,N_43265);
xnor U44470 (N_44470,N_43356,N_43570);
or U44471 (N_44471,N_42261,N_43953);
or U44472 (N_44472,N_43086,N_43574);
xor U44473 (N_44473,N_42190,N_43677);
xor U44474 (N_44474,N_43892,N_42008);
nand U44475 (N_44475,N_42983,N_42074);
nor U44476 (N_44476,N_42904,N_43016);
nor U44477 (N_44477,N_43125,N_43566);
xnor U44478 (N_44478,N_43646,N_43069);
nand U44479 (N_44479,N_43684,N_42617);
xnor U44480 (N_44480,N_42902,N_42742);
xor U44481 (N_44481,N_42118,N_42364);
or U44482 (N_44482,N_42929,N_43205);
and U44483 (N_44483,N_42974,N_43558);
nor U44484 (N_44484,N_43463,N_43666);
or U44485 (N_44485,N_42311,N_42240);
xor U44486 (N_44486,N_43691,N_43403);
nor U44487 (N_44487,N_42763,N_42678);
xor U44488 (N_44488,N_42173,N_43997);
nor U44489 (N_44489,N_43325,N_42076);
xor U44490 (N_44490,N_43713,N_43057);
nor U44491 (N_44491,N_42395,N_42489);
nor U44492 (N_44492,N_43848,N_43871);
nand U44493 (N_44493,N_43277,N_42402);
or U44494 (N_44494,N_43002,N_42733);
nor U44495 (N_44495,N_42414,N_42053);
or U44496 (N_44496,N_42558,N_43384);
nand U44497 (N_44497,N_42841,N_43749);
or U44498 (N_44498,N_42237,N_42797);
and U44499 (N_44499,N_42755,N_43306);
and U44500 (N_44500,N_43681,N_43019);
nand U44501 (N_44501,N_42705,N_42954);
and U44502 (N_44502,N_43222,N_43453);
xnor U44503 (N_44503,N_43577,N_43702);
or U44504 (N_44504,N_42809,N_42032);
or U44505 (N_44505,N_43424,N_43441);
nand U44506 (N_44506,N_43136,N_42342);
and U44507 (N_44507,N_43786,N_42391);
nor U44508 (N_44508,N_43225,N_42963);
nand U44509 (N_44509,N_43951,N_42221);
nor U44510 (N_44510,N_43588,N_43242);
or U44511 (N_44511,N_42256,N_42186);
and U44512 (N_44512,N_42647,N_42431);
and U44513 (N_44513,N_43029,N_42885);
nand U44514 (N_44514,N_43859,N_43281);
xor U44515 (N_44515,N_42549,N_42254);
nand U44516 (N_44516,N_43288,N_43500);
and U44517 (N_44517,N_42157,N_42867);
xor U44518 (N_44518,N_43938,N_42505);
nor U44519 (N_44519,N_42837,N_43949);
nand U44520 (N_44520,N_42426,N_43778);
nor U44521 (N_44521,N_43939,N_42353);
nor U44522 (N_44522,N_42958,N_43762);
nor U44523 (N_44523,N_42299,N_42058);
or U44524 (N_44524,N_42649,N_42056);
or U44525 (N_44525,N_42329,N_42286);
and U44526 (N_44526,N_43503,N_43665);
or U44527 (N_44527,N_42443,N_42613);
or U44528 (N_44528,N_43616,N_43630);
or U44529 (N_44529,N_43793,N_43518);
and U44530 (N_44530,N_42844,N_42943);
or U44531 (N_44531,N_42986,N_42175);
nand U44532 (N_44532,N_43755,N_42897);
xnor U44533 (N_44533,N_43756,N_43870);
nand U44534 (N_44534,N_43552,N_43105);
nand U44535 (N_44535,N_43091,N_42694);
nor U44536 (N_44536,N_42557,N_42176);
nand U44537 (N_44537,N_43511,N_42971);
and U44538 (N_44538,N_42140,N_42915);
nand U44539 (N_44539,N_42044,N_42903);
nor U44540 (N_44540,N_43011,N_42464);
or U44541 (N_44541,N_43992,N_43831);
or U44542 (N_44542,N_42612,N_43656);
or U44543 (N_44543,N_42289,N_42439);
nand U44544 (N_44544,N_43374,N_43680);
xnor U44545 (N_44545,N_42820,N_42787);
nor U44546 (N_44546,N_42033,N_42014);
nand U44547 (N_44547,N_43773,N_43669);
nor U44548 (N_44548,N_42834,N_43107);
xnor U44549 (N_44549,N_43640,N_43435);
nand U44550 (N_44550,N_42073,N_42846);
nor U44551 (N_44551,N_42434,N_43950);
nor U44552 (N_44552,N_42422,N_42813);
and U44553 (N_44553,N_43822,N_42734);
nand U44554 (N_44554,N_43323,N_43967);
nand U44555 (N_44555,N_43167,N_43559);
and U44556 (N_44556,N_42265,N_43720);
nor U44557 (N_44557,N_43137,N_43337);
and U44558 (N_44558,N_42015,N_43479);
or U44559 (N_44559,N_43979,N_43620);
and U44560 (N_44560,N_43119,N_42997);
or U44561 (N_44561,N_43537,N_43383);
and U44562 (N_44562,N_43077,N_42788);
nand U44563 (N_44563,N_42899,N_43780);
or U44564 (N_44564,N_42587,N_43546);
nand U44565 (N_44565,N_42239,N_42367);
and U44566 (N_44566,N_42436,N_43707);
nand U44567 (N_44567,N_43168,N_42982);
or U44568 (N_44568,N_43103,N_42840);
xnor U44569 (N_44569,N_42538,N_42021);
nor U44570 (N_44570,N_42398,N_43501);
xnor U44571 (N_44571,N_42243,N_42127);
nor U44572 (N_44572,N_43724,N_43847);
nand U44573 (N_44573,N_42799,N_42197);
nor U44574 (N_44574,N_43679,N_42675);
nand U44575 (N_44575,N_43159,N_43809);
or U44576 (N_44576,N_42623,N_42611);
or U44577 (N_44577,N_43569,N_43726);
or U44578 (N_44578,N_42306,N_43902);
xnor U44579 (N_44579,N_42832,N_43079);
or U44580 (N_44580,N_43839,N_43133);
and U44581 (N_44581,N_42401,N_43273);
nor U44582 (N_44582,N_43868,N_43431);
nand U44583 (N_44583,N_43063,N_43585);
or U44584 (N_44584,N_42459,N_43194);
nand U44585 (N_44585,N_42663,N_43528);
nor U44586 (N_44586,N_43657,N_42783);
xnor U44587 (N_44587,N_43776,N_42765);
or U44588 (N_44588,N_42296,N_43805);
or U44589 (N_44589,N_43746,N_42901);
nor U44590 (N_44590,N_42718,N_43587);
and U44591 (N_44591,N_43999,N_43985);
xnor U44592 (N_44592,N_43700,N_43033);
xnor U44593 (N_44593,N_42775,N_43021);
or U44594 (N_44594,N_43532,N_43451);
xnor U44595 (N_44595,N_43026,N_43409);
xor U44596 (N_44596,N_42034,N_42372);
or U44597 (N_44597,N_42596,N_43885);
xnor U44598 (N_44598,N_42894,N_42092);
and U44599 (N_44599,N_43605,N_43719);
or U44600 (N_44600,N_43987,N_43548);
nor U44601 (N_44601,N_43722,N_42412);
or U44602 (N_44602,N_42479,N_42644);
and U44603 (N_44603,N_42334,N_42757);
and U44604 (N_44604,N_43948,N_42491);
and U44605 (N_44605,N_43196,N_42279);
nand U44606 (N_44606,N_42744,N_43833);
and U44607 (N_44607,N_43246,N_43353);
nor U44608 (N_44608,N_43676,N_43637);
xnor U44609 (N_44609,N_42444,N_42916);
and U44610 (N_44610,N_42096,N_42521);
nand U44611 (N_44611,N_43301,N_42192);
nand U44612 (N_44612,N_42203,N_42283);
nor U44613 (N_44613,N_43343,N_42191);
nor U44614 (N_44614,N_42241,N_42732);
nand U44615 (N_44615,N_43887,N_42585);
and U44616 (N_44616,N_43652,N_43214);
nand U44617 (N_44617,N_42860,N_43432);
or U44618 (N_44618,N_42269,N_43413);
nand U44619 (N_44619,N_42523,N_43519);
nand U44620 (N_44620,N_42251,N_42149);
xor U44621 (N_44621,N_43898,N_43710);
nor U44622 (N_44622,N_42953,N_43729);
nor U44623 (N_44623,N_43098,N_42347);
or U44624 (N_44624,N_42448,N_43437);
or U44625 (N_44625,N_43642,N_43050);
nor U44626 (N_44626,N_43028,N_43644);
or U44627 (N_44627,N_42068,N_43255);
or U44628 (N_44628,N_43764,N_43791);
or U44629 (N_44629,N_42378,N_42650);
and U44630 (N_44630,N_42994,N_42553);
xor U44631 (N_44631,N_42394,N_42051);
xor U44632 (N_44632,N_43481,N_42771);
nand U44633 (N_44633,N_42031,N_42770);
xnor U44634 (N_44634,N_42007,N_43889);
xnor U44635 (N_44635,N_42121,N_43492);
nand U44636 (N_44636,N_42244,N_43653);
nor U44637 (N_44637,N_43373,N_42411);
or U44638 (N_44638,N_42938,N_42330);
or U44639 (N_44639,N_43627,N_43739);
or U44640 (N_44640,N_42136,N_43043);
nor U44641 (N_44641,N_42779,N_42515);
xnor U44642 (N_44642,N_43454,N_42964);
and U44643 (N_44643,N_42308,N_43709);
nor U44644 (N_44644,N_43975,N_43211);
or U44645 (N_44645,N_43825,N_43836);
or U44646 (N_44646,N_42572,N_43561);
nand U44647 (N_44647,N_43483,N_42657);
nand U44648 (N_44648,N_43708,N_42785);
or U44649 (N_44649,N_43765,N_43568);
and U44650 (N_44650,N_42879,N_42802);
or U44651 (N_44651,N_43796,N_42278);
and U44652 (N_44652,N_43024,N_43256);
or U44653 (N_44653,N_42934,N_43664);
or U44654 (N_44654,N_42972,N_42970);
nor U44655 (N_44655,N_42108,N_43816);
nor U44656 (N_44656,N_42936,N_42696);
nand U44657 (N_44657,N_43414,N_42499);
and U44658 (N_44658,N_43506,N_42036);
or U44659 (N_44659,N_43108,N_43264);
or U44660 (N_44660,N_42654,N_43121);
and U44661 (N_44661,N_42721,N_42466);
nand U44662 (N_44662,N_43427,N_43564);
nor U44663 (N_44663,N_42284,N_42736);
or U44664 (N_44664,N_43259,N_42161);
or U44665 (N_44665,N_43741,N_43138);
or U44666 (N_44666,N_42724,N_42409);
xor U44667 (N_44667,N_42776,N_43185);
or U44668 (N_44668,N_42354,N_43697);
nor U44669 (N_44669,N_43408,N_42598);
nand U44670 (N_44670,N_42951,N_42125);
nor U44671 (N_44671,N_43248,N_42680);
nor U44672 (N_44672,N_42282,N_43497);
and U44673 (N_44673,N_43296,N_43928);
nand U44674 (N_44674,N_43678,N_42691);
nand U44675 (N_44675,N_43283,N_42798);
nand U44676 (N_44676,N_43976,N_42335);
and U44677 (N_44677,N_43804,N_42417);
nor U44678 (N_44678,N_43467,N_43539);
nor U44679 (N_44679,N_43388,N_43770);
xor U44680 (N_44680,N_42104,N_43698);
nand U44681 (N_44681,N_42925,N_43813);
and U44682 (N_44682,N_42026,N_42300);
or U44683 (N_44683,N_43294,N_43386);
nor U44684 (N_44684,N_42041,N_42356);
nand U44685 (N_44685,N_42216,N_43580);
or U44686 (N_44686,N_43267,N_43230);
and U44687 (N_44687,N_42061,N_42518);
and U44688 (N_44688,N_43295,N_42035);
nor U44689 (N_44689,N_43271,N_43310);
and U44690 (N_44690,N_43080,N_43738);
nor U44691 (N_44691,N_43361,N_43404);
or U44692 (N_44692,N_43307,N_43457);
nand U44693 (N_44693,N_42920,N_43480);
or U44694 (N_44694,N_42001,N_43563);
and U44695 (N_44695,N_42510,N_42360);
nand U44696 (N_44696,N_43416,N_42552);
xnor U44697 (N_44697,N_43840,N_42923);
xnor U44698 (N_44698,N_43041,N_42653);
or U44699 (N_44699,N_42658,N_42119);
nor U44700 (N_44700,N_42165,N_42706);
nand U44701 (N_44701,N_42253,N_42821);
nand U44702 (N_44702,N_42124,N_43320);
or U44703 (N_44703,N_43104,N_43188);
or U44704 (N_44704,N_43866,N_42326);
xor U44705 (N_44705,N_43841,N_42807);
xnor U44706 (N_44706,N_43797,N_42445);
nor U44707 (N_44707,N_43912,N_42927);
xnor U44708 (N_44708,N_42786,N_43161);
nand U44709 (N_44709,N_43176,N_42493);
or U44710 (N_44710,N_43462,N_43247);
or U44711 (N_44711,N_42517,N_43685);
and U44712 (N_44712,N_42302,N_42248);
and U44713 (N_44713,N_43812,N_43659);
xnor U44714 (N_44714,N_43235,N_43406);
nand U44715 (N_44715,N_42497,N_42194);
nand U44716 (N_44716,N_42531,N_42390);
xor U44717 (N_44717,N_42377,N_43970);
nand U44718 (N_44718,N_43358,N_43591);
nand U44719 (N_44719,N_42453,N_43801);
nor U44720 (N_44720,N_43352,N_42599);
nor U44721 (N_44721,N_42942,N_43540);
xor U44722 (N_44722,N_42050,N_43827);
or U44723 (N_44723,N_43012,N_42926);
nor U44724 (N_44724,N_42796,N_42078);
xnor U44725 (N_44725,N_43172,N_43655);
nand U44726 (N_44726,N_43428,N_43735);
nand U44727 (N_44727,N_42548,N_43978);
and U44728 (N_44728,N_42527,N_42424);
nand U44729 (N_44729,N_42848,N_43111);
and U44730 (N_44730,N_42978,N_43129);
nand U44731 (N_44731,N_42627,N_43318);
nor U44732 (N_44732,N_43036,N_42703);
and U44733 (N_44733,N_42737,N_42002);
nor U44734 (N_44734,N_43212,N_43760);
or U44735 (N_44735,N_42564,N_42973);
nor U44736 (N_44736,N_43461,N_42047);
xor U44737 (N_44737,N_43191,N_43171);
or U44738 (N_44738,N_43370,N_43219);
nand U44739 (N_44739,N_43900,N_43556);
xnor U44740 (N_44740,N_42998,N_43943);
nor U44741 (N_44741,N_42532,N_42615);
nand U44742 (N_44742,N_43712,N_42463);
xor U44743 (N_44743,N_43959,N_43195);
nand U44744 (N_44744,N_43331,N_42473);
and U44745 (N_44745,N_42550,N_42293);
nand U44746 (N_44746,N_43199,N_42522);
and U44747 (N_44747,N_42725,N_42569);
or U44748 (N_44748,N_42432,N_43488);
nand U44749 (N_44749,N_43761,N_43154);
nand U44750 (N_44750,N_42132,N_43078);
and U44751 (N_44751,N_43759,N_43823);
nand U44752 (N_44752,N_42413,N_42710);
xnor U44753 (N_44753,N_42534,N_42825);
nor U44754 (N_44754,N_42333,N_42645);
or U44755 (N_44755,N_43706,N_42155);
nor U44756 (N_44756,N_43008,N_42651);
nand U44757 (N_44757,N_43915,N_42331);
nand U44758 (N_44758,N_43648,N_43253);
xnor U44759 (N_44759,N_43251,N_42156);
xnor U44760 (N_44760,N_42446,N_42152);
nor U44761 (N_44761,N_43330,N_42917);
nand U44762 (N_44762,N_42975,N_43302);
xor U44763 (N_44763,N_43662,N_43298);
nor U44764 (N_44764,N_43923,N_43990);
and U44765 (N_44765,N_43830,N_42573);
xor U44766 (N_44766,N_43986,N_42593);
xnor U44767 (N_44767,N_43769,N_43475);
and U44768 (N_44768,N_43144,N_42374);
nand U44769 (N_44769,N_43197,N_43270);
xnor U44770 (N_44770,N_42811,N_42343);
xor U44771 (N_44771,N_42625,N_43683);
nand U44772 (N_44772,N_43216,N_43065);
nand U44773 (N_44773,N_42425,N_42543);
or U44774 (N_44774,N_42154,N_42702);
or U44775 (N_44775,N_43489,N_42672);
and U44776 (N_44776,N_42632,N_43166);
or U44777 (N_44777,N_42064,N_43633);
xor U44778 (N_44778,N_43052,N_43327);
xnor U44779 (N_44779,N_42072,N_42891);
or U44780 (N_44780,N_42849,N_43844);
and U44781 (N_44781,N_43203,N_42815);
and U44782 (N_44782,N_42812,N_42423);
xor U44783 (N_44783,N_43808,N_43508);
nor U44784 (N_44784,N_43886,N_42297);
or U44785 (N_44785,N_43879,N_42712);
and U44786 (N_44786,N_42666,N_42633);
nand U44787 (N_44787,N_42222,N_43850);
and U44788 (N_44788,N_42407,N_42116);
nand U44789 (N_44789,N_43156,N_42634);
and U44790 (N_44790,N_42853,N_42430);
nor U44791 (N_44791,N_42877,N_42018);
xor U44792 (N_44792,N_43792,N_42348);
nor U44793 (N_44793,N_42016,N_42315);
nor U44794 (N_44794,N_42452,N_42214);
nor U44795 (N_44795,N_42681,N_42267);
and U44796 (N_44796,N_42114,N_42144);
xor U44797 (N_44797,N_43649,N_42322);
and U44798 (N_44798,N_43621,N_42913);
xor U44799 (N_44799,N_42150,N_43874);
and U44800 (N_44800,N_43037,N_43226);
xor U44801 (N_44801,N_43747,N_43799);
nor U44802 (N_44802,N_42454,N_42492);
nand U44803 (N_44803,N_43258,N_43821);
and U44804 (N_44804,N_43357,N_43775);
nand U44805 (N_44805,N_43890,N_43148);
nand U44806 (N_44806,N_43579,N_43183);
and U44807 (N_44807,N_43650,N_43785);
or U44808 (N_44808,N_42418,N_43907);
or U44809 (N_44809,N_42693,N_42313);
nand U44810 (N_44810,N_42912,N_43278);
and U44811 (N_44811,N_42379,N_42359);
or U44812 (N_44812,N_42490,N_42690);
xnor U44813 (N_44813,N_43751,N_42094);
nand U44814 (N_44814,N_42246,N_42588);
nand U44815 (N_44815,N_43860,N_43541);
or U44816 (N_44816,N_43047,N_43400);
nor U44817 (N_44817,N_42778,N_43682);
or U44818 (N_44818,N_43152,N_43328);
nor U44819 (N_44819,N_43170,N_43916);
xor U44820 (N_44820,N_43618,N_42081);
and U44821 (N_44821,N_43198,N_42610);
xor U44822 (N_44822,N_43097,N_42172);
nand U44823 (N_44823,N_43186,N_43845);
nand U44824 (N_44824,N_42890,N_43459);
nor U44825 (N_44825,N_42352,N_42122);
or U44826 (N_44826,N_43285,N_42560);
or U44827 (N_44827,N_42110,N_42999);
xnor U44828 (N_44828,N_43829,N_43937);
xor U44829 (N_44829,N_43127,N_42817);
xnor U44830 (N_44830,N_43334,N_43261);
nand U44831 (N_44831,N_42544,N_43894);
or U44832 (N_44832,N_43465,N_42164);
xnor U44833 (N_44833,N_42921,N_43607);
nand U44834 (N_44834,N_42833,N_43802);
nand U44835 (N_44835,N_42408,N_42945);
or U44836 (N_44836,N_43187,N_42085);
nor U44837 (N_44837,N_43316,N_43704);
or U44838 (N_44838,N_42946,N_42637);
nor U44839 (N_44839,N_43661,N_43317);
and U44840 (N_44840,N_43933,N_43929);
and U44841 (N_44841,N_43075,N_42563);
or U44842 (N_44842,N_42831,N_42000);
or U44843 (N_44843,N_43355,N_42158);
xnor U44844 (N_44844,N_42485,N_42969);
and U44845 (N_44845,N_42556,N_42767);
and U44846 (N_44846,N_43365,N_43303);
or U44847 (N_44847,N_43366,N_43795);
xnor U44848 (N_44848,N_43499,N_43947);
and U44849 (N_44849,N_43297,N_42055);
and U44850 (N_44850,N_43843,N_42160);
or U44851 (N_44851,N_42562,N_42823);
and U44852 (N_44852,N_42178,N_43737);
nand U44853 (N_44853,N_42181,N_42766);
xor U44854 (N_44854,N_42472,N_43602);
nor U44855 (N_44855,N_43192,N_43576);
xor U44856 (N_44856,N_43132,N_43308);
or U44857 (N_44857,N_42295,N_43102);
nand U44858 (N_44858,N_43824,N_43023);
nor U44859 (N_44859,N_42985,N_43407);
and U44860 (N_44860,N_42208,N_42328);
nand U44861 (N_44861,N_42907,N_42609);
xnor U44862 (N_44862,N_43287,N_43354);
and U44863 (N_44863,N_43151,N_42276);
or U44864 (N_44864,N_43567,N_43596);
xor U44865 (N_44865,N_43904,N_42695);
nand U44866 (N_44866,N_43730,N_43493);
or U44867 (N_44867,N_43964,N_43391);
xnor U44868 (N_44868,N_43876,N_43789);
xnor U44869 (N_44869,N_42758,N_43007);
or U44870 (N_44870,N_42042,N_42271);
and U44871 (N_44871,N_43969,N_43529);
xnor U44872 (N_44872,N_42447,N_43449);
nand U44873 (N_44873,N_43696,N_43234);
nand U44874 (N_44874,N_43592,N_42806);
xnor U44875 (N_44875,N_43430,N_43145);
and U44876 (N_44876,N_43022,N_43895);
nand U44877 (N_44877,N_43232,N_42528);
or U44878 (N_44878,N_43645,N_43066);
xnor U44879 (N_44879,N_43380,N_42039);
nor U44880 (N_44880,N_42385,N_43903);
nor U44881 (N_44881,N_42373,N_42003);
and U44882 (N_44882,N_43445,N_42745);
nor U44883 (N_44883,N_43758,N_42312);
or U44884 (N_44884,N_43858,N_42782);
and U44885 (N_44885,N_43982,N_42465);
or U44886 (N_44886,N_42516,N_42198);
nor U44887 (N_44887,N_42597,N_42838);
and U44888 (N_44888,N_42218,N_43955);
or U44889 (N_44889,N_42746,N_43333);
or U44890 (N_44890,N_42461,N_43734);
and U44891 (N_44891,N_43074,N_43593);
or U44892 (N_44892,N_42743,N_42168);
and U44893 (N_44893,N_42870,N_42575);
xnor U44894 (N_44894,N_43502,N_42567);
or U44895 (N_44895,N_43911,N_43639);
nor U44896 (N_44896,N_42487,N_42065);
nor U44897 (N_44897,N_42803,N_42707);
or U44898 (N_44898,N_42361,N_42079);
and U44899 (N_44899,N_42314,N_43433);
and U44900 (N_44900,N_43173,N_42405);
xor U44901 (N_44901,N_42720,N_43393);
or U44902 (N_44902,N_43983,N_42368);
nand U44903 (N_44903,N_43555,N_42052);
xnor U44904 (N_44904,N_43184,N_42595);
nor U44905 (N_44905,N_42868,N_43060);
nand U44906 (N_44906,N_43299,N_43861);
and U44907 (N_44907,N_43486,N_43477);
nor U44908 (N_44908,N_42483,N_43731);
and U44909 (N_44909,N_42363,N_42750);
nand U44910 (N_44910,N_43973,N_42135);
nand U44911 (N_44911,N_43390,N_43114);
xnor U44912 (N_44912,N_43286,N_42561);
nand U44913 (N_44913,N_43174,N_43010);
xor U44914 (N_44914,N_42930,N_42655);
or U44915 (N_44915,N_42380,N_43243);
nor U44916 (N_44916,N_43856,N_42949);
nor U44917 (N_44917,N_42980,N_43954);
nor U44918 (N_44918,N_43141,N_43134);
nand U44919 (N_44919,N_42226,N_43632);
or U44920 (N_44920,N_42388,N_42950);
nor U44921 (N_44921,N_43068,N_42301);
xor U44922 (N_44922,N_43153,N_42435);
nor U44923 (N_44923,N_42905,N_42514);
or U44924 (N_44924,N_43660,N_43181);
and U44925 (N_44925,N_42498,N_43818);
xnor U44926 (N_44926,N_43614,N_42098);
nand U44927 (N_44927,N_42570,N_43351);
or U44928 (N_44928,N_42540,N_42231);
nor U44929 (N_44929,N_42699,N_42207);
xor U44930 (N_44930,N_42262,N_42685);
and U44931 (N_44931,N_43315,N_42211);
nand U44932 (N_44932,N_42387,N_42869);
and U44933 (N_44933,N_43507,N_42400);
nand U44934 (N_44934,N_42566,N_43864);
or U44935 (N_44935,N_42084,N_42668);
xnor U44936 (N_44936,N_43763,N_43375);
nor U44937 (N_44937,N_43941,N_42661);
and U44938 (N_44938,N_42397,N_42496);
nand U44939 (N_44939,N_43921,N_42111);
nor U44940 (N_44940,N_43599,N_43971);
xnor U44941 (N_44941,N_43834,N_42677);
nand U44942 (N_44942,N_43118,N_42235);
and U44943 (N_44943,N_42648,N_43425);
or U44944 (N_44944,N_42888,N_43473);
nand U44945 (N_44945,N_43359,N_43070);
nor U44946 (N_44946,N_42861,N_42177);
and U44947 (N_44947,N_42346,N_43832);
or U44948 (N_44948,N_42620,N_42457);
and U44949 (N_44949,N_43515,N_42238);
or U44950 (N_44950,N_42684,N_43115);
and U44951 (N_44951,N_42526,N_42227);
nand U44952 (N_44952,N_43732,N_43304);
nand U44953 (N_44953,N_43658,N_42169);
or U44954 (N_44954,N_43006,N_43628);
and U44955 (N_44955,N_43842,N_43000);
nand U44956 (N_44956,N_42759,N_42641);
xor U44957 (N_44957,N_43940,N_43863);
nand U44958 (N_44958,N_42659,N_42881);
nor U44959 (N_44959,N_43757,N_43263);
and U44960 (N_44960,N_42507,N_43444);
nand U44961 (N_44961,N_42576,N_42873);
or U44962 (N_44962,N_42875,N_43249);
nand U44963 (N_44963,N_43623,N_43420);
nor U44964 (N_44964,N_42474,N_42206);
and U44965 (N_44965,N_43798,N_43031);
or U44966 (N_44966,N_43339,N_43217);
nor U44967 (N_44967,N_42735,N_42180);
nor U44968 (N_44968,N_43855,N_42059);
nand U44969 (N_44969,N_42428,N_42371);
and U44970 (N_44970,N_42476,N_42652);
or U44971 (N_44971,N_42129,N_42773);
nor U44972 (N_44972,N_43456,N_42349);
nand U44973 (N_44973,N_43157,N_42624);
xor U44974 (N_44974,N_42145,N_43061);
and U44975 (N_44975,N_43624,N_42589);
xnor U44976 (N_44976,N_42049,N_42280);
or U44977 (N_44977,N_43865,N_43405);
xor U44978 (N_44978,N_43046,N_43321);
and U44979 (N_44979,N_43629,N_42924);
nor U44980 (N_44980,N_42332,N_43631);
or U44981 (N_44981,N_43617,N_43945);
or U44982 (N_44982,N_42449,N_42298);
and U44983 (N_44983,N_43784,N_43787);
nand U44984 (N_44984,N_42607,N_43452);
xnor U44985 (N_44985,N_42740,N_43504);
xor U44986 (N_44986,N_43750,N_43671);
nand U44987 (N_44987,N_42341,N_42580);
nand U44988 (N_44988,N_42965,N_42010);
xnor U44989 (N_44989,N_42469,N_43622);
and U44990 (N_44990,N_43553,N_42006);
and U44991 (N_44991,N_43589,N_43854);
nand U44992 (N_44992,N_42143,N_42303);
nor U44993 (N_44993,N_43725,N_42247);
xnor U44994 (N_44994,N_42382,N_43647);
or U44995 (N_44995,N_43130,N_42674);
nor U44996 (N_44996,N_42028,N_43906);
or U44997 (N_44997,N_43027,N_42202);
and U44998 (N_44998,N_43914,N_42664);
nor U44999 (N_44999,N_42880,N_43535);
and U45000 (N_45000,N_42210,N_42190);
nand U45001 (N_45001,N_42754,N_42908);
nor U45002 (N_45002,N_43617,N_42173);
or U45003 (N_45003,N_42081,N_43976);
or U45004 (N_45004,N_42506,N_42357);
nor U45005 (N_45005,N_42274,N_43530);
and U45006 (N_45006,N_43743,N_43127);
nor U45007 (N_45007,N_42165,N_43839);
xnor U45008 (N_45008,N_42655,N_43049);
and U45009 (N_45009,N_42408,N_42190);
nor U45010 (N_45010,N_42708,N_42900);
or U45011 (N_45011,N_42269,N_42113);
nor U45012 (N_45012,N_42576,N_42864);
and U45013 (N_45013,N_43442,N_42269);
and U45014 (N_45014,N_43181,N_42722);
nand U45015 (N_45015,N_42098,N_42863);
or U45016 (N_45016,N_42474,N_42083);
nand U45017 (N_45017,N_42461,N_42262);
nand U45018 (N_45018,N_42750,N_42758);
or U45019 (N_45019,N_43499,N_43760);
xor U45020 (N_45020,N_42960,N_42201);
nand U45021 (N_45021,N_43558,N_42724);
and U45022 (N_45022,N_42054,N_43323);
nand U45023 (N_45023,N_43290,N_43585);
or U45024 (N_45024,N_42252,N_43000);
or U45025 (N_45025,N_43950,N_42166);
xor U45026 (N_45026,N_43893,N_42415);
and U45027 (N_45027,N_43603,N_43118);
nor U45028 (N_45028,N_43618,N_42961);
and U45029 (N_45029,N_42994,N_43674);
nor U45030 (N_45030,N_43452,N_42758);
nor U45031 (N_45031,N_43691,N_43445);
nor U45032 (N_45032,N_43571,N_43327);
or U45033 (N_45033,N_42869,N_43176);
nor U45034 (N_45034,N_43632,N_43039);
and U45035 (N_45035,N_42350,N_43441);
or U45036 (N_45036,N_43080,N_42518);
nand U45037 (N_45037,N_42410,N_43006);
or U45038 (N_45038,N_43750,N_42613);
nor U45039 (N_45039,N_43192,N_43320);
and U45040 (N_45040,N_43702,N_43443);
nand U45041 (N_45041,N_42613,N_42549);
xor U45042 (N_45042,N_42501,N_42094);
xor U45043 (N_45043,N_42266,N_43415);
nand U45044 (N_45044,N_42852,N_42744);
nand U45045 (N_45045,N_43540,N_42364);
nor U45046 (N_45046,N_43008,N_43748);
nor U45047 (N_45047,N_43509,N_42902);
or U45048 (N_45048,N_43846,N_43851);
nand U45049 (N_45049,N_42021,N_43425);
or U45050 (N_45050,N_43013,N_42697);
nand U45051 (N_45051,N_42122,N_43885);
and U45052 (N_45052,N_43227,N_43075);
nor U45053 (N_45053,N_42401,N_42483);
nand U45054 (N_45054,N_43823,N_43077);
or U45055 (N_45055,N_43552,N_43907);
nor U45056 (N_45056,N_42969,N_42886);
nand U45057 (N_45057,N_42049,N_43282);
or U45058 (N_45058,N_42929,N_42739);
or U45059 (N_45059,N_43239,N_42922);
nand U45060 (N_45060,N_42017,N_43757);
xor U45061 (N_45061,N_43170,N_43104);
nand U45062 (N_45062,N_43483,N_42770);
and U45063 (N_45063,N_42719,N_43285);
xor U45064 (N_45064,N_43277,N_43616);
xnor U45065 (N_45065,N_42213,N_43651);
xor U45066 (N_45066,N_42647,N_43896);
or U45067 (N_45067,N_43146,N_42135);
nor U45068 (N_45068,N_42639,N_43146);
or U45069 (N_45069,N_42958,N_42599);
nand U45070 (N_45070,N_43346,N_43097);
nand U45071 (N_45071,N_43364,N_42930);
xnor U45072 (N_45072,N_43376,N_42973);
nor U45073 (N_45073,N_42866,N_43086);
nand U45074 (N_45074,N_42843,N_42734);
and U45075 (N_45075,N_42083,N_43366);
or U45076 (N_45076,N_42632,N_42832);
or U45077 (N_45077,N_43777,N_42564);
or U45078 (N_45078,N_42670,N_43489);
xnor U45079 (N_45079,N_42420,N_42398);
or U45080 (N_45080,N_42560,N_43694);
nor U45081 (N_45081,N_42831,N_43164);
or U45082 (N_45082,N_42256,N_43473);
or U45083 (N_45083,N_42792,N_42111);
nor U45084 (N_45084,N_43739,N_42439);
nand U45085 (N_45085,N_43574,N_43351);
nor U45086 (N_45086,N_42384,N_42429);
nand U45087 (N_45087,N_43958,N_42910);
xor U45088 (N_45088,N_42975,N_42230);
nor U45089 (N_45089,N_42638,N_43862);
xor U45090 (N_45090,N_42675,N_43736);
and U45091 (N_45091,N_42608,N_42196);
or U45092 (N_45092,N_43624,N_43961);
and U45093 (N_45093,N_42929,N_42188);
xnor U45094 (N_45094,N_42243,N_43729);
nand U45095 (N_45095,N_43072,N_43525);
nor U45096 (N_45096,N_43970,N_43566);
and U45097 (N_45097,N_42963,N_43243);
nand U45098 (N_45098,N_42471,N_43383);
nand U45099 (N_45099,N_43795,N_42792);
nand U45100 (N_45100,N_42895,N_43025);
nand U45101 (N_45101,N_43722,N_42000);
nand U45102 (N_45102,N_43537,N_42970);
nor U45103 (N_45103,N_43414,N_42990);
or U45104 (N_45104,N_43419,N_43254);
nand U45105 (N_45105,N_43407,N_43566);
or U45106 (N_45106,N_43088,N_43936);
nor U45107 (N_45107,N_42218,N_43566);
and U45108 (N_45108,N_42027,N_43446);
xor U45109 (N_45109,N_43559,N_43921);
or U45110 (N_45110,N_42995,N_42189);
xor U45111 (N_45111,N_42458,N_43074);
nand U45112 (N_45112,N_43264,N_43502);
nand U45113 (N_45113,N_43722,N_42915);
nor U45114 (N_45114,N_43839,N_43769);
nand U45115 (N_45115,N_42919,N_43660);
xnor U45116 (N_45116,N_43231,N_42696);
or U45117 (N_45117,N_43087,N_43419);
xnor U45118 (N_45118,N_42912,N_43977);
nand U45119 (N_45119,N_42598,N_43668);
nor U45120 (N_45120,N_43245,N_43476);
xor U45121 (N_45121,N_43653,N_43252);
and U45122 (N_45122,N_43403,N_43314);
xor U45123 (N_45123,N_42992,N_42865);
or U45124 (N_45124,N_42979,N_42881);
nand U45125 (N_45125,N_42577,N_43631);
or U45126 (N_45126,N_42751,N_43758);
nor U45127 (N_45127,N_43538,N_43559);
or U45128 (N_45128,N_43984,N_43050);
and U45129 (N_45129,N_43594,N_42390);
nand U45130 (N_45130,N_43300,N_42897);
and U45131 (N_45131,N_43219,N_43116);
and U45132 (N_45132,N_43888,N_43393);
nor U45133 (N_45133,N_43199,N_42449);
and U45134 (N_45134,N_42254,N_43754);
xnor U45135 (N_45135,N_42570,N_43209);
nand U45136 (N_45136,N_43391,N_42018);
and U45137 (N_45137,N_42494,N_42534);
and U45138 (N_45138,N_42030,N_43781);
nor U45139 (N_45139,N_43135,N_42122);
nand U45140 (N_45140,N_43389,N_43851);
or U45141 (N_45141,N_43811,N_42526);
nor U45142 (N_45142,N_42137,N_43465);
xor U45143 (N_45143,N_42950,N_42288);
nor U45144 (N_45144,N_43051,N_42836);
xnor U45145 (N_45145,N_42085,N_42173);
xnor U45146 (N_45146,N_42908,N_42827);
and U45147 (N_45147,N_42501,N_42500);
nand U45148 (N_45148,N_42893,N_43409);
or U45149 (N_45149,N_43668,N_43485);
nor U45150 (N_45150,N_42034,N_43151);
nand U45151 (N_45151,N_43471,N_43447);
xor U45152 (N_45152,N_43894,N_43719);
and U45153 (N_45153,N_42587,N_42812);
and U45154 (N_45154,N_42154,N_43555);
nand U45155 (N_45155,N_42340,N_42966);
nor U45156 (N_45156,N_43499,N_43548);
and U45157 (N_45157,N_42417,N_42350);
xnor U45158 (N_45158,N_43727,N_42560);
nand U45159 (N_45159,N_42104,N_43411);
nor U45160 (N_45160,N_42954,N_43792);
and U45161 (N_45161,N_43757,N_43180);
nand U45162 (N_45162,N_43172,N_43953);
nor U45163 (N_45163,N_42962,N_43520);
or U45164 (N_45164,N_43958,N_43266);
or U45165 (N_45165,N_43282,N_42523);
or U45166 (N_45166,N_43093,N_42419);
nor U45167 (N_45167,N_43313,N_43662);
or U45168 (N_45168,N_42340,N_42382);
nand U45169 (N_45169,N_43715,N_43765);
xor U45170 (N_45170,N_43090,N_42035);
xnor U45171 (N_45171,N_43970,N_43588);
and U45172 (N_45172,N_43308,N_42909);
nor U45173 (N_45173,N_43398,N_43282);
nor U45174 (N_45174,N_42055,N_42540);
nand U45175 (N_45175,N_42696,N_42028);
nor U45176 (N_45176,N_42331,N_43718);
and U45177 (N_45177,N_42152,N_43353);
nand U45178 (N_45178,N_42561,N_42602);
and U45179 (N_45179,N_42825,N_43770);
nand U45180 (N_45180,N_43410,N_43901);
xor U45181 (N_45181,N_42522,N_43987);
xor U45182 (N_45182,N_42842,N_42172);
nand U45183 (N_45183,N_42498,N_42172);
and U45184 (N_45184,N_43233,N_42787);
and U45185 (N_45185,N_42833,N_43173);
or U45186 (N_45186,N_43406,N_43307);
nor U45187 (N_45187,N_43145,N_42606);
xnor U45188 (N_45188,N_43920,N_43417);
nand U45189 (N_45189,N_43028,N_43203);
nand U45190 (N_45190,N_42124,N_43578);
nor U45191 (N_45191,N_42370,N_42125);
nor U45192 (N_45192,N_42037,N_43697);
xor U45193 (N_45193,N_43248,N_42809);
xnor U45194 (N_45194,N_42552,N_43972);
nor U45195 (N_45195,N_42665,N_42438);
nand U45196 (N_45196,N_43348,N_42811);
nor U45197 (N_45197,N_43362,N_43931);
xnor U45198 (N_45198,N_42483,N_43907);
nor U45199 (N_45199,N_43727,N_43154);
and U45200 (N_45200,N_43155,N_43544);
xor U45201 (N_45201,N_43985,N_42480);
or U45202 (N_45202,N_43339,N_43777);
or U45203 (N_45203,N_43545,N_43286);
nand U45204 (N_45204,N_43606,N_43598);
or U45205 (N_45205,N_43232,N_43550);
or U45206 (N_45206,N_43385,N_42255);
nand U45207 (N_45207,N_43287,N_42621);
nand U45208 (N_45208,N_42160,N_43537);
or U45209 (N_45209,N_43304,N_42225);
xor U45210 (N_45210,N_43518,N_43116);
xnor U45211 (N_45211,N_42785,N_42059);
nor U45212 (N_45212,N_43081,N_42156);
and U45213 (N_45213,N_43158,N_42406);
and U45214 (N_45214,N_42521,N_43995);
and U45215 (N_45215,N_42678,N_42101);
nand U45216 (N_45216,N_43306,N_43763);
or U45217 (N_45217,N_42044,N_43662);
nor U45218 (N_45218,N_42014,N_43911);
nand U45219 (N_45219,N_43056,N_42713);
nor U45220 (N_45220,N_43213,N_43584);
xnor U45221 (N_45221,N_42896,N_42488);
nor U45222 (N_45222,N_43631,N_43503);
and U45223 (N_45223,N_42125,N_42208);
or U45224 (N_45224,N_42921,N_43599);
nand U45225 (N_45225,N_43085,N_42875);
xor U45226 (N_45226,N_43192,N_43480);
and U45227 (N_45227,N_42763,N_42101);
nand U45228 (N_45228,N_43750,N_43954);
or U45229 (N_45229,N_43856,N_42522);
xor U45230 (N_45230,N_42439,N_42050);
nand U45231 (N_45231,N_42799,N_42552);
nor U45232 (N_45232,N_43981,N_42603);
nand U45233 (N_45233,N_42186,N_42894);
nor U45234 (N_45234,N_43410,N_43623);
nor U45235 (N_45235,N_43903,N_42309);
and U45236 (N_45236,N_43498,N_42753);
or U45237 (N_45237,N_42981,N_42170);
and U45238 (N_45238,N_42772,N_42228);
nand U45239 (N_45239,N_43762,N_43770);
and U45240 (N_45240,N_42192,N_43386);
xor U45241 (N_45241,N_43453,N_43090);
or U45242 (N_45242,N_42781,N_42993);
or U45243 (N_45243,N_42959,N_43688);
nand U45244 (N_45244,N_43607,N_42675);
and U45245 (N_45245,N_43714,N_43007);
nor U45246 (N_45246,N_43428,N_43920);
nor U45247 (N_45247,N_43022,N_42708);
nand U45248 (N_45248,N_42847,N_42652);
nor U45249 (N_45249,N_42646,N_42002);
nand U45250 (N_45250,N_43247,N_42853);
xnor U45251 (N_45251,N_43662,N_42160);
nand U45252 (N_45252,N_42889,N_43089);
xor U45253 (N_45253,N_42490,N_43890);
xnor U45254 (N_45254,N_42758,N_42039);
nor U45255 (N_45255,N_42363,N_42038);
xor U45256 (N_45256,N_43630,N_43754);
nor U45257 (N_45257,N_43181,N_43155);
nand U45258 (N_45258,N_42996,N_43632);
or U45259 (N_45259,N_43273,N_43243);
and U45260 (N_45260,N_42120,N_42184);
xor U45261 (N_45261,N_43372,N_43475);
or U45262 (N_45262,N_43255,N_43132);
and U45263 (N_45263,N_43824,N_42999);
xor U45264 (N_45264,N_43851,N_42126);
or U45265 (N_45265,N_43547,N_42229);
and U45266 (N_45266,N_42522,N_42578);
xnor U45267 (N_45267,N_43847,N_42246);
or U45268 (N_45268,N_42331,N_43283);
xor U45269 (N_45269,N_43448,N_43355);
and U45270 (N_45270,N_42216,N_42686);
and U45271 (N_45271,N_43098,N_43997);
nand U45272 (N_45272,N_42173,N_43446);
and U45273 (N_45273,N_42829,N_42818);
and U45274 (N_45274,N_43574,N_42352);
nand U45275 (N_45275,N_43912,N_43313);
nor U45276 (N_45276,N_43366,N_43425);
and U45277 (N_45277,N_42935,N_43367);
and U45278 (N_45278,N_42840,N_43836);
xor U45279 (N_45279,N_43111,N_42329);
nand U45280 (N_45280,N_42466,N_42281);
or U45281 (N_45281,N_42543,N_43409);
xor U45282 (N_45282,N_42903,N_43876);
nand U45283 (N_45283,N_43866,N_43809);
nor U45284 (N_45284,N_42903,N_42323);
and U45285 (N_45285,N_43235,N_42436);
xor U45286 (N_45286,N_43673,N_42969);
xnor U45287 (N_45287,N_43209,N_43406);
or U45288 (N_45288,N_42539,N_42024);
nand U45289 (N_45289,N_43650,N_42429);
or U45290 (N_45290,N_42618,N_42704);
nand U45291 (N_45291,N_43618,N_43418);
and U45292 (N_45292,N_43560,N_42123);
and U45293 (N_45293,N_43751,N_43117);
nor U45294 (N_45294,N_42119,N_42762);
nor U45295 (N_45295,N_43628,N_42504);
and U45296 (N_45296,N_42070,N_43239);
nand U45297 (N_45297,N_43654,N_43671);
or U45298 (N_45298,N_43333,N_42204);
nor U45299 (N_45299,N_42145,N_42692);
and U45300 (N_45300,N_42072,N_43576);
or U45301 (N_45301,N_42663,N_42333);
or U45302 (N_45302,N_42051,N_43250);
xor U45303 (N_45303,N_42009,N_42793);
or U45304 (N_45304,N_42527,N_43916);
xnor U45305 (N_45305,N_43109,N_42260);
and U45306 (N_45306,N_42567,N_43478);
nand U45307 (N_45307,N_42026,N_43409);
xnor U45308 (N_45308,N_42345,N_42934);
or U45309 (N_45309,N_43688,N_43500);
xor U45310 (N_45310,N_43070,N_42047);
nand U45311 (N_45311,N_43265,N_42674);
and U45312 (N_45312,N_42181,N_43194);
nand U45313 (N_45313,N_42227,N_43855);
nor U45314 (N_45314,N_43049,N_42585);
nand U45315 (N_45315,N_42330,N_42967);
nor U45316 (N_45316,N_43661,N_42532);
nand U45317 (N_45317,N_43035,N_43858);
nand U45318 (N_45318,N_42206,N_42305);
xor U45319 (N_45319,N_42429,N_43795);
nor U45320 (N_45320,N_42899,N_43797);
or U45321 (N_45321,N_43263,N_42707);
nand U45322 (N_45322,N_42977,N_42514);
and U45323 (N_45323,N_42123,N_42734);
nand U45324 (N_45324,N_43746,N_43925);
and U45325 (N_45325,N_42779,N_43440);
and U45326 (N_45326,N_43782,N_43800);
xor U45327 (N_45327,N_43648,N_42922);
or U45328 (N_45328,N_43472,N_43277);
nor U45329 (N_45329,N_43177,N_42094);
or U45330 (N_45330,N_42473,N_43799);
nand U45331 (N_45331,N_42546,N_42628);
or U45332 (N_45332,N_43724,N_43999);
nor U45333 (N_45333,N_43343,N_43036);
nand U45334 (N_45334,N_43111,N_42204);
nor U45335 (N_45335,N_43408,N_43264);
or U45336 (N_45336,N_42492,N_43611);
xnor U45337 (N_45337,N_42710,N_42988);
nand U45338 (N_45338,N_43163,N_42054);
or U45339 (N_45339,N_43888,N_42717);
and U45340 (N_45340,N_43188,N_42338);
nand U45341 (N_45341,N_43205,N_42674);
xnor U45342 (N_45342,N_43615,N_43321);
xnor U45343 (N_45343,N_43722,N_43294);
nor U45344 (N_45344,N_43428,N_43349);
or U45345 (N_45345,N_43709,N_43759);
and U45346 (N_45346,N_43981,N_42719);
or U45347 (N_45347,N_42630,N_42790);
and U45348 (N_45348,N_43356,N_42456);
nor U45349 (N_45349,N_42422,N_42571);
or U45350 (N_45350,N_43293,N_43639);
nand U45351 (N_45351,N_42480,N_42283);
xnor U45352 (N_45352,N_43779,N_43719);
nand U45353 (N_45353,N_43764,N_42304);
or U45354 (N_45354,N_42479,N_42170);
nand U45355 (N_45355,N_43606,N_43447);
or U45356 (N_45356,N_42716,N_43641);
or U45357 (N_45357,N_42951,N_42890);
and U45358 (N_45358,N_42628,N_42853);
or U45359 (N_45359,N_42627,N_42575);
or U45360 (N_45360,N_42378,N_42481);
or U45361 (N_45361,N_43224,N_42931);
nor U45362 (N_45362,N_43316,N_43218);
or U45363 (N_45363,N_43141,N_43241);
and U45364 (N_45364,N_42638,N_42222);
and U45365 (N_45365,N_42628,N_43984);
nor U45366 (N_45366,N_42363,N_43866);
or U45367 (N_45367,N_42723,N_42058);
nand U45368 (N_45368,N_43803,N_42443);
xor U45369 (N_45369,N_43634,N_42008);
and U45370 (N_45370,N_42667,N_43521);
and U45371 (N_45371,N_42864,N_42616);
nor U45372 (N_45372,N_43108,N_43360);
and U45373 (N_45373,N_43642,N_43140);
nor U45374 (N_45374,N_43229,N_42669);
nand U45375 (N_45375,N_43529,N_42103);
nor U45376 (N_45376,N_43417,N_43955);
and U45377 (N_45377,N_42813,N_43660);
xnor U45378 (N_45378,N_42771,N_43336);
xor U45379 (N_45379,N_42646,N_42966);
and U45380 (N_45380,N_43661,N_42923);
nor U45381 (N_45381,N_42032,N_42292);
xor U45382 (N_45382,N_42731,N_43012);
and U45383 (N_45383,N_43971,N_43598);
or U45384 (N_45384,N_42242,N_42004);
nor U45385 (N_45385,N_43603,N_42457);
nor U45386 (N_45386,N_43051,N_42130);
nand U45387 (N_45387,N_42075,N_43839);
and U45388 (N_45388,N_42984,N_43104);
xor U45389 (N_45389,N_43194,N_42532);
or U45390 (N_45390,N_42779,N_43545);
xnor U45391 (N_45391,N_42305,N_42817);
nand U45392 (N_45392,N_42674,N_42696);
nor U45393 (N_45393,N_43703,N_43179);
nand U45394 (N_45394,N_42180,N_43212);
xnor U45395 (N_45395,N_43137,N_43957);
nor U45396 (N_45396,N_42680,N_42884);
or U45397 (N_45397,N_43796,N_42309);
or U45398 (N_45398,N_42220,N_43526);
and U45399 (N_45399,N_43471,N_43005);
nand U45400 (N_45400,N_43336,N_43034);
nor U45401 (N_45401,N_43693,N_42097);
or U45402 (N_45402,N_43828,N_43172);
nand U45403 (N_45403,N_42977,N_42108);
xor U45404 (N_45404,N_43544,N_42859);
nand U45405 (N_45405,N_43073,N_43531);
nand U45406 (N_45406,N_42868,N_43045);
xor U45407 (N_45407,N_42808,N_43374);
or U45408 (N_45408,N_42289,N_43618);
nand U45409 (N_45409,N_43781,N_43039);
nand U45410 (N_45410,N_42967,N_43627);
or U45411 (N_45411,N_42270,N_43682);
nor U45412 (N_45412,N_42553,N_43488);
and U45413 (N_45413,N_42557,N_43640);
xnor U45414 (N_45414,N_43436,N_42010);
and U45415 (N_45415,N_43318,N_42821);
nand U45416 (N_45416,N_43659,N_43611);
and U45417 (N_45417,N_43239,N_42493);
xnor U45418 (N_45418,N_42343,N_43215);
or U45419 (N_45419,N_43146,N_43504);
nand U45420 (N_45420,N_42034,N_42808);
nor U45421 (N_45421,N_43550,N_43617);
nand U45422 (N_45422,N_43793,N_42181);
and U45423 (N_45423,N_42259,N_43465);
xnor U45424 (N_45424,N_42405,N_42112);
or U45425 (N_45425,N_43644,N_43660);
nand U45426 (N_45426,N_43470,N_42309);
and U45427 (N_45427,N_43659,N_42037);
nor U45428 (N_45428,N_43632,N_43907);
xnor U45429 (N_45429,N_43553,N_43686);
nor U45430 (N_45430,N_43842,N_43174);
or U45431 (N_45431,N_43242,N_42727);
nand U45432 (N_45432,N_42015,N_43859);
and U45433 (N_45433,N_43976,N_43471);
nand U45434 (N_45434,N_43549,N_43884);
nand U45435 (N_45435,N_43027,N_42612);
xor U45436 (N_45436,N_42825,N_43425);
nor U45437 (N_45437,N_42755,N_43120);
nor U45438 (N_45438,N_43237,N_43481);
nor U45439 (N_45439,N_43410,N_42564);
nor U45440 (N_45440,N_43052,N_43681);
nor U45441 (N_45441,N_42453,N_43645);
nand U45442 (N_45442,N_43038,N_43435);
and U45443 (N_45443,N_42398,N_42721);
or U45444 (N_45444,N_42526,N_43423);
nor U45445 (N_45445,N_43476,N_42031);
xor U45446 (N_45446,N_42417,N_42603);
nor U45447 (N_45447,N_42191,N_43262);
nor U45448 (N_45448,N_43397,N_42810);
or U45449 (N_45449,N_43223,N_43621);
xor U45450 (N_45450,N_42999,N_42759);
and U45451 (N_45451,N_42387,N_42923);
and U45452 (N_45452,N_42547,N_42085);
nor U45453 (N_45453,N_43920,N_42900);
and U45454 (N_45454,N_42914,N_43346);
or U45455 (N_45455,N_42359,N_42946);
nand U45456 (N_45456,N_43061,N_43462);
nand U45457 (N_45457,N_43671,N_42900);
nand U45458 (N_45458,N_42400,N_42274);
and U45459 (N_45459,N_42697,N_43104);
and U45460 (N_45460,N_43816,N_43818);
xnor U45461 (N_45461,N_42738,N_43074);
xnor U45462 (N_45462,N_42537,N_42694);
or U45463 (N_45463,N_42630,N_43120);
xnor U45464 (N_45464,N_42197,N_42573);
nor U45465 (N_45465,N_42223,N_43020);
nor U45466 (N_45466,N_43435,N_42284);
nor U45467 (N_45467,N_43855,N_42753);
and U45468 (N_45468,N_42624,N_42233);
nand U45469 (N_45469,N_43107,N_42115);
nor U45470 (N_45470,N_43783,N_42897);
nand U45471 (N_45471,N_43633,N_43332);
and U45472 (N_45472,N_43864,N_43144);
and U45473 (N_45473,N_42319,N_43600);
and U45474 (N_45474,N_43614,N_43861);
or U45475 (N_45475,N_42036,N_43481);
xnor U45476 (N_45476,N_42336,N_42021);
xnor U45477 (N_45477,N_42121,N_43647);
nand U45478 (N_45478,N_42620,N_42386);
and U45479 (N_45479,N_43497,N_42575);
and U45480 (N_45480,N_42334,N_43306);
or U45481 (N_45481,N_43836,N_43978);
nand U45482 (N_45482,N_42419,N_42455);
nor U45483 (N_45483,N_42502,N_42899);
and U45484 (N_45484,N_42118,N_43914);
or U45485 (N_45485,N_42461,N_42121);
xnor U45486 (N_45486,N_42414,N_42395);
and U45487 (N_45487,N_43814,N_42964);
nand U45488 (N_45488,N_43403,N_43185);
or U45489 (N_45489,N_43065,N_43372);
or U45490 (N_45490,N_43048,N_42983);
nand U45491 (N_45491,N_42735,N_43222);
xor U45492 (N_45492,N_42793,N_43614);
or U45493 (N_45493,N_43197,N_43744);
and U45494 (N_45494,N_43969,N_42371);
nand U45495 (N_45495,N_42581,N_42699);
xnor U45496 (N_45496,N_42739,N_42772);
nor U45497 (N_45497,N_43836,N_43528);
nand U45498 (N_45498,N_43424,N_42138);
nand U45499 (N_45499,N_43919,N_42110);
nor U45500 (N_45500,N_43031,N_42146);
nand U45501 (N_45501,N_43056,N_43261);
xor U45502 (N_45502,N_43143,N_43569);
or U45503 (N_45503,N_43906,N_42504);
nand U45504 (N_45504,N_42767,N_42834);
or U45505 (N_45505,N_42897,N_43387);
nand U45506 (N_45506,N_42960,N_43422);
and U45507 (N_45507,N_43681,N_42528);
or U45508 (N_45508,N_42227,N_42579);
nor U45509 (N_45509,N_42072,N_43363);
nand U45510 (N_45510,N_43581,N_43025);
and U45511 (N_45511,N_42476,N_42186);
or U45512 (N_45512,N_43964,N_42668);
or U45513 (N_45513,N_42278,N_42914);
nor U45514 (N_45514,N_43058,N_43426);
nand U45515 (N_45515,N_42323,N_42530);
nor U45516 (N_45516,N_42169,N_43804);
nor U45517 (N_45517,N_43673,N_42905);
or U45518 (N_45518,N_42784,N_43675);
or U45519 (N_45519,N_43697,N_43919);
nand U45520 (N_45520,N_43147,N_42560);
or U45521 (N_45521,N_43277,N_43704);
xor U45522 (N_45522,N_42393,N_43636);
and U45523 (N_45523,N_42424,N_42396);
nand U45524 (N_45524,N_43683,N_42093);
nor U45525 (N_45525,N_43164,N_42764);
and U45526 (N_45526,N_42377,N_42149);
or U45527 (N_45527,N_42421,N_42570);
and U45528 (N_45528,N_42666,N_42752);
nor U45529 (N_45529,N_42427,N_42657);
xor U45530 (N_45530,N_43834,N_43476);
or U45531 (N_45531,N_43144,N_43507);
xnor U45532 (N_45532,N_43758,N_42713);
nand U45533 (N_45533,N_42364,N_42447);
nand U45534 (N_45534,N_43987,N_43990);
xor U45535 (N_45535,N_42973,N_43212);
nand U45536 (N_45536,N_43741,N_43363);
nand U45537 (N_45537,N_42277,N_42315);
nor U45538 (N_45538,N_42718,N_42236);
xor U45539 (N_45539,N_42322,N_42280);
nand U45540 (N_45540,N_43257,N_43056);
nor U45541 (N_45541,N_42978,N_43390);
and U45542 (N_45542,N_43722,N_43264);
and U45543 (N_45543,N_43060,N_43196);
xor U45544 (N_45544,N_43354,N_42820);
nand U45545 (N_45545,N_42476,N_43797);
and U45546 (N_45546,N_42153,N_43230);
and U45547 (N_45547,N_43567,N_43580);
and U45548 (N_45548,N_43194,N_43331);
and U45549 (N_45549,N_42463,N_42526);
nand U45550 (N_45550,N_43004,N_42073);
or U45551 (N_45551,N_43839,N_43235);
or U45552 (N_45552,N_42313,N_42194);
xor U45553 (N_45553,N_42864,N_43090);
nor U45554 (N_45554,N_43218,N_42091);
xnor U45555 (N_45555,N_43128,N_43893);
and U45556 (N_45556,N_43222,N_43499);
nor U45557 (N_45557,N_42071,N_43555);
and U45558 (N_45558,N_42368,N_43506);
xnor U45559 (N_45559,N_42786,N_42544);
xor U45560 (N_45560,N_43778,N_43766);
or U45561 (N_45561,N_43000,N_42421);
nand U45562 (N_45562,N_43889,N_43466);
xnor U45563 (N_45563,N_42388,N_42012);
and U45564 (N_45564,N_43726,N_43426);
nor U45565 (N_45565,N_43970,N_42967);
and U45566 (N_45566,N_43655,N_43985);
and U45567 (N_45567,N_43239,N_43993);
nor U45568 (N_45568,N_42656,N_43970);
nor U45569 (N_45569,N_42968,N_43029);
nand U45570 (N_45570,N_42601,N_43906);
nand U45571 (N_45571,N_42230,N_43251);
nor U45572 (N_45572,N_42325,N_43269);
nand U45573 (N_45573,N_43440,N_42412);
nand U45574 (N_45574,N_42235,N_42966);
xnor U45575 (N_45575,N_43591,N_43708);
xor U45576 (N_45576,N_43262,N_42691);
or U45577 (N_45577,N_43073,N_42846);
or U45578 (N_45578,N_42863,N_42747);
nor U45579 (N_45579,N_42129,N_42030);
nor U45580 (N_45580,N_42323,N_43348);
and U45581 (N_45581,N_43220,N_43454);
nand U45582 (N_45582,N_43575,N_43010);
and U45583 (N_45583,N_42501,N_42016);
nand U45584 (N_45584,N_42746,N_42144);
xnor U45585 (N_45585,N_43654,N_43760);
or U45586 (N_45586,N_42536,N_43278);
xnor U45587 (N_45587,N_43807,N_42404);
xor U45588 (N_45588,N_42272,N_42971);
and U45589 (N_45589,N_43770,N_43910);
or U45590 (N_45590,N_42857,N_43301);
nand U45591 (N_45591,N_42711,N_43165);
or U45592 (N_45592,N_42720,N_42121);
or U45593 (N_45593,N_43410,N_43462);
xor U45594 (N_45594,N_42727,N_42134);
nand U45595 (N_45595,N_43570,N_43949);
or U45596 (N_45596,N_43180,N_43401);
nor U45597 (N_45597,N_43399,N_43371);
and U45598 (N_45598,N_43440,N_42501);
nand U45599 (N_45599,N_43541,N_42916);
nand U45600 (N_45600,N_43809,N_42726);
xnor U45601 (N_45601,N_42950,N_42928);
xnor U45602 (N_45602,N_42103,N_43217);
nand U45603 (N_45603,N_42205,N_43404);
nand U45604 (N_45604,N_42114,N_43976);
or U45605 (N_45605,N_42845,N_42372);
xor U45606 (N_45606,N_42315,N_42963);
xnor U45607 (N_45607,N_43152,N_43362);
and U45608 (N_45608,N_42438,N_43946);
xnor U45609 (N_45609,N_43994,N_42082);
nand U45610 (N_45610,N_42879,N_42936);
or U45611 (N_45611,N_42328,N_42378);
xnor U45612 (N_45612,N_42244,N_42514);
or U45613 (N_45613,N_43309,N_42118);
and U45614 (N_45614,N_43658,N_43451);
xnor U45615 (N_45615,N_42180,N_42947);
and U45616 (N_45616,N_43064,N_42411);
and U45617 (N_45617,N_43895,N_43615);
nor U45618 (N_45618,N_43136,N_42863);
nand U45619 (N_45619,N_42530,N_43718);
or U45620 (N_45620,N_42074,N_42162);
or U45621 (N_45621,N_43650,N_43230);
xnor U45622 (N_45622,N_43173,N_43948);
nand U45623 (N_45623,N_43802,N_43181);
nor U45624 (N_45624,N_43694,N_43183);
or U45625 (N_45625,N_43778,N_42501);
and U45626 (N_45626,N_42613,N_42420);
and U45627 (N_45627,N_42082,N_42772);
and U45628 (N_45628,N_43375,N_43427);
xnor U45629 (N_45629,N_43770,N_43248);
and U45630 (N_45630,N_42581,N_42016);
xnor U45631 (N_45631,N_43658,N_43560);
or U45632 (N_45632,N_43920,N_43103);
nor U45633 (N_45633,N_42339,N_42240);
nor U45634 (N_45634,N_43545,N_42582);
xor U45635 (N_45635,N_42241,N_42154);
and U45636 (N_45636,N_43894,N_42260);
and U45637 (N_45637,N_43356,N_42842);
nand U45638 (N_45638,N_43128,N_43415);
and U45639 (N_45639,N_42020,N_42539);
nor U45640 (N_45640,N_42486,N_43112);
and U45641 (N_45641,N_42698,N_42232);
nor U45642 (N_45642,N_43754,N_43733);
xor U45643 (N_45643,N_42846,N_42255);
or U45644 (N_45644,N_42657,N_43546);
or U45645 (N_45645,N_43538,N_43542);
nand U45646 (N_45646,N_43613,N_43094);
nand U45647 (N_45647,N_42027,N_42977);
or U45648 (N_45648,N_42015,N_43142);
nand U45649 (N_45649,N_42389,N_43698);
or U45650 (N_45650,N_42587,N_43082);
xor U45651 (N_45651,N_42079,N_42263);
nand U45652 (N_45652,N_43965,N_43414);
nor U45653 (N_45653,N_42483,N_42172);
nand U45654 (N_45654,N_43643,N_42869);
nand U45655 (N_45655,N_42932,N_42000);
nand U45656 (N_45656,N_43015,N_43811);
or U45657 (N_45657,N_43412,N_43220);
or U45658 (N_45658,N_43240,N_42177);
nor U45659 (N_45659,N_42915,N_43738);
nand U45660 (N_45660,N_43099,N_43443);
or U45661 (N_45661,N_42926,N_42413);
nor U45662 (N_45662,N_43722,N_43695);
nor U45663 (N_45663,N_42652,N_42202);
xor U45664 (N_45664,N_42413,N_43057);
and U45665 (N_45665,N_43882,N_42670);
xnor U45666 (N_45666,N_42550,N_42405);
nor U45667 (N_45667,N_42594,N_42353);
and U45668 (N_45668,N_42552,N_43223);
or U45669 (N_45669,N_43002,N_43983);
nor U45670 (N_45670,N_43510,N_42067);
xor U45671 (N_45671,N_42408,N_42857);
nand U45672 (N_45672,N_42058,N_42742);
and U45673 (N_45673,N_42183,N_43725);
nor U45674 (N_45674,N_42670,N_42939);
or U45675 (N_45675,N_43365,N_42109);
xor U45676 (N_45676,N_43270,N_43590);
nand U45677 (N_45677,N_43411,N_42574);
and U45678 (N_45678,N_43661,N_43227);
and U45679 (N_45679,N_43387,N_43925);
xnor U45680 (N_45680,N_43944,N_42625);
or U45681 (N_45681,N_43748,N_42492);
or U45682 (N_45682,N_42758,N_42285);
or U45683 (N_45683,N_43904,N_42758);
nor U45684 (N_45684,N_42590,N_42015);
and U45685 (N_45685,N_42827,N_42757);
or U45686 (N_45686,N_43152,N_43993);
nand U45687 (N_45687,N_43373,N_43870);
nand U45688 (N_45688,N_43503,N_43880);
or U45689 (N_45689,N_42278,N_42858);
nor U45690 (N_45690,N_43469,N_42691);
or U45691 (N_45691,N_42362,N_42575);
nand U45692 (N_45692,N_42391,N_43039);
and U45693 (N_45693,N_42407,N_42388);
or U45694 (N_45694,N_42938,N_42423);
and U45695 (N_45695,N_43456,N_42078);
xnor U45696 (N_45696,N_42243,N_43052);
or U45697 (N_45697,N_42417,N_43963);
nor U45698 (N_45698,N_43822,N_42820);
nor U45699 (N_45699,N_42567,N_42572);
xor U45700 (N_45700,N_43253,N_43297);
nor U45701 (N_45701,N_43224,N_43488);
or U45702 (N_45702,N_42887,N_42206);
or U45703 (N_45703,N_43918,N_43799);
nor U45704 (N_45704,N_43117,N_42916);
xor U45705 (N_45705,N_42683,N_42941);
or U45706 (N_45706,N_42934,N_43082);
and U45707 (N_45707,N_43615,N_43998);
xor U45708 (N_45708,N_43621,N_42487);
xor U45709 (N_45709,N_42498,N_43755);
or U45710 (N_45710,N_42449,N_43249);
xor U45711 (N_45711,N_42898,N_42328);
xnor U45712 (N_45712,N_43343,N_43663);
xor U45713 (N_45713,N_43006,N_43255);
nor U45714 (N_45714,N_43944,N_43629);
and U45715 (N_45715,N_42870,N_42911);
nand U45716 (N_45716,N_43544,N_43899);
and U45717 (N_45717,N_42478,N_43945);
nor U45718 (N_45718,N_42410,N_42796);
nor U45719 (N_45719,N_42014,N_42230);
or U45720 (N_45720,N_42723,N_43689);
or U45721 (N_45721,N_42799,N_42794);
nand U45722 (N_45722,N_42637,N_42108);
nand U45723 (N_45723,N_43886,N_42079);
nor U45724 (N_45724,N_43054,N_42415);
or U45725 (N_45725,N_42558,N_42163);
and U45726 (N_45726,N_42530,N_42079);
nor U45727 (N_45727,N_43076,N_42996);
nand U45728 (N_45728,N_42009,N_43851);
nand U45729 (N_45729,N_43203,N_43431);
nand U45730 (N_45730,N_43564,N_42918);
nor U45731 (N_45731,N_42466,N_43354);
nor U45732 (N_45732,N_42545,N_42291);
nor U45733 (N_45733,N_42732,N_43494);
or U45734 (N_45734,N_43199,N_43481);
nand U45735 (N_45735,N_42370,N_42092);
xnor U45736 (N_45736,N_43869,N_42254);
nor U45737 (N_45737,N_42633,N_42230);
xor U45738 (N_45738,N_42905,N_43672);
and U45739 (N_45739,N_43162,N_43006);
nor U45740 (N_45740,N_43687,N_43066);
and U45741 (N_45741,N_43226,N_43104);
nor U45742 (N_45742,N_42845,N_42394);
nand U45743 (N_45743,N_42414,N_43009);
nor U45744 (N_45744,N_43918,N_42751);
nor U45745 (N_45745,N_42556,N_43286);
xnor U45746 (N_45746,N_43145,N_43648);
and U45747 (N_45747,N_42091,N_42274);
or U45748 (N_45748,N_42843,N_43190);
nand U45749 (N_45749,N_43908,N_43289);
nor U45750 (N_45750,N_43734,N_42446);
xnor U45751 (N_45751,N_43051,N_43099);
nand U45752 (N_45752,N_43229,N_42322);
nor U45753 (N_45753,N_42862,N_42347);
nor U45754 (N_45754,N_42591,N_43038);
nor U45755 (N_45755,N_42350,N_43059);
nor U45756 (N_45756,N_42980,N_42440);
xor U45757 (N_45757,N_43888,N_42042);
or U45758 (N_45758,N_43026,N_42934);
nand U45759 (N_45759,N_43195,N_42267);
xor U45760 (N_45760,N_42052,N_43242);
xor U45761 (N_45761,N_42739,N_42079);
xor U45762 (N_45762,N_42887,N_42525);
and U45763 (N_45763,N_43774,N_43012);
and U45764 (N_45764,N_43431,N_43957);
nor U45765 (N_45765,N_43273,N_42120);
and U45766 (N_45766,N_43538,N_43406);
and U45767 (N_45767,N_42770,N_43760);
or U45768 (N_45768,N_42648,N_43414);
or U45769 (N_45769,N_43224,N_42517);
or U45770 (N_45770,N_43998,N_43777);
nand U45771 (N_45771,N_42563,N_42295);
nor U45772 (N_45772,N_43634,N_42873);
nand U45773 (N_45773,N_42509,N_42027);
nor U45774 (N_45774,N_42600,N_43299);
nor U45775 (N_45775,N_43569,N_43196);
or U45776 (N_45776,N_42098,N_42892);
nor U45777 (N_45777,N_43954,N_43272);
and U45778 (N_45778,N_42905,N_42821);
nand U45779 (N_45779,N_42759,N_42401);
nor U45780 (N_45780,N_43412,N_42325);
or U45781 (N_45781,N_42649,N_43293);
and U45782 (N_45782,N_42449,N_43613);
xor U45783 (N_45783,N_43711,N_42830);
or U45784 (N_45784,N_42732,N_42365);
xor U45785 (N_45785,N_42761,N_43921);
nand U45786 (N_45786,N_43310,N_43784);
nand U45787 (N_45787,N_42334,N_43793);
nor U45788 (N_45788,N_43088,N_43541);
xor U45789 (N_45789,N_43992,N_43051);
nand U45790 (N_45790,N_42789,N_42658);
nor U45791 (N_45791,N_42561,N_42634);
nand U45792 (N_45792,N_43034,N_43424);
or U45793 (N_45793,N_43164,N_42469);
xor U45794 (N_45794,N_42311,N_42044);
nor U45795 (N_45795,N_43514,N_42031);
or U45796 (N_45796,N_43282,N_42572);
and U45797 (N_45797,N_42093,N_42847);
or U45798 (N_45798,N_42838,N_43171);
nand U45799 (N_45799,N_43672,N_42907);
xor U45800 (N_45800,N_43374,N_43712);
and U45801 (N_45801,N_43037,N_42858);
nand U45802 (N_45802,N_42808,N_42839);
xor U45803 (N_45803,N_43993,N_43704);
or U45804 (N_45804,N_42609,N_42537);
or U45805 (N_45805,N_43904,N_43136);
nor U45806 (N_45806,N_42623,N_42859);
nor U45807 (N_45807,N_42505,N_42333);
or U45808 (N_45808,N_43490,N_43737);
and U45809 (N_45809,N_42359,N_43415);
xnor U45810 (N_45810,N_43750,N_43071);
xor U45811 (N_45811,N_43711,N_42103);
xor U45812 (N_45812,N_42589,N_42022);
nor U45813 (N_45813,N_43208,N_43813);
or U45814 (N_45814,N_43106,N_43639);
nor U45815 (N_45815,N_43061,N_42380);
and U45816 (N_45816,N_42514,N_43032);
and U45817 (N_45817,N_43025,N_42356);
nand U45818 (N_45818,N_43371,N_42659);
xnor U45819 (N_45819,N_43336,N_43868);
or U45820 (N_45820,N_42262,N_42290);
nor U45821 (N_45821,N_43324,N_43021);
or U45822 (N_45822,N_43964,N_43559);
or U45823 (N_45823,N_43318,N_43596);
nand U45824 (N_45824,N_43169,N_42229);
and U45825 (N_45825,N_42115,N_42326);
xor U45826 (N_45826,N_42396,N_42765);
nor U45827 (N_45827,N_42582,N_42671);
nand U45828 (N_45828,N_42560,N_43778);
nand U45829 (N_45829,N_42007,N_42335);
nand U45830 (N_45830,N_43537,N_43544);
nand U45831 (N_45831,N_43085,N_42503);
or U45832 (N_45832,N_43934,N_43710);
nor U45833 (N_45833,N_42467,N_42862);
nand U45834 (N_45834,N_42448,N_43332);
nand U45835 (N_45835,N_42001,N_43183);
and U45836 (N_45836,N_42017,N_43819);
nand U45837 (N_45837,N_43944,N_42544);
xor U45838 (N_45838,N_43732,N_43263);
or U45839 (N_45839,N_43938,N_43555);
or U45840 (N_45840,N_43805,N_42512);
xnor U45841 (N_45841,N_42678,N_43505);
xnor U45842 (N_45842,N_42383,N_42451);
xnor U45843 (N_45843,N_42277,N_43203);
xor U45844 (N_45844,N_43094,N_43612);
and U45845 (N_45845,N_42162,N_42595);
nor U45846 (N_45846,N_43309,N_43117);
xnor U45847 (N_45847,N_42174,N_43904);
nand U45848 (N_45848,N_42691,N_42746);
nor U45849 (N_45849,N_42872,N_43117);
nand U45850 (N_45850,N_43585,N_42909);
nor U45851 (N_45851,N_42616,N_42931);
xnor U45852 (N_45852,N_42709,N_42862);
nand U45853 (N_45853,N_42296,N_43410);
xor U45854 (N_45854,N_43025,N_42144);
or U45855 (N_45855,N_42959,N_42276);
xor U45856 (N_45856,N_42493,N_42851);
xor U45857 (N_45857,N_43944,N_42058);
nor U45858 (N_45858,N_43898,N_43220);
xnor U45859 (N_45859,N_42270,N_43169);
nand U45860 (N_45860,N_42984,N_43691);
and U45861 (N_45861,N_42569,N_43360);
or U45862 (N_45862,N_42486,N_42447);
and U45863 (N_45863,N_43305,N_43376);
and U45864 (N_45864,N_42793,N_42063);
or U45865 (N_45865,N_42660,N_43366);
nand U45866 (N_45866,N_42772,N_43557);
or U45867 (N_45867,N_43301,N_42974);
nor U45868 (N_45868,N_42506,N_43597);
or U45869 (N_45869,N_42604,N_42490);
nor U45870 (N_45870,N_43147,N_43157);
xor U45871 (N_45871,N_43195,N_42542);
and U45872 (N_45872,N_42700,N_43944);
and U45873 (N_45873,N_43087,N_43347);
or U45874 (N_45874,N_42617,N_42420);
xor U45875 (N_45875,N_42167,N_43058);
nor U45876 (N_45876,N_42258,N_42405);
and U45877 (N_45877,N_42348,N_43611);
or U45878 (N_45878,N_42805,N_42385);
nand U45879 (N_45879,N_42872,N_42475);
nor U45880 (N_45880,N_42243,N_43935);
xor U45881 (N_45881,N_43347,N_43486);
nor U45882 (N_45882,N_43125,N_43664);
nor U45883 (N_45883,N_43283,N_43921);
or U45884 (N_45884,N_43727,N_43434);
and U45885 (N_45885,N_43774,N_43105);
xor U45886 (N_45886,N_43701,N_43044);
or U45887 (N_45887,N_43588,N_43827);
xor U45888 (N_45888,N_42010,N_43648);
xnor U45889 (N_45889,N_43434,N_43892);
nand U45890 (N_45890,N_42106,N_43708);
nand U45891 (N_45891,N_43165,N_43197);
xor U45892 (N_45892,N_42306,N_42183);
nand U45893 (N_45893,N_43479,N_42420);
xnor U45894 (N_45894,N_43197,N_43797);
xnor U45895 (N_45895,N_42760,N_42092);
nand U45896 (N_45896,N_42029,N_42538);
or U45897 (N_45897,N_42092,N_43038);
nand U45898 (N_45898,N_42124,N_42681);
nor U45899 (N_45899,N_42182,N_43536);
nor U45900 (N_45900,N_42002,N_42530);
nand U45901 (N_45901,N_43276,N_42931);
or U45902 (N_45902,N_43084,N_42680);
nor U45903 (N_45903,N_43473,N_43747);
xnor U45904 (N_45904,N_43512,N_42553);
nand U45905 (N_45905,N_42181,N_42254);
and U45906 (N_45906,N_42452,N_43123);
xnor U45907 (N_45907,N_43089,N_43094);
and U45908 (N_45908,N_43857,N_43172);
nand U45909 (N_45909,N_43678,N_42705);
nand U45910 (N_45910,N_42557,N_42632);
and U45911 (N_45911,N_43026,N_42348);
xor U45912 (N_45912,N_43445,N_43203);
or U45913 (N_45913,N_42930,N_43629);
nor U45914 (N_45914,N_42243,N_43349);
nor U45915 (N_45915,N_43720,N_42394);
or U45916 (N_45916,N_43957,N_42869);
nand U45917 (N_45917,N_43643,N_43897);
nor U45918 (N_45918,N_43524,N_43863);
and U45919 (N_45919,N_43351,N_42468);
nor U45920 (N_45920,N_42813,N_43986);
and U45921 (N_45921,N_42750,N_43570);
nor U45922 (N_45922,N_42181,N_43924);
xnor U45923 (N_45923,N_43959,N_42584);
xnor U45924 (N_45924,N_43833,N_42323);
nand U45925 (N_45925,N_42721,N_43572);
nor U45926 (N_45926,N_43468,N_43067);
nor U45927 (N_45927,N_42527,N_42474);
nor U45928 (N_45928,N_42208,N_42970);
xor U45929 (N_45929,N_43242,N_43740);
nand U45930 (N_45930,N_42945,N_43594);
xor U45931 (N_45931,N_43312,N_43359);
or U45932 (N_45932,N_43006,N_43674);
nand U45933 (N_45933,N_42860,N_43022);
nor U45934 (N_45934,N_42086,N_43059);
nor U45935 (N_45935,N_43504,N_43531);
nand U45936 (N_45936,N_42721,N_42486);
nand U45937 (N_45937,N_43234,N_43745);
or U45938 (N_45938,N_42914,N_43766);
and U45939 (N_45939,N_43705,N_43110);
nand U45940 (N_45940,N_42061,N_43505);
xor U45941 (N_45941,N_42334,N_43935);
or U45942 (N_45942,N_43401,N_43015);
xnor U45943 (N_45943,N_43209,N_43893);
xor U45944 (N_45944,N_42497,N_43230);
and U45945 (N_45945,N_42886,N_43134);
or U45946 (N_45946,N_42715,N_42306);
or U45947 (N_45947,N_43356,N_42156);
or U45948 (N_45948,N_43261,N_43211);
xor U45949 (N_45949,N_43468,N_42840);
and U45950 (N_45950,N_42622,N_42603);
and U45951 (N_45951,N_42180,N_43110);
or U45952 (N_45952,N_42815,N_43605);
xnor U45953 (N_45953,N_43854,N_43239);
nand U45954 (N_45954,N_42080,N_43436);
xnor U45955 (N_45955,N_42966,N_42175);
and U45956 (N_45956,N_43324,N_43159);
nor U45957 (N_45957,N_43593,N_43236);
and U45958 (N_45958,N_42462,N_43353);
nor U45959 (N_45959,N_43185,N_42953);
or U45960 (N_45960,N_43845,N_43239);
xor U45961 (N_45961,N_43701,N_43728);
and U45962 (N_45962,N_42162,N_42307);
nand U45963 (N_45963,N_43857,N_43940);
and U45964 (N_45964,N_43544,N_42725);
nand U45965 (N_45965,N_42363,N_42526);
xnor U45966 (N_45966,N_42104,N_42599);
xnor U45967 (N_45967,N_43956,N_42283);
nor U45968 (N_45968,N_42083,N_43494);
or U45969 (N_45969,N_42846,N_42911);
nor U45970 (N_45970,N_43131,N_43386);
and U45971 (N_45971,N_42515,N_43828);
nand U45972 (N_45972,N_43156,N_43815);
or U45973 (N_45973,N_43812,N_43597);
xor U45974 (N_45974,N_42377,N_43780);
or U45975 (N_45975,N_42926,N_42780);
xnor U45976 (N_45976,N_42379,N_43787);
xor U45977 (N_45977,N_42997,N_42877);
or U45978 (N_45978,N_42889,N_43365);
nand U45979 (N_45979,N_42367,N_43331);
nor U45980 (N_45980,N_42130,N_43417);
or U45981 (N_45981,N_42830,N_42773);
xor U45982 (N_45982,N_42194,N_43514);
and U45983 (N_45983,N_42527,N_43417);
and U45984 (N_45984,N_43872,N_42193);
and U45985 (N_45985,N_43251,N_42516);
nor U45986 (N_45986,N_42357,N_42261);
and U45987 (N_45987,N_42631,N_43695);
and U45988 (N_45988,N_42049,N_42556);
or U45989 (N_45989,N_42955,N_42317);
xnor U45990 (N_45990,N_42470,N_43093);
and U45991 (N_45991,N_42864,N_42454);
xor U45992 (N_45992,N_43513,N_43853);
nand U45993 (N_45993,N_42998,N_42721);
and U45994 (N_45994,N_43646,N_42943);
and U45995 (N_45995,N_42305,N_43565);
nand U45996 (N_45996,N_42066,N_42198);
xor U45997 (N_45997,N_42181,N_43056);
or U45998 (N_45998,N_43090,N_42439);
xnor U45999 (N_45999,N_43027,N_43072);
nor U46000 (N_46000,N_45982,N_44983);
nor U46001 (N_46001,N_44783,N_44234);
xnor U46002 (N_46002,N_45471,N_44526);
nor U46003 (N_46003,N_44292,N_44589);
and U46004 (N_46004,N_44464,N_44148);
and U46005 (N_46005,N_45367,N_45707);
nand U46006 (N_46006,N_45320,N_44987);
nor U46007 (N_46007,N_45242,N_45805);
or U46008 (N_46008,N_45675,N_44721);
nor U46009 (N_46009,N_44326,N_45840);
nor U46010 (N_46010,N_44800,N_45610);
xor U46011 (N_46011,N_44053,N_44193);
nor U46012 (N_46012,N_44533,N_45773);
nor U46013 (N_46013,N_45767,N_44633);
nor U46014 (N_46014,N_45094,N_44830);
xnor U46015 (N_46015,N_44417,N_45299);
and U46016 (N_46016,N_45928,N_45657);
and U46017 (N_46017,N_44584,N_44873);
nand U46018 (N_46018,N_44444,N_45683);
or U46019 (N_46019,N_44974,N_44263);
nor U46020 (N_46020,N_44261,N_45969);
and U46021 (N_46021,N_45131,N_45075);
or U46022 (N_46022,N_45182,N_44018);
and U46023 (N_46023,N_45578,N_45852);
xnor U46024 (N_46024,N_44970,N_45209);
xnor U46025 (N_46025,N_44542,N_44063);
and U46026 (N_46026,N_45240,N_45561);
or U46027 (N_46027,N_45785,N_45487);
and U46028 (N_46028,N_45725,N_44335);
nor U46029 (N_46029,N_44502,N_44070);
and U46030 (N_46030,N_44937,N_44095);
nor U46031 (N_46031,N_45863,N_44620);
and U46032 (N_46032,N_45992,N_44511);
and U46033 (N_46033,N_44043,N_45125);
nor U46034 (N_46034,N_45964,N_45690);
and U46035 (N_46035,N_45359,N_45078);
nand U46036 (N_46036,N_45967,N_44075);
and U46037 (N_46037,N_45113,N_45894);
nand U46038 (N_46038,N_45495,N_44534);
and U46039 (N_46039,N_44808,N_45744);
nand U46040 (N_46040,N_44553,N_45274);
and U46041 (N_46041,N_44792,N_45458);
and U46042 (N_46042,N_44400,N_45331);
xor U46043 (N_46043,N_45574,N_45736);
or U46044 (N_46044,N_44210,N_44097);
nor U46045 (N_46045,N_44878,N_44723);
xnor U46046 (N_46046,N_45181,N_45018);
xnor U46047 (N_46047,N_44732,N_44863);
nand U46048 (N_46048,N_45356,N_45721);
and U46049 (N_46049,N_44154,N_44136);
nor U46050 (N_46050,N_44009,N_44952);
nand U46051 (N_46051,N_45454,N_45919);
xnor U46052 (N_46052,N_44169,N_44551);
nand U46053 (N_46053,N_44538,N_45842);
xor U46054 (N_46054,N_45255,N_44806);
nand U46055 (N_46055,N_45634,N_44085);
xor U46056 (N_46056,N_44494,N_45552);
or U46057 (N_46057,N_45210,N_44254);
xnor U46058 (N_46058,N_45243,N_45850);
xor U46059 (N_46059,N_45269,N_45778);
or U46060 (N_46060,N_44157,N_45271);
nand U46061 (N_46061,N_44113,N_45765);
xor U46062 (N_46062,N_44879,N_44159);
or U46063 (N_46063,N_44885,N_44945);
or U46064 (N_46064,N_45074,N_45195);
xor U46065 (N_46065,N_44177,N_45038);
or U46066 (N_46066,N_45710,N_44977);
nor U46067 (N_46067,N_45046,N_44675);
nor U46068 (N_46068,N_44237,N_45317);
or U46069 (N_46069,N_44574,N_45731);
and U46070 (N_46070,N_45417,N_44601);
nor U46071 (N_46071,N_45579,N_45005);
and U46072 (N_46072,N_45792,N_44373);
and U46073 (N_46073,N_45449,N_45508);
and U46074 (N_46074,N_45739,N_44065);
and U46075 (N_46075,N_44356,N_44605);
nor U46076 (N_46076,N_45564,N_45685);
and U46077 (N_46077,N_45387,N_44936);
nand U46078 (N_46078,N_45830,N_45577);
or U46079 (N_46079,N_44299,N_45039);
and U46080 (N_46080,N_44365,N_45238);
nor U46081 (N_46081,N_45073,N_44120);
and U46082 (N_46082,N_45581,N_44669);
nand U46083 (N_46083,N_44837,N_44378);
and U46084 (N_46084,N_44190,N_45627);
or U46085 (N_46085,N_45162,N_45312);
xnor U46086 (N_46086,N_45745,N_45455);
or U46087 (N_46087,N_45839,N_44349);
or U46088 (N_46088,N_44985,N_45213);
nand U46089 (N_46089,N_44214,N_44765);
or U46090 (N_46090,N_45793,N_45343);
nand U46091 (N_46091,N_45434,N_44414);
nor U46092 (N_46092,N_45396,N_45165);
xnor U46093 (N_46093,N_44036,N_44647);
and U46094 (N_46094,N_44957,N_45545);
xor U46095 (N_46095,N_44745,N_45229);
nor U46096 (N_46096,N_45931,N_44026);
nor U46097 (N_46097,N_44390,N_45522);
nor U46098 (N_46098,N_44173,N_44433);
xnor U46099 (N_46099,N_45045,N_44333);
and U46100 (N_46100,N_45953,N_45712);
xnor U46101 (N_46101,N_44838,N_45918);
nor U46102 (N_46102,N_44933,N_45171);
and U46103 (N_46103,N_44215,N_44908);
nor U46104 (N_46104,N_45788,N_44962);
or U46105 (N_46105,N_45965,N_45147);
or U46106 (N_46106,N_45499,N_45787);
xor U46107 (N_46107,N_45247,N_45491);
xor U46108 (N_46108,N_44849,N_45349);
or U46109 (N_46109,N_45813,N_44602);
nor U46110 (N_46110,N_44858,N_45479);
and U46111 (N_46111,N_45470,N_44920);
or U46112 (N_46112,N_44692,N_44258);
nand U46113 (N_46113,N_44662,N_44896);
nor U46114 (N_46114,N_45511,N_44304);
or U46115 (N_46115,N_45058,N_45060);
nor U46116 (N_46116,N_45207,N_44743);
nand U46117 (N_46117,N_44519,N_44324);
xnor U46118 (N_46118,N_45847,N_45421);
xnor U46119 (N_46119,N_44245,N_45093);
nor U46120 (N_46120,N_44344,N_44430);
nand U46121 (N_46121,N_45538,N_44803);
xor U46122 (N_46122,N_45007,N_44242);
nand U46123 (N_46123,N_44541,N_45228);
and U46124 (N_46124,N_44413,N_45310);
nor U46125 (N_46125,N_45733,N_45700);
or U46126 (N_46126,N_45987,N_45883);
xor U46127 (N_46127,N_44603,N_45889);
xor U46128 (N_46128,N_45670,N_45400);
nand U46129 (N_46129,N_45020,N_45150);
nand U46130 (N_46130,N_44906,N_44833);
xnor U46131 (N_46131,N_45880,N_45302);
or U46132 (N_46132,N_45430,N_44068);
nand U46133 (N_46133,N_44687,N_44932);
nor U46134 (N_46134,N_45697,N_44663);
nand U46135 (N_46135,N_45693,N_44066);
or U46136 (N_46136,N_44883,N_45701);
nand U46137 (N_46137,N_45630,N_45703);
nand U46138 (N_46138,N_45659,N_44161);
xnor U46139 (N_46139,N_44124,N_45575);
nor U46140 (N_46140,N_44203,N_44489);
or U46141 (N_46141,N_44999,N_45085);
xor U46142 (N_46142,N_45504,N_44287);
or U46143 (N_46143,N_45319,N_44546);
nor U46144 (N_46144,N_45122,N_45900);
nor U46145 (N_46145,N_44090,N_45107);
nand U46146 (N_46146,N_45542,N_44008);
xnor U46147 (N_46147,N_45071,N_44392);
and U46148 (N_46148,N_45993,N_44853);
or U46149 (N_46149,N_45591,N_45775);
nand U46150 (N_46150,N_45485,N_45891);
nand U46151 (N_46151,N_44290,N_44456);
and U46152 (N_46152,N_45724,N_44402);
xor U46153 (N_46153,N_45270,N_45300);
and U46154 (N_46154,N_45565,N_44831);
xnor U46155 (N_46155,N_45509,N_44967);
and U46156 (N_46156,N_45585,N_45451);
and U46157 (N_46157,N_44894,N_44088);
and U46158 (N_46158,N_44924,N_44485);
nand U46159 (N_46159,N_45617,N_45194);
xor U46160 (N_46160,N_44360,N_45087);
or U46161 (N_46161,N_44342,N_45002);
nor U46162 (N_46162,N_44825,N_44006);
xor U46163 (N_46163,N_45338,N_44865);
or U46164 (N_46164,N_44488,N_44102);
and U46165 (N_46165,N_44082,N_44828);
nor U46166 (N_46166,N_45407,N_45408);
and U46167 (N_46167,N_45374,N_45977);
nor U46168 (N_46168,N_44050,N_44595);
nand U46169 (N_46169,N_44320,N_45711);
and U46170 (N_46170,N_45594,N_44759);
and U46171 (N_46171,N_44752,N_44575);
and U46172 (N_46172,N_45111,N_45602);
xnor U46173 (N_46173,N_44802,N_44505);
nand U46174 (N_46174,N_45163,N_45426);
xor U46175 (N_46175,N_44766,N_44637);
and U46176 (N_46176,N_44117,N_45570);
and U46177 (N_46177,N_45436,N_45937);
and U46178 (N_46178,N_44507,N_45676);
nor U46179 (N_46179,N_45906,N_44612);
xnor U46180 (N_46180,N_44618,N_45480);
and U46181 (N_46181,N_44701,N_44656);
and U46182 (N_46182,N_45280,N_44998);
xor U46183 (N_46183,N_45867,N_44267);
and U46184 (N_46184,N_45829,N_44958);
nor U46185 (N_46185,N_44420,N_44517);
xor U46186 (N_46186,N_45529,N_45326);
or U46187 (N_46187,N_44121,N_45445);
and U46188 (N_46188,N_44561,N_44138);
xnor U46189 (N_46189,N_44953,N_45203);
xnor U46190 (N_46190,N_44416,N_45996);
nand U46191 (N_46191,N_45835,N_45029);
nor U46192 (N_46192,N_44409,N_44529);
or U46193 (N_46193,N_45998,N_45789);
xnor U46194 (N_46194,N_45492,N_44573);
nor U46195 (N_46195,N_45248,N_44524);
xor U46196 (N_46196,N_44316,N_45216);
or U46197 (N_46197,N_44588,N_44549);
and U46198 (N_46198,N_44297,N_44330);
nand U46199 (N_46199,N_44576,N_44798);
nand U46200 (N_46200,N_44727,N_44221);
and U46201 (N_46201,N_45862,N_44498);
nor U46202 (N_46202,N_45208,N_44740);
nand U46203 (N_46203,N_44126,N_45489);
xnor U46204 (N_46204,N_45502,N_44702);
or U46205 (N_46205,N_45102,N_45348);
xnor U46206 (N_46206,N_44199,N_44988);
xnor U46207 (N_46207,N_45358,N_45422);
or U46208 (N_46208,N_45366,N_44426);
nand U46209 (N_46209,N_45249,N_45266);
nand U46210 (N_46210,N_45772,N_44799);
and U46211 (N_46211,N_44239,N_45878);
xnor U46212 (N_46212,N_45418,N_44415);
nor U46213 (N_46213,N_45346,N_45121);
xnor U46214 (N_46214,N_44518,N_44790);
or U46215 (N_46215,N_44216,N_44145);
nor U46216 (N_46216,N_44904,N_44364);
and U46217 (N_46217,N_45682,N_45447);
nor U46218 (N_46218,N_44722,N_45006);
or U46219 (N_46219,N_45469,N_45934);
and U46220 (N_46220,N_45315,N_45543);
and U46221 (N_46221,N_45339,N_45450);
or U46222 (N_46222,N_44657,N_44112);
or U46223 (N_46223,N_44171,N_45554);
and U46224 (N_46224,N_44593,N_44391);
xnor U46225 (N_46225,N_45428,N_44230);
nand U46226 (N_46226,N_45179,N_44566);
nor U46227 (N_46227,N_45301,N_44389);
nand U46228 (N_46228,N_44064,N_45737);
and U46229 (N_46229,N_44341,N_45606);
and U46230 (N_46230,N_45369,N_44613);
or U46231 (N_46231,N_44960,N_45800);
or U46232 (N_46232,N_44011,N_44891);
or U46233 (N_46233,N_44086,N_44107);
and U46234 (N_46234,N_44362,N_44812);
or U46235 (N_46235,N_45373,N_44055);
or U46236 (N_46236,N_45140,N_44291);
nand U46237 (N_46237,N_45921,N_44981);
and U46238 (N_46238,N_44581,N_44950);
nor U46239 (N_46239,N_44910,N_45905);
and U46240 (N_46240,N_45128,N_45875);
nand U46241 (N_46241,N_44461,N_44471);
nand U46242 (N_46242,N_45652,N_45233);
nor U46243 (N_46243,N_44959,N_44616);
nor U46244 (N_46244,N_44038,N_44965);
and U46245 (N_46245,N_44582,N_44513);
or U46246 (N_46246,N_44580,N_44770);
or U46247 (N_46247,N_44228,N_45943);
xnor U46248 (N_46248,N_45753,N_44516);
or U46249 (N_46249,N_45599,N_44841);
nor U46250 (N_46250,N_45086,N_44673);
and U46251 (N_46251,N_45528,N_44836);
xnor U46252 (N_46252,N_44919,N_44668);
nand U46253 (N_46253,N_45215,N_45569);
nand U46254 (N_46254,N_44087,N_45580);
xnor U46255 (N_46255,N_45156,N_44811);
nor U46256 (N_46256,N_44822,N_45160);
and U46257 (N_46257,N_44226,N_45353);
nand U46258 (N_46258,N_44321,N_44104);
xnor U46259 (N_46259,N_45371,N_44590);
and U46260 (N_46260,N_44013,N_45549);
and U46261 (N_46261,N_44984,N_45858);
nor U46262 (N_46262,N_45911,N_45719);
nand U46263 (N_46263,N_44949,N_44780);
nand U46264 (N_46264,N_45292,N_44846);
nand U46265 (N_46265,N_44788,N_45566);
or U46266 (N_46266,N_45152,N_45596);
nor U46267 (N_46267,N_45028,N_44467);
nand U46268 (N_46268,N_45516,N_45443);
nand U46269 (N_46269,N_44719,N_45226);
xnor U46270 (N_46270,N_44938,N_44346);
xor U46271 (N_46271,N_45350,N_44544);
nand U46272 (N_46272,N_44583,N_44108);
nand U46273 (N_46273,N_44659,N_44751);
nor U46274 (N_46274,N_44850,N_45572);
xnor U46275 (N_46275,N_45362,N_44961);
xnor U46276 (N_46276,N_45077,N_44394);
nand U46277 (N_46277,N_45754,N_45391);
nor U46278 (N_46278,N_45730,N_44127);
nor U46279 (N_46279,N_45132,N_45275);
xnor U46280 (N_46280,N_45024,N_44144);
or U46281 (N_46281,N_44698,N_45735);
and U46282 (N_46282,N_44223,N_45896);
and U46283 (N_46283,N_45063,N_45424);
nand U46284 (N_46284,N_44852,N_45397);
and U46285 (N_46285,N_45611,N_45457);
nand U46286 (N_46286,N_45000,N_44405);
nor U46287 (N_46287,N_45468,N_45877);
nor U46288 (N_46288,N_45604,N_44654);
or U46289 (N_46289,N_44057,N_44617);
or U46290 (N_46290,N_45115,N_44328);
and U46291 (N_46291,N_44632,N_45419);
nand U46292 (N_46292,N_45250,N_44243);
or U46293 (N_46293,N_45833,N_45493);
xnor U46294 (N_46294,N_45717,N_44285);
and U46295 (N_46295,N_44480,N_45022);
nor U46296 (N_46296,N_45971,N_45874);
nor U46297 (N_46297,N_44492,N_45649);
nor U46298 (N_46298,N_45645,N_44074);
xnor U46299 (N_46299,N_45047,N_44619);
and U46300 (N_46300,N_44652,N_45536);
xor U46301 (N_46301,N_44046,N_44474);
nand U46302 (N_46302,N_44220,N_45101);
xnor U46303 (N_46303,N_45395,N_45674);
xor U46304 (N_46304,N_45819,N_45042);
or U46305 (N_46305,N_45429,N_44855);
xnor U46306 (N_46306,N_45756,N_45145);
and U46307 (N_46307,N_45855,N_44479);
nand U46308 (N_46308,N_45154,N_45252);
and U46309 (N_46309,N_45178,N_44458);
nand U46310 (N_46310,N_45550,N_44911);
or U46311 (N_46311,N_45861,N_44401);
or U46312 (N_46312,N_44880,N_45755);
and U46313 (N_46313,N_45589,N_45925);
or U46314 (N_46314,N_45036,N_44775);
nor U46315 (N_46315,N_44343,N_45081);
or U46316 (N_46316,N_45263,N_45054);
and U46317 (N_46317,N_44991,N_44350);
or U46318 (N_46318,N_44928,N_44528);
or U46319 (N_46319,N_45806,N_44579);
nand U46320 (N_46320,N_44639,N_44412);
and U46321 (N_46321,N_44556,N_45282);
nand U46322 (N_46322,N_44403,N_45378);
xnor U46323 (N_46323,N_44969,N_44867);
xor U46324 (N_46324,N_45605,N_44591);
or U46325 (N_46325,N_44315,N_45211);
nand U46326 (N_46326,N_44168,N_45206);
and U46327 (N_46327,N_44866,N_44348);
or U46328 (N_46328,N_44178,N_45390);
or U46329 (N_46329,N_45625,N_44819);
or U46330 (N_46330,N_44739,N_45979);
nor U46331 (N_46331,N_45278,N_44062);
and U46332 (N_46332,N_45963,N_44164);
nor U46333 (N_46333,N_45435,N_44441);
nand U46334 (N_46334,N_44882,N_44303);
and U46335 (N_46335,N_44889,N_44979);
or U46336 (N_46336,N_45968,N_44163);
and U46337 (N_46337,N_45313,N_45523);
nand U46338 (N_46338,N_45116,N_45986);
or U46339 (N_46339,N_45377,N_45403);
or U46340 (N_46340,N_44700,N_44381);
and U46341 (N_46341,N_44020,N_44678);
xor U46342 (N_46342,N_45665,N_45836);
nand U46343 (N_46343,N_44964,N_45540);
and U46344 (N_46344,N_44995,N_45118);
and U46345 (N_46345,N_45482,N_44302);
xor U46346 (N_46346,N_45595,N_45960);
nor U46347 (N_46347,N_45853,N_45709);
and U46348 (N_46348,N_45167,N_45288);
nand U46349 (N_46349,N_44207,N_45751);
nor U46350 (N_46350,N_45053,N_45794);
xnor U46351 (N_46351,N_44366,N_44897);
nand U46352 (N_46352,N_44472,N_44249);
xor U46353 (N_46353,N_45548,N_45886);
and U46354 (N_46354,N_44826,N_44101);
xnor U46355 (N_46355,N_45831,N_45032);
nor U46356 (N_46356,N_44531,N_45679);
nor U46357 (N_46357,N_45316,N_44729);
or U46358 (N_46358,N_45671,N_45644);
xor U46359 (N_46359,N_45234,N_45512);
and U46360 (N_46360,N_45563,N_45948);
or U46361 (N_46361,N_45926,N_45791);
nand U46362 (N_46362,N_45957,N_45825);
or U46363 (N_46363,N_45049,N_44925);
nand U46364 (N_46364,N_44629,N_45622);
xor U46365 (N_46365,N_45412,N_44829);
and U46366 (N_46366,N_44111,N_44329);
xor U46367 (N_46367,N_45342,N_44468);
nor U46368 (N_46368,N_45385,N_45108);
xnor U46369 (N_46369,N_45587,N_44670);
nor U46370 (N_46370,N_44737,N_44103);
and U46371 (N_46371,N_45083,N_45914);
nor U46372 (N_46372,N_44848,N_45534);
and U46373 (N_46373,N_45654,N_44437);
and U46374 (N_46374,N_44109,N_44080);
nand U46375 (N_46375,N_45868,N_44396);
and U46376 (N_46376,N_44259,N_45205);
xor U46377 (N_46377,N_44040,N_45218);
or U46378 (N_46378,N_44515,N_45064);
nor U46379 (N_46379,N_45030,N_45220);
nand U46380 (N_46380,N_44240,N_44487);
and U46381 (N_46381,N_44886,N_45786);
nand U46382 (N_46382,N_44547,N_44017);
xnor U46383 (N_46383,N_44359,N_45956);
or U46384 (N_46384,N_44311,N_45025);
nor U46385 (N_46385,N_45734,N_45603);
and U46386 (N_46386,N_44247,N_45533);
nor U46387 (N_46387,N_44715,N_44338);
or U46388 (N_46388,N_44310,N_45438);
nand U46389 (N_46389,N_44083,N_45881);
and U46390 (N_46390,N_45783,N_45808);
nand U46391 (N_46391,N_44093,N_44625);
xor U46392 (N_46392,N_44817,N_44921);
nand U46393 (N_46393,N_45376,N_44874);
xor U46394 (N_46394,N_45461,N_45192);
and U46395 (N_46395,N_45647,N_44160);
nand U46396 (N_46396,N_44809,N_44973);
and U46397 (N_46397,N_44913,N_44607);
or U46398 (N_46398,N_44695,N_44682);
xnor U46399 (N_46399,N_44621,N_45388);
nor U46400 (N_46400,N_45498,N_44918);
xor U46401 (N_46401,N_44369,N_44351);
nand U46402 (N_46402,N_45807,N_45866);
xnor U46403 (N_46403,N_45834,N_45272);
nor U46404 (N_46404,N_44915,N_45695);
or U46405 (N_46405,N_45660,N_45198);
nor U46406 (N_46406,N_45096,N_44931);
xor U46407 (N_46407,N_45202,N_44030);
or U46408 (N_46408,N_45537,N_44674);
or U46409 (N_46409,N_45084,N_45884);
xor U46410 (N_46410,N_45583,N_45651);
xnor U46411 (N_46411,N_45506,N_45157);
nand U46412 (N_46412,N_44149,N_45547);
nand U46413 (N_46413,N_44832,N_44100);
or U46414 (N_46414,N_44184,N_44514);
and U46415 (N_46415,N_44917,N_44246);
xor U46416 (N_46416,N_44767,N_44250);
xnor U46417 (N_46417,N_44231,N_44992);
xor U46418 (N_46418,N_44643,N_45974);
nor U46419 (N_46419,N_44035,N_45802);
xnor U46420 (N_46420,N_44422,N_44717);
or U46421 (N_46421,N_45091,N_44522);
and U46422 (N_46422,N_45100,N_44587);
xor U46423 (N_46423,N_44312,N_44888);
xor U46424 (N_46424,N_44916,N_44060);
nand U46425 (N_46425,N_44548,N_44379);
and U46426 (N_46426,N_45155,N_45988);
nand U46427 (N_46427,N_44861,N_45409);
xor U46428 (N_46428,N_44693,N_45513);
nor U46429 (N_46429,N_44476,N_45507);
nor U46430 (N_46430,N_44265,N_45262);
nand U46431 (N_46431,N_44747,N_44694);
nand U46432 (N_46432,N_44843,N_44902);
and U46433 (N_46433,N_44345,N_45483);
nor U46434 (N_46434,N_45246,N_44976);
nand U46435 (N_46435,N_45056,N_44777);
nor U46436 (N_46436,N_44372,N_45556);
nand U46437 (N_46437,N_44470,N_44881);
nor U46438 (N_46438,N_45464,N_45311);
and U46439 (N_46439,N_44434,N_44890);
xor U46440 (N_46440,N_44056,N_45927);
xor U46441 (N_46441,N_44705,N_44398);
nor U46442 (N_46442,N_45991,N_44382);
or U46443 (N_46443,N_45954,N_44114);
xor U46444 (N_46444,N_44432,N_45285);
or U46445 (N_46445,N_45031,N_45441);
xor U46446 (N_46446,N_45917,N_45559);
nor U46447 (N_46447,N_44651,N_44450);
nand U46448 (N_46448,N_45505,N_44182);
or U46449 (N_46449,N_44624,N_44001);
nand U46450 (N_46450,N_45909,N_44034);
and U46451 (N_46451,N_44762,N_44596);
nand U46452 (N_46452,N_44971,N_44418);
and U46453 (N_46453,N_45539,N_44189);
xor U46454 (N_46454,N_45609,N_45187);
xnor U46455 (N_46455,N_45328,N_45244);
nor U46456 (N_46456,N_45144,N_44857);
and U46457 (N_46457,N_45729,N_45224);
nand U46458 (N_46458,N_44684,N_45851);
nand U46459 (N_46459,N_44264,N_45279);
xnor U46460 (N_46460,N_44380,N_45392);
nor U46461 (N_46461,N_44209,N_44640);
or U46462 (N_46462,N_45713,N_44443);
or U46463 (N_46463,N_45932,N_45955);
nor U46464 (N_46464,N_45055,N_44776);
nor U46465 (N_46465,N_44997,N_44758);
xnor U46466 (N_46466,N_44248,N_44763);
and U46467 (N_46467,N_45336,N_45427);
and U46468 (N_46468,N_44367,N_44340);
nand U46469 (N_46469,N_45771,N_44482);
nand U46470 (N_46470,N_44045,N_44731);
xnor U46471 (N_46471,N_45066,N_45614);
or U46472 (N_46472,N_44054,N_44165);
xnor U46473 (N_46473,N_44914,N_44205);
nand U46474 (N_46474,N_44115,N_44336);
nor U46475 (N_46475,N_45360,N_45531);
and U46476 (N_46476,N_44069,N_45696);
or U46477 (N_46477,N_44294,N_45462);
or U46478 (N_46478,N_44804,N_45079);
nand U46479 (N_46479,N_44130,N_44211);
and U46480 (N_46480,N_45801,N_45290);
nand U46481 (N_46481,N_44842,N_45832);
and U46482 (N_46482,N_44005,N_45615);
or U46483 (N_46483,N_45325,N_44665);
nor U46484 (N_46484,N_45557,N_44608);
xnor U46485 (N_46485,N_44194,N_44941);
or U46486 (N_46486,N_45620,N_45260);
nand U46487 (N_46487,N_44975,N_45902);
nand U46488 (N_46488,N_44787,N_45624);
xnor U46489 (N_46489,N_45639,N_45673);
nand U46490 (N_46490,N_44404,N_44644);
nor U46491 (N_46491,N_45766,N_45026);
or U46492 (N_46492,N_44993,N_45009);
nand U46493 (N_46493,N_45947,N_44172);
or U46494 (N_46494,N_44688,N_44152);
or U46495 (N_46495,N_45404,N_44972);
nand U46496 (N_46496,N_45920,N_45626);
xnor U46497 (N_46497,N_45985,N_45173);
or U46498 (N_46498,N_45294,N_44483);
or U46499 (N_46499,N_45465,N_45318);
and U46500 (N_46500,N_45658,N_45929);
or U46501 (N_46501,N_45017,N_44142);
xor U46502 (N_46502,N_44135,N_44658);
nand U46503 (N_46503,N_45551,N_44820);
xnor U46504 (N_46504,N_45183,N_44307);
nand U46505 (N_46505,N_45705,N_44845);
xnor U46506 (N_46506,N_44730,N_44834);
and U46507 (N_46507,N_45437,N_44509);
xor U46508 (N_46508,N_45068,N_44206);
and U46509 (N_46509,N_45037,N_45139);
nand U46510 (N_46510,N_44314,N_44597);
nor U46511 (N_46511,N_44884,N_44912);
xnor U46512 (N_46512,N_44823,N_45264);
nor U46513 (N_46513,N_45860,N_45959);
nor U46514 (N_46514,N_44718,N_45910);
or U46515 (N_46515,N_45488,N_45432);
nand U46516 (N_46516,N_45520,N_44375);
nand U46517 (N_46517,N_45161,N_44810);
xnor U46518 (N_46518,N_45824,N_45268);
nor U46519 (N_46519,N_45386,N_45568);
nor U46520 (N_46520,N_45251,N_45646);
xnor U46521 (N_46521,N_45567,N_45095);
nand U46522 (N_46522,N_45341,N_45584);
or U46523 (N_46523,N_44195,N_45699);
or U46524 (N_46524,N_44929,N_44754);
nand U46525 (N_46525,N_45558,N_45780);
xnor U46526 (N_46526,N_45923,N_45981);
nor U46527 (N_46527,N_45003,N_45307);
nor U46528 (N_46528,N_44061,N_44847);
and U46529 (N_46529,N_45306,N_45184);
nor U46530 (N_46530,N_45650,N_44094);
nor U46531 (N_46531,N_45484,N_44934);
nand U46532 (N_46532,N_45526,N_45398);
xor U46533 (N_46533,N_45126,N_45916);
xor U46534 (N_46534,N_44623,N_44253);
or U46535 (N_46535,N_45219,N_44671);
nor U46536 (N_46536,N_45001,N_45277);
or U46537 (N_46537,N_44746,N_44477);
nor U46538 (N_46538,N_45798,N_45888);
or U46539 (N_46539,N_44497,N_44262);
nand U46540 (N_46540,N_45621,N_44681);
nor U46541 (N_46541,N_45854,N_45907);
nor U46542 (N_46542,N_44501,N_44646);
nand U46543 (N_46543,N_45689,N_45303);
nor U46544 (N_46544,N_45327,N_44044);
xor U46545 (N_46545,N_45466,N_44630);
nor U46546 (N_46546,N_44308,N_44286);
nor U46547 (N_46547,N_45221,N_44436);
nand U46548 (N_46548,N_44703,N_45930);
nor U46549 (N_46549,N_44188,N_45966);
or U46550 (N_46550,N_45678,N_44990);
nand U46551 (N_46551,N_44058,N_44019);
and U46552 (N_46552,N_44276,N_44406);
nand U46553 (N_46553,N_44923,N_44930);
nand U46554 (N_46554,N_44429,N_45628);
nand U46555 (N_46555,N_45490,N_45431);
and U46556 (N_46556,N_44004,N_44224);
xor U46557 (N_46557,N_44217,N_44181);
nor U46558 (N_46558,N_45159,N_44720);
or U46559 (N_46559,N_44000,N_44134);
and U46560 (N_46560,N_45692,N_44503);
and U46561 (N_46561,N_44555,N_45876);
xnor U46562 (N_46562,N_44563,N_44773);
nor U46563 (N_46563,N_44741,N_45663);
nor U46564 (N_46564,N_45448,N_44893);
and U46565 (N_46565,N_45571,N_44504);
and U46566 (N_46566,N_45414,N_45080);
and U46567 (N_46567,N_45681,N_44162);
and U46568 (N_46568,N_44385,N_45815);
nand U46569 (N_46569,N_45476,N_45023);
and U46570 (N_46570,N_45297,N_44905);
xnor U46571 (N_46571,N_45158,N_44284);
or U46572 (N_46572,N_44774,N_44014);
nor U46573 (N_46573,N_44175,N_45130);
or U46574 (N_46574,N_45241,N_45401);
nor U46575 (N_46575,N_45899,N_44872);
nand U46576 (N_46576,N_44235,N_44868);
xor U46577 (N_46577,N_44645,N_44192);
nand U46578 (N_46578,N_44685,N_44447);
nand U46579 (N_46579,N_45393,N_44072);
nand U46580 (N_46580,N_44572,N_44023);
nor U46581 (N_46581,N_45460,N_45134);
or U46582 (N_46582,N_45687,N_45496);
nand U46583 (N_46583,N_45185,N_45164);
and U46584 (N_46584,N_44092,N_44636);
xnor U46585 (N_46585,N_45997,N_45012);
and U46586 (N_46586,N_44185,N_45239);
and U46587 (N_46587,N_44465,N_45295);
xnor U46588 (N_46588,N_44676,N_44793);
and U46589 (N_46589,N_44951,N_44252);
and U46590 (N_46590,N_45291,N_44313);
and U46591 (N_46591,N_44059,N_44559);
nand U46592 (N_46592,N_44594,N_44073);
or U46593 (N_46593,N_45669,N_44183);
and U46594 (N_46594,N_45382,N_45746);
or U46595 (N_46595,N_44395,N_44028);
nand U46596 (N_46596,N_45694,N_45276);
nand U46597 (N_46597,N_44530,N_44728);
and U46598 (N_46598,N_45892,N_44523);
nand U46599 (N_46599,N_44196,N_44296);
nand U46600 (N_46600,N_44491,N_45843);
nand U46601 (N_46601,N_45738,N_44273);
and U46602 (N_46602,N_44600,N_45612);
nand U46603 (N_46603,N_45304,N_44560);
nor U46604 (N_46604,N_44438,N_44900);
nor U46605 (N_46605,N_44493,N_44212);
and U46606 (N_46606,N_44105,N_44421);
nor U46607 (N_46607,N_44564,N_44047);
nor U46608 (N_46608,N_44550,N_44578);
xor U46609 (N_46609,N_45763,N_45330);
and U46610 (N_46610,N_45636,N_45072);
nand U46611 (N_46611,N_44478,N_44186);
xnor U46612 (N_46612,N_44940,N_44358);
nor U46613 (N_46613,N_45517,N_45527);
xor U46614 (N_46614,N_45261,N_44821);
and U46615 (N_46615,N_45718,N_44269);
and U46616 (N_46616,N_44448,N_44948);
nand U46617 (N_46617,N_44796,N_45433);
nand U46618 (N_46618,N_44251,N_45057);
xnor U46619 (N_46619,N_45944,N_45972);
or U46620 (N_46620,N_44714,N_45950);
or U46621 (N_46621,N_45347,N_44814);
nand U46622 (N_46622,N_44048,N_45231);
nand U46623 (N_46623,N_45010,N_44219);
xnor U46624 (N_46624,N_44944,N_45089);
nor U46625 (N_46625,N_44052,N_44764);
or U46626 (N_46626,N_44197,N_44143);
nand U46627 (N_46627,N_44734,N_44986);
or U46628 (N_46628,N_45015,N_44554);
and U46629 (N_46629,N_45642,N_45643);
nand U46630 (N_46630,N_44318,N_44151);
xnor U46631 (N_46631,N_45553,N_45051);
or U46632 (N_46632,N_44091,N_45667);
or U46633 (N_46633,N_44892,N_45416);
and U46634 (N_46634,N_44610,N_44445);
nand U46635 (N_46635,N_45973,N_45329);
xor U46636 (N_46636,N_44225,N_45013);
and U46637 (N_46637,N_44994,N_45090);
nor U46638 (N_46638,N_44446,N_45641);
and U46639 (N_46639,N_44824,N_44903);
nor U46640 (N_46640,N_44325,N_44510);
nor U46641 (N_46641,N_45857,N_45980);
nand U46642 (N_46642,N_44167,N_44577);
nand U46643 (N_46643,N_44407,N_45782);
and U46644 (N_46644,N_45344,N_44760);
and U46645 (N_46645,N_45335,N_44462);
nor U46646 (N_46646,N_45473,N_45804);
or U46647 (N_46647,N_45105,N_44078);
or U46648 (N_46648,N_45518,N_44860);
or U46649 (N_46649,N_45514,N_45871);
and U46650 (N_46650,N_45702,N_44795);
nor U46651 (N_46651,N_45873,N_44208);
or U46652 (N_46652,N_44508,N_45014);
or U46653 (N_46653,N_45357,N_45174);
and U46654 (N_46654,N_44012,N_44966);
nor U46655 (N_46655,N_44386,N_44805);
nand U46656 (N_46656,N_44327,N_44496);
or U46657 (N_46657,N_44761,N_44558);
and U46658 (N_46658,N_44634,N_45812);
nand U46659 (N_46659,N_45668,N_44033);
or U46660 (N_46660,N_44704,N_44411);
xnor U46661 (N_46661,N_44042,N_45287);
nand U46662 (N_46662,N_45760,N_44757);
nand U46663 (N_46663,N_44779,N_45922);
or U46664 (N_46664,N_45859,N_44927);
and U46665 (N_46665,N_44631,N_44031);
nor U46666 (N_46666,N_45097,N_45592);
and U46667 (N_46667,N_45535,N_45364);
and U46668 (N_46668,N_44281,N_44106);
and U46669 (N_46669,N_45799,N_45481);
xnor U46670 (N_46670,N_44486,N_45501);
and U46671 (N_46671,N_44679,N_44453);
and U46672 (N_46672,N_45774,N_44628);
nand U46673 (N_46673,N_45380,N_44037);
and U46674 (N_46674,N_45935,N_44955);
nor U46675 (N_46675,N_45474,N_45779);
nor U46676 (N_46676,N_45334,N_45904);
nor U46677 (N_46677,N_45375,N_45758);
xnor U46678 (N_46678,N_44568,N_44641);
nor U46679 (N_46679,N_45016,N_45176);
or U46680 (N_46680,N_44536,N_44869);
nor U46681 (N_46681,N_44233,N_45440);
or U46682 (N_46682,N_44870,N_45989);
nand U46683 (N_46683,N_44425,N_45666);
and U46684 (N_46684,N_45684,N_45008);
and U46685 (N_46685,N_45257,N_45406);
nor U46686 (N_46686,N_45999,N_45608);
nor U46687 (N_46687,N_44374,N_45816);
and U46688 (N_46688,N_45796,N_44778);
nand U46689 (N_46689,N_44614,N_45245);
or U46690 (N_46690,N_44270,N_45811);
or U46691 (N_46691,N_45648,N_45354);
and U46692 (N_46692,N_44785,N_44440);
nand U46693 (N_46693,N_44709,N_44110);
nor U46694 (N_46694,N_44352,N_44331);
nor U46695 (N_46695,N_44282,N_45764);
nand U46696 (N_46696,N_45759,N_45882);
or U46697 (N_46697,N_44238,N_45059);
nand U46698 (N_46698,N_45913,N_44570);
or U46699 (N_46699,N_45170,N_44939);
xnor U46700 (N_46700,N_45041,N_44604);
nand U46701 (N_46701,N_45142,N_44586);
xor U46702 (N_46702,N_45453,N_44025);
xor U46703 (N_46703,N_45938,N_45237);
nor U46704 (N_46704,N_45446,N_44089);
or U46705 (N_46705,N_44909,N_44410);
nor U46706 (N_46706,N_45510,N_44125);
and U46707 (N_46707,N_44289,N_44495);
and U46708 (N_46708,N_44655,N_44213);
nor U46709 (N_46709,N_44689,N_44801);
and U46710 (N_46710,N_45352,N_45732);
nand U46711 (N_46711,N_45452,N_44255);
nand U46712 (N_46712,N_45688,N_44525);
or U46713 (N_46713,N_44187,N_45826);
or U46714 (N_46714,N_45112,N_45340);
nor U46715 (N_46715,N_44690,N_44371);
xor U46716 (N_46716,N_44419,N_44439);
nor U46717 (N_46717,N_44898,N_44424);
xor U46718 (N_46718,N_44332,N_45915);
nand U46719 (N_46719,N_44609,N_44027);
nand U46720 (N_46720,N_45048,N_44899);
xor U46721 (N_46721,N_44781,N_45444);
nand U46722 (N_46722,N_44653,N_44660);
or U46723 (N_46723,N_44840,N_45828);
nand U46724 (N_46724,N_44552,N_44545);
nor U46725 (N_46725,N_45515,N_45214);
and U46726 (N_46726,N_44611,N_44922);
or U46727 (N_46727,N_44260,N_44935);
nor U46728 (N_46728,N_44140,N_45477);
xor U46729 (N_46729,N_44543,N_45573);
and U46730 (N_46730,N_45752,N_45321);
nand U46731 (N_46731,N_44098,N_44334);
nor U46732 (N_46732,N_44506,N_44672);
nand U46733 (N_46733,N_44361,N_44191);
nor U46734 (N_46734,N_44275,N_44039);
nor U46735 (N_46735,N_44010,N_45769);
and U46736 (N_46736,N_44648,N_45503);
nand U46737 (N_46737,N_45995,N_44024);
and U46738 (N_46738,N_45151,N_44750);
or U46739 (N_46739,N_45590,N_45706);
xnor U46740 (N_46740,N_45727,N_45781);
and U46741 (N_46741,N_44096,N_45332);
and U46742 (N_46742,N_44428,N_45472);
nor U46743 (N_46743,N_44677,N_45052);
and U46744 (N_46744,N_44711,N_45936);
xnor U46745 (N_46745,N_45741,N_45912);
nor U46746 (N_46746,N_45521,N_45757);
nor U46747 (N_46747,N_45399,N_44650);
or U46748 (N_46748,N_44003,N_45704);
nand U46749 (N_46749,N_44851,N_45337);
or U46750 (N_46750,N_44499,N_44738);
or U46751 (N_46751,N_45146,N_44535);
or U46752 (N_46752,N_44129,N_45716);
or U46753 (N_46753,N_44166,N_45402);
and U46754 (N_46754,N_44642,N_44946);
nor U46755 (N_46755,N_44298,N_44733);
nor U46756 (N_46756,N_44756,N_44141);
and U46757 (N_46757,N_45740,N_44512);
and U46758 (N_46758,N_44022,N_45143);
nor U46759 (N_46759,N_44753,N_45136);
xor U46760 (N_46760,N_45166,N_45761);
nand U46761 (N_46761,N_44393,N_45137);
or U46762 (N_46762,N_45821,N_44696);
or U46763 (N_46763,N_45803,N_44076);
nand U46764 (N_46764,N_45175,N_44980);
xor U46765 (N_46765,N_44452,N_45661);
xor U46766 (N_46766,N_45410,N_44854);
nand U46767 (N_46767,N_44132,N_45662);
xor U46768 (N_46768,N_44427,N_45289);
nand U46769 (N_46769,N_44475,N_45177);
nand U46770 (N_46770,N_44707,N_44638);
nor U46771 (N_46771,N_44887,N_45562);
and U46772 (N_46772,N_45762,N_44201);
and U46773 (N_46773,N_44271,N_45893);
or U46774 (N_46774,N_44399,N_44856);
or U46775 (N_46775,N_44963,N_45864);
xnor U46776 (N_46776,N_45281,N_45777);
nor U46777 (N_46777,N_44691,N_44520);
and U46778 (N_46778,N_44002,N_44481);
nor U46779 (N_46779,N_45099,N_45486);
xnor U46780 (N_46780,N_45286,N_45225);
nor U46781 (N_46781,N_45619,N_45784);
and U46782 (N_46782,N_44202,N_45728);
and U46783 (N_46783,N_45305,N_45749);
or U46784 (N_46784,N_44744,N_44435);
nand U46785 (N_46785,N_44569,N_44791);
xnor U46786 (N_46786,N_45838,N_45379);
nor U46787 (N_46787,N_44442,N_45961);
and U46788 (N_46788,N_45588,N_45949);
or U46789 (N_46789,N_45070,N_44768);
nor U46790 (N_46790,N_44278,N_44716);
or U46791 (N_46791,N_44323,N_45691);
and U46792 (N_46792,N_44968,N_44724);
or U46793 (N_46793,N_45817,N_44521);
or U46794 (N_46794,N_45168,N_44454);
xor U46795 (N_46795,N_44844,N_44697);
nor U46796 (N_46796,N_45033,N_44954);
nand U46797 (N_46797,N_44943,N_45940);
xor U46798 (N_46798,N_45976,N_45411);
and U46799 (N_46799,N_44277,N_44119);
nand U46800 (N_46800,N_44128,N_45990);
nand U46801 (N_46801,N_44769,N_45984);
nor U46802 (N_46802,N_45200,N_45308);
xor U46803 (N_46803,N_45631,N_45942);
nor U46804 (N_46804,N_45872,N_44322);
or U46805 (N_46805,N_44079,N_45459);
xnor U46806 (N_46806,N_45952,N_44626);
and U46807 (N_46807,N_44875,N_44354);
and U46808 (N_46808,N_45903,N_44713);
and U46809 (N_46809,N_45361,N_45153);
nand U46810 (N_46810,N_44664,N_44712);
nand U46811 (N_46811,N_44978,N_44680);
xor U46812 (N_46812,N_44500,N_45750);
nand U46813 (N_46813,N_44490,N_44667);
and U46814 (N_46814,N_45082,N_45365);
nor U46815 (N_46815,N_45519,N_45885);
and U46816 (N_46816,N_44782,N_45050);
nand U46817 (N_46817,N_44532,N_45616);
nor U46818 (N_46818,N_45129,N_45869);
and U46819 (N_46819,N_45284,N_45887);
xnor U46820 (N_46820,N_45098,N_45188);
or U46821 (N_46821,N_44131,N_44748);
xor U46822 (N_46822,N_45597,N_44431);
nor U46823 (N_46823,N_45941,N_45598);
or U46824 (N_46824,N_44032,N_45525);
xor U46825 (N_46825,N_45546,N_44942);
nand U46826 (N_46826,N_44982,N_44585);
or U46827 (N_46827,N_45823,N_44571);
nor U46828 (N_46828,N_44071,N_44179);
xor U46829 (N_46829,N_45363,N_44726);
nor U46830 (N_46830,N_45124,N_45296);
xor U46831 (N_46831,N_44139,N_45848);
and U46832 (N_46832,N_45708,N_45790);
and U46833 (N_46833,N_44562,N_45672);
nor U46834 (N_46834,N_44133,N_45664);
or U46835 (N_46835,N_44029,N_45415);
and U46836 (N_46836,N_45743,N_45629);
or U46837 (N_46837,N_45267,N_44592);
nand U46838 (N_46838,N_44257,N_44473);
and U46839 (N_46839,N_45370,N_44947);
and U46840 (N_46840,N_45235,N_45653);
nor U46841 (N_46841,N_44353,N_44827);
and U46842 (N_46842,N_44339,N_45497);
or U46843 (N_46843,N_44606,N_44084);
xor U46844 (N_46844,N_45092,N_44540);
xnor U46845 (N_46845,N_44864,N_44384);
nand U46846 (N_46846,N_45962,N_45897);
nand U46847 (N_46847,N_44236,N_44859);
or U46848 (N_46848,N_44147,N_45405);
nor U46849 (N_46849,N_45467,N_45413);
and U46850 (N_46850,N_44683,N_45635);
nor U46851 (N_46851,N_45582,N_45822);
nor U46852 (N_46852,N_44784,N_44241);
nand U46853 (N_46853,N_44710,N_44118);
nor U46854 (N_46854,N_45895,N_44725);
nand U46855 (N_46855,N_44368,N_45062);
and U46856 (N_46856,N_44081,N_45714);
nor U46857 (N_46857,N_44174,N_45768);
or U46858 (N_46858,N_44355,N_44789);
xor U46859 (N_46859,N_44137,N_45637);
or U46860 (N_46860,N_44295,N_45109);
or U46861 (N_46861,N_44176,N_45439);
nand U46862 (N_46862,N_45169,N_45524);
nor U46863 (N_46863,N_45827,N_44268);
nor U46864 (N_46864,N_45879,N_45994);
or U46865 (N_46865,N_44895,N_44300);
nor U46866 (N_46866,N_45946,N_45172);
or U46867 (N_46867,N_45463,N_44622);
xor U46868 (N_46868,N_45975,N_45809);
and U46869 (N_46869,N_45227,N_45655);
or U46870 (N_46870,N_45541,N_45600);
nand U46871 (N_46871,N_45067,N_45500);
nor U46872 (N_46872,N_44484,N_45283);
nor U46873 (N_46873,N_45607,N_45958);
and U46874 (N_46874,N_45898,N_45846);
nand U46875 (N_46875,N_44408,N_45069);
nor U46876 (N_46876,N_44123,N_44772);
nor U46877 (N_46877,N_44227,N_44067);
and U46878 (N_46878,N_44317,N_45381);
nor U46879 (N_46879,N_45199,N_44686);
or U46880 (N_46880,N_45638,N_44016);
xnor U46881 (N_46881,N_45389,N_45747);
nor U46882 (N_46882,N_44288,N_45222);
xnor U46883 (N_46883,N_45019,N_44153);
xor U46884 (N_46884,N_44598,N_45256);
or U46885 (N_46885,N_45383,N_45236);
nor U46886 (N_46886,N_44347,N_44021);
xor U46887 (N_46887,N_45530,N_44170);
nand U46888 (N_46888,N_44835,N_44749);
nand U46889 (N_46889,N_45795,N_45742);
or U46890 (N_46890,N_45196,N_44198);
and U46891 (N_46891,N_45908,N_45722);
xor U46892 (N_46892,N_44871,N_45135);
and U46893 (N_46893,N_44742,N_45127);
nand U46894 (N_46894,N_44615,N_45223);
nand U46895 (N_46895,N_45820,N_45021);
xnor U46896 (N_46896,N_44256,N_44309);
nand U46897 (N_46897,N_45456,N_44319);
and U46898 (N_46898,N_44661,N_45027);
nand U46899 (N_46899,N_45273,N_45837);
nor U46900 (N_46900,N_44363,N_45970);
and U46901 (N_46901,N_45201,N_44244);
or U46902 (N_46902,N_44807,N_45141);
nand U46903 (N_46903,N_45939,N_44229);
xnor U46904 (N_46904,N_45104,N_45686);
xor U46905 (N_46905,N_45044,N_45217);
xnor U46906 (N_46906,N_44150,N_44699);
or U46907 (N_46907,N_45117,N_45043);
xor U46908 (N_46908,N_45841,N_44649);
nand U46909 (N_46909,N_45204,N_44280);
xor U46910 (N_46910,N_44877,N_44049);
or U46911 (N_46911,N_44459,N_44155);
nor U46912 (N_46912,N_45355,N_45114);
and U46913 (N_46913,N_44463,N_45983);
nor U46914 (N_46914,N_45230,N_44989);
and U46915 (N_46915,N_45814,N_44666);
xor U46916 (N_46916,N_44077,N_44451);
and U46917 (N_46917,N_44771,N_45698);
xnor U46918 (N_46918,N_44301,N_45120);
nor U46919 (N_46919,N_44218,N_44706);
xor U46920 (N_46920,N_45845,N_45586);
nor U46921 (N_46921,N_44539,N_44293);
or U46922 (N_46922,N_45776,N_44736);
and U46923 (N_46923,N_44423,N_44815);
xor U46924 (N_46924,N_45040,N_44794);
xor U46925 (N_46925,N_45309,N_45011);
or U46926 (N_46926,N_44567,N_44370);
and U46927 (N_46927,N_44306,N_45945);
and U46928 (N_46928,N_45924,N_44527);
or U46929 (N_46929,N_44627,N_45333);
nor U46930 (N_46930,N_45193,N_44305);
nand U46931 (N_46931,N_45818,N_45191);
nand U46932 (N_46932,N_44337,N_45656);
and U46933 (N_46933,N_45123,N_44274);
and U46934 (N_46934,N_45560,N_45555);
xor U46935 (N_46935,N_45265,N_45601);
xor U46936 (N_46936,N_45632,N_45425);
or U46937 (N_46937,N_44839,N_45061);
nand U46938 (N_46938,N_45901,N_44397);
nor U46939 (N_46939,N_44926,N_45715);
nand U46940 (N_46940,N_44457,N_44122);
and U46941 (N_46941,N_45232,N_45103);
and U46942 (N_46942,N_44051,N_44449);
and U46943 (N_46943,N_45726,N_45314);
nand U46944 (N_46944,N_45368,N_44279);
or U46945 (N_46945,N_44146,N_44755);
and U46946 (N_46946,N_45324,N_45186);
and U46947 (N_46947,N_45189,N_44388);
and U46948 (N_46948,N_44469,N_44599);
and U46949 (N_46949,N_45797,N_44266);
or U46950 (N_46950,N_45076,N_45197);
nor U46951 (N_46951,N_44180,N_45106);
xor U46952 (N_46952,N_44156,N_45258);
nand U46953 (N_46953,N_45322,N_44797);
and U46954 (N_46954,N_45394,N_45475);
nor U46955 (N_46955,N_44907,N_44455);
nor U46956 (N_46956,N_45351,N_45613);
nor U46957 (N_46957,N_45856,N_44565);
nand U46958 (N_46958,N_45148,N_44357);
xnor U46959 (N_46959,N_45119,N_45034);
or U46960 (N_46960,N_45494,N_45180);
nand U46961 (N_46961,N_44786,N_45933);
nor U46962 (N_46962,N_45384,N_44007);
xor U46963 (N_46963,N_45442,N_45423);
or U46964 (N_46964,N_45680,N_44015);
or U46965 (N_46965,N_44818,N_45870);
or U46966 (N_46966,N_45190,N_45133);
or U46967 (N_46967,N_45544,N_44222);
xnor U46968 (N_46968,N_45633,N_45254);
and U46969 (N_46969,N_44635,N_45110);
and U46970 (N_46970,N_44376,N_44813);
nand U46971 (N_46971,N_44116,N_44557);
xnor U46972 (N_46972,N_45951,N_44158);
xnor U46973 (N_46973,N_44996,N_45372);
nand U46974 (N_46974,N_45004,N_44041);
nor U46975 (N_46975,N_45253,N_44232);
and U46976 (N_46976,N_45532,N_45576);
nor U46977 (N_46977,N_45810,N_45478);
and U46978 (N_46978,N_45978,N_44708);
nand U46979 (N_46979,N_44901,N_45323);
or U46980 (N_46980,N_45259,N_44099);
or U46981 (N_46981,N_45593,N_44537);
nor U46982 (N_46982,N_44200,N_45298);
nand U46983 (N_46983,N_44816,N_45748);
nand U46984 (N_46984,N_44956,N_45212);
or U46985 (N_46985,N_45640,N_44466);
and U46986 (N_46986,N_45618,N_44204);
nand U46987 (N_46987,N_45149,N_44272);
xor U46988 (N_46988,N_45720,N_44460);
and U46989 (N_46989,N_45677,N_44283);
or U46990 (N_46990,N_45890,N_45420);
nand U46991 (N_46991,N_45723,N_44876);
or U46992 (N_46992,N_44735,N_45035);
or U46993 (N_46993,N_44377,N_45770);
nor U46994 (N_46994,N_45849,N_44862);
and U46995 (N_46995,N_44387,N_45088);
and U46996 (N_46996,N_45138,N_45065);
or U46997 (N_46997,N_45345,N_45623);
or U46998 (N_46998,N_45293,N_45844);
or U46999 (N_46999,N_45865,N_44383);
nor U47000 (N_47000,N_45646,N_45655);
nor U47001 (N_47001,N_44207,N_45538);
and U47002 (N_47002,N_44017,N_45810);
nor U47003 (N_47003,N_45614,N_45096);
or U47004 (N_47004,N_45141,N_45012);
nor U47005 (N_47005,N_45091,N_45863);
xnor U47006 (N_47006,N_45694,N_45126);
or U47007 (N_47007,N_45951,N_44041);
xor U47008 (N_47008,N_45420,N_45341);
or U47009 (N_47009,N_44527,N_45255);
or U47010 (N_47010,N_44414,N_44299);
or U47011 (N_47011,N_44169,N_44483);
xnor U47012 (N_47012,N_45030,N_44441);
nor U47013 (N_47013,N_45484,N_45704);
and U47014 (N_47014,N_45604,N_44993);
xor U47015 (N_47015,N_45737,N_45315);
xnor U47016 (N_47016,N_44290,N_45168);
and U47017 (N_47017,N_44840,N_44464);
and U47018 (N_47018,N_45040,N_44755);
nor U47019 (N_47019,N_45152,N_45658);
xor U47020 (N_47020,N_45578,N_45860);
xor U47021 (N_47021,N_44640,N_45889);
nor U47022 (N_47022,N_45850,N_45844);
nor U47023 (N_47023,N_44719,N_44505);
or U47024 (N_47024,N_45666,N_44572);
or U47025 (N_47025,N_44196,N_44412);
nor U47026 (N_47026,N_44218,N_45740);
or U47027 (N_47027,N_45879,N_44997);
or U47028 (N_47028,N_45011,N_45394);
nand U47029 (N_47029,N_44617,N_45522);
xor U47030 (N_47030,N_45195,N_45250);
xnor U47031 (N_47031,N_45991,N_44136);
xor U47032 (N_47032,N_44050,N_45272);
nand U47033 (N_47033,N_44539,N_44402);
or U47034 (N_47034,N_45921,N_45077);
nor U47035 (N_47035,N_44696,N_44166);
nor U47036 (N_47036,N_44232,N_44188);
or U47037 (N_47037,N_45974,N_44250);
xnor U47038 (N_47038,N_45371,N_44610);
and U47039 (N_47039,N_45575,N_45065);
and U47040 (N_47040,N_44195,N_44089);
and U47041 (N_47041,N_44131,N_45231);
and U47042 (N_47042,N_45761,N_44071);
and U47043 (N_47043,N_44769,N_45122);
nor U47044 (N_47044,N_44448,N_45462);
or U47045 (N_47045,N_45170,N_44738);
nand U47046 (N_47046,N_45286,N_45193);
nor U47047 (N_47047,N_44546,N_44440);
nand U47048 (N_47048,N_45534,N_44843);
nor U47049 (N_47049,N_45373,N_44537);
and U47050 (N_47050,N_45502,N_44299);
xor U47051 (N_47051,N_44685,N_45360);
and U47052 (N_47052,N_44359,N_45583);
nor U47053 (N_47053,N_44636,N_45199);
and U47054 (N_47054,N_45630,N_45654);
and U47055 (N_47055,N_44322,N_44428);
nor U47056 (N_47056,N_44825,N_45952);
or U47057 (N_47057,N_44598,N_45835);
nand U47058 (N_47058,N_45215,N_44697);
xor U47059 (N_47059,N_44156,N_44121);
nand U47060 (N_47060,N_45108,N_44430);
nor U47061 (N_47061,N_45017,N_44002);
xnor U47062 (N_47062,N_44620,N_45265);
xnor U47063 (N_47063,N_45183,N_44420);
nand U47064 (N_47064,N_44208,N_44480);
or U47065 (N_47065,N_44473,N_44586);
nor U47066 (N_47066,N_44803,N_45967);
nand U47067 (N_47067,N_45868,N_45727);
nor U47068 (N_47068,N_44536,N_44416);
nand U47069 (N_47069,N_44266,N_44307);
nand U47070 (N_47070,N_44468,N_45869);
and U47071 (N_47071,N_45189,N_45366);
or U47072 (N_47072,N_44678,N_45024);
nand U47073 (N_47073,N_44485,N_45496);
nor U47074 (N_47074,N_44460,N_44560);
nor U47075 (N_47075,N_44630,N_45828);
nand U47076 (N_47076,N_45550,N_45167);
and U47077 (N_47077,N_44441,N_45176);
or U47078 (N_47078,N_44330,N_44795);
nor U47079 (N_47079,N_44650,N_44840);
or U47080 (N_47080,N_45148,N_45683);
nand U47081 (N_47081,N_44980,N_45586);
nor U47082 (N_47082,N_45023,N_44789);
or U47083 (N_47083,N_44784,N_44838);
xnor U47084 (N_47084,N_44857,N_44806);
nor U47085 (N_47085,N_45893,N_44316);
nor U47086 (N_47086,N_44817,N_44207);
or U47087 (N_47087,N_44805,N_45959);
nor U47088 (N_47088,N_45063,N_45240);
nand U47089 (N_47089,N_44039,N_44657);
nand U47090 (N_47090,N_44294,N_45005);
xnor U47091 (N_47091,N_44545,N_44866);
xor U47092 (N_47092,N_45891,N_45988);
and U47093 (N_47093,N_44387,N_45620);
xnor U47094 (N_47094,N_44901,N_44212);
or U47095 (N_47095,N_44979,N_45661);
and U47096 (N_47096,N_45940,N_44537);
nand U47097 (N_47097,N_44259,N_45097);
xnor U47098 (N_47098,N_44137,N_44264);
or U47099 (N_47099,N_44852,N_45550);
or U47100 (N_47100,N_45707,N_45804);
and U47101 (N_47101,N_45390,N_45497);
xor U47102 (N_47102,N_44364,N_45389);
or U47103 (N_47103,N_45024,N_45198);
nand U47104 (N_47104,N_45941,N_44041);
and U47105 (N_47105,N_45860,N_44189);
or U47106 (N_47106,N_44967,N_44958);
nor U47107 (N_47107,N_45370,N_44884);
nor U47108 (N_47108,N_44767,N_45996);
xnor U47109 (N_47109,N_45635,N_45588);
or U47110 (N_47110,N_44807,N_45289);
and U47111 (N_47111,N_44521,N_45010);
nor U47112 (N_47112,N_45961,N_45130);
xor U47113 (N_47113,N_45194,N_44723);
or U47114 (N_47114,N_44591,N_45301);
nand U47115 (N_47115,N_44009,N_44925);
and U47116 (N_47116,N_44679,N_44590);
and U47117 (N_47117,N_45168,N_45506);
nor U47118 (N_47118,N_44970,N_44940);
nand U47119 (N_47119,N_45473,N_45557);
xor U47120 (N_47120,N_44054,N_45400);
and U47121 (N_47121,N_45802,N_44270);
nand U47122 (N_47122,N_45541,N_44200);
or U47123 (N_47123,N_45339,N_44188);
nor U47124 (N_47124,N_45794,N_45581);
and U47125 (N_47125,N_44744,N_44557);
or U47126 (N_47126,N_44626,N_45913);
nor U47127 (N_47127,N_44316,N_44229);
and U47128 (N_47128,N_45360,N_45650);
and U47129 (N_47129,N_44752,N_44286);
nand U47130 (N_47130,N_45019,N_45797);
nor U47131 (N_47131,N_45719,N_44434);
and U47132 (N_47132,N_45356,N_44734);
xor U47133 (N_47133,N_44603,N_44154);
and U47134 (N_47134,N_45355,N_44430);
xor U47135 (N_47135,N_44527,N_44485);
xor U47136 (N_47136,N_44545,N_44651);
xnor U47137 (N_47137,N_45303,N_44433);
nor U47138 (N_47138,N_45428,N_44507);
or U47139 (N_47139,N_45039,N_44326);
nand U47140 (N_47140,N_45403,N_45112);
nor U47141 (N_47141,N_44697,N_45445);
nand U47142 (N_47142,N_45363,N_44455);
or U47143 (N_47143,N_44599,N_45498);
and U47144 (N_47144,N_45840,N_44576);
nand U47145 (N_47145,N_44048,N_44880);
and U47146 (N_47146,N_45839,N_44657);
or U47147 (N_47147,N_44166,N_44595);
nor U47148 (N_47148,N_45962,N_44603);
and U47149 (N_47149,N_44166,N_44107);
and U47150 (N_47150,N_45711,N_44897);
nand U47151 (N_47151,N_45525,N_44451);
nand U47152 (N_47152,N_45813,N_45506);
nand U47153 (N_47153,N_45821,N_45516);
or U47154 (N_47154,N_45039,N_45029);
or U47155 (N_47155,N_44014,N_45541);
nand U47156 (N_47156,N_44354,N_45467);
xnor U47157 (N_47157,N_44174,N_45671);
or U47158 (N_47158,N_45468,N_45151);
nand U47159 (N_47159,N_44461,N_45003);
nand U47160 (N_47160,N_45681,N_44069);
or U47161 (N_47161,N_45347,N_45377);
nor U47162 (N_47162,N_44844,N_45124);
nand U47163 (N_47163,N_44495,N_44339);
and U47164 (N_47164,N_44673,N_44885);
and U47165 (N_47165,N_44011,N_45068);
xnor U47166 (N_47166,N_45961,N_45014);
or U47167 (N_47167,N_45379,N_44737);
nand U47168 (N_47168,N_44596,N_45769);
and U47169 (N_47169,N_44315,N_45414);
or U47170 (N_47170,N_44503,N_44528);
xor U47171 (N_47171,N_44616,N_44343);
xor U47172 (N_47172,N_44857,N_44737);
and U47173 (N_47173,N_44940,N_44926);
xnor U47174 (N_47174,N_44929,N_44418);
nor U47175 (N_47175,N_45747,N_45958);
and U47176 (N_47176,N_44981,N_44685);
or U47177 (N_47177,N_45548,N_44533);
and U47178 (N_47178,N_45599,N_44815);
nand U47179 (N_47179,N_44160,N_44062);
xnor U47180 (N_47180,N_44931,N_44555);
and U47181 (N_47181,N_45073,N_45928);
or U47182 (N_47182,N_45037,N_44723);
or U47183 (N_47183,N_44074,N_45363);
or U47184 (N_47184,N_45647,N_44832);
xnor U47185 (N_47185,N_45381,N_45044);
xor U47186 (N_47186,N_45015,N_45083);
nand U47187 (N_47187,N_44869,N_45142);
xnor U47188 (N_47188,N_45701,N_45812);
nand U47189 (N_47189,N_44329,N_45830);
nor U47190 (N_47190,N_45287,N_45372);
nor U47191 (N_47191,N_44023,N_45379);
or U47192 (N_47192,N_45976,N_44216);
nand U47193 (N_47193,N_45873,N_44018);
xor U47194 (N_47194,N_44871,N_44997);
xnor U47195 (N_47195,N_45457,N_44281);
or U47196 (N_47196,N_44535,N_44104);
or U47197 (N_47197,N_45023,N_45722);
nor U47198 (N_47198,N_44964,N_45681);
xnor U47199 (N_47199,N_45408,N_45779);
xnor U47200 (N_47200,N_45730,N_44753);
nor U47201 (N_47201,N_45899,N_44752);
nand U47202 (N_47202,N_44389,N_45640);
or U47203 (N_47203,N_45946,N_45109);
xnor U47204 (N_47204,N_45866,N_44659);
nor U47205 (N_47205,N_44331,N_44637);
nor U47206 (N_47206,N_44331,N_45257);
xnor U47207 (N_47207,N_44954,N_44300);
nand U47208 (N_47208,N_44079,N_45469);
xor U47209 (N_47209,N_45867,N_45539);
and U47210 (N_47210,N_44876,N_45832);
xor U47211 (N_47211,N_45920,N_44064);
nand U47212 (N_47212,N_45852,N_45219);
nand U47213 (N_47213,N_44871,N_45356);
or U47214 (N_47214,N_45444,N_44172);
xor U47215 (N_47215,N_44550,N_44687);
nor U47216 (N_47216,N_45693,N_44549);
xnor U47217 (N_47217,N_45083,N_44887);
nor U47218 (N_47218,N_45533,N_44908);
nor U47219 (N_47219,N_44742,N_45014);
and U47220 (N_47220,N_44816,N_45347);
nor U47221 (N_47221,N_44711,N_44607);
nand U47222 (N_47222,N_44909,N_45442);
nand U47223 (N_47223,N_45586,N_44713);
nor U47224 (N_47224,N_44625,N_44388);
xor U47225 (N_47225,N_45492,N_45647);
nor U47226 (N_47226,N_45853,N_44077);
or U47227 (N_47227,N_45766,N_44543);
or U47228 (N_47228,N_45509,N_45459);
nor U47229 (N_47229,N_45567,N_45301);
nor U47230 (N_47230,N_44653,N_45730);
or U47231 (N_47231,N_45132,N_45429);
nor U47232 (N_47232,N_44208,N_45281);
or U47233 (N_47233,N_45664,N_44794);
nor U47234 (N_47234,N_45189,N_44343);
or U47235 (N_47235,N_44979,N_45880);
nor U47236 (N_47236,N_44531,N_45669);
nand U47237 (N_47237,N_45246,N_45103);
and U47238 (N_47238,N_44982,N_45549);
or U47239 (N_47239,N_45651,N_45749);
nand U47240 (N_47240,N_45326,N_45799);
nor U47241 (N_47241,N_44937,N_44204);
xor U47242 (N_47242,N_45370,N_44177);
and U47243 (N_47243,N_45201,N_45027);
xor U47244 (N_47244,N_45572,N_45730);
nand U47245 (N_47245,N_44935,N_45384);
or U47246 (N_47246,N_44259,N_45945);
or U47247 (N_47247,N_45719,N_45430);
nand U47248 (N_47248,N_44194,N_45975);
nor U47249 (N_47249,N_45402,N_44210);
or U47250 (N_47250,N_44249,N_44845);
xnor U47251 (N_47251,N_45341,N_44102);
or U47252 (N_47252,N_45825,N_45262);
nand U47253 (N_47253,N_45268,N_44978);
xnor U47254 (N_47254,N_45804,N_44684);
and U47255 (N_47255,N_45327,N_45810);
and U47256 (N_47256,N_45100,N_45514);
xor U47257 (N_47257,N_44241,N_44910);
nand U47258 (N_47258,N_45597,N_45300);
xor U47259 (N_47259,N_44582,N_44018);
xor U47260 (N_47260,N_45039,N_44033);
or U47261 (N_47261,N_44114,N_44689);
or U47262 (N_47262,N_44246,N_45659);
xor U47263 (N_47263,N_45501,N_44286);
nor U47264 (N_47264,N_44918,N_45958);
nand U47265 (N_47265,N_45410,N_44797);
or U47266 (N_47266,N_44249,N_45408);
or U47267 (N_47267,N_44461,N_45409);
nand U47268 (N_47268,N_45293,N_44172);
nand U47269 (N_47269,N_45434,N_45265);
and U47270 (N_47270,N_45852,N_44377);
or U47271 (N_47271,N_45777,N_44930);
xnor U47272 (N_47272,N_44852,N_45539);
nor U47273 (N_47273,N_44801,N_44699);
xnor U47274 (N_47274,N_45213,N_44191);
nand U47275 (N_47275,N_45606,N_45201);
nand U47276 (N_47276,N_44901,N_44887);
or U47277 (N_47277,N_44445,N_45922);
or U47278 (N_47278,N_44799,N_44277);
nand U47279 (N_47279,N_44901,N_44545);
nor U47280 (N_47280,N_44195,N_44269);
or U47281 (N_47281,N_45807,N_44448);
or U47282 (N_47282,N_45125,N_45382);
and U47283 (N_47283,N_45251,N_45519);
nand U47284 (N_47284,N_44989,N_45572);
or U47285 (N_47285,N_45044,N_45814);
or U47286 (N_47286,N_44844,N_45987);
nand U47287 (N_47287,N_44535,N_44314);
nand U47288 (N_47288,N_45875,N_44542);
xnor U47289 (N_47289,N_44713,N_45217);
nor U47290 (N_47290,N_45798,N_45119);
nand U47291 (N_47291,N_45981,N_44960);
and U47292 (N_47292,N_44572,N_44618);
nor U47293 (N_47293,N_44681,N_45182);
or U47294 (N_47294,N_45082,N_44282);
nor U47295 (N_47295,N_44996,N_44671);
or U47296 (N_47296,N_45144,N_45594);
xnor U47297 (N_47297,N_45286,N_45518);
xnor U47298 (N_47298,N_45467,N_45401);
and U47299 (N_47299,N_45339,N_44590);
xor U47300 (N_47300,N_45467,N_45000);
or U47301 (N_47301,N_45696,N_44980);
nand U47302 (N_47302,N_44467,N_44312);
nand U47303 (N_47303,N_45612,N_44337);
or U47304 (N_47304,N_44276,N_45693);
or U47305 (N_47305,N_44927,N_44347);
nand U47306 (N_47306,N_45727,N_44953);
xnor U47307 (N_47307,N_44431,N_45888);
xnor U47308 (N_47308,N_44434,N_44897);
or U47309 (N_47309,N_44607,N_45950);
or U47310 (N_47310,N_45419,N_44986);
nor U47311 (N_47311,N_45703,N_45414);
and U47312 (N_47312,N_44787,N_44119);
xor U47313 (N_47313,N_44418,N_45813);
nor U47314 (N_47314,N_44756,N_45579);
nor U47315 (N_47315,N_45826,N_44605);
and U47316 (N_47316,N_44874,N_44305);
nor U47317 (N_47317,N_45935,N_45222);
and U47318 (N_47318,N_44558,N_45311);
nand U47319 (N_47319,N_45903,N_45808);
or U47320 (N_47320,N_44573,N_45118);
nand U47321 (N_47321,N_44380,N_45099);
and U47322 (N_47322,N_45010,N_45133);
and U47323 (N_47323,N_44363,N_44385);
and U47324 (N_47324,N_45431,N_45517);
nor U47325 (N_47325,N_45852,N_44852);
xor U47326 (N_47326,N_44762,N_44694);
xor U47327 (N_47327,N_45089,N_45592);
and U47328 (N_47328,N_44057,N_44491);
and U47329 (N_47329,N_45373,N_45096);
xnor U47330 (N_47330,N_45747,N_45482);
nor U47331 (N_47331,N_45758,N_44998);
and U47332 (N_47332,N_45848,N_45496);
xnor U47333 (N_47333,N_44573,N_45802);
nand U47334 (N_47334,N_44077,N_45586);
nor U47335 (N_47335,N_45926,N_44691);
nor U47336 (N_47336,N_45137,N_44807);
nor U47337 (N_47337,N_45102,N_45676);
or U47338 (N_47338,N_44952,N_44263);
or U47339 (N_47339,N_44161,N_45639);
and U47340 (N_47340,N_45590,N_44408);
nand U47341 (N_47341,N_45191,N_44740);
or U47342 (N_47342,N_44089,N_45305);
or U47343 (N_47343,N_44327,N_44407);
xnor U47344 (N_47344,N_45131,N_45173);
and U47345 (N_47345,N_44646,N_45767);
nand U47346 (N_47346,N_44391,N_45165);
nand U47347 (N_47347,N_45750,N_45195);
or U47348 (N_47348,N_45152,N_44333);
nand U47349 (N_47349,N_44209,N_45688);
nor U47350 (N_47350,N_45318,N_45029);
nand U47351 (N_47351,N_44905,N_44217);
xnor U47352 (N_47352,N_45305,N_44553);
nor U47353 (N_47353,N_45768,N_44325);
and U47354 (N_47354,N_44358,N_44657);
nor U47355 (N_47355,N_45696,N_45364);
nor U47356 (N_47356,N_45177,N_45828);
and U47357 (N_47357,N_45759,N_44449);
nor U47358 (N_47358,N_44072,N_44568);
xnor U47359 (N_47359,N_45144,N_45434);
nand U47360 (N_47360,N_45920,N_45812);
xor U47361 (N_47361,N_44342,N_44494);
and U47362 (N_47362,N_45648,N_45755);
or U47363 (N_47363,N_45608,N_44347);
or U47364 (N_47364,N_45910,N_44811);
and U47365 (N_47365,N_45310,N_44514);
and U47366 (N_47366,N_44023,N_45154);
nand U47367 (N_47367,N_44935,N_44528);
or U47368 (N_47368,N_44190,N_44788);
nand U47369 (N_47369,N_44547,N_44721);
nor U47370 (N_47370,N_44774,N_45322);
or U47371 (N_47371,N_44407,N_45179);
nor U47372 (N_47372,N_45258,N_45223);
and U47373 (N_47373,N_44694,N_45527);
nand U47374 (N_47374,N_45560,N_44821);
nand U47375 (N_47375,N_44994,N_45066);
nor U47376 (N_47376,N_45508,N_44232);
xor U47377 (N_47377,N_45463,N_44150);
or U47378 (N_47378,N_44425,N_44989);
nor U47379 (N_47379,N_44293,N_45634);
nand U47380 (N_47380,N_45307,N_45164);
nor U47381 (N_47381,N_45260,N_45785);
and U47382 (N_47382,N_45237,N_44392);
and U47383 (N_47383,N_44508,N_45373);
and U47384 (N_47384,N_45130,N_44922);
xnor U47385 (N_47385,N_44539,N_44890);
or U47386 (N_47386,N_44451,N_45950);
nand U47387 (N_47387,N_45193,N_45179);
nand U47388 (N_47388,N_44558,N_44315);
xnor U47389 (N_47389,N_45162,N_44727);
nand U47390 (N_47390,N_44610,N_44419);
nand U47391 (N_47391,N_45628,N_45047);
or U47392 (N_47392,N_45978,N_44210);
nor U47393 (N_47393,N_44251,N_44750);
xnor U47394 (N_47394,N_44026,N_45996);
and U47395 (N_47395,N_45467,N_44511);
nor U47396 (N_47396,N_44647,N_45573);
nand U47397 (N_47397,N_45942,N_44175);
and U47398 (N_47398,N_45370,N_44510);
nor U47399 (N_47399,N_45149,N_45320);
nor U47400 (N_47400,N_45084,N_45225);
nand U47401 (N_47401,N_45980,N_44805);
and U47402 (N_47402,N_44830,N_45596);
and U47403 (N_47403,N_45049,N_45206);
nand U47404 (N_47404,N_44900,N_44754);
or U47405 (N_47405,N_44348,N_45787);
and U47406 (N_47406,N_44644,N_44445);
or U47407 (N_47407,N_45243,N_45603);
xnor U47408 (N_47408,N_44885,N_45746);
or U47409 (N_47409,N_44064,N_44417);
nor U47410 (N_47410,N_45630,N_44748);
and U47411 (N_47411,N_44515,N_44064);
xnor U47412 (N_47412,N_45586,N_45339);
nand U47413 (N_47413,N_44955,N_45610);
nor U47414 (N_47414,N_45964,N_45888);
nor U47415 (N_47415,N_44930,N_45364);
nand U47416 (N_47416,N_45131,N_45034);
and U47417 (N_47417,N_44203,N_44182);
nor U47418 (N_47418,N_45755,N_45705);
nand U47419 (N_47419,N_44181,N_44737);
nand U47420 (N_47420,N_45316,N_44272);
nand U47421 (N_47421,N_45707,N_45320);
xnor U47422 (N_47422,N_44890,N_44626);
or U47423 (N_47423,N_44826,N_44415);
nor U47424 (N_47424,N_44857,N_44282);
nand U47425 (N_47425,N_45849,N_45600);
nand U47426 (N_47426,N_44978,N_45508);
nor U47427 (N_47427,N_45705,N_44902);
nand U47428 (N_47428,N_44991,N_44475);
nand U47429 (N_47429,N_44875,N_44346);
nand U47430 (N_47430,N_44609,N_45511);
xnor U47431 (N_47431,N_45244,N_45279);
nand U47432 (N_47432,N_45835,N_45385);
and U47433 (N_47433,N_44396,N_45345);
or U47434 (N_47434,N_44497,N_45682);
and U47435 (N_47435,N_44483,N_44165);
nor U47436 (N_47436,N_45400,N_45499);
or U47437 (N_47437,N_45245,N_44353);
and U47438 (N_47438,N_44106,N_44502);
nor U47439 (N_47439,N_44662,N_45723);
or U47440 (N_47440,N_44336,N_44249);
and U47441 (N_47441,N_45749,N_45338);
nand U47442 (N_47442,N_45393,N_44742);
and U47443 (N_47443,N_44991,N_45198);
nand U47444 (N_47444,N_44005,N_44033);
nor U47445 (N_47445,N_44656,N_44661);
nand U47446 (N_47446,N_45818,N_44604);
nor U47447 (N_47447,N_45062,N_44958);
and U47448 (N_47448,N_44496,N_44726);
and U47449 (N_47449,N_44260,N_45628);
nand U47450 (N_47450,N_44646,N_44309);
or U47451 (N_47451,N_44124,N_45790);
xnor U47452 (N_47452,N_44537,N_45849);
and U47453 (N_47453,N_44820,N_44307);
and U47454 (N_47454,N_44107,N_45831);
xnor U47455 (N_47455,N_45300,N_45808);
nor U47456 (N_47456,N_44524,N_45715);
xor U47457 (N_47457,N_44752,N_44536);
nand U47458 (N_47458,N_45506,N_44044);
xor U47459 (N_47459,N_44992,N_45079);
nor U47460 (N_47460,N_45290,N_44372);
or U47461 (N_47461,N_44563,N_45735);
nand U47462 (N_47462,N_44686,N_45514);
and U47463 (N_47463,N_45728,N_44194);
nor U47464 (N_47464,N_44722,N_45657);
and U47465 (N_47465,N_44219,N_45862);
nand U47466 (N_47466,N_45069,N_44792);
nor U47467 (N_47467,N_44911,N_45056);
or U47468 (N_47468,N_44075,N_44790);
nand U47469 (N_47469,N_45379,N_45773);
and U47470 (N_47470,N_45243,N_44579);
nand U47471 (N_47471,N_44297,N_45349);
nor U47472 (N_47472,N_45795,N_45977);
and U47473 (N_47473,N_44471,N_44270);
nor U47474 (N_47474,N_44026,N_45148);
xnor U47475 (N_47475,N_44695,N_45632);
and U47476 (N_47476,N_45358,N_44953);
and U47477 (N_47477,N_45324,N_44843);
or U47478 (N_47478,N_44522,N_45656);
xor U47479 (N_47479,N_44279,N_44335);
nand U47480 (N_47480,N_45071,N_45487);
nand U47481 (N_47481,N_45663,N_44817);
and U47482 (N_47482,N_44185,N_44270);
nor U47483 (N_47483,N_45521,N_44869);
nor U47484 (N_47484,N_44995,N_44526);
nand U47485 (N_47485,N_45157,N_44486);
and U47486 (N_47486,N_45242,N_44047);
nor U47487 (N_47487,N_44136,N_44358);
or U47488 (N_47488,N_44164,N_44294);
xnor U47489 (N_47489,N_44372,N_44475);
nand U47490 (N_47490,N_44486,N_44883);
nand U47491 (N_47491,N_44618,N_45845);
and U47492 (N_47492,N_45378,N_45014);
or U47493 (N_47493,N_44863,N_45407);
nand U47494 (N_47494,N_44223,N_45439);
and U47495 (N_47495,N_44127,N_44976);
nand U47496 (N_47496,N_45375,N_45968);
and U47497 (N_47497,N_44580,N_45931);
nand U47498 (N_47498,N_45943,N_45582);
xor U47499 (N_47499,N_44492,N_45255);
nand U47500 (N_47500,N_45783,N_45544);
or U47501 (N_47501,N_45124,N_44988);
and U47502 (N_47502,N_45819,N_44186);
and U47503 (N_47503,N_44113,N_44706);
or U47504 (N_47504,N_45070,N_44771);
xor U47505 (N_47505,N_45128,N_44264);
xnor U47506 (N_47506,N_45996,N_45497);
or U47507 (N_47507,N_44605,N_45586);
nand U47508 (N_47508,N_44975,N_44963);
nand U47509 (N_47509,N_45344,N_45064);
or U47510 (N_47510,N_45135,N_45716);
nor U47511 (N_47511,N_45836,N_44142);
or U47512 (N_47512,N_44460,N_44862);
xnor U47513 (N_47513,N_45246,N_45660);
nor U47514 (N_47514,N_45535,N_44554);
and U47515 (N_47515,N_45251,N_45146);
or U47516 (N_47516,N_45757,N_44357);
xor U47517 (N_47517,N_44631,N_45899);
and U47518 (N_47518,N_45609,N_44770);
and U47519 (N_47519,N_45868,N_44218);
or U47520 (N_47520,N_44798,N_44930);
nand U47521 (N_47521,N_44622,N_45412);
xor U47522 (N_47522,N_44267,N_45645);
nand U47523 (N_47523,N_45867,N_45141);
xor U47524 (N_47524,N_45557,N_45326);
nand U47525 (N_47525,N_45133,N_44567);
nor U47526 (N_47526,N_44143,N_44850);
and U47527 (N_47527,N_45060,N_45314);
nor U47528 (N_47528,N_45072,N_45195);
xnor U47529 (N_47529,N_44366,N_44364);
nand U47530 (N_47530,N_44465,N_44450);
nand U47531 (N_47531,N_45161,N_45936);
nand U47532 (N_47532,N_44399,N_45278);
or U47533 (N_47533,N_45718,N_44550);
nand U47534 (N_47534,N_44302,N_45047);
nand U47535 (N_47535,N_44732,N_45771);
or U47536 (N_47536,N_45430,N_44084);
xnor U47537 (N_47537,N_45128,N_44113);
xor U47538 (N_47538,N_45616,N_45335);
or U47539 (N_47539,N_44767,N_45325);
nor U47540 (N_47540,N_44444,N_44691);
nor U47541 (N_47541,N_44423,N_44641);
nor U47542 (N_47542,N_45690,N_45867);
and U47543 (N_47543,N_45295,N_45251);
nand U47544 (N_47544,N_44148,N_44362);
nand U47545 (N_47545,N_45767,N_44328);
nor U47546 (N_47546,N_45113,N_44005);
and U47547 (N_47547,N_45062,N_45636);
or U47548 (N_47548,N_45274,N_45877);
and U47549 (N_47549,N_45681,N_44255);
or U47550 (N_47550,N_45429,N_45755);
and U47551 (N_47551,N_45635,N_44694);
and U47552 (N_47552,N_44141,N_44463);
nor U47553 (N_47553,N_44156,N_44909);
nor U47554 (N_47554,N_44314,N_45667);
and U47555 (N_47555,N_45951,N_44822);
nand U47556 (N_47556,N_45665,N_45167);
xor U47557 (N_47557,N_45137,N_45889);
nor U47558 (N_47558,N_45140,N_44758);
and U47559 (N_47559,N_45120,N_44675);
or U47560 (N_47560,N_45016,N_44544);
nand U47561 (N_47561,N_44413,N_44018);
xor U47562 (N_47562,N_45144,N_44159);
or U47563 (N_47563,N_44805,N_45536);
nand U47564 (N_47564,N_45166,N_44041);
nand U47565 (N_47565,N_45304,N_45887);
and U47566 (N_47566,N_45889,N_45863);
xnor U47567 (N_47567,N_44629,N_44031);
or U47568 (N_47568,N_45217,N_44778);
nand U47569 (N_47569,N_44851,N_45294);
xnor U47570 (N_47570,N_45505,N_44619);
nand U47571 (N_47571,N_44735,N_45328);
and U47572 (N_47572,N_45577,N_45029);
or U47573 (N_47573,N_44904,N_44166);
nand U47574 (N_47574,N_44265,N_44486);
nand U47575 (N_47575,N_44038,N_45755);
nand U47576 (N_47576,N_44059,N_45222);
xor U47577 (N_47577,N_45966,N_45069);
or U47578 (N_47578,N_45495,N_44992);
or U47579 (N_47579,N_44325,N_44060);
or U47580 (N_47580,N_44828,N_44942);
nor U47581 (N_47581,N_44488,N_44967);
nor U47582 (N_47582,N_45355,N_44834);
xnor U47583 (N_47583,N_45777,N_45999);
or U47584 (N_47584,N_44360,N_45319);
nor U47585 (N_47585,N_44228,N_45790);
or U47586 (N_47586,N_44725,N_45541);
and U47587 (N_47587,N_45577,N_44893);
nor U47588 (N_47588,N_45156,N_45843);
nor U47589 (N_47589,N_45999,N_45585);
xor U47590 (N_47590,N_45859,N_44795);
nand U47591 (N_47591,N_44070,N_45144);
and U47592 (N_47592,N_44017,N_44298);
and U47593 (N_47593,N_45545,N_45650);
xor U47594 (N_47594,N_45007,N_45126);
or U47595 (N_47595,N_44575,N_44299);
nor U47596 (N_47596,N_44629,N_44345);
nor U47597 (N_47597,N_45383,N_45899);
nand U47598 (N_47598,N_44179,N_44473);
and U47599 (N_47599,N_44013,N_45351);
nand U47600 (N_47600,N_44145,N_45756);
or U47601 (N_47601,N_45035,N_45027);
xnor U47602 (N_47602,N_44282,N_45653);
nand U47603 (N_47603,N_45282,N_45091);
nor U47604 (N_47604,N_45088,N_45803);
or U47605 (N_47605,N_45319,N_45146);
nand U47606 (N_47606,N_45596,N_45972);
or U47607 (N_47607,N_44036,N_45705);
xor U47608 (N_47608,N_44198,N_45819);
or U47609 (N_47609,N_44607,N_44946);
nor U47610 (N_47610,N_45307,N_45017);
or U47611 (N_47611,N_44853,N_45630);
and U47612 (N_47612,N_44101,N_44034);
or U47613 (N_47613,N_44704,N_45874);
nor U47614 (N_47614,N_45391,N_45300);
nand U47615 (N_47615,N_45762,N_45867);
or U47616 (N_47616,N_45435,N_45226);
and U47617 (N_47617,N_45045,N_44078);
nand U47618 (N_47618,N_44470,N_45301);
xnor U47619 (N_47619,N_45273,N_44898);
nor U47620 (N_47620,N_44161,N_44192);
nor U47621 (N_47621,N_45795,N_45926);
or U47622 (N_47622,N_44162,N_44315);
nor U47623 (N_47623,N_45430,N_44043);
and U47624 (N_47624,N_45350,N_44953);
and U47625 (N_47625,N_44912,N_44115);
or U47626 (N_47626,N_45088,N_45685);
nand U47627 (N_47627,N_44375,N_45802);
and U47628 (N_47628,N_44926,N_44624);
nand U47629 (N_47629,N_45647,N_45196);
xor U47630 (N_47630,N_45628,N_45145);
and U47631 (N_47631,N_45182,N_44676);
nor U47632 (N_47632,N_45970,N_44085);
nand U47633 (N_47633,N_44952,N_44157);
xnor U47634 (N_47634,N_45294,N_45638);
or U47635 (N_47635,N_45473,N_45405);
nor U47636 (N_47636,N_45042,N_44564);
and U47637 (N_47637,N_45387,N_44620);
nand U47638 (N_47638,N_44395,N_45055);
and U47639 (N_47639,N_45799,N_44313);
nand U47640 (N_47640,N_45124,N_44374);
xnor U47641 (N_47641,N_45036,N_45572);
xnor U47642 (N_47642,N_45459,N_44509);
or U47643 (N_47643,N_44877,N_44618);
or U47644 (N_47644,N_44575,N_44208);
xnor U47645 (N_47645,N_44449,N_44221);
and U47646 (N_47646,N_44077,N_45145);
nor U47647 (N_47647,N_44440,N_44010);
and U47648 (N_47648,N_45966,N_44936);
xnor U47649 (N_47649,N_44175,N_44790);
nand U47650 (N_47650,N_44406,N_45579);
nand U47651 (N_47651,N_44814,N_45676);
nor U47652 (N_47652,N_44433,N_44008);
xnor U47653 (N_47653,N_44850,N_45627);
nor U47654 (N_47654,N_45635,N_45027);
nor U47655 (N_47655,N_45329,N_44380);
nand U47656 (N_47656,N_45095,N_45029);
or U47657 (N_47657,N_44273,N_44901);
and U47658 (N_47658,N_44320,N_44717);
nand U47659 (N_47659,N_45595,N_44041);
nand U47660 (N_47660,N_44979,N_45558);
or U47661 (N_47661,N_44143,N_45993);
or U47662 (N_47662,N_44166,N_45230);
and U47663 (N_47663,N_44087,N_45270);
and U47664 (N_47664,N_45817,N_45622);
and U47665 (N_47665,N_45774,N_45986);
and U47666 (N_47666,N_45036,N_45759);
or U47667 (N_47667,N_45727,N_44907);
and U47668 (N_47668,N_44951,N_45959);
or U47669 (N_47669,N_44281,N_45455);
and U47670 (N_47670,N_45914,N_45645);
nor U47671 (N_47671,N_44767,N_44859);
and U47672 (N_47672,N_45196,N_45071);
xor U47673 (N_47673,N_44186,N_44796);
nor U47674 (N_47674,N_45195,N_44796);
or U47675 (N_47675,N_44882,N_44714);
nor U47676 (N_47676,N_45563,N_44385);
nor U47677 (N_47677,N_45149,N_44900);
nor U47678 (N_47678,N_45760,N_45670);
or U47679 (N_47679,N_44199,N_45936);
nor U47680 (N_47680,N_44835,N_45191);
and U47681 (N_47681,N_45023,N_44087);
xor U47682 (N_47682,N_45017,N_45234);
nand U47683 (N_47683,N_44163,N_45687);
xnor U47684 (N_47684,N_45975,N_44579);
and U47685 (N_47685,N_44313,N_45085);
xor U47686 (N_47686,N_44372,N_44134);
or U47687 (N_47687,N_45512,N_45004);
xnor U47688 (N_47688,N_44349,N_45196);
nand U47689 (N_47689,N_45513,N_44264);
nor U47690 (N_47690,N_45638,N_45941);
or U47691 (N_47691,N_44580,N_44961);
or U47692 (N_47692,N_44468,N_45134);
nand U47693 (N_47693,N_45563,N_44504);
and U47694 (N_47694,N_44744,N_44354);
xor U47695 (N_47695,N_44497,N_44619);
and U47696 (N_47696,N_44037,N_45775);
or U47697 (N_47697,N_44350,N_44424);
or U47698 (N_47698,N_45124,N_44483);
nand U47699 (N_47699,N_44250,N_44567);
nand U47700 (N_47700,N_44810,N_44015);
nand U47701 (N_47701,N_45191,N_44446);
xnor U47702 (N_47702,N_45840,N_45284);
nand U47703 (N_47703,N_44324,N_44554);
and U47704 (N_47704,N_45610,N_44410);
xor U47705 (N_47705,N_45690,N_44497);
or U47706 (N_47706,N_45485,N_45864);
nand U47707 (N_47707,N_44996,N_44333);
xnor U47708 (N_47708,N_45786,N_45868);
nand U47709 (N_47709,N_44659,N_44179);
nor U47710 (N_47710,N_45098,N_44886);
or U47711 (N_47711,N_44056,N_44357);
nand U47712 (N_47712,N_45981,N_45960);
and U47713 (N_47713,N_45527,N_44271);
nor U47714 (N_47714,N_45540,N_45951);
and U47715 (N_47715,N_45941,N_44168);
and U47716 (N_47716,N_45492,N_45963);
nor U47717 (N_47717,N_45363,N_44316);
nand U47718 (N_47718,N_45235,N_45861);
and U47719 (N_47719,N_44897,N_44054);
nor U47720 (N_47720,N_44001,N_45268);
xor U47721 (N_47721,N_44454,N_44214);
nand U47722 (N_47722,N_44637,N_45747);
nand U47723 (N_47723,N_44232,N_45211);
and U47724 (N_47724,N_45494,N_44742);
and U47725 (N_47725,N_44444,N_44579);
and U47726 (N_47726,N_44023,N_44392);
and U47727 (N_47727,N_45935,N_44399);
xor U47728 (N_47728,N_44940,N_45095);
xnor U47729 (N_47729,N_44981,N_44585);
or U47730 (N_47730,N_44402,N_45232);
xnor U47731 (N_47731,N_45981,N_44076);
xnor U47732 (N_47732,N_45233,N_45439);
nand U47733 (N_47733,N_45566,N_44560);
or U47734 (N_47734,N_44912,N_45576);
xnor U47735 (N_47735,N_44841,N_44255);
and U47736 (N_47736,N_45565,N_45166);
nand U47737 (N_47737,N_45019,N_45923);
xnor U47738 (N_47738,N_44127,N_44346);
nand U47739 (N_47739,N_44614,N_45667);
or U47740 (N_47740,N_44999,N_45116);
nor U47741 (N_47741,N_44541,N_45093);
nor U47742 (N_47742,N_44644,N_45002);
nand U47743 (N_47743,N_45194,N_44616);
or U47744 (N_47744,N_44262,N_45822);
nand U47745 (N_47745,N_44902,N_45936);
or U47746 (N_47746,N_44392,N_45589);
or U47747 (N_47747,N_44577,N_44859);
or U47748 (N_47748,N_45633,N_45321);
and U47749 (N_47749,N_45675,N_44042);
nand U47750 (N_47750,N_44402,N_44183);
xnor U47751 (N_47751,N_44816,N_44840);
xor U47752 (N_47752,N_45814,N_45099);
and U47753 (N_47753,N_45039,N_44579);
or U47754 (N_47754,N_44096,N_45307);
or U47755 (N_47755,N_45913,N_45230);
nor U47756 (N_47756,N_44926,N_45534);
xor U47757 (N_47757,N_44628,N_44762);
nand U47758 (N_47758,N_45583,N_45134);
xnor U47759 (N_47759,N_45141,N_44267);
nor U47760 (N_47760,N_44804,N_45345);
nand U47761 (N_47761,N_44154,N_44552);
or U47762 (N_47762,N_44503,N_44161);
and U47763 (N_47763,N_45121,N_45791);
and U47764 (N_47764,N_45034,N_45890);
nor U47765 (N_47765,N_44244,N_44807);
and U47766 (N_47766,N_44370,N_44687);
nor U47767 (N_47767,N_45209,N_44817);
nor U47768 (N_47768,N_44109,N_45512);
and U47769 (N_47769,N_44561,N_45238);
and U47770 (N_47770,N_45874,N_44976);
or U47771 (N_47771,N_44229,N_45802);
nor U47772 (N_47772,N_44648,N_44267);
or U47773 (N_47773,N_45949,N_45750);
and U47774 (N_47774,N_45399,N_44486);
nand U47775 (N_47775,N_45327,N_45343);
nand U47776 (N_47776,N_44362,N_45936);
nor U47777 (N_47777,N_44278,N_44916);
xor U47778 (N_47778,N_45362,N_44599);
nor U47779 (N_47779,N_45584,N_45863);
and U47780 (N_47780,N_45071,N_45942);
nand U47781 (N_47781,N_45137,N_44748);
or U47782 (N_47782,N_45852,N_45027);
xor U47783 (N_47783,N_45637,N_44526);
nand U47784 (N_47784,N_45065,N_44336);
xnor U47785 (N_47785,N_44015,N_44808);
nor U47786 (N_47786,N_45445,N_44932);
nand U47787 (N_47787,N_44039,N_44341);
xor U47788 (N_47788,N_45816,N_44791);
and U47789 (N_47789,N_44411,N_45726);
nand U47790 (N_47790,N_44026,N_45907);
xnor U47791 (N_47791,N_44135,N_44913);
or U47792 (N_47792,N_45423,N_44032);
and U47793 (N_47793,N_44956,N_45034);
nor U47794 (N_47794,N_45788,N_44897);
nor U47795 (N_47795,N_45021,N_44021);
and U47796 (N_47796,N_45368,N_44746);
xnor U47797 (N_47797,N_44029,N_44345);
or U47798 (N_47798,N_45926,N_44892);
or U47799 (N_47799,N_45896,N_45930);
nand U47800 (N_47800,N_44475,N_44146);
nand U47801 (N_47801,N_45632,N_44143);
xor U47802 (N_47802,N_44678,N_44606);
and U47803 (N_47803,N_44028,N_44772);
nor U47804 (N_47804,N_45662,N_44609);
nand U47805 (N_47805,N_45121,N_45013);
or U47806 (N_47806,N_44892,N_45472);
xor U47807 (N_47807,N_44123,N_45191);
nand U47808 (N_47808,N_45504,N_45556);
nand U47809 (N_47809,N_45257,N_44975);
nand U47810 (N_47810,N_44608,N_44876);
and U47811 (N_47811,N_45067,N_44013);
and U47812 (N_47812,N_45734,N_45394);
and U47813 (N_47813,N_45138,N_44347);
nor U47814 (N_47814,N_45102,N_45072);
or U47815 (N_47815,N_44045,N_44687);
xor U47816 (N_47816,N_45253,N_45021);
and U47817 (N_47817,N_44564,N_45757);
xnor U47818 (N_47818,N_45901,N_44704);
or U47819 (N_47819,N_45146,N_45991);
and U47820 (N_47820,N_44553,N_44539);
xor U47821 (N_47821,N_44346,N_45731);
and U47822 (N_47822,N_45701,N_44531);
xor U47823 (N_47823,N_44847,N_44868);
xnor U47824 (N_47824,N_44386,N_44095);
and U47825 (N_47825,N_45875,N_44889);
nor U47826 (N_47826,N_45503,N_44571);
nand U47827 (N_47827,N_44352,N_44656);
and U47828 (N_47828,N_44280,N_44318);
nor U47829 (N_47829,N_45156,N_44828);
or U47830 (N_47830,N_44910,N_45264);
nand U47831 (N_47831,N_45259,N_44374);
nor U47832 (N_47832,N_44757,N_44158);
xnor U47833 (N_47833,N_45793,N_44009);
and U47834 (N_47834,N_45471,N_44406);
xnor U47835 (N_47835,N_44423,N_44382);
nand U47836 (N_47836,N_44296,N_45192);
or U47837 (N_47837,N_44259,N_44219);
or U47838 (N_47838,N_44862,N_45485);
xnor U47839 (N_47839,N_44677,N_44870);
and U47840 (N_47840,N_44120,N_44099);
nand U47841 (N_47841,N_45618,N_45517);
xnor U47842 (N_47842,N_44225,N_44400);
or U47843 (N_47843,N_44796,N_45872);
nand U47844 (N_47844,N_45565,N_44354);
and U47845 (N_47845,N_44610,N_44699);
and U47846 (N_47846,N_44139,N_45277);
xor U47847 (N_47847,N_44159,N_45620);
nand U47848 (N_47848,N_45342,N_44469);
or U47849 (N_47849,N_44409,N_45394);
nand U47850 (N_47850,N_45177,N_45960);
nand U47851 (N_47851,N_44539,N_44242);
xnor U47852 (N_47852,N_44085,N_45135);
nor U47853 (N_47853,N_44439,N_44143);
nand U47854 (N_47854,N_44504,N_44394);
nor U47855 (N_47855,N_44665,N_44060);
nand U47856 (N_47856,N_45103,N_45455);
or U47857 (N_47857,N_44988,N_45438);
xnor U47858 (N_47858,N_45206,N_44880);
or U47859 (N_47859,N_45905,N_44760);
nand U47860 (N_47860,N_45041,N_44919);
nor U47861 (N_47861,N_44988,N_44533);
and U47862 (N_47862,N_44353,N_45178);
xor U47863 (N_47863,N_44303,N_44913);
and U47864 (N_47864,N_44493,N_45401);
nor U47865 (N_47865,N_44299,N_45101);
nand U47866 (N_47866,N_44989,N_44217);
nor U47867 (N_47867,N_44436,N_44343);
and U47868 (N_47868,N_44631,N_44197);
or U47869 (N_47869,N_45575,N_45217);
or U47870 (N_47870,N_44231,N_44087);
nand U47871 (N_47871,N_45329,N_44997);
nand U47872 (N_47872,N_45804,N_44192);
or U47873 (N_47873,N_45459,N_44595);
or U47874 (N_47874,N_44959,N_45266);
xnor U47875 (N_47875,N_44115,N_45038);
nand U47876 (N_47876,N_44845,N_44705);
nor U47877 (N_47877,N_44248,N_45004);
xor U47878 (N_47878,N_44848,N_45714);
nand U47879 (N_47879,N_45939,N_45003);
nand U47880 (N_47880,N_44610,N_44014);
xor U47881 (N_47881,N_44906,N_44330);
nor U47882 (N_47882,N_44544,N_44545);
nand U47883 (N_47883,N_45230,N_44533);
nand U47884 (N_47884,N_44597,N_44906);
and U47885 (N_47885,N_45138,N_45333);
and U47886 (N_47886,N_45428,N_44347);
nor U47887 (N_47887,N_44475,N_45879);
or U47888 (N_47888,N_44432,N_44461);
nand U47889 (N_47889,N_44591,N_45978);
and U47890 (N_47890,N_44697,N_45425);
and U47891 (N_47891,N_45789,N_44795);
or U47892 (N_47892,N_44492,N_44605);
xor U47893 (N_47893,N_44382,N_44038);
xor U47894 (N_47894,N_44409,N_45419);
nand U47895 (N_47895,N_45870,N_44278);
xnor U47896 (N_47896,N_45729,N_44678);
and U47897 (N_47897,N_44964,N_45238);
nand U47898 (N_47898,N_45461,N_45142);
nand U47899 (N_47899,N_45480,N_45511);
nand U47900 (N_47900,N_45528,N_45052);
nor U47901 (N_47901,N_44545,N_45238);
nand U47902 (N_47902,N_44594,N_44094);
and U47903 (N_47903,N_44949,N_44813);
or U47904 (N_47904,N_45493,N_44572);
and U47905 (N_47905,N_44834,N_44433);
nand U47906 (N_47906,N_44092,N_44741);
or U47907 (N_47907,N_44606,N_44457);
or U47908 (N_47908,N_44260,N_45019);
nand U47909 (N_47909,N_45900,N_44469);
or U47910 (N_47910,N_45029,N_45393);
or U47911 (N_47911,N_45087,N_44215);
nand U47912 (N_47912,N_44151,N_44707);
or U47913 (N_47913,N_45115,N_45344);
and U47914 (N_47914,N_44368,N_44884);
nand U47915 (N_47915,N_45283,N_44086);
or U47916 (N_47916,N_45964,N_45780);
nand U47917 (N_47917,N_44598,N_45523);
nand U47918 (N_47918,N_44774,N_44933);
nor U47919 (N_47919,N_45279,N_45966);
xnor U47920 (N_47920,N_44817,N_45180);
nor U47921 (N_47921,N_45749,N_44274);
and U47922 (N_47922,N_44503,N_44633);
and U47923 (N_47923,N_45020,N_44979);
xnor U47924 (N_47924,N_45672,N_44973);
and U47925 (N_47925,N_44724,N_44489);
xnor U47926 (N_47926,N_45095,N_44284);
nor U47927 (N_47927,N_44813,N_44265);
and U47928 (N_47928,N_45852,N_44959);
nor U47929 (N_47929,N_45572,N_44895);
or U47930 (N_47930,N_44881,N_45573);
and U47931 (N_47931,N_44309,N_44505);
nor U47932 (N_47932,N_44256,N_44630);
or U47933 (N_47933,N_44888,N_44036);
or U47934 (N_47934,N_45239,N_45897);
nor U47935 (N_47935,N_45408,N_45196);
nor U47936 (N_47936,N_45546,N_44714);
and U47937 (N_47937,N_45248,N_44096);
xnor U47938 (N_47938,N_44394,N_44573);
and U47939 (N_47939,N_44913,N_44131);
xnor U47940 (N_47940,N_44608,N_44620);
or U47941 (N_47941,N_45703,N_44959);
xnor U47942 (N_47942,N_45611,N_44086);
xor U47943 (N_47943,N_44067,N_44959);
or U47944 (N_47944,N_44491,N_44715);
nor U47945 (N_47945,N_45666,N_45979);
nand U47946 (N_47946,N_44091,N_45859);
and U47947 (N_47947,N_44726,N_44147);
nand U47948 (N_47948,N_44562,N_45031);
xor U47949 (N_47949,N_45547,N_44815);
and U47950 (N_47950,N_44304,N_45561);
nand U47951 (N_47951,N_45514,N_45621);
or U47952 (N_47952,N_45061,N_45711);
and U47953 (N_47953,N_45001,N_44564);
or U47954 (N_47954,N_44300,N_45293);
nor U47955 (N_47955,N_45351,N_45686);
xor U47956 (N_47956,N_44524,N_44256);
xor U47957 (N_47957,N_44555,N_44425);
nand U47958 (N_47958,N_45473,N_44991);
nand U47959 (N_47959,N_45871,N_44056);
nand U47960 (N_47960,N_45276,N_45432);
and U47961 (N_47961,N_45941,N_44560);
nand U47962 (N_47962,N_45769,N_44503);
or U47963 (N_47963,N_44540,N_44209);
nand U47964 (N_47964,N_45944,N_45659);
and U47965 (N_47965,N_44566,N_45024);
or U47966 (N_47966,N_44100,N_45376);
nor U47967 (N_47967,N_45779,N_45493);
xor U47968 (N_47968,N_45386,N_44134);
and U47969 (N_47969,N_44522,N_45065);
or U47970 (N_47970,N_45735,N_44553);
or U47971 (N_47971,N_44889,N_44248);
and U47972 (N_47972,N_45825,N_45811);
and U47973 (N_47973,N_44595,N_44370);
and U47974 (N_47974,N_45172,N_45416);
and U47975 (N_47975,N_45464,N_45160);
and U47976 (N_47976,N_44498,N_44247);
xor U47977 (N_47977,N_44218,N_44961);
nor U47978 (N_47978,N_45250,N_44627);
xor U47979 (N_47979,N_44857,N_45052);
nor U47980 (N_47980,N_44202,N_44168);
xor U47981 (N_47981,N_45699,N_44165);
and U47982 (N_47982,N_45020,N_44127);
nor U47983 (N_47983,N_44769,N_45780);
nand U47984 (N_47984,N_45872,N_44611);
xor U47985 (N_47985,N_45780,N_44334);
xnor U47986 (N_47986,N_44209,N_45051);
xnor U47987 (N_47987,N_45151,N_45383);
xnor U47988 (N_47988,N_44433,N_45898);
and U47989 (N_47989,N_45072,N_45421);
nor U47990 (N_47990,N_45948,N_45876);
xor U47991 (N_47991,N_45391,N_44145);
or U47992 (N_47992,N_44056,N_44342);
nor U47993 (N_47993,N_45684,N_44711);
or U47994 (N_47994,N_44526,N_45372);
or U47995 (N_47995,N_45841,N_44714);
nand U47996 (N_47996,N_44554,N_44372);
xnor U47997 (N_47997,N_44630,N_45469);
and U47998 (N_47998,N_44330,N_44879);
nor U47999 (N_47999,N_44982,N_44767);
nor U48000 (N_48000,N_46435,N_46255);
or U48001 (N_48001,N_47488,N_47023);
nor U48002 (N_48002,N_47882,N_47081);
and U48003 (N_48003,N_46431,N_46711);
xor U48004 (N_48004,N_47096,N_47753);
nor U48005 (N_48005,N_47506,N_46437);
and U48006 (N_48006,N_46706,N_47251);
or U48007 (N_48007,N_46519,N_46951);
nor U48008 (N_48008,N_46566,N_47189);
or U48009 (N_48009,N_47627,N_46544);
nand U48010 (N_48010,N_47881,N_46683);
or U48011 (N_48011,N_46997,N_47870);
nand U48012 (N_48012,N_47325,N_47712);
and U48013 (N_48013,N_46295,N_47643);
and U48014 (N_48014,N_46841,N_47873);
nor U48015 (N_48015,N_47697,N_46629);
nand U48016 (N_48016,N_46491,N_47232);
and U48017 (N_48017,N_47938,N_47138);
and U48018 (N_48018,N_47581,N_47006);
xnor U48019 (N_48019,N_46622,N_47367);
or U48020 (N_48020,N_46274,N_47743);
and U48021 (N_48021,N_47310,N_46845);
xnor U48022 (N_48022,N_46085,N_47242);
nor U48023 (N_48023,N_46869,N_47534);
or U48024 (N_48024,N_46318,N_46773);
or U48025 (N_48025,N_47469,N_46385);
or U48026 (N_48026,N_46679,N_46176);
nor U48027 (N_48027,N_46228,N_46852);
or U48028 (N_48028,N_47767,N_46775);
xor U48029 (N_48029,N_46463,N_46363);
nor U48030 (N_48030,N_46858,N_47246);
xor U48031 (N_48031,N_47227,N_46734);
nand U48032 (N_48032,N_46304,N_47719);
nand U48033 (N_48033,N_47253,N_47164);
nor U48034 (N_48034,N_47760,N_47680);
xor U48035 (N_48035,N_46696,N_47048);
nor U48036 (N_48036,N_46210,N_47957);
or U48037 (N_48037,N_46292,N_47517);
and U48038 (N_48038,N_46795,N_46614);
xnor U48039 (N_48039,N_46698,N_47705);
nor U48040 (N_48040,N_47336,N_47306);
nor U48041 (N_48041,N_46344,N_46301);
or U48042 (N_48042,N_46330,N_46296);
or U48043 (N_48043,N_46727,N_47279);
nand U48044 (N_48044,N_47054,N_47405);
xor U48045 (N_48045,N_46461,N_46187);
xor U48046 (N_48046,N_46764,N_47772);
nand U48047 (N_48047,N_46045,N_46066);
and U48048 (N_48048,N_47004,N_47028);
nand U48049 (N_48049,N_47585,N_46827);
nand U48050 (N_48050,N_46032,N_47852);
nor U48051 (N_48051,N_46074,N_46523);
nand U48052 (N_48052,N_46139,N_46443);
nand U48053 (N_48053,N_47731,N_46648);
nor U48054 (N_48054,N_47612,N_47710);
or U48055 (N_48055,N_47777,N_46645);
or U48056 (N_48056,N_47039,N_47605);
or U48057 (N_48057,N_47747,N_46810);
nand U48058 (N_48058,N_47518,N_47036);
nand U48059 (N_48059,N_46597,N_46105);
nor U48060 (N_48060,N_47502,N_46678);
or U48061 (N_48061,N_47830,N_46005);
xor U48062 (N_48062,N_47298,N_47897);
xnor U48063 (N_48063,N_47713,N_47633);
xnor U48064 (N_48064,N_46901,N_47443);
nor U48065 (N_48065,N_47442,N_46140);
xnor U48066 (N_48066,N_46244,N_47959);
xor U48067 (N_48067,N_46427,N_47569);
nor U48068 (N_48068,N_46532,N_46320);
and U48069 (N_48069,N_46753,N_47451);
or U48070 (N_48070,N_46424,N_46023);
and U48071 (N_48071,N_47616,N_47821);
nor U48072 (N_48072,N_46536,N_46169);
nand U48073 (N_48073,N_46831,N_46932);
or U48074 (N_48074,N_46230,N_47171);
or U48075 (N_48075,N_47812,N_47018);
xnor U48076 (N_48076,N_46127,N_47920);
xnor U48077 (N_48077,N_46952,N_46580);
nor U48078 (N_48078,N_47807,N_47066);
or U48079 (N_48079,N_47464,N_46325);
nor U48080 (N_48080,N_46560,N_47531);
nor U48081 (N_48081,N_47218,N_46197);
xor U48082 (N_48082,N_47009,N_46028);
xor U48083 (N_48083,N_46910,N_46487);
nor U48084 (N_48084,N_47369,N_46546);
xor U48085 (N_48085,N_46259,N_46785);
nor U48086 (N_48086,N_47259,N_46986);
nor U48087 (N_48087,N_46989,N_46552);
xnor U48088 (N_48088,N_47343,N_46660);
and U48089 (N_48089,N_47528,N_47049);
or U48090 (N_48090,N_46243,N_47941);
nor U48091 (N_48091,N_46293,N_47472);
xnor U48092 (N_48092,N_47931,N_46843);
xnor U48093 (N_48093,N_46403,N_47780);
and U48094 (N_48094,N_46089,N_47674);
or U48095 (N_48095,N_46913,N_47571);
nand U48096 (N_48096,N_47149,N_46113);
nor U48097 (N_48097,N_46441,N_47480);
and U48098 (N_48098,N_46788,N_47094);
or U48099 (N_48099,N_46680,N_47683);
nand U48100 (N_48100,N_47085,N_47117);
and U48101 (N_48101,N_47474,N_46053);
xnor U48102 (N_48102,N_47965,N_46885);
nand U48103 (N_48103,N_47043,N_46490);
nand U48104 (N_48104,N_47435,N_46774);
or U48105 (N_48105,N_47623,N_47338);
nand U48106 (N_48106,N_46413,N_46149);
or U48107 (N_48107,N_47496,N_47476);
nand U48108 (N_48108,N_46075,N_47110);
nand U48109 (N_48109,N_47864,N_46218);
and U48110 (N_48110,N_46043,N_46505);
and U48111 (N_48111,N_47930,N_47078);
or U48112 (N_48112,N_46763,N_46656);
nand U48113 (N_48113,N_47391,N_46055);
and U48114 (N_48114,N_46836,N_46057);
and U48115 (N_48115,N_47204,N_46077);
and U48116 (N_48116,N_46368,N_46609);
and U48117 (N_48117,N_46486,N_46062);
or U48118 (N_48118,N_47748,N_46960);
and U48119 (N_48119,N_47077,N_47910);
and U48120 (N_48120,N_47255,N_47907);
xnor U48121 (N_48121,N_46954,N_47046);
xor U48122 (N_48122,N_47704,N_46452);
nor U48123 (N_48123,N_47254,N_46011);
and U48124 (N_48124,N_47814,N_47419);
and U48125 (N_48125,N_47217,N_46610);
nand U48126 (N_48126,N_47438,N_47083);
nor U48127 (N_48127,N_46496,N_47354);
or U48128 (N_48128,N_47877,N_47996);
nor U48129 (N_48129,N_46006,N_46022);
nor U48130 (N_48130,N_47459,N_46971);
and U48131 (N_48131,N_46762,N_46359);
xor U48132 (N_48132,N_47434,N_46959);
nand U48133 (N_48133,N_46334,N_46765);
and U48134 (N_48134,N_47590,N_47266);
and U48135 (N_48135,N_47188,N_46751);
nor U48136 (N_48136,N_47422,N_46829);
or U48137 (N_48137,N_47105,N_46094);
xnor U48138 (N_48138,N_47408,N_47762);
nor U48139 (N_48139,N_47535,N_47826);
nand U48140 (N_48140,N_47076,N_47484);
and U48141 (N_48141,N_47103,N_47655);
nor U48142 (N_48142,N_47221,N_47979);
or U48143 (N_48143,N_47681,N_47308);
or U48144 (N_48144,N_46002,N_47832);
nand U48145 (N_48145,N_47774,N_46111);
or U48146 (N_48146,N_46689,N_47113);
or U48147 (N_48147,N_46850,N_47545);
xor U48148 (N_48148,N_47170,N_47924);
or U48149 (N_48149,N_47328,N_47948);
xnor U48150 (N_48150,N_46444,N_47470);
xor U48151 (N_48151,N_47026,N_47498);
nor U48152 (N_48152,N_47027,N_46647);
nor U48153 (N_48153,N_47896,N_46256);
nand U48154 (N_48154,N_47178,N_46034);
and U48155 (N_48155,N_47257,N_47146);
or U48156 (N_48156,N_47387,N_46803);
nand U48157 (N_48157,N_46958,N_47904);
and U48158 (N_48158,N_46786,N_46950);
xnor U48159 (N_48159,N_46341,N_47406);
xnor U48160 (N_48160,N_46721,N_46746);
or U48161 (N_48161,N_46839,N_46524);
and U48162 (N_48162,N_46048,N_47234);
and U48163 (N_48163,N_46464,N_47166);
and U48164 (N_48164,N_47946,N_46020);
xor U48165 (N_48165,N_47603,N_47925);
nand U48166 (N_48166,N_47733,N_47879);
nand U48167 (N_48167,N_46134,N_47558);
nand U48168 (N_48168,N_47745,N_46927);
and U48169 (N_48169,N_47521,N_46287);
nand U48170 (N_48170,N_46966,N_46137);
and U48171 (N_48171,N_47566,N_46965);
nor U48172 (N_48172,N_47044,N_46429);
and U48173 (N_48173,N_47889,N_46088);
nand U48174 (N_48174,N_47417,N_47237);
nand U48175 (N_48175,N_46981,N_47557);
and U48176 (N_48176,N_47431,N_47143);
or U48177 (N_48177,N_46905,N_47876);
nor U48178 (N_48178,N_46453,N_47764);
or U48179 (N_48179,N_47332,N_46426);
nand U48180 (N_48180,N_47104,N_46970);
xor U48181 (N_48181,N_46717,N_46240);
nand U48182 (N_48182,N_47329,N_46151);
and U48183 (N_48183,N_47903,N_47766);
xnor U48184 (N_48184,N_47967,N_46940);
xnor U48185 (N_48185,N_47202,N_46015);
or U48186 (N_48186,N_46922,N_47447);
nor U48187 (N_48187,N_46097,N_47849);
xnor U48188 (N_48188,N_47144,N_47586);
xor U48189 (N_48189,N_47231,N_46783);
and U48190 (N_48190,N_47583,N_46107);
and U48191 (N_48191,N_47060,N_47124);
or U48192 (N_48192,N_47892,N_46818);
or U48193 (N_48193,N_47444,N_46136);
or U48194 (N_48194,N_47527,N_47019);
xor U48195 (N_48195,N_46608,N_47723);
nor U48196 (N_48196,N_46191,N_47159);
or U48197 (N_48197,N_46714,N_47185);
and U48198 (N_48198,N_46628,N_46733);
or U48199 (N_48199,N_46147,N_47000);
or U48200 (N_48200,N_46277,N_47454);
and U48201 (N_48201,N_47787,N_47993);
nor U48202 (N_48202,N_46939,N_47935);
nand U48203 (N_48203,N_46090,N_46216);
and U48204 (N_48204,N_46779,N_47005);
or U48205 (N_48205,N_47186,N_47837);
or U48206 (N_48206,N_47450,N_46564);
nor U48207 (N_48207,N_46931,N_46510);
and U48208 (N_48208,N_46572,N_46725);
and U48209 (N_48209,N_47779,N_47543);
nor U48210 (N_48210,N_46911,N_47089);
and U48211 (N_48211,N_46548,N_46348);
nand U48212 (N_48212,N_47515,N_46898);
nand U48213 (N_48213,N_47230,N_47548);
xnor U48214 (N_48214,N_46438,N_47858);
nand U48215 (N_48215,N_47183,N_47647);
xor U48216 (N_48216,N_46029,N_47030);
or U48217 (N_48217,N_46848,N_47735);
nand U48218 (N_48218,N_47510,N_47884);
and U48219 (N_48219,N_47906,N_46967);
xnor U48220 (N_48220,N_46578,N_47778);
or U48221 (N_48221,N_47715,N_47768);
and U48222 (N_48222,N_46367,N_47172);
or U48223 (N_48223,N_47269,N_46943);
nand U48224 (N_48224,N_47866,N_47639);
nor U48225 (N_48225,N_46484,N_46161);
nand U48226 (N_48226,N_47233,N_46157);
nand U48227 (N_48227,N_46881,N_46448);
nand U48228 (N_48228,N_47785,N_47642);
xor U48229 (N_48229,N_47148,N_46815);
xnor U48230 (N_48230,N_47592,N_46104);
xnor U48231 (N_48231,N_46709,N_46868);
and U48232 (N_48232,N_46719,N_46076);
nor U48233 (N_48233,N_46442,N_47716);
or U48234 (N_48234,N_46565,N_47372);
nand U48235 (N_48235,N_46875,N_46902);
and U48236 (N_48236,N_46518,N_47120);
nand U48237 (N_48237,N_47893,N_47669);
nand U48238 (N_48238,N_46313,N_46621);
xnor U48239 (N_48239,N_46419,N_47532);
nor U48240 (N_48240,N_46677,N_46808);
or U48241 (N_48241,N_46480,N_47071);
xnor U48242 (N_48242,N_46471,N_46623);
or U48243 (N_48243,N_47195,N_46878);
or U48244 (N_48244,N_47205,N_46364);
nand U48245 (N_48245,N_47694,N_47987);
or U48246 (N_48246,N_46846,N_47102);
xnor U48247 (N_48247,N_47667,N_46771);
nor U48248 (N_48248,N_46856,N_46106);
nor U48249 (N_48249,N_47839,N_47564);
nor U48250 (N_48250,N_46953,N_47756);
nand U48251 (N_48251,N_47173,N_47370);
or U48252 (N_48252,N_46099,N_46286);
and U48253 (N_48253,N_46477,N_47389);
and U48254 (N_48254,N_46498,N_46626);
xor U48255 (N_48255,N_46227,N_47657);
or U48256 (N_48256,N_47206,N_47074);
or U48257 (N_48257,N_46404,N_47176);
nor U48258 (N_48258,N_46204,N_46279);
nand U48259 (N_48259,N_47666,N_47806);
nand U48260 (N_48260,N_47093,N_46805);
nor U48261 (N_48261,N_47795,N_47810);
and U48262 (N_48262,N_46945,N_46353);
or U48263 (N_48263,N_47182,N_46635);
and U48264 (N_48264,N_47670,N_46947);
and U48265 (N_48265,N_46782,N_47289);
nor U48266 (N_48266,N_46221,N_47047);
or U48267 (N_48267,N_47374,N_46874);
and U48268 (N_48268,N_46824,N_46143);
or U48269 (N_48269,N_46352,N_47828);
or U48270 (N_48270,N_47200,N_47033);
nand U48271 (N_48271,N_46562,N_46963);
nand U48272 (N_48272,N_47499,N_47818);
or U48273 (N_48273,N_47158,N_46234);
or U48274 (N_48274,N_46417,N_47942);
nand U48275 (N_48275,N_46754,N_46924);
nor U48276 (N_48276,N_46466,N_47703);
xnor U48277 (N_48277,N_46633,N_46616);
and U48278 (N_48278,N_46619,N_47652);
and U48279 (N_48279,N_46766,N_47483);
or U48280 (N_48280,N_47923,N_47540);
or U48281 (N_48281,N_47114,N_47356);
xor U48282 (N_48282,N_47561,N_47707);
nand U48283 (N_48283,N_46072,N_47128);
nor U48284 (N_48284,N_47448,N_47915);
nor U48285 (N_48285,N_47177,N_46718);
and U48286 (N_48286,N_46550,N_46863);
xor U48287 (N_48287,N_46772,N_47692);
xnor U48288 (N_48288,N_47458,N_46702);
nor U48289 (N_48289,N_46957,N_46035);
xnor U48290 (N_48290,N_47111,N_46125);
and U48291 (N_48291,N_47600,N_47512);
nor U48292 (N_48292,N_47956,N_47212);
and U48293 (N_48293,N_47478,N_46820);
nand U48294 (N_48294,N_46728,N_46668);
xnor U48295 (N_48295,N_47265,N_46472);
nor U48296 (N_48296,N_47416,N_46280);
xor U48297 (N_48297,N_46847,N_47880);
xnor U48298 (N_48298,N_46509,N_47210);
nor U48299 (N_48299,N_46968,N_47950);
nand U48300 (N_48300,N_46687,N_47929);
and U48301 (N_48301,N_47580,N_46246);
or U48302 (N_48302,N_47396,N_47998);
nor U48303 (N_48303,N_46308,N_47127);
and U48304 (N_48304,N_46613,N_46081);
nor U48305 (N_48305,N_47816,N_46270);
xor U48306 (N_48306,N_47501,N_46690);
xnor U48307 (N_48307,N_47167,N_47939);
nand U48308 (N_48308,N_47746,N_46693);
nor U48309 (N_48309,N_47944,N_46411);
nor U48310 (N_48310,N_46908,N_46790);
or U48311 (N_48311,N_47366,N_47211);
nand U48312 (N_48312,N_46082,N_47736);
nor U48313 (N_48313,N_47015,N_47365);
and U48314 (N_48314,N_47091,N_47485);
nand U48315 (N_48315,N_47622,N_47701);
or U48316 (N_48316,N_47181,N_47399);
nand U48317 (N_48317,N_46167,N_47437);
nor U48318 (N_48318,N_46569,N_46675);
and U48319 (N_48319,N_47150,N_47058);
nor U48320 (N_48320,N_47522,N_46671);
and U48321 (N_48321,N_46384,N_47722);
or U48322 (N_48322,N_46041,N_46064);
nand U48323 (N_48323,N_47514,N_46337);
and U48324 (N_48324,N_47426,N_47902);
and U48325 (N_48325,N_47773,N_46439);
nand U48326 (N_48326,N_47471,N_46080);
nor U48327 (N_48327,N_47021,N_46716);
xnor U48328 (N_48328,N_47115,N_46316);
nand U48329 (N_48329,N_47052,N_46252);
xnor U48330 (N_48330,N_47313,N_47525);
nand U48331 (N_48331,N_47985,N_47793);
xor U48332 (N_48332,N_47125,N_46695);
or U48333 (N_48333,N_46059,N_46380);
nor U48334 (N_48334,N_46067,N_47608);
and U48335 (N_48335,N_46755,N_47554);
and U48336 (N_48336,N_46872,N_46225);
xnor U48337 (N_48337,N_47260,N_47943);
and U48338 (N_48338,N_47358,N_47840);
and U48339 (N_48339,N_47546,N_47862);
xor U48340 (N_48340,N_46310,N_47653);
xnor U48341 (N_48341,N_46837,N_46640);
or U48342 (N_48342,N_46642,N_46712);
and U48343 (N_48343,N_47686,N_46520);
nor U48344 (N_48344,N_47154,N_47126);
nand U48345 (N_48345,N_47098,N_47314);
nor U48346 (N_48346,N_46456,N_46573);
nor U48347 (N_48347,N_47988,N_46261);
xor U48348 (N_48348,N_46575,N_47216);
nand U48349 (N_48349,N_47981,N_46079);
nand U48350 (N_48350,N_47890,N_47595);
and U48351 (N_48351,N_46311,N_47755);
nor U48352 (N_48352,N_46084,N_46199);
and U48353 (N_48353,N_46811,N_47520);
nand U48354 (N_48354,N_46145,N_47481);
nand U48355 (N_48355,N_47045,N_47994);
nor U48356 (N_48356,N_47055,N_47861);
xor U48357 (N_48357,N_46302,N_46052);
nor U48358 (N_48358,N_47371,N_46465);
and U48359 (N_48359,N_46993,N_47721);
nor U48360 (N_48360,N_46912,N_46242);
or U48361 (N_48361,N_47162,N_46585);
and U48362 (N_48362,N_46796,N_46665);
xor U48363 (N_48363,N_47403,N_46738);
xnor U48364 (N_48364,N_46859,N_47174);
xor U48365 (N_48365,N_47562,N_47057);
or U48366 (N_48366,N_46909,N_46156);
and U48367 (N_48367,N_47349,N_46389);
and U48368 (N_48368,N_47610,N_46589);
and U48369 (N_48369,N_46402,N_47636);
or U48370 (N_48370,N_46899,N_47345);
nand U48371 (N_48371,N_46867,N_47741);
nand U48372 (N_48372,N_46605,N_47491);
nor U48373 (N_48373,N_46984,N_46676);
nor U48374 (N_48374,N_46071,N_47397);
xnor U48375 (N_48375,N_46667,N_46258);
and U48376 (N_48376,N_46780,N_47754);
and U48377 (N_48377,N_46688,N_47913);
and U48378 (N_48378,N_46339,N_46305);
nand U48379 (N_48379,N_47990,N_47958);
xnor U48380 (N_48380,N_46001,N_46594);
xnor U48381 (N_48381,N_46861,N_47850);
nor U48382 (N_48382,N_46030,N_46345);
nor U48383 (N_48383,N_47671,N_46710);
nor U48384 (N_48384,N_46567,N_47051);
or U48385 (N_48385,N_47119,N_47385);
and U48386 (N_48386,N_46659,N_46864);
nand U48387 (N_48387,N_46990,N_47771);
xor U48388 (N_48388,N_47799,N_46723);
nand U48389 (N_48389,N_47468,N_46294);
and U48390 (N_48390,N_47794,N_46663);
nor U48391 (N_48391,N_47516,N_46529);
nand U48392 (N_48392,N_47805,N_46956);
nand U48393 (N_48393,N_47637,N_46459);
nand U48394 (N_48394,N_46525,N_47236);
nand U48395 (N_48395,N_47107,N_46322);
nor U48396 (N_48396,N_47827,N_47219);
or U48397 (N_48397,N_47673,N_47281);
and U48398 (N_48398,N_46778,N_47068);
or U48399 (N_48399,N_46154,N_47157);
nand U48400 (N_48400,N_46355,N_46114);
and U48401 (N_48401,N_46893,N_47577);
nor U48402 (N_48402,N_47949,N_46271);
nor U48403 (N_48403,N_46425,N_47953);
nor U48404 (N_48404,N_46661,N_47654);
nand U48405 (N_48405,N_46365,N_47373);
or U48406 (N_48406,N_47305,N_46941);
xnor U48407 (N_48407,N_46324,N_47191);
or U48408 (N_48408,N_46944,N_46307);
and U48409 (N_48409,N_46581,N_46237);
xnor U48410 (N_48410,N_46896,N_46146);
nand U48411 (N_48411,N_47035,N_46350);
nand U48412 (N_48412,N_47410,N_46724);
xor U48413 (N_48413,N_46101,N_47213);
or U48414 (N_48414,N_46631,N_46599);
nor U48415 (N_48415,N_47808,N_47738);
or U48416 (N_48416,N_46888,N_46691);
nor U48417 (N_48417,N_46574,N_47082);
or U48418 (N_48418,N_47108,N_47368);
nand U48419 (N_48419,N_46282,N_47473);
or U48420 (N_48420,N_46329,N_46933);
xnor U48421 (N_48421,N_47180,N_46112);
or U48422 (N_48422,N_46326,N_47696);
nor U48423 (N_48423,N_47252,N_46806);
or U48424 (N_48424,N_46999,N_46207);
nor U48425 (N_48425,N_47591,N_46422);
xnor U48426 (N_48426,N_46272,N_47393);
nand U48427 (N_48427,N_47918,N_47802);
nor U48428 (N_48428,N_47198,N_46376);
xor U48429 (N_48429,N_47765,N_46200);
and U48430 (N_48430,N_47224,N_46078);
nand U48431 (N_48431,N_47582,N_46587);
nand U48432 (N_48432,N_47286,N_47040);
xor U48433 (N_48433,N_46317,N_47615);
xor U48434 (N_48434,N_46705,N_47782);
or U48435 (N_48435,N_46853,N_47337);
nor U48436 (N_48436,N_46184,N_46460);
nor U48437 (N_48437,N_47197,N_47309);
xnor U48438 (N_48438,N_47155,N_46070);
nand U48439 (N_48439,N_47318,N_46331);
and U48440 (N_48440,N_46602,N_46387);
nand U48441 (N_48441,N_47646,N_47572);
xor U48442 (N_48442,N_47282,N_46974);
or U48443 (N_48443,N_47971,N_47065);
or U48444 (N_48444,N_46787,N_46886);
xor U48445 (N_48445,N_46281,N_47689);
nor U48446 (N_48446,N_47168,N_47874);
xor U48447 (N_48447,N_46361,N_47169);
nand U48448 (N_48448,N_46547,N_46876);
nand U48449 (N_48449,N_47092,N_46423);
xnor U48450 (N_48450,N_47334,N_46467);
and U48451 (N_48451,N_47095,N_47479);
xor U48452 (N_48452,N_47436,N_47982);
xnor U48453 (N_48453,N_46333,N_46290);
and U48454 (N_48454,N_46982,N_46248);
or U48455 (N_48455,N_46217,N_46500);
nand U48456 (N_48456,N_46636,N_47969);
nor U48457 (N_48457,N_47507,N_47433);
nand U48458 (N_48458,N_46319,N_47863);
or U48459 (N_48459,N_47460,N_46297);
xor U48460 (N_48460,N_47868,N_46674);
and U48461 (N_48461,N_47594,N_47151);
or U48462 (N_48462,N_47263,N_46735);
and U48463 (N_48463,N_46087,N_47576);
nor U48464 (N_48464,N_47829,N_46390);
xnor U48465 (N_48465,N_47720,N_47222);
xor U48466 (N_48466,N_46926,N_47539);
and U48467 (N_48467,N_47031,N_47857);
xnor U48468 (N_48468,N_46314,N_47070);
xor U48469 (N_48469,N_46854,N_46979);
nor U48470 (N_48470,N_47611,N_47729);
or U48471 (N_48471,N_47340,N_46205);
xnor U48472 (N_48472,N_46269,N_46065);
or U48473 (N_48473,N_46995,N_46285);
and U48474 (N_48474,N_46516,N_46637);
nor U48475 (N_48475,N_47734,N_47037);
or U48476 (N_48476,N_47599,N_47718);
and U48477 (N_48477,N_47661,N_46494);
nor U48478 (N_48478,N_47175,N_46421);
or U48479 (N_48479,N_46284,N_46468);
and U48480 (N_48480,N_46434,N_47482);
and U48481 (N_48481,N_47977,N_46701);
nor U48482 (N_48482,N_46857,N_47872);
nand U48483 (N_48483,N_46478,N_47511);
nor U48484 (N_48484,N_46684,N_47088);
and U48485 (N_48485,N_46262,N_46817);
nor U48486 (N_48486,N_47384,N_46312);
and U48487 (N_48487,N_46485,N_47109);
and U48488 (N_48488,N_46483,N_46508);
xor U48489 (N_48489,N_47609,N_46741);
and U48490 (N_48490,N_47463,N_46356);
nor U48491 (N_48491,N_46177,N_46155);
nand U48492 (N_48492,N_46975,N_47871);
nor U48493 (N_48493,N_47392,N_47725);
xor U48494 (N_48494,N_46770,N_46238);
nor U48495 (N_48495,N_46503,N_47201);
or U48496 (N_48496,N_46533,N_46887);
nand U48497 (N_48497,N_46489,N_46056);
nor U48498 (N_48498,N_46634,N_47834);
xor U48499 (N_48499,N_46215,N_47307);
and U48500 (N_48500,N_46730,N_46542);
nor U48501 (N_48501,N_46162,N_47714);
and U48502 (N_48502,N_46394,N_47311);
nand U48503 (N_48503,N_47280,N_46593);
xor U48504 (N_48504,N_46354,N_46937);
xnor U48505 (N_48505,N_47847,N_47856);
or U48506 (N_48506,N_47823,N_47432);
or U48507 (N_48507,N_46653,N_46923);
and U48508 (N_48508,N_46054,N_47800);
xor U48509 (N_48509,N_46031,N_46499);
xnor U48510 (N_48510,N_47934,N_47819);
or U48511 (N_48511,N_47208,N_47156);
nand U48512 (N_48512,N_47508,N_46405);
or U48513 (N_48513,N_46268,N_47798);
xnor U48514 (N_48514,N_47740,N_47625);
or U48515 (N_48515,N_47226,N_47976);
nand U48516 (N_48516,N_46540,N_46530);
nor U48517 (N_48517,N_46880,N_47376);
xnor U48518 (N_48518,N_47602,N_46729);
and U48519 (N_48519,N_46700,N_46039);
and U48520 (N_48520,N_46291,N_47813);
xnor U48521 (N_48521,N_47898,N_47842);
nand U48522 (N_48522,N_47122,N_46583);
and U48523 (N_48523,N_46208,N_47415);
nand U48524 (N_48524,N_46198,N_46807);
or U48525 (N_48525,N_46512,N_47342);
nor U48526 (N_48526,N_46809,N_46357);
nor U48527 (N_48527,N_46929,N_47228);
xnor U48528 (N_48528,N_46432,N_47732);
and U48529 (N_48529,N_46577,N_46832);
or U48530 (N_48530,N_47455,N_46193);
nor U48531 (N_48531,N_46697,N_46388);
nand U48532 (N_48532,N_46935,N_46016);
and U48533 (N_48533,N_47691,N_46784);
xor U48534 (N_48534,N_46860,N_46555);
or U48535 (N_48535,N_47456,N_47817);
or U48536 (N_48536,N_47901,N_47775);
nor U48537 (N_48537,N_47249,N_47769);
or U48538 (N_48538,N_47875,N_46794);
or U48539 (N_48539,N_46890,N_46206);
xnor U48540 (N_48540,N_46985,N_47025);
or U48541 (N_48541,N_47631,N_47853);
xor U48542 (N_48542,N_47220,N_47300);
nor U48543 (N_48543,N_46681,N_47140);
nor U48544 (N_48544,N_46158,N_46142);
xor U48545 (N_48545,N_46328,N_47940);
xor U48546 (N_48546,N_47656,N_46050);
xor U48547 (N_48547,N_47549,N_47029);
nand U48548 (N_48548,N_47295,N_47317);
nand U48549 (N_48549,N_46372,N_46915);
and U48550 (N_48550,N_47811,N_47560);
or U48551 (N_48551,N_47118,N_46692);
nand U48552 (N_48552,N_47351,N_46250);
and U48553 (N_48553,N_46415,N_47493);
or U48554 (N_48554,N_46152,N_47770);
nor U48555 (N_48555,N_46983,N_46220);
or U48556 (N_48556,N_46233,N_47524);
or U48557 (N_48557,N_47624,N_46495);
and U48558 (N_48558,N_47632,N_47293);
nand U48559 (N_48559,N_46083,N_47536);
nor U48560 (N_48560,N_47256,N_47014);
nor U48561 (N_48561,N_46414,N_47955);
or U48562 (N_48562,N_46347,N_46116);
and U48563 (N_48563,N_47398,N_47975);
or U48564 (N_48564,N_47225,N_46748);
nand U48565 (N_48565,N_46232,N_46186);
nor U48566 (N_48566,N_46196,N_47537);
nand U48567 (N_48567,N_47848,N_47352);
nor U48568 (N_48568,N_47597,N_47291);
xnor U48569 (N_48569,N_47270,N_46511);
or U48570 (N_48570,N_46842,N_46655);
nor U48571 (N_48571,N_46247,N_47665);
nand U48572 (N_48572,N_47382,N_47621);
xor U48573 (N_48573,N_47316,N_47388);
or U48574 (N_48574,N_47843,N_46907);
and U48575 (N_48575,N_46096,N_46446);
or U48576 (N_48576,N_46264,N_47084);
or U48577 (N_48577,N_46744,N_47968);
nor U48578 (N_48578,N_47017,N_46482);
nor U48579 (N_48579,N_46801,N_47888);
and U48580 (N_48580,N_47620,N_46895);
nor U48581 (N_48581,N_47355,N_46804);
nand U48582 (N_48582,N_47509,N_47584);
or U48583 (N_48583,N_46672,N_47394);
nand U48584 (N_48584,N_46033,N_47290);
nand U48585 (N_48585,N_46479,N_47983);
nand U48586 (N_48586,N_47908,N_47917);
nand U48587 (N_48587,N_47424,N_46362);
xor U48588 (N_48588,N_46825,N_47695);
nand U48589 (N_48589,N_46571,N_47601);
or U48590 (N_48590,N_46037,N_46666);
nor U48591 (N_48591,N_46288,N_47012);
and U48592 (N_48592,N_46517,N_47932);
xor U48593 (N_48593,N_47886,N_47739);
or U48594 (N_48594,N_46792,N_47744);
and U48595 (N_48595,N_47038,N_47430);
nor U48596 (N_48596,N_46473,N_46018);
nor U48597 (N_48597,N_46369,N_46936);
and U48598 (N_48598,N_47261,N_46408);
nand U48599 (N_48599,N_47836,N_46061);
or U48600 (N_48600,N_46998,N_46992);
nor U48601 (N_48601,N_46165,N_46450);
or U48602 (N_48602,N_47073,N_46747);
or U48603 (N_48603,N_46584,N_46192);
or U48604 (N_48604,N_47786,N_46260);
and U48605 (N_48605,N_46526,N_47693);
xnor U48606 (N_48606,N_46235,N_47331);
nand U48607 (N_48607,N_47467,N_47190);
or U48608 (N_48608,N_47556,N_46664);
nor U48609 (N_48609,N_47663,N_46188);
and U48610 (N_48610,N_46172,N_46175);
or U48611 (N_48611,N_46254,N_47687);
xnor U48612 (N_48612,N_46879,N_47137);
nand U48613 (N_48613,N_46527,N_46004);
or U48614 (N_48614,N_47947,N_47412);
nand U48615 (N_48615,N_47954,N_47333);
nand U48616 (N_48616,N_47682,N_47960);
xnor U48617 (N_48617,N_46420,N_46009);
nor U48618 (N_48618,N_47867,N_46366);
and U48619 (N_48619,N_47179,N_47792);
or U48620 (N_48620,N_46761,N_46126);
xnor U48621 (N_48621,N_46699,N_47007);
or U48622 (N_48622,N_47123,N_47321);
xor U48623 (N_48623,N_47660,N_47320);
xnor U48624 (N_48624,N_47427,N_46802);
and U48625 (N_48625,N_46513,N_47075);
nand U48626 (N_48626,N_46793,N_46000);
nor U48627 (N_48627,N_47377,N_46019);
or U48628 (N_48628,N_47809,N_46013);
and U48629 (N_48629,N_46726,N_46551);
nor U48630 (N_48630,N_46507,N_47303);
nand U48631 (N_48631,N_46430,N_46159);
nor U48632 (N_48632,N_46739,N_47010);
and U48633 (N_48633,N_47086,N_46643);
nor U48634 (N_48634,N_46181,N_47523);
or U48635 (N_48635,N_46391,N_46769);
nor U48636 (N_48636,N_46654,N_46743);
nand U48637 (N_48637,N_46814,N_46166);
xor U48638 (N_48638,N_47492,N_47750);
or U48639 (N_48639,N_46449,N_47783);
or U48640 (N_48640,N_47761,N_46873);
nand U48641 (N_48641,N_46556,N_47239);
nand U48642 (N_48642,N_46436,N_47820);
or U48643 (N_48643,N_47184,N_47678);
or U48644 (N_48644,N_47133,N_46327);
nor U48645 (N_48645,N_47490,N_46212);
or U48646 (N_48646,N_46737,N_47383);
or U48647 (N_48647,N_47992,N_47899);
or U48648 (N_48648,N_47297,N_46275);
nor U48649 (N_48649,N_46917,N_47063);
and U48650 (N_48650,N_46042,N_46060);
and U48651 (N_48651,N_47995,N_46949);
and U48652 (N_48652,N_46299,N_47072);
nand U48653 (N_48653,N_47453,N_46504);
nor U48654 (N_48654,N_47519,N_47267);
nor U48655 (N_48655,N_46393,N_47165);
xnor U48656 (N_48656,N_46554,N_47613);
nor U48657 (N_48657,N_46014,N_47440);
nor U48658 (N_48658,N_47796,N_46171);
and U48659 (N_48659,N_46289,N_46251);
nor U48660 (N_48660,N_47804,N_47292);
or U48661 (N_48661,N_46838,N_46144);
nand U48662 (N_48662,N_46229,N_47749);
or U48663 (N_48663,N_46194,N_46124);
and U48664 (N_48664,N_46007,N_46994);
or U48665 (N_48665,N_46025,N_46068);
and U48666 (N_48666,N_47784,N_46646);
nor U48667 (N_48667,N_47244,N_46100);
or U48668 (N_48668,N_46195,N_46987);
and U48669 (N_48669,N_46749,N_47241);
xor U48670 (N_48670,N_46179,N_47553);
nand U48671 (N_48671,N_47390,N_46445);
and U48672 (N_48672,N_46767,N_46759);
and U48673 (N_48673,N_46226,N_47937);
nand U48674 (N_48674,N_47003,N_46713);
nand U48675 (N_48675,N_46036,N_46742);
and U48676 (N_48676,N_47672,N_47142);
or U48677 (N_48677,N_46374,N_47542);
nor U48678 (N_48678,N_47550,N_47596);
xnor U48679 (N_48679,N_47147,N_46026);
xor U48680 (N_48680,N_46934,N_47379);
and U48681 (N_48681,N_46835,N_47626);
xor U48682 (N_48682,N_46501,N_46492);
and U48683 (N_48683,N_46851,N_47855);
nand U48684 (N_48684,N_47250,N_46410);
xnor U48685 (N_48685,N_46570,N_47700);
xor U48686 (N_48686,N_47100,N_46791);
and U48687 (N_48687,N_46185,N_47428);
and U48688 (N_48688,N_47664,N_47315);
nor U48689 (N_48689,N_47423,N_47997);
and U48690 (N_48690,N_46283,N_47452);
xor U48691 (N_48691,N_47262,N_46916);
or U48692 (N_48692,N_47851,N_46378);
nor U48693 (N_48693,N_47344,N_47758);
nand U48694 (N_48694,N_46920,N_46224);
and U48695 (N_48695,N_46148,N_46174);
nand U48696 (N_48696,N_47132,N_46141);
nor U48697 (N_48697,N_46826,N_46703);
nor U48698 (N_48698,N_46046,N_47008);
xnor U48699 (N_48699,N_47675,N_47963);
nor U48700 (N_48700,N_47573,N_47011);
and U48701 (N_48701,N_47970,N_46153);
nand U48702 (N_48702,N_47776,N_46371);
and U48703 (N_48703,N_47445,N_47363);
nor U48704 (N_48704,N_47989,N_47914);
nand U48705 (N_48705,N_46756,N_47991);
nor U48706 (N_48706,N_46298,N_46973);
nor U48707 (N_48707,N_47090,N_46253);
and U48708 (N_48708,N_47619,N_46412);
xor U48709 (N_48709,N_46118,N_47651);
xnor U48710 (N_48710,N_46024,N_46855);
nor U48711 (N_48711,N_47822,N_46607);
nor U48712 (N_48712,N_46182,N_47024);
xor U48713 (N_48713,N_47276,N_46758);
nand U48714 (N_48714,N_46816,N_47248);
or U48715 (N_48715,N_47559,N_47457);
nand U48716 (N_48716,N_46561,N_46543);
and U48717 (N_48717,N_47544,N_47702);
nand U48718 (N_48718,N_47141,N_47698);
xnor U48719 (N_48719,N_46889,N_47688);
xor U48720 (N_48720,N_46704,N_46190);
or U48721 (N_48721,N_46265,N_46715);
or U48722 (N_48722,N_47984,N_46740);
nand U48723 (N_48723,N_47353,N_46092);
xor U48724 (N_48724,N_46946,N_46919);
or U48725 (N_48725,N_46406,N_46969);
and U48726 (N_48726,N_46914,N_46563);
xor U48727 (N_48727,N_47418,N_47844);
or U48728 (N_48728,N_47339,N_47964);
nor U48729 (N_48729,N_46458,N_46732);
nor U48730 (N_48730,N_46267,N_46418);
or U48731 (N_48731,N_47214,N_46731);
or U48732 (N_48732,N_47278,N_47494);
or U48733 (N_48733,N_47709,N_46183);
xor U48734 (N_48734,N_46757,N_46720);
nand U48735 (N_48735,N_47130,N_46133);
nand U48736 (N_48736,N_47587,N_46822);
nand U48737 (N_48737,N_46948,N_46428);
nand U48738 (N_48738,N_46349,N_46095);
xor U48739 (N_48739,N_47414,N_47644);
or U48740 (N_48740,N_46844,N_47294);
nor U48741 (N_48741,N_47726,N_46401);
xor U48742 (N_48742,N_46638,N_46866);
and U48743 (N_48743,N_47101,N_47579);
or U48744 (N_48744,N_47420,N_47706);
or U48745 (N_48745,N_47360,N_47951);
nand U48746 (N_48746,N_46163,N_46799);
nand U48747 (N_48747,N_46649,N_46395);
or U48748 (N_48748,N_47803,N_47163);
xor U48749 (N_48749,N_46469,N_46601);
nor U48750 (N_48750,N_46455,N_47737);
nand U48751 (N_48751,N_46604,N_47972);
or U48752 (N_48752,N_46038,N_46211);
nand U48753 (N_48753,N_47357,N_47883);
xor U48754 (N_48754,N_47860,N_46214);
and U48755 (N_48755,N_47801,N_47962);
or U48756 (N_48756,N_47022,N_46120);
and U48757 (N_48757,N_46870,N_46351);
nor U48758 (N_48758,N_47825,N_46073);
or U48759 (N_48759,N_46338,N_46877);
and U48760 (N_48760,N_47894,N_46828);
nor U48761 (N_48761,N_47529,N_46538);
nor U48762 (N_48762,N_47676,N_46800);
nor U48763 (N_48763,N_47752,N_47302);
and U48764 (N_48764,N_46164,N_46620);
or U48765 (N_48765,N_47489,N_47900);
or U48766 (N_48766,N_47690,N_47304);
xor U48767 (N_48767,N_46416,N_47116);
and U48768 (N_48768,N_46454,N_46972);
or U48769 (N_48769,N_47402,N_47645);
and U48770 (N_48770,N_47223,N_47324);
nor U48771 (N_48771,N_46612,N_47364);
nand U48772 (N_48772,N_47927,N_47727);
xnor U48773 (N_48773,N_46209,N_46093);
nor U48774 (N_48774,N_47961,N_46624);
and U48775 (N_48775,N_46760,N_46377);
xor U48776 (N_48776,N_47504,N_47854);
and U48777 (N_48777,N_47475,N_47288);
and U48778 (N_48778,N_47966,N_47346);
or U48779 (N_48779,N_46650,N_46502);
xor U48780 (N_48780,N_46682,N_47662);
nand U48781 (N_48781,N_47912,N_47973);
xor U48782 (N_48782,N_47824,N_46223);
nor U48783 (N_48783,N_46962,N_46976);
nand U48784 (N_48784,N_46938,N_46475);
and U48785 (N_48785,N_46058,N_46119);
nor U48786 (N_48786,N_46231,N_47153);
nor U48787 (N_48787,N_47386,N_47034);
nand U48788 (N_48788,N_46399,N_47032);
xor U48789 (N_48789,N_46892,N_47598);
or U48790 (N_48790,N_46882,N_46219);
nand U48791 (N_48791,N_46370,N_46470);
and U48792 (N_48792,N_46625,N_46980);
xnor U48793 (N_48793,N_46553,N_46644);
nor U48794 (N_48794,N_47650,N_46522);
nand U48795 (N_48795,N_46122,N_47717);
nor U48796 (N_48796,N_47243,N_47002);
nand U48797 (N_48797,N_47129,N_46440);
xor U48798 (N_48798,N_47411,N_46300);
and U48799 (N_48799,N_46481,N_46178);
nand U48800 (N_48800,N_46603,N_47497);
and U48801 (N_48801,N_47618,N_47845);
or U48802 (N_48802,N_47699,N_46925);
or U48803 (N_48803,N_47607,N_46245);
xnor U48804 (N_48804,N_46708,N_46834);
and U48805 (N_48805,N_47588,N_46303);
nand U48806 (N_48806,N_46545,N_46988);
xor U48807 (N_48807,N_46996,N_47042);
xor U48808 (N_48808,N_46833,N_47277);
nand U48809 (N_48809,N_47495,N_47952);
nand U48810 (N_48810,N_47563,N_47916);
nor U48811 (N_48811,N_46273,N_46170);
nand U48812 (N_48812,N_46476,N_46652);
nor U48813 (N_48813,N_47194,N_47640);
nand U48814 (N_48814,N_46618,N_47878);
nand U48815 (N_48815,N_47831,N_46918);
nand U48816 (N_48816,N_46798,N_47268);
or U48817 (N_48817,N_46150,N_46883);
or U48818 (N_48818,N_46884,N_47513);
and U48819 (N_48819,N_47350,N_47199);
nor U48820 (N_48820,N_47578,N_47551);
or U48821 (N_48821,N_46202,N_46309);
and U48822 (N_48822,N_46121,N_47781);
and U48823 (N_48823,N_47835,N_47685);
nand U48824 (N_48824,N_46928,N_47909);
xnor U48825 (N_48825,N_47617,N_46457);
nor U48826 (N_48826,N_46849,N_46375);
and U48827 (N_48827,N_47503,N_47135);
nor U48828 (N_48828,N_47161,N_47284);
xor U48829 (N_48829,N_46462,N_46110);
or U48830 (N_48830,N_47299,N_46263);
nand U48831 (N_48831,N_46360,N_47887);
nor U48832 (N_48832,N_47533,N_46669);
or U48833 (N_48833,N_46213,N_46600);
nand U48834 (N_48834,N_47160,N_46978);
nand U48835 (N_48835,N_47099,N_47441);
and U48836 (N_48836,N_47013,N_46346);
nor U48837 (N_48837,N_46558,N_47323);
nor U48838 (N_48838,N_47381,N_46736);
or U48839 (N_48839,N_47378,N_47604);
nor U48840 (N_48840,N_46123,N_47069);
xnor U48841 (N_48841,N_46051,N_46955);
nand U48842 (N_48842,N_46108,N_46109);
xnor U48843 (N_48843,N_46904,N_46131);
and U48844 (N_48844,N_47283,N_47921);
nand U48845 (N_48845,N_47649,N_47409);
xnor U48846 (N_48846,N_46017,N_46752);
xnor U48847 (N_48847,N_46400,N_47347);
nor U48848 (N_48848,N_47192,N_47425);
nor U48849 (N_48849,N_46559,N_47446);
xor U48850 (N_48850,N_46789,N_46750);
nand U48851 (N_48851,N_46128,N_47319);
xnor U48852 (N_48852,N_46894,N_47429);
or U48853 (N_48853,N_46535,N_46098);
xnor U48854 (N_48854,N_47933,N_46398);
or U48855 (N_48855,N_46813,N_46332);
xor U48856 (N_48856,N_46008,N_46497);
or U48857 (N_48857,N_47742,N_46611);
and U48858 (N_48858,N_46797,N_46433);
and U48859 (N_48859,N_47538,N_47846);
nand U48860 (N_48860,N_47790,N_46903);
or U48861 (N_48861,N_47570,N_46694);
or U48862 (N_48862,N_47885,N_47145);
nand U48863 (N_48863,N_46396,N_47421);
or U48864 (N_48864,N_46386,N_46606);
nor U48865 (N_48865,N_46871,N_46541);
and U48866 (N_48866,N_46630,N_47978);
xor U48867 (N_48867,N_46383,N_47575);
and U48868 (N_48868,N_47629,N_47209);
nand U48869 (N_48869,N_46840,N_46222);
and U48870 (N_48870,N_47628,N_47287);
and U48871 (N_48871,N_47449,N_47020);
xor U48872 (N_48872,N_46673,N_46707);
nor U48873 (N_48873,N_46539,N_47067);
and U48874 (N_48874,N_46044,N_46323);
or U48875 (N_48875,N_46160,N_47606);
nor U48876 (N_48876,N_47797,N_47547);
xor U48877 (N_48877,N_47757,N_47203);
or U48878 (N_48878,N_47050,N_47728);
nand U48879 (N_48879,N_47833,N_47348);
xnor U48880 (N_48880,N_46239,N_47895);
nand U48881 (N_48881,N_47919,N_47327);
nor U48882 (N_48882,N_47152,N_47359);
nand U48883 (N_48883,N_46641,N_46130);
nand U48884 (N_48884,N_47684,N_46379);
or U48885 (N_48885,N_47593,N_47891);
or U48886 (N_48886,N_46627,N_47574);
or U48887 (N_48887,N_47567,N_46407);
nand U48888 (N_48888,N_46381,N_46549);
and U48889 (N_48889,N_46091,N_46047);
xnor U48890 (N_48890,N_47751,N_47926);
or U48891 (N_48891,N_46135,N_46315);
nor U48892 (N_48892,N_46168,N_46819);
and U48893 (N_48893,N_46537,N_47361);
and U48894 (N_48894,N_47838,N_46906);
nor U48895 (N_48895,N_47275,N_47677);
xor U48896 (N_48896,N_47062,N_46812);
nand U48897 (N_48897,N_46409,N_47648);
xnor U48898 (N_48898,N_46662,N_47465);
nand U48899 (N_48899,N_47059,N_46010);
xnor U48900 (N_48900,N_46138,N_46777);
nor U48901 (N_48901,N_47439,N_46474);
xnor U48902 (N_48902,N_47080,N_46977);
or U48903 (N_48903,N_47134,N_47296);
xnor U48904 (N_48904,N_47273,N_47658);
or U48905 (N_48905,N_46897,N_46257);
and U48906 (N_48906,N_46278,N_46768);
and U48907 (N_48907,N_46639,N_47196);
xor U48908 (N_48908,N_46241,N_47335);
nand U48909 (N_48909,N_47530,N_47400);
or U48910 (N_48910,N_46249,N_47112);
and U48911 (N_48911,N_47614,N_47708);
nand U48912 (N_48912,N_46040,N_47541);
xor U48913 (N_48913,N_46528,N_46063);
or U48914 (N_48914,N_46745,N_47788);
or U48915 (N_48915,N_46189,N_46865);
or U48916 (N_48916,N_47841,N_46579);
xor U48917 (N_48917,N_47815,N_46336);
xnor U48918 (N_48918,N_47341,N_46201);
xnor U48919 (N_48919,N_47945,N_46557);
nand U48920 (N_48920,N_46722,N_47922);
nor U48921 (N_48921,N_46514,N_46343);
xnor U48922 (N_48922,N_47097,N_47974);
xor U48923 (N_48923,N_47375,N_47312);
nand U48924 (N_48924,N_47079,N_46781);
nand U48925 (N_48925,N_47106,N_47730);
xor U48926 (N_48926,N_47635,N_47053);
and U48927 (N_48927,N_46340,N_46576);
nand U48928 (N_48928,N_46588,N_46964);
nor U48929 (N_48929,N_47789,N_47285);
nand U48930 (N_48930,N_47395,N_46027);
xnor U48931 (N_48931,N_47235,N_47568);
nand U48932 (N_48932,N_47087,N_47131);
and U48933 (N_48933,N_46921,N_47064);
xnor U48934 (N_48934,N_47980,N_46129);
nor U48935 (N_48935,N_47911,N_47240);
and U48936 (N_48936,N_47928,N_47301);
and U48937 (N_48937,N_47001,N_46830);
nor U48938 (N_48938,N_47193,N_47487);
and U48939 (N_48939,N_46651,N_47271);
nor U48940 (N_48940,N_46596,N_46657);
and U48941 (N_48941,N_46069,N_47061);
nand U48942 (N_48942,N_47362,N_46615);
xor U48943 (N_48943,N_46991,N_46686);
nor U48944 (N_48944,N_47016,N_46488);
xnor U48945 (N_48945,N_46236,N_47526);
or U48946 (N_48946,N_47207,N_47215);
nand U48947 (N_48947,N_46617,N_46173);
nor U48948 (N_48948,N_46891,N_47859);
nor U48949 (N_48949,N_47401,N_46521);
or U48950 (N_48950,N_46930,N_46595);
xnor U48951 (N_48951,N_47404,N_46900);
and U48952 (N_48952,N_47634,N_46862);
xor U48953 (N_48953,N_46534,N_47555);
or U48954 (N_48954,N_46086,N_47668);
xnor U48955 (N_48955,N_47462,N_47711);
and U48956 (N_48956,N_46823,N_47486);
nor U48957 (N_48957,N_47986,N_46515);
nor U48958 (N_48958,N_46531,N_46392);
xor U48959 (N_48959,N_47380,N_46821);
or U48960 (N_48960,N_47865,N_47589);
nand U48961 (N_48961,N_46942,N_46103);
xnor U48962 (N_48962,N_47679,N_46658);
nand U48963 (N_48963,N_46493,N_47659);
or U48964 (N_48964,N_47264,N_46115);
nor U48965 (N_48965,N_46203,N_47139);
and U48966 (N_48966,N_47187,N_46342);
xor U48967 (N_48967,N_46586,N_46632);
and U48968 (N_48968,N_47466,N_46592);
xnor U48969 (N_48969,N_47247,N_46373);
nor U48970 (N_48970,N_46506,N_47330);
xor U48971 (N_48971,N_46102,N_46266);
xor U48972 (N_48972,N_46276,N_46321);
or U48973 (N_48973,N_47272,N_47999);
nor U48974 (N_48974,N_47500,N_46021);
nor U48975 (N_48975,N_46382,N_46598);
nand U48976 (N_48976,N_47245,N_47461);
nor U48977 (N_48977,N_47322,N_47630);
xor U48978 (N_48978,N_47477,N_47136);
xor U48979 (N_48979,N_46582,N_47791);
and U48980 (N_48980,N_47936,N_46961);
xnor U48981 (N_48981,N_46590,N_46132);
or U48982 (N_48982,N_47407,N_46003);
or U48983 (N_48983,N_47565,N_46180);
xnor U48984 (N_48984,N_47724,N_46397);
nand U48985 (N_48985,N_47869,N_47238);
xor U48986 (N_48986,N_47413,N_47763);
and U48987 (N_48987,N_47326,N_46591);
xor U48988 (N_48988,N_46049,N_46568);
nor U48989 (N_48989,N_46451,N_47056);
nor U48990 (N_48990,N_47759,N_47041);
and U48991 (N_48991,N_47229,N_47638);
or U48992 (N_48992,N_47274,N_46335);
nand U48993 (N_48993,N_46776,N_46685);
nor U48994 (N_48994,N_47552,N_47641);
nor U48995 (N_48995,N_46012,N_47121);
xnor U48996 (N_48996,N_47905,N_46358);
nor U48997 (N_48997,N_46447,N_46117);
and U48998 (N_48998,N_47258,N_46306);
nand U48999 (N_48999,N_47505,N_46670);
or U49000 (N_49000,N_47337,N_47597);
xnor U49001 (N_49001,N_46666,N_46294);
or U49002 (N_49002,N_47768,N_46382);
nor U49003 (N_49003,N_47046,N_46825);
xnor U49004 (N_49004,N_47896,N_46543);
xor U49005 (N_49005,N_47344,N_46539);
xnor U49006 (N_49006,N_47195,N_47761);
or U49007 (N_49007,N_46896,N_47863);
and U49008 (N_49008,N_47655,N_47712);
or U49009 (N_49009,N_47046,N_47112);
or U49010 (N_49010,N_46505,N_46163);
and U49011 (N_49011,N_47889,N_46376);
nor U49012 (N_49012,N_46502,N_46848);
xor U49013 (N_49013,N_46300,N_47871);
nor U49014 (N_49014,N_46538,N_46921);
xor U49015 (N_49015,N_46198,N_46856);
or U49016 (N_49016,N_46618,N_47207);
nand U49017 (N_49017,N_47295,N_47035);
xor U49018 (N_49018,N_47492,N_46763);
nand U49019 (N_49019,N_46049,N_47589);
or U49020 (N_49020,N_47045,N_47064);
nand U49021 (N_49021,N_47949,N_46862);
nor U49022 (N_49022,N_47520,N_46660);
xor U49023 (N_49023,N_47022,N_47631);
nand U49024 (N_49024,N_47473,N_47308);
or U49025 (N_49025,N_46428,N_46616);
and U49026 (N_49026,N_46142,N_46745);
nor U49027 (N_49027,N_46775,N_46854);
xnor U49028 (N_49028,N_46759,N_47032);
nor U49029 (N_49029,N_46332,N_47093);
nand U49030 (N_49030,N_46938,N_47872);
xnor U49031 (N_49031,N_47760,N_47735);
or U49032 (N_49032,N_47868,N_46401);
and U49033 (N_49033,N_47784,N_46123);
xor U49034 (N_49034,N_46710,N_46757);
nor U49035 (N_49035,N_46707,N_47833);
or U49036 (N_49036,N_47800,N_47671);
or U49037 (N_49037,N_47748,N_47363);
or U49038 (N_49038,N_47846,N_47039);
and U49039 (N_49039,N_46744,N_46134);
nor U49040 (N_49040,N_46545,N_46063);
or U49041 (N_49041,N_47247,N_47303);
nand U49042 (N_49042,N_47782,N_47230);
xor U49043 (N_49043,N_46913,N_46013);
nor U49044 (N_49044,N_47931,N_47664);
and U49045 (N_49045,N_46561,N_46187);
or U49046 (N_49046,N_47478,N_47739);
nand U49047 (N_49047,N_46315,N_47355);
or U49048 (N_49048,N_46803,N_46107);
or U49049 (N_49049,N_47763,N_47876);
nor U49050 (N_49050,N_46134,N_46323);
nor U49051 (N_49051,N_46542,N_47668);
xor U49052 (N_49052,N_46354,N_46211);
and U49053 (N_49053,N_47010,N_46214);
nor U49054 (N_49054,N_47197,N_46520);
nor U49055 (N_49055,N_46726,N_46056);
nand U49056 (N_49056,N_47087,N_46169);
or U49057 (N_49057,N_47851,N_47176);
or U49058 (N_49058,N_46480,N_47097);
and U49059 (N_49059,N_47215,N_46827);
and U49060 (N_49060,N_46431,N_46835);
nand U49061 (N_49061,N_46526,N_47772);
and U49062 (N_49062,N_47627,N_46077);
and U49063 (N_49063,N_46307,N_46561);
or U49064 (N_49064,N_47220,N_47085);
xnor U49065 (N_49065,N_46876,N_47921);
xor U49066 (N_49066,N_47004,N_46408);
or U49067 (N_49067,N_46416,N_46360);
nand U49068 (N_49068,N_47271,N_47808);
and U49069 (N_49069,N_46350,N_46267);
xnor U49070 (N_49070,N_46689,N_46286);
nand U49071 (N_49071,N_47800,N_47255);
xor U49072 (N_49072,N_46022,N_46930);
nor U49073 (N_49073,N_46753,N_47984);
or U49074 (N_49074,N_47243,N_47261);
nor U49075 (N_49075,N_46785,N_46438);
or U49076 (N_49076,N_47500,N_46896);
and U49077 (N_49077,N_46268,N_47288);
xor U49078 (N_49078,N_46520,N_46714);
nor U49079 (N_49079,N_47622,N_46302);
or U49080 (N_49080,N_47034,N_46036);
nand U49081 (N_49081,N_46079,N_47428);
or U49082 (N_49082,N_47075,N_47094);
nor U49083 (N_49083,N_46987,N_46775);
nor U49084 (N_49084,N_47566,N_46156);
nor U49085 (N_49085,N_47808,N_47004);
nor U49086 (N_49086,N_46691,N_47174);
nor U49087 (N_49087,N_46289,N_46099);
nand U49088 (N_49088,N_47778,N_46562);
xnor U49089 (N_49089,N_46073,N_47301);
and U49090 (N_49090,N_47330,N_46239);
and U49091 (N_49091,N_46246,N_47755);
nand U49092 (N_49092,N_46347,N_46230);
xor U49093 (N_49093,N_46667,N_47743);
and U49094 (N_49094,N_47625,N_46307);
and U49095 (N_49095,N_47065,N_47570);
and U49096 (N_49096,N_46639,N_47925);
nand U49097 (N_49097,N_46679,N_47354);
nor U49098 (N_49098,N_46116,N_46734);
nor U49099 (N_49099,N_46048,N_47322);
or U49100 (N_49100,N_47890,N_46905);
and U49101 (N_49101,N_47045,N_46051);
nor U49102 (N_49102,N_47168,N_47348);
nand U49103 (N_49103,N_46767,N_47452);
nor U49104 (N_49104,N_47987,N_46353);
nand U49105 (N_49105,N_46044,N_47452);
xnor U49106 (N_49106,N_47411,N_46832);
nand U49107 (N_49107,N_47305,N_46893);
or U49108 (N_49108,N_46676,N_46741);
nand U49109 (N_49109,N_46896,N_46500);
nor U49110 (N_49110,N_47081,N_47184);
xnor U49111 (N_49111,N_47682,N_47592);
nor U49112 (N_49112,N_46499,N_46500);
or U49113 (N_49113,N_46014,N_46019);
nor U49114 (N_49114,N_46830,N_46035);
and U49115 (N_49115,N_46664,N_46965);
nor U49116 (N_49116,N_47598,N_46883);
nand U49117 (N_49117,N_47645,N_47233);
and U49118 (N_49118,N_47017,N_47362);
or U49119 (N_49119,N_46131,N_47390);
nand U49120 (N_49120,N_46657,N_46059);
xor U49121 (N_49121,N_47932,N_46088);
xor U49122 (N_49122,N_46237,N_47188);
or U49123 (N_49123,N_47762,N_47301);
xnor U49124 (N_49124,N_46334,N_46793);
nand U49125 (N_49125,N_46707,N_47217);
nor U49126 (N_49126,N_46193,N_46147);
nor U49127 (N_49127,N_47528,N_47037);
xor U49128 (N_49128,N_46388,N_47217);
nand U49129 (N_49129,N_47205,N_47641);
xor U49130 (N_49130,N_46242,N_46862);
or U49131 (N_49131,N_46231,N_46303);
nand U49132 (N_49132,N_46177,N_47920);
xor U49133 (N_49133,N_47693,N_46677);
nor U49134 (N_49134,N_46990,N_46698);
nor U49135 (N_49135,N_47032,N_47935);
and U49136 (N_49136,N_46010,N_46571);
nand U49137 (N_49137,N_46228,N_46458);
nor U49138 (N_49138,N_46086,N_47247);
or U49139 (N_49139,N_47923,N_46807);
xnor U49140 (N_49140,N_47646,N_46659);
or U49141 (N_49141,N_47638,N_47396);
xnor U49142 (N_49142,N_47374,N_46822);
or U49143 (N_49143,N_46681,N_47912);
xnor U49144 (N_49144,N_46870,N_47618);
and U49145 (N_49145,N_46819,N_46531);
nor U49146 (N_49146,N_46054,N_47339);
nor U49147 (N_49147,N_47388,N_46494);
and U49148 (N_49148,N_47641,N_47795);
and U49149 (N_49149,N_46335,N_47228);
and U49150 (N_49150,N_47399,N_46973);
nor U49151 (N_49151,N_46144,N_46768);
xor U49152 (N_49152,N_47630,N_47440);
and U49153 (N_49153,N_46512,N_46985);
xor U49154 (N_49154,N_46764,N_47891);
xnor U49155 (N_49155,N_47884,N_46565);
xor U49156 (N_49156,N_47770,N_46070);
xnor U49157 (N_49157,N_47138,N_47261);
xnor U49158 (N_49158,N_46796,N_46939);
nand U49159 (N_49159,N_46914,N_47621);
and U49160 (N_49160,N_46753,N_46953);
nor U49161 (N_49161,N_46086,N_47352);
nand U49162 (N_49162,N_47093,N_47833);
xor U49163 (N_49163,N_46497,N_47105);
and U49164 (N_49164,N_46145,N_46943);
nor U49165 (N_49165,N_46884,N_47982);
xnor U49166 (N_49166,N_46051,N_46859);
nor U49167 (N_49167,N_47011,N_46923);
nand U49168 (N_49168,N_47408,N_46008);
or U49169 (N_49169,N_47219,N_47270);
nand U49170 (N_49170,N_47597,N_47452);
and U49171 (N_49171,N_47841,N_47265);
or U49172 (N_49172,N_47056,N_47265);
nor U49173 (N_49173,N_46486,N_46663);
nor U49174 (N_49174,N_47105,N_47179);
nor U49175 (N_49175,N_47826,N_46175);
nor U49176 (N_49176,N_47490,N_46045);
or U49177 (N_49177,N_46783,N_47447);
nor U49178 (N_49178,N_47356,N_46633);
or U49179 (N_49179,N_46772,N_47648);
xnor U49180 (N_49180,N_46376,N_47822);
nand U49181 (N_49181,N_47417,N_47752);
xnor U49182 (N_49182,N_46587,N_46094);
or U49183 (N_49183,N_47901,N_46609);
nand U49184 (N_49184,N_46796,N_47575);
and U49185 (N_49185,N_47615,N_46451);
nand U49186 (N_49186,N_46068,N_47381);
or U49187 (N_49187,N_46302,N_47199);
and U49188 (N_49188,N_46003,N_47911);
nand U49189 (N_49189,N_46711,N_46679);
nor U49190 (N_49190,N_47915,N_46705);
nand U49191 (N_49191,N_47086,N_46361);
and U49192 (N_49192,N_46793,N_46514);
and U49193 (N_49193,N_47927,N_47393);
or U49194 (N_49194,N_47332,N_47879);
and U49195 (N_49195,N_47617,N_46869);
or U49196 (N_49196,N_47902,N_46445);
nor U49197 (N_49197,N_46881,N_47972);
xor U49198 (N_49198,N_46195,N_46491);
nand U49199 (N_49199,N_47442,N_47127);
and U49200 (N_49200,N_46038,N_46515);
nand U49201 (N_49201,N_47558,N_46189);
nor U49202 (N_49202,N_47350,N_47936);
or U49203 (N_49203,N_46424,N_47082);
nor U49204 (N_49204,N_46753,N_47569);
xnor U49205 (N_49205,N_47141,N_47541);
nor U49206 (N_49206,N_46788,N_47530);
nor U49207 (N_49207,N_47122,N_46168);
nor U49208 (N_49208,N_46874,N_47147);
and U49209 (N_49209,N_46333,N_47315);
or U49210 (N_49210,N_46772,N_47707);
nand U49211 (N_49211,N_47928,N_46154);
nor U49212 (N_49212,N_47073,N_46306);
nand U49213 (N_49213,N_47429,N_47363);
and U49214 (N_49214,N_47245,N_46267);
xnor U49215 (N_49215,N_46248,N_46136);
nor U49216 (N_49216,N_46519,N_47968);
nand U49217 (N_49217,N_46073,N_46017);
xor U49218 (N_49218,N_47370,N_46098);
xnor U49219 (N_49219,N_46671,N_46715);
or U49220 (N_49220,N_46183,N_46523);
nand U49221 (N_49221,N_47582,N_47875);
nand U49222 (N_49222,N_47209,N_47884);
or U49223 (N_49223,N_46700,N_47724);
or U49224 (N_49224,N_46743,N_46227);
xor U49225 (N_49225,N_46764,N_46878);
and U49226 (N_49226,N_47011,N_46730);
nand U49227 (N_49227,N_47144,N_47046);
or U49228 (N_49228,N_46145,N_47714);
xor U49229 (N_49229,N_47868,N_46495);
or U49230 (N_49230,N_46501,N_46818);
or U49231 (N_49231,N_47656,N_47740);
nor U49232 (N_49232,N_47448,N_46944);
nor U49233 (N_49233,N_46708,N_47715);
xnor U49234 (N_49234,N_46873,N_47740);
xnor U49235 (N_49235,N_46331,N_46668);
and U49236 (N_49236,N_47694,N_47228);
xnor U49237 (N_49237,N_46815,N_47806);
nand U49238 (N_49238,N_47927,N_47066);
or U49239 (N_49239,N_47220,N_47959);
and U49240 (N_49240,N_47966,N_46394);
or U49241 (N_49241,N_47770,N_46690);
xnor U49242 (N_49242,N_46120,N_46453);
or U49243 (N_49243,N_46337,N_47958);
nor U49244 (N_49244,N_46365,N_47828);
nor U49245 (N_49245,N_46160,N_46166);
nand U49246 (N_49246,N_47757,N_47258);
nor U49247 (N_49247,N_46505,N_46698);
xor U49248 (N_49248,N_46142,N_46850);
or U49249 (N_49249,N_47951,N_46931);
nand U49250 (N_49250,N_47111,N_47533);
or U49251 (N_49251,N_47932,N_46285);
or U49252 (N_49252,N_47093,N_47726);
nor U49253 (N_49253,N_46782,N_46663);
nor U49254 (N_49254,N_47677,N_47466);
nor U49255 (N_49255,N_47535,N_47245);
or U49256 (N_49256,N_46178,N_47991);
nor U49257 (N_49257,N_47895,N_47456);
xor U49258 (N_49258,N_46590,N_46265);
nor U49259 (N_49259,N_47652,N_47359);
and U49260 (N_49260,N_47206,N_47716);
and U49261 (N_49261,N_46847,N_47294);
nor U49262 (N_49262,N_47801,N_47177);
xor U49263 (N_49263,N_46730,N_47295);
xnor U49264 (N_49264,N_46726,N_46080);
xor U49265 (N_49265,N_46210,N_47149);
xnor U49266 (N_49266,N_46912,N_47810);
nor U49267 (N_49267,N_47348,N_47587);
nor U49268 (N_49268,N_46759,N_46197);
or U49269 (N_49269,N_46042,N_46979);
and U49270 (N_49270,N_47380,N_46678);
and U49271 (N_49271,N_47073,N_46896);
and U49272 (N_49272,N_46687,N_47308);
nand U49273 (N_49273,N_46067,N_47954);
or U49274 (N_49274,N_46844,N_47831);
or U49275 (N_49275,N_46528,N_46703);
and U49276 (N_49276,N_47099,N_47145);
nand U49277 (N_49277,N_46926,N_46585);
nand U49278 (N_49278,N_46054,N_47400);
nor U49279 (N_49279,N_47047,N_47915);
or U49280 (N_49280,N_47470,N_46101);
nand U49281 (N_49281,N_47370,N_46023);
xor U49282 (N_49282,N_47763,N_46171);
nand U49283 (N_49283,N_46907,N_47139);
nand U49284 (N_49284,N_46190,N_46074);
nor U49285 (N_49285,N_47191,N_46809);
nor U49286 (N_49286,N_46266,N_46882);
and U49287 (N_49287,N_47929,N_47040);
and U49288 (N_49288,N_46580,N_47555);
or U49289 (N_49289,N_47485,N_47835);
xor U49290 (N_49290,N_46308,N_47970);
nor U49291 (N_49291,N_46310,N_46118);
and U49292 (N_49292,N_46758,N_46597);
and U49293 (N_49293,N_47024,N_47045);
nand U49294 (N_49294,N_46737,N_46239);
xor U49295 (N_49295,N_47052,N_46842);
or U49296 (N_49296,N_47547,N_47270);
xnor U49297 (N_49297,N_47360,N_47435);
and U49298 (N_49298,N_46543,N_46147);
nand U49299 (N_49299,N_47881,N_46417);
and U49300 (N_49300,N_46033,N_47973);
xor U49301 (N_49301,N_47155,N_46705);
nand U49302 (N_49302,N_47199,N_47707);
xor U49303 (N_49303,N_47736,N_46503);
nor U49304 (N_49304,N_47549,N_46128);
nor U49305 (N_49305,N_46440,N_47155);
nor U49306 (N_49306,N_46644,N_46114);
xor U49307 (N_49307,N_46428,N_47426);
or U49308 (N_49308,N_46283,N_46551);
or U49309 (N_49309,N_46837,N_47122);
nand U49310 (N_49310,N_47865,N_47209);
xor U49311 (N_49311,N_47887,N_46311);
and U49312 (N_49312,N_47121,N_47475);
nor U49313 (N_49313,N_47790,N_46822);
nor U49314 (N_49314,N_47091,N_47076);
nand U49315 (N_49315,N_47953,N_47970);
or U49316 (N_49316,N_46245,N_47176);
xnor U49317 (N_49317,N_46623,N_46825);
and U49318 (N_49318,N_46568,N_46898);
and U49319 (N_49319,N_47363,N_46010);
nand U49320 (N_49320,N_47815,N_47131);
or U49321 (N_49321,N_46483,N_47041);
and U49322 (N_49322,N_46782,N_47821);
xnor U49323 (N_49323,N_46354,N_46877);
nor U49324 (N_49324,N_46093,N_47058);
nor U49325 (N_49325,N_47002,N_47515);
or U49326 (N_49326,N_47254,N_47736);
or U49327 (N_49327,N_46939,N_47721);
nand U49328 (N_49328,N_46178,N_47637);
or U49329 (N_49329,N_46043,N_46914);
xnor U49330 (N_49330,N_46346,N_47760);
and U49331 (N_49331,N_47618,N_47005);
xor U49332 (N_49332,N_47742,N_46254);
and U49333 (N_49333,N_47812,N_47438);
nand U49334 (N_49334,N_47058,N_46762);
nor U49335 (N_49335,N_47770,N_46090);
and U49336 (N_49336,N_47616,N_46531);
and U49337 (N_49337,N_46965,N_47208);
nor U49338 (N_49338,N_46645,N_46812);
or U49339 (N_49339,N_46481,N_47052);
nor U49340 (N_49340,N_46348,N_47279);
xnor U49341 (N_49341,N_46899,N_46455);
xnor U49342 (N_49342,N_47265,N_47718);
or U49343 (N_49343,N_46880,N_46554);
nand U49344 (N_49344,N_46220,N_47348);
nand U49345 (N_49345,N_47970,N_47309);
and U49346 (N_49346,N_47791,N_47674);
xnor U49347 (N_49347,N_47356,N_47563);
nor U49348 (N_49348,N_47116,N_46639);
xnor U49349 (N_49349,N_47971,N_46521);
xor U49350 (N_49350,N_46604,N_47123);
and U49351 (N_49351,N_46379,N_47516);
or U49352 (N_49352,N_47433,N_47686);
xor U49353 (N_49353,N_47638,N_46721);
or U49354 (N_49354,N_47689,N_46583);
xor U49355 (N_49355,N_46633,N_46733);
nand U49356 (N_49356,N_46154,N_47814);
nand U49357 (N_49357,N_46824,N_46404);
nand U49358 (N_49358,N_46509,N_46890);
nand U49359 (N_49359,N_46521,N_47600);
xor U49360 (N_49360,N_47318,N_46859);
or U49361 (N_49361,N_47235,N_47278);
and U49362 (N_49362,N_46540,N_46074);
and U49363 (N_49363,N_46780,N_47611);
nor U49364 (N_49364,N_47955,N_46361);
nor U49365 (N_49365,N_47496,N_47660);
or U49366 (N_49366,N_47436,N_47178);
nand U49367 (N_49367,N_47014,N_47686);
and U49368 (N_49368,N_46937,N_47570);
xnor U49369 (N_49369,N_47057,N_46288);
and U49370 (N_49370,N_46708,N_47017);
nor U49371 (N_49371,N_46495,N_47987);
nor U49372 (N_49372,N_46247,N_47715);
nor U49373 (N_49373,N_46612,N_47436);
xor U49374 (N_49374,N_46664,N_46673);
xor U49375 (N_49375,N_47993,N_47556);
or U49376 (N_49376,N_47347,N_46559);
nand U49377 (N_49377,N_46465,N_47669);
or U49378 (N_49378,N_47745,N_47238);
and U49379 (N_49379,N_47777,N_47130);
nor U49380 (N_49380,N_47341,N_47780);
and U49381 (N_49381,N_47536,N_47203);
or U49382 (N_49382,N_47448,N_47606);
nor U49383 (N_49383,N_47010,N_46563);
xnor U49384 (N_49384,N_47787,N_47544);
nor U49385 (N_49385,N_47900,N_47143);
nand U49386 (N_49386,N_47136,N_46810);
xnor U49387 (N_49387,N_47593,N_47913);
nor U49388 (N_49388,N_46217,N_46834);
or U49389 (N_49389,N_46995,N_46858);
and U49390 (N_49390,N_47864,N_47197);
or U49391 (N_49391,N_46056,N_46856);
nand U49392 (N_49392,N_47505,N_46346);
or U49393 (N_49393,N_47040,N_46067);
xnor U49394 (N_49394,N_47868,N_46429);
or U49395 (N_49395,N_47211,N_47286);
xor U49396 (N_49396,N_46556,N_47366);
xnor U49397 (N_49397,N_46122,N_47255);
or U49398 (N_49398,N_46453,N_46800);
xor U49399 (N_49399,N_47547,N_47070);
or U49400 (N_49400,N_47565,N_47598);
nand U49401 (N_49401,N_46924,N_47318);
or U49402 (N_49402,N_47971,N_46885);
xnor U49403 (N_49403,N_47098,N_46205);
or U49404 (N_49404,N_46784,N_47714);
nand U49405 (N_49405,N_47681,N_47801);
nand U49406 (N_49406,N_47883,N_46986);
or U49407 (N_49407,N_46803,N_46800);
nor U49408 (N_49408,N_46228,N_47312);
nor U49409 (N_49409,N_47179,N_47437);
nor U49410 (N_49410,N_46337,N_47814);
or U49411 (N_49411,N_46920,N_46586);
or U49412 (N_49412,N_47389,N_46405);
nor U49413 (N_49413,N_46444,N_46793);
xnor U49414 (N_49414,N_46480,N_47480);
nand U49415 (N_49415,N_46809,N_46063);
or U49416 (N_49416,N_46168,N_47519);
and U49417 (N_49417,N_46148,N_46060);
xnor U49418 (N_49418,N_47837,N_46715);
nor U49419 (N_49419,N_46615,N_46587);
xnor U49420 (N_49420,N_46026,N_46354);
nor U49421 (N_49421,N_46011,N_47643);
nand U49422 (N_49422,N_46250,N_46016);
xnor U49423 (N_49423,N_47110,N_47157);
xor U49424 (N_49424,N_46057,N_46134);
or U49425 (N_49425,N_46146,N_46974);
and U49426 (N_49426,N_46820,N_46604);
nand U49427 (N_49427,N_46232,N_46557);
nand U49428 (N_49428,N_47799,N_46526);
xor U49429 (N_49429,N_46274,N_47119);
nor U49430 (N_49430,N_47867,N_47906);
xor U49431 (N_49431,N_47570,N_47829);
nand U49432 (N_49432,N_47932,N_46008);
nor U49433 (N_49433,N_46126,N_47358);
or U49434 (N_49434,N_46896,N_47561);
nand U49435 (N_49435,N_46904,N_47799);
or U49436 (N_49436,N_47641,N_46004);
or U49437 (N_49437,N_46795,N_46686);
nand U49438 (N_49438,N_46783,N_47296);
xnor U49439 (N_49439,N_46268,N_46547);
xor U49440 (N_49440,N_47258,N_46920);
and U49441 (N_49441,N_46365,N_47389);
nor U49442 (N_49442,N_47903,N_47642);
or U49443 (N_49443,N_46868,N_46507);
nor U49444 (N_49444,N_46790,N_47269);
nor U49445 (N_49445,N_46329,N_47200);
nand U49446 (N_49446,N_46457,N_46831);
xnor U49447 (N_49447,N_47031,N_47631);
xnor U49448 (N_49448,N_47382,N_47379);
and U49449 (N_49449,N_46134,N_46804);
or U49450 (N_49450,N_47996,N_47031);
xnor U49451 (N_49451,N_46806,N_46593);
nor U49452 (N_49452,N_46440,N_46782);
or U49453 (N_49453,N_46954,N_46951);
nor U49454 (N_49454,N_46099,N_47870);
or U49455 (N_49455,N_47591,N_46035);
xor U49456 (N_49456,N_47528,N_46967);
nand U49457 (N_49457,N_46320,N_47989);
or U49458 (N_49458,N_46361,N_46883);
nor U49459 (N_49459,N_47219,N_46874);
xor U49460 (N_49460,N_46771,N_46496);
nor U49461 (N_49461,N_47998,N_46549);
xnor U49462 (N_49462,N_47127,N_47712);
xor U49463 (N_49463,N_47676,N_46248);
nor U49464 (N_49464,N_47741,N_46016);
or U49465 (N_49465,N_46548,N_47339);
xnor U49466 (N_49466,N_46430,N_46963);
nor U49467 (N_49467,N_47284,N_46809);
and U49468 (N_49468,N_47400,N_46107);
xnor U49469 (N_49469,N_46411,N_46711);
nand U49470 (N_49470,N_47214,N_47044);
or U49471 (N_49471,N_47781,N_46338);
xor U49472 (N_49472,N_46479,N_47240);
xor U49473 (N_49473,N_47830,N_46298);
nand U49474 (N_49474,N_47746,N_46953);
nor U49475 (N_49475,N_46283,N_46229);
nand U49476 (N_49476,N_47798,N_46217);
nor U49477 (N_49477,N_46973,N_47027);
and U49478 (N_49478,N_46570,N_46545);
nor U49479 (N_49479,N_46710,N_46688);
nand U49480 (N_49480,N_47642,N_46442);
nand U49481 (N_49481,N_46250,N_46756);
or U49482 (N_49482,N_46309,N_47065);
xor U49483 (N_49483,N_47851,N_47429);
xnor U49484 (N_49484,N_47533,N_47428);
nand U49485 (N_49485,N_47800,N_47403);
nand U49486 (N_49486,N_47345,N_46391);
nand U49487 (N_49487,N_47122,N_46068);
nand U49488 (N_49488,N_46400,N_47217);
or U49489 (N_49489,N_47806,N_47487);
or U49490 (N_49490,N_47219,N_46251);
nand U49491 (N_49491,N_47402,N_47149);
and U49492 (N_49492,N_47665,N_46384);
or U49493 (N_49493,N_46822,N_47679);
nor U49494 (N_49494,N_46666,N_46286);
or U49495 (N_49495,N_47214,N_46242);
xor U49496 (N_49496,N_47037,N_46081);
nor U49497 (N_49497,N_46791,N_46998);
or U49498 (N_49498,N_46240,N_47132);
nor U49499 (N_49499,N_47590,N_47938);
or U49500 (N_49500,N_47319,N_46140);
nor U49501 (N_49501,N_47340,N_46930);
nand U49502 (N_49502,N_47892,N_46030);
nor U49503 (N_49503,N_46814,N_46746);
or U49504 (N_49504,N_46287,N_46546);
nand U49505 (N_49505,N_47576,N_46183);
or U49506 (N_49506,N_47825,N_47414);
or U49507 (N_49507,N_47076,N_46506);
nand U49508 (N_49508,N_47090,N_46972);
xnor U49509 (N_49509,N_47460,N_47905);
nor U49510 (N_49510,N_46100,N_47191);
or U49511 (N_49511,N_47724,N_47601);
nor U49512 (N_49512,N_47505,N_47969);
xnor U49513 (N_49513,N_47216,N_46127);
nand U49514 (N_49514,N_46760,N_47936);
nor U49515 (N_49515,N_47067,N_46780);
xnor U49516 (N_49516,N_46802,N_47755);
nand U49517 (N_49517,N_46873,N_46659);
xor U49518 (N_49518,N_47235,N_46290);
nor U49519 (N_49519,N_47384,N_47165);
xor U49520 (N_49520,N_47985,N_46916);
nand U49521 (N_49521,N_46882,N_46716);
nand U49522 (N_49522,N_47466,N_46933);
nor U49523 (N_49523,N_46956,N_46162);
and U49524 (N_49524,N_46818,N_46308);
nor U49525 (N_49525,N_47959,N_47498);
nor U49526 (N_49526,N_47167,N_46459);
or U49527 (N_49527,N_47385,N_47086);
nand U49528 (N_49528,N_47547,N_46516);
xor U49529 (N_49529,N_47850,N_47969);
and U49530 (N_49530,N_47712,N_47241);
nand U49531 (N_49531,N_46088,N_46585);
xor U49532 (N_49532,N_46791,N_46207);
and U49533 (N_49533,N_46672,N_47460);
xnor U49534 (N_49534,N_47949,N_47864);
xor U49535 (N_49535,N_47201,N_47503);
nand U49536 (N_49536,N_47179,N_46126);
nor U49537 (N_49537,N_46622,N_46570);
and U49538 (N_49538,N_47001,N_46255);
xnor U49539 (N_49539,N_47644,N_46229);
nor U49540 (N_49540,N_46206,N_46930);
xor U49541 (N_49541,N_47626,N_46495);
xnor U49542 (N_49542,N_46542,N_47589);
nor U49543 (N_49543,N_46804,N_46050);
nor U49544 (N_49544,N_47307,N_46292);
or U49545 (N_49545,N_47606,N_47308);
and U49546 (N_49546,N_47237,N_47299);
or U49547 (N_49547,N_46667,N_47647);
nor U49548 (N_49548,N_46142,N_47992);
nand U49549 (N_49549,N_47702,N_46939);
or U49550 (N_49550,N_47072,N_46937);
nand U49551 (N_49551,N_47807,N_47826);
nor U49552 (N_49552,N_46939,N_46326);
nand U49553 (N_49553,N_47488,N_46949);
xnor U49554 (N_49554,N_47475,N_47847);
and U49555 (N_49555,N_47236,N_47498);
nor U49556 (N_49556,N_46836,N_47752);
or U49557 (N_49557,N_47825,N_46946);
or U49558 (N_49558,N_47241,N_46327);
nor U49559 (N_49559,N_46681,N_46111);
nand U49560 (N_49560,N_47855,N_47838);
nor U49561 (N_49561,N_46801,N_46709);
nand U49562 (N_49562,N_47687,N_47327);
xnor U49563 (N_49563,N_46629,N_46079);
nor U49564 (N_49564,N_46886,N_47132);
or U49565 (N_49565,N_46360,N_47054);
xnor U49566 (N_49566,N_47046,N_46556);
and U49567 (N_49567,N_47067,N_46246);
nor U49568 (N_49568,N_46620,N_47978);
or U49569 (N_49569,N_46392,N_47638);
nor U49570 (N_49570,N_47129,N_46710);
nand U49571 (N_49571,N_47117,N_46544);
nand U49572 (N_49572,N_47534,N_46421);
xnor U49573 (N_49573,N_47810,N_47163);
nor U49574 (N_49574,N_47605,N_47887);
nor U49575 (N_49575,N_47484,N_46401);
xor U49576 (N_49576,N_46409,N_46050);
and U49577 (N_49577,N_47183,N_47656);
xor U49578 (N_49578,N_46576,N_47821);
and U49579 (N_49579,N_47794,N_46621);
xnor U49580 (N_49580,N_47134,N_47849);
or U49581 (N_49581,N_47992,N_47575);
or U49582 (N_49582,N_47180,N_47256);
xnor U49583 (N_49583,N_46905,N_47747);
and U49584 (N_49584,N_46491,N_47875);
nor U49585 (N_49585,N_47585,N_47201);
or U49586 (N_49586,N_46995,N_47258);
and U49587 (N_49587,N_47290,N_47579);
nor U49588 (N_49588,N_46269,N_46592);
xnor U49589 (N_49589,N_46207,N_46309);
or U49590 (N_49590,N_46987,N_47519);
or U49591 (N_49591,N_47204,N_47148);
and U49592 (N_49592,N_47616,N_47666);
xnor U49593 (N_49593,N_46745,N_46395);
nor U49594 (N_49594,N_47516,N_46474);
nand U49595 (N_49595,N_47206,N_47117);
nand U49596 (N_49596,N_47138,N_46630);
nor U49597 (N_49597,N_46161,N_46691);
xnor U49598 (N_49598,N_46685,N_47182);
or U49599 (N_49599,N_47442,N_47829);
nand U49600 (N_49600,N_47880,N_46829);
or U49601 (N_49601,N_46244,N_47519);
or U49602 (N_49602,N_47531,N_46748);
and U49603 (N_49603,N_46870,N_47701);
xnor U49604 (N_49604,N_47697,N_47965);
and U49605 (N_49605,N_47164,N_46674);
xor U49606 (N_49606,N_47401,N_46438);
or U49607 (N_49607,N_46364,N_47881);
or U49608 (N_49608,N_47333,N_47409);
and U49609 (N_49609,N_47442,N_46194);
nand U49610 (N_49610,N_47588,N_47528);
nand U49611 (N_49611,N_47038,N_47768);
or U49612 (N_49612,N_46312,N_47010);
nand U49613 (N_49613,N_47154,N_47543);
nor U49614 (N_49614,N_47637,N_47066);
nand U49615 (N_49615,N_46471,N_47976);
xnor U49616 (N_49616,N_47071,N_46961);
nor U49617 (N_49617,N_47379,N_46527);
or U49618 (N_49618,N_46420,N_46162);
or U49619 (N_49619,N_46943,N_47088);
nor U49620 (N_49620,N_47748,N_47485);
nor U49621 (N_49621,N_46673,N_47210);
xnor U49622 (N_49622,N_46252,N_47284);
nand U49623 (N_49623,N_47321,N_47792);
nor U49624 (N_49624,N_46086,N_46571);
or U49625 (N_49625,N_47463,N_46644);
nand U49626 (N_49626,N_46256,N_47085);
xor U49627 (N_49627,N_46356,N_46184);
or U49628 (N_49628,N_47492,N_46941);
nand U49629 (N_49629,N_47842,N_47697);
xor U49630 (N_49630,N_47498,N_46403);
or U49631 (N_49631,N_47289,N_47520);
and U49632 (N_49632,N_47887,N_47017);
nor U49633 (N_49633,N_47521,N_46435);
nor U49634 (N_49634,N_47262,N_46067);
nor U49635 (N_49635,N_47400,N_47554);
or U49636 (N_49636,N_46809,N_47438);
or U49637 (N_49637,N_47546,N_46849);
nor U49638 (N_49638,N_46765,N_46706);
and U49639 (N_49639,N_46128,N_47042);
and U49640 (N_49640,N_46588,N_46098);
xor U49641 (N_49641,N_47726,N_47196);
nor U49642 (N_49642,N_46627,N_46495);
nand U49643 (N_49643,N_46672,N_47716);
or U49644 (N_49644,N_46776,N_47635);
or U49645 (N_49645,N_47473,N_47488);
nor U49646 (N_49646,N_46306,N_47279);
nor U49647 (N_49647,N_46144,N_46690);
xnor U49648 (N_49648,N_47246,N_46017);
and U49649 (N_49649,N_46448,N_47469);
xor U49650 (N_49650,N_47680,N_47659);
and U49651 (N_49651,N_47190,N_47188);
nand U49652 (N_49652,N_47083,N_47224);
nand U49653 (N_49653,N_47215,N_47033);
or U49654 (N_49654,N_47718,N_47487);
and U49655 (N_49655,N_47128,N_46318);
or U49656 (N_49656,N_46559,N_47770);
or U49657 (N_49657,N_47946,N_46839);
xor U49658 (N_49658,N_46359,N_46027);
nor U49659 (N_49659,N_46352,N_46684);
nand U49660 (N_49660,N_46948,N_46778);
xnor U49661 (N_49661,N_46804,N_46178);
xor U49662 (N_49662,N_47704,N_46090);
nand U49663 (N_49663,N_47277,N_46411);
nor U49664 (N_49664,N_46780,N_47805);
nand U49665 (N_49665,N_47769,N_47785);
and U49666 (N_49666,N_46397,N_46890);
and U49667 (N_49667,N_47128,N_46810);
and U49668 (N_49668,N_47650,N_47882);
or U49669 (N_49669,N_46273,N_47541);
or U49670 (N_49670,N_47540,N_47182);
xor U49671 (N_49671,N_47823,N_47300);
and U49672 (N_49672,N_46238,N_47313);
and U49673 (N_49673,N_46845,N_46561);
nand U49674 (N_49674,N_47637,N_46133);
or U49675 (N_49675,N_47431,N_47890);
nor U49676 (N_49676,N_46128,N_46576);
and U49677 (N_49677,N_47443,N_47024);
nand U49678 (N_49678,N_47337,N_47632);
nor U49679 (N_49679,N_46777,N_46184);
nor U49680 (N_49680,N_46832,N_46239);
nor U49681 (N_49681,N_46704,N_47624);
nor U49682 (N_49682,N_46851,N_46075);
or U49683 (N_49683,N_47366,N_47407);
xnor U49684 (N_49684,N_46427,N_46958);
or U49685 (N_49685,N_46867,N_46298);
and U49686 (N_49686,N_46312,N_46540);
or U49687 (N_49687,N_47984,N_46990);
or U49688 (N_49688,N_47515,N_46092);
xnor U49689 (N_49689,N_47735,N_46399);
nor U49690 (N_49690,N_46045,N_46061);
xnor U49691 (N_49691,N_47069,N_47330);
or U49692 (N_49692,N_47640,N_46271);
nand U49693 (N_49693,N_46065,N_47034);
or U49694 (N_49694,N_47295,N_47116);
and U49695 (N_49695,N_46753,N_47523);
or U49696 (N_49696,N_46474,N_46510);
xnor U49697 (N_49697,N_46251,N_46677);
and U49698 (N_49698,N_46618,N_46557);
nor U49699 (N_49699,N_47094,N_46252);
nor U49700 (N_49700,N_46565,N_46864);
nor U49701 (N_49701,N_46219,N_47098);
xnor U49702 (N_49702,N_46792,N_46557);
or U49703 (N_49703,N_47847,N_47146);
and U49704 (N_49704,N_46534,N_47889);
nor U49705 (N_49705,N_46594,N_47778);
or U49706 (N_49706,N_47538,N_46525);
and U49707 (N_49707,N_47901,N_47322);
nor U49708 (N_49708,N_47668,N_47308);
or U49709 (N_49709,N_47711,N_46860);
nand U49710 (N_49710,N_46075,N_46035);
nand U49711 (N_49711,N_47801,N_46257);
and U49712 (N_49712,N_47160,N_46755);
or U49713 (N_49713,N_47050,N_47804);
xor U49714 (N_49714,N_46433,N_47369);
or U49715 (N_49715,N_46531,N_46305);
nand U49716 (N_49716,N_47019,N_47692);
or U49717 (N_49717,N_46966,N_46954);
or U49718 (N_49718,N_46217,N_46742);
xnor U49719 (N_49719,N_47337,N_47445);
xnor U49720 (N_49720,N_46997,N_47168);
nor U49721 (N_49721,N_46094,N_47062);
xor U49722 (N_49722,N_46233,N_46929);
xnor U49723 (N_49723,N_46152,N_46991);
nand U49724 (N_49724,N_46834,N_47033);
nor U49725 (N_49725,N_46769,N_46559);
nand U49726 (N_49726,N_46763,N_46193);
or U49727 (N_49727,N_46909,N_47555);
nand U49728 (N_49728,N_47980,N_46555);
xnor U49729 (N_49729,N_47457,N_47981);
and U49730 (N_49730,N_46867,N_47621);
nand U49731 (N_49731,N_47500,N_47757);
or U49732 (N_49732,N_47616,N_46607);
or U49733 (N_49733,N_47247,N_47033);
nor U49734 (N_49734,N_47169,N_46559);
nor U49735 (N_49735,N_46333,N_47283);
xor U49736 (N_49736,N_46526,N_47471);
nand U49737 (N_49737,N_46332,N_47600);
nor U49738 (N_49738,N_47486,N_47985);
nor U49739 (N_49739,N_47399,N_47193);
xor U49740 (N_49740,N_46634,N_47145);
xor U49741 (N_49741,N_46767,N_46246);
nor U49742 (N_49742,N_47231,N_46963);
nor U49743 (N_49743,N_46091,N_47057);
or U49744 (N_49744,N_46036,N_47406);
nand U49745 (N_49745,N_47117,N_46919);
nor U49746 (N_49746,N_46505,N_46583);
and U49747 (N_49747,N_47827,N_46129);
or U49748 (N_49748,N_47632,N_46119);
xnor U49749 (N_49749,N_47608,N_47989);
or U49750 (N_49750,N_46589,N_46477);
nor U49751 (N_49751,N_47550,N_47599);
xor U49752 (N_49752,N_46032,N_46583);
nand U49753 (N_49753,N_47891,N_46569);
or U49754 (N_49754,N_47607,N_47198);
xor U49755 (N_49755,N_46746,N_47476);
nor U49756 (N_49756,N_47409,N_47279);
or U49757 (N_49757,N_46114,N_47435);
and U49758 (N_49758,N_47292,N_46741);
xor U49759 (N_49759,N_47141,N_47705);
or U49760 (N_49760,N_46965,N_47124);
nor U49761 (N_49761,N_46238,N_47030);
nor U49762 (N_49762,N_47360,N_47810);
xnor U49763 (N_49763,N_46344,N_46790);
nand U49764 (N_49764,N_46919,N_47834);
nor U49765 (N_49765,N_46381,N_46715);
xor U49766 (N_49766,N_47788,N_47060);
nor U49767 (N_49767,N_46726,N_47618);
and U49768 (N_49768,N_46915,N_47274);
or U49769 (N_49769,N_47731,N_46342);
nand U49770 (N_49770,N_46399,N_47988);
or U49771 (N_49771,N_46576,N_47518);
or U49772 (N_49772,N_47264,N_46671);
nand U49773 (N_49773,N_46918,N_46188);
and U49774 (N_49774,N_47605,N_46020);
and U49775 (N_49775,N_46340,N_47680);
or U49776 (N_49776,N_47525,N_47789);
and U49777 (N_49777,N_47354,N_47919);
or U49778 (N_49778,N_46634,N_46769);
nor U49779 (N_49779,N_47431,N_46895);
and U49780 (N_49780,N_47066,N_47572);
and U49781 (N_49781,N_47338,N_47745);
xnor U49782 (N_49782,N_47321,N_46926);
and U49783 (N_49783,N_46620,N_47383);
nor U49784 (N_49784,N_46374,N_46465);
nor U49785 (N_49785,N_46023,N_47485);
xor U49786 (N_49786,N_47166,N_47109);
nand U49787 (N_49787,N_47851,N_47645);
or U49788 (N_49788,N_47423,N_47251);
nor U49789 (N_49789,N_46144,N_46999);
nand U49790 (N_49790,N_46613,N_47160);
nor U49791 (N_49791,N_47621,N_47187);
nor U49792 (N_49792,N_46106,N_46318);
xnor U49793 (N_49793,N_46320,N_47890);
nor U49794 (N_49794,N_47533,N_47019);
or U49795 (N_49795,N_47863,N_46371);
nor U49796 (N_49796,N_47033,N_47498);
xnor U49797 (N_49797,N_46988,N_47475);
and U49798 (N_49798,N_46565,N_46934);
and U49799 (N_49799,N_47950,N_47871);
or U49800 (N_49800,N_46785,N_46243);
or U49801 (N_49801,N_47823,N_47596);
nand U49802 (N_49802,N_46325,N_46806);
or U49803 (N_49803,N_46426,N_46762);
nor U49804 (N_49804,N_46341,N_47323);
or U49805 (N_49805,N_46485,N_46984);
nand U49806 (N_49806,N_46217,N_47421);
nor U49807 (N_49807,N_46874,N_47824);
and U49808 (N_49808,N_46412,N_47442);
nand U49809 (N_49809,N_46258,N_47834);
and U49810 (N_49810,N_46561,N_46620);
or U49811 (N_49811,N_47378,N_47705);
nor U49812 (N_49812,N_47840,N_47016);
or U49813 (N_49813,N_46779,N_47473);
xor U49814 (N_49814,N_46071,N_46148);
nor U49815 (N_49815,N_47155,N_46182);
or U49816 (N_49816,N_46947,N_47780);
and U49817 (N_49817,N_47415,N_46278);
nor U49818 (N_49818,N_46825,N_47960);
nor U49819 (N_49819,N_47230,N_46665);
or U49820 (N_49820,N_46765,N_47948);
and U49821 (N_49821,N_47288,N_47496);
and U49822 (N_49822,N_47889,N_47691);
nand U49823 (N_49823,N_47443,N_46079);
nor U49824 (N_49824,N_47982,N_47760);
and U49825 (N_49825,N_46279,N_47728);
and U49826 (N_49826,N_46274,N_46525);
xnor U49827 (N_49827,N_47125,N_47938);
xor U49828 (N_49828,N_46883,N_46363);
nor U49829 (N_49829,N_46229,N_47326);
or U49830 (N_49830,N_47203,N_46336);
nand U49831 (N_49831,N_46880,N_46591);
and U49832 (N_49832,N_46435,N_46549);
nand U49833 (N_49833,N_47170,N_46605);
or U49834 (N_49834,N_46441,N_47754);
nand U49835 (N_49835,N_46088,N_47518);
and U49836 (N_49836,N_47476,N_46461);
xnor U49837 (N_49837,N_46552,N_47176);
or U49838 (N_49838,N_47318,N_47069);
or U49839 (N_49839,N_46307,N_46074);
nand U49840 (N_49840,N_46635,N_46268);
and U49841 (N_49841,N_47402,N_46972);
or U49842 (N_49842,N_47390,N_46316);
nand U49843 (N_49843,N_46765,N_46512);
nand U49844 (N_49844,N_47556,N_46782);
nand U49845 (N_49845,N_46561,N_47864);
or U49846 (N_49846,N_47449,N_46780);
xor U49847 (N_49847,N_46559,N_46350);
nand U49848 (N_49848,N_46654,N_47239);
xnor U49849 (N_49849,N_46754,N_46337);
or U49850 (N_49850,N_47430,N_46215);
and U49851 (N_49851,N_46158,N_46913);
and U49852 (N_49852,N_46021,N_47243);
nand U49853 (N_49853,N_46804,N_46373);
and U49854 (N_49854,N_47539,N_47742);
or U49855 (N_49855,N_47030,N_47412);
or U49856 (N_49856,N_47629,N_47088);
or U49857 (N_49857,N_46789,N_47592);
or U49858 (N_49858,N_46800,N_46994);
xor U49859 (N_49859,N_46715,N_46450);
and U49860 (N_49860,N_47584,N_46813);
xnor U49861 (N_49861,N_47627,N_46307);
xnor U49862 (N_49862,N_47530,N_46116);
and U49863 (N_49863,N_47492,N_47692);
nand U49864 (N_49864,N_47104,N_46561);
and U49865 (N_49865,N_47309,N_46806);
or U49866 (N_49866,N_47210,N_46391);
and U49867 (N_49867,N_47172,N_47641);
and U49868 (N_49868,N_47704,N_46874);
nand U49869 (N_49869,N_47286,N_47096);
xnor U49870 (N_49870,N_46613,N_47013);
nand U49871 (N_49871,N_47799,N_47821);
and U49872 (N_49872,N_46898,N_47605);
nor U49873 (N_49873,N_47639,N_46204);
nand U49874 (N_49874,N_46419,N_46128);
xor U49875 (N_49875,N_47224,N_46074);
and U49876 (N_49876,N_47947,N_47958);
nor U49877 (N_49877,N_46203,N_47396);
xor U49878 (N_49878,N_46432,N_46139);
or U49879 (N_49879,N_47321,N_47900);
nand U49880 (N_49880,N_47009,N_46149);
xnor U49881 (N_49881,N_46369,N_46949);
nand U49882 (N_49882,N_47967,N_47425);
and U49883 (N_49883,N_47405,N_46764);
xor U49884 (N_49884,N_46128,N_47130);
nand U49885 (N_49885,N_47801,N_46883);
nand U49886 (N_49886,N_46019,N_46704);
nand U49887 (N_49887,N_46235,N_46431);
and U49888 (N_49888,N_46805,N_47506);
and U49889 (N_49889,N_46301,N_46573);
and U49890 (N_49890,N_47537,N_47535);
nand U49891 (N_49891,N_47675,N_47577);
nor U49892 (N_49892,N_46864,N_46664);
xnor U49893 (N_49893,N_46569,N_46376);
nor U49894 (N_49894,N_46645,N_46244);
nand U49895 (N_49895,N_46153,N_47903);
xnor U49896 (N_49896,N_46904,N_47711);
nand U49897 (N_49897,N_46131,N_46574);
nor U49898 (N_49898,N_47855,N_47066);
and U49899 (N_49899,N_46936,N_47887);
or U49900 (N_49900,N_46199,N_47496);
nor U49901 (N_49901,N_47890,N_47641);
xnor U49902 (N_49902,N_47515,N_47493);
xor U49903 (N_49903,N_47243,N_47038);
and U49904 (N_49904,N_46427,N_47108);
nor U49905 (N_49905,N_47038,N_47227);
nor U49906 (N_49906,N_46442,N_47926);
nand U49907 (N_49907,N_47647,N_47595);
nand U49908 (N_49908,N_47408,N_47174);
nor U49909 (N_49909,N_46554,N_46091);
and U49910 (N_49910,N_47340,N_46256);
nand U49911 (N_49911,N_47542,N_47204);
nand U49912 (N_49912,N_47943,N_47249);
nor U49913 (N_49913,N_47828,N_46213);
nor U49914 (N_49914,N_47878,N_47820);
xnor U49915 (N_49915,N_46186,N_46046);
or U49916 (N_49916,N_46678,N_47081);
and U49917 (N_49917,N_47180,N_46355);
nand U49918 (N_49918,N_47539,N_46810);
or U49919 (N_49919,N_46891,N_46442);
nand U49920 (N_49920,N_47952,N_46794);
xor U49921 (N_49921,N_46697,N_46514);
xnor U49922 (N_49922,N_46581,N_46583);
nor U49923 (N_49923,N_47565,N_47094);
or U49924 (N_49924,N_47001,N_47886);
xor U49925 (N_49925,N_46628,N_47727);
xor U49926 (N_49926,N_47821,N_47178);
and U49927 (N_49927,N_47996,N_47804);
nor U49928 (N_49928,N_47269,N_46672);
nand U49929 (N_49929,N_47048,N_47778);
nand U49930 (N_49930,N_47487,N_47920);
nor U49931 (N_49931,N_46282,N_46017);
nand U49932 (N_49932,N_47188,N_46123);
xnor U49933 (N_49933,N_47861,N_46550);
nand U49934 (N_49934,N_47325,N_46205);
or U49935 (N_49935,N_47671,N_46357);
or U49936 (N_49936,N_47415,N_47432);
and U49937 (N_49937,N_46438,N_47575);
nand U49938 (N_49938,N_46305,N_47311);
xor U49939 (N_49939,N_46641,N_46605);
nor U49940 (N_49940,N_47354,N_46993);
xor U49941 (N_49941,N_47700,N_47386);
or U49942 (N_49942,N_46938,N_47272);
or U49943 (N_49943,N_47346,N_46329);
or U49944 (N_49944,N_46568,N_46944);
nand U49945 (N_49945,N_47173,N_46026);
or U49946 (N_49946,N_46972,N_47481);
xnor U49947 (N_49947,N_46462,N_47034);
nand U49948 (N_49948,N_47374,N_47593);
or U49949 (N_49949,N_46967,N_46995);
xor U49950 (N_49950,N_46771,N_47517);
or U49951 (N_49951,N_46776,N_46286);
and U49952 (N_49952,N_46835,N_46674);
nor U49953 (N_49953,N_46322,N_46589);
or U49954 (N_49954,N_46406,N_47102);
or U49955 (N_49955,N_46871,N_47675);
or U49956 (N_49956,N_47766,N_46375);
nor U49957 (N_49957,N_47987,N_46347);
xor U49958 (N_49958,N_47751,N_46684);
or U49959 (N_49959,N_46558,N_47511);
and U49960 (N_49960,N_47075,N_46448);
or U49961 (N_49961,N_46782,N_46641);
nand U49962 (N_49962,N_47764,N_47734);
or U49963 (N_49963,N_46437,N_46115);
and U49964 (N_49964,N_47678,N_46534);
xor U49965 (N_49965,N_46483,N_47933);
nor U49966 (N_49966,N_46483,N_46542);
nand U49967 (N_49967,N_46413,N_47402);
xnor U49968 (N_49968,N_46502,N_46209);
nand U49969 (N_49969,N_46439,N_46537);
nand U49970 (N_49970,N_47097,N_47584);
nor U49971 (N_49971,N_47418,N_47877);
nand U49972 (N_49972,N_46439,N_46997);
nor U49973 (N_49973,N_47143,N_47683);
and U49974 (N_49974,N_47254,N_46295);
or U49975 (N_49975,N_46297,N_47146);
or U49976 (N_49976,N_47032,N_46317);
xnor U49977 (N_49977,N_46962,N_47215);
nand U49978 (N_49978,N_47023,N_47492);
xor U49979 (N_49979,N_47930,N_47330);
nand U49980 (N_49980,N_46794,N_47526);
and U49981 (N_49981,N_47852,N_47142);
or U49982 (N_49982,N_46346,N_47391);
and U49983 (N_49983,N_47084,N_47550);
nor U49984 (N_49984,N_46185,N_46770);
nor U49985 (N_49985,N_47697,N_46149);
xor U49986 (N_49986,N_47468,N_46779);
nand U49987 (N_49987,N_47088,N_46331);
nor U49988 (N_49988,N_46465,N_47921);
or U49989 (N_49989,N_47703,N_47118);
nor U49990 (N_49990,N_46500,N_47752);
and U49991 (N_49991,N_47093,N_47572);
nor U49992 (N_49992,N_46139,N_46740);
nor U49993 (N_49993,N_47623,N_47598);
or U49994 (N_49994,N_47804,N_46410);
nand U49995 (N_49995,N_47261,N_46970);
nor U49996 (N_49996,N_46853,N_47664);
nor U49997 (N_49997,N_46676,N_46851);
xor U49998 (N_49998,N_46845,N_47193);
and U49999 (N_49999,N_46982,N_47872);
and UO_0 (O_0,N_48468,N_49147);
nand UO_1 (O_1,N_48480,N_49710);
and UO_2 (O_2,N_49428,N_48065);
or UO_3 (O_3,N_49963,N_49016);
nand UO_4 (O_4,N_49469,N_49881);
and UO_5 (O_5,N_48129,N_48971);
and UO_6 (O_6,N_48484,N_48584);
and UO_7 (O_7,N_48016,N_48115);
and UO_8 (O_8,N_48314,N_48061);
nor UO_9 (O_9,N_48378,N_48824);
and UO_10 (O_10,N_48083,N_49411);
and UO_11 (O_11,N_48560,N_48652);
nand UO_12 (O_12,N_48568,N_48268);
xnor UO_13 (O_13,N_48470,N_48659);
and UO_14 (O_14,N_48991,N_49993);
xor UO_15 (O_15,N_48842,N_49707);
nor UO_16 (O_16,N_49197,N_49533);
or UO_17 (O_17,N_49778,N_49483);
or UO_18 (O_18,N_49275,N_48998);
nand UO_19 (O_19,N_49874,N_49090);
or UO_20 (O_20,N_48757,N_49613);
xnor UO_21 (O_21,N_49142,N_49986);
nor UO_22 (O_22,N_48653,N_49006);
and UO_23 (O_23,N_49797,N_48644);
nor UO_24 (O_24,N_49671,N_49500);
or UO_25 (O_25,N_49798,N_48994);
or UO_26 (O_26,N_49954,N_48098);
and UO_27 (O_27,N_48395,N_48849);
xnor UO_28 (O_28,N_49650,N_48218);
xnor UO_29 (O_29,N_49265,N_48202);
and UO_30 (O_30,N_48615,N_48368);
nor UO_31 (O_31,N_49601,N_48388);
and UO_32 (O_32,N_48566,N_49154);
nor UO_33 (O_33,N_48467,N_49890);
xor UO_34 (O_34,N_49549,N_48352);
xor UO_35 (O_35,N_48785,N_48015);
nand UO_36 (O_36,N_48908,N_48794);
nand UO_37 (O_37,N_49043,N_49784);
nor UO_38 (O_38,N_48465,N_48239);
xnor UO_39 (O_39,N_49834,N_49193);
and UO_40 (O_40,N_49464,N_49634);
nand UO_41 (O_41,N_49564,N_49025);
xor UO_42 (O_42,N_48204,N_49860);
xnor UO_43 (O_43,N_48157,N_48125);
and UO_44 (O_44,N_49290,N_48214);
xor UO_45 (O_45,N_49139,N_49839);
nand UO_46 (O_46,N_48198,N_49855);
nor UO_47 (O_47,N_49746,N_49900);
and UO_48 (O_48,N_49218,N_49427);
and UO_49 (O_49,N_49442,N_48542);
or UO_50 (O_50,N_48285,N_49737);
or UO_51 (O_51,N_49050,N_49165);
nor UO_52 (O_52,N_48851,N_48443);
or UO_53 (O_53,N_48071,N_49921);
or UO_54 (O_54,N_49096,N_48739);
nor UO_55 (O_55,N_48775,N_49271);
nor UO_56 (O_56,N_48509,N_49135);
and UO_57 (O_57,N_49308,N_49024);
or UO_58 (O_58,N_48183,N_49272);
or UO_59 (O_59,N_48654,N_48563);
nand UO_60 (O_60,N_49934,N_49786);
nand UO_61 (O_61,N_49131,N_49748);
nor UO_62 (O_62,N_48657,N_48505);
nand UO_63 (O_63,N_49882,N_49527);
and UO_64 (O_64,N_49468,N_48992);
nor UO_65 (O_65,N_48689,N_49976);
or UO_66 (O_66,N_48028,N_49978);
nor UO_67 (O_67,N_48860,N_48397);
or UO_68 (O_68,N_48551,N_48034);
or UO_69 (O_69,N_48105,N_49597);
nand UO_70 (O_70,N_49371,N_48738);
and UO_71 (O_71,N_48338,N_48651);
and UO_72 (O_72,N_48940,N_48411);
xnor UO_73 (O_73,N_49719,N_49917);
nor UO_74 (O_74,N_49312,N_48730);
or UO_75 (O_75,N_49941,N_49665);
and UO_76 (O_76,N_49156,N_48255);
nor UO_77 (O_77,N_48629,N_49823);
and UO_78 (O_78,N_48697,N_49962);
nand UO_79 (O_79,N_49432,N_48166);
nand UO_80 (O_80,N_49568,N_48773);
xor UO_81 (O_81,N_48458,N_49875);
nand UO_82 (O_82,N_49261,N_48164);
nand UO_83 (O_83,N_48791,N_49158);
and UO_84 (O_84,N_49037,N_49221);
nand UO_85 (O_85,N_48799,N_49883);
or UO_86 (O_86,N_49658,N_49583);
nor UO_87 (O_87,N_49887,N_48062);
or UO_88 (O_88,N_49967,N_48171);
nand UO_89 (O_89,N_48847,N_49945);
xor UO_90 (O_90,N_48007,N_49414);
nor UO_91 (O_91,N_48891,N_49393);
nand UO_92 (O_92,N_49950,N_49578);
xor UO_93 (O_93,N_49287,N_49582);
nand UO_94 (O_94,N_49970,N_48391);
or UO_95 (O_95,N_48237,N_48752);
xnor UO_96 (O_96,N_49576,N_49998);
and UO_97 (O_97,N_48017,N_48506);
or UO_98 (O_98,N_49063,N_48769);
or UO_99 (O_99,N_49447,N_48390);
nor UO_100 (O_100,N_48173,N_49920);
nor UO_101 (O_101,N_48309,N_49231);
nand UO_102 (O_102,N_49350,N_48887);
nor UO_103 (O_103,N_49132,N_49808);
nand UO_104 (O_104,N_48628,N_49421);
xor UO_105 (O_105,N_48511,N_48302);
nor UO_106 (O_106,N_48611,N_49189);
nand UO_107 (O_107,N_49383,N_49529);
and UO_108 (O_108,N_49083,N_48503);
xor UO_109 (O_109,N_48996,N_49675);
xor UO_110 (O_110,N_48608,N_48777);
nor UO_111 (O_111,N_48333,N_48369);
nand UO_112 (O_112,N_49289,N_49669);
or UO_113 (O_113,N_49773,N_48723);
nor UO_114 (O_114,N_49078,N_49636);
nand UO_115 (O_115,N_48937,N_49944);
nor UO_116 (O_116,N_49622,N_48481);
xnor UO_117 (O_117,N_48939,N_48363);
xor UO_118 (O_118,N_49355,N_48052);
nand UO_119 (O_119,N_48492,N_48528);
nor UO_120 (O_120,N_49942,N_49047);
and UO_121 (O_121,N_48732,N_49007);
and UO_122 (O_122,N_49870,N_49930);
or UO_123 (O_123,N_49792,N_48848);
or UO_124 (O_124,N_48792,N_49559);
nor UO_125 (O_125,N_49143,N_48488);
nand UO_126 (O_126,N_48328,N_49562);
or UO_127 (O_127,N_49466,N_48721);
xnor UO_128 (O_128,N_48261,N_48120);
nor UO_129 (O_129,N_49424,N_48002);
nor UO_130 (O_130,N_48864,N_49984);
and UO_131 (O_131,N_48347,N_49357);
xnor UO_132 (O_132,N_49817,N_48962);
xnor UO_133 (O_133,N_49170,N_48916);
nor UO_134 (O_134,N_48189,N_49150);
xor UO_135 (O_135,N_49535,N_48206);
xnor UO_136 (O_136,N_48946,N_48057);
or UO_137 (O_137,N_48463,N_49129);
and UO_138 (O_138,N_48473,N_49459);
nand UO_139 (O_139,N_49159,N_48857);
nor UO_140 (O_140,N_48854,N_48485);
or UO_141 (O_141,N_49988,N_48696);
nor UO_142 (O_142,N_48784,N_48605);
or UO_143 (O_143,N_48232,N_49865);
and UO_144 (O_144,N_48288,N_49401);
xor UO_145 (O_145,N_49045,N_48330);
and UO_146 (O_146,N_48987,N_48925);
xor UO_147 (O_147,N_49715,N_48523);
nand UO_148 (O_148,N_48903,N_49240);
and UO_149 (O_149,N_49761,N_49062);
or UO_150 (O_150,N_48574,N_49926);
or UO_151 (O_151,N_48744,N_48260);
xor UO_152 (O_152,N_49588,N_49082);
xnor UO_153 (O_153,N_48695,N_49811);
and UO_154 (O_154,N_48095,N_48922);
or UO_155 (O_155,N_49276,N_48627);
nand UO_156 (O_156,N_48444,N_49364);
xor UO_157 (O_157,N_48043,N_48290);
or UO_158 (O_158,N_49434,N_49462);
xor UO_159 (O_159,N_49619,N_48068);
and UO_160 (O_160,N_48085,N_49035);
xor UO_161 (O_161,N_49463,N_49630);
or UO_162 (O_162,N_49450,N_49845);
nor UO_163 (O_163,N_49281,N_49028);
nor UO_164 (O_164,N_49819,N_49736);
xor UO_165 (O_165,N_49708,N_48911);
nor UO_166 (O_166,N_49638,N_48673);
nor UO_167 (O_167,N_49124,N_49895);
nand UO_168 (O_168,N_49136,N_48241);
and UO_169 (O_169,N_49661,N_48907);
xor UO_170 (O_170,N_48975,N_49435);
and UO_171 (O_171,N_48222,N_49904);
nand UO_172 (O_172,N_48094,N_49893);
nor UO_173 (O_173,N_49964,N_48945);
nand UO_174 (O_174,N_49932,N_48275);
xor UO_175 (O_175,N_49596,N_48949);
or UO_176 (O_176,N_48393,N_48895);
xor UO_177 (O_177,N_48195,N_49418);
xor UO_178 (O_178,N_48631,N_48455);
xnor UO_179 (O_179,N_48549,N_48459);
xnor UO_180 (O_180,N_48672,N_48519);
or UO_181 (O_181,N_49347,N_49186);
nor UO_182 (O_182,N_49117,N_49426);
nor UO_183 (O_183,N_49734,N_48958);
and UO_184 (O_184,N_49627,N_49064);
nand UO_185 (O_185,N_49612,N_48176);
and UO_186 (O_186,N_48576,N_48306);
or UO_187 (O_187,N_48893,N_49258);
nand UO_188 (O_188,N_48131,N_48543);
or UO_189 (O_189,N_49948,N_49381);
xor UO_190 (O_190,N_49239,N_49451);
nor UO_191 (O_191,N_49455,N_49031);
xnor UO_192 (O_192,N_49115,N_49825);
xor UO_193 (O_193,N_48335,N_48491);
and UO_194 (O_194,N_49810,N_48558);
nand UO_195 (O_195,N_49252,N_49949);
or UO_196 (O_196,N_48165,N_48639);
and UO_197 (O_197,N_48296,N_48741);
or UO_198 (O_198,N_48929,N_48985);
and UO_199 (O_199,N_49779,N_49125);
or UO_200 (O_200,N_48538,N_48064);
nor UO_201 (O_201,N_48595,N_49927);
or UO_202 (O_202,N_48342,N_49595);
or UO_203 (O_203,N_48282,N_48984);
nand UO_204 (O_204,N_48587,N_49718);
and UO_205 (O_205,N_48039,N_49303);
and UO_206 (O_206,N_48927,N_49742);
and UO_207 (O_207,N_48196,N_48554);
xor UO_208 (O_208,N_48529,N_48321);
nor UO_209 (O_209,N_48399,N_48827);
xnor UO_210 (O_210,N_48797,N_49781);
nor UO_211 (O_211,N_48240,N_49645);
or UO_212 (O_212,N_48426,N_49524);
and UO_213 (O_213,N_48955,N_48731);
xor UO_214 (O_214,N_48546,N_48771);
xnor UO_215 (O_215,N_49586,N_48515);
and UO_216 (O_216,N_48942,N_49306);
or UO_217 (O_217,N_48802,N_49332);
nand UO_218 (O_218,N_49759,N_48194);
nand UO_219 (O_219,N_48358,N_48601);
nand UO_220 (O_220,N_49858,N_49351);
nand UO_221 (O_221,N_48216,N_49333);
xnor UO_222 (O_222,N_48295,N_49548);
nand UO_223 (O_223,N_48570,N_49345);
or UO_224 (O_224,N_48318,N_48320);
nor UO_225 (O_225,N_49104,N_48990);
xnor UO_226 (O_226,N_48266,N_49841);
xnor UO_227 (O_227,N_48316,N_48759);
xor UO_228 (O_228,N_49471,N_48155);
nand UO_229 (O_229,N_48966,N_48346);
nand UO_230 (O_230,N_48425,N_48339);
nand UO_231 (O_231,N_49387,N_49722);
and UO_232 (O_232,N_48960,N_48223);
nand UO_233 (O_233,N_49668,N_48906);
and UO_234 (O_234,N_48040,N_48361);
nor UO_235 (O_235,N_49696,N_49423);
and UO_236 (O_236,N_49906,N_48385);
xor UO_237 (O_237,N_49752,N_49461);
nor UO_238 (O_238,N_49727,N_49829);
and UO_239 (O_239,N_48508,N_49913);
or UO_240 (O_240,N_49151,N_49251);
and UO_241 (O_241,N_48109,N_48021);
and UO_242 (O_242,N_48379,N_48038);
and UO_243 (O_243,N_49687,N_49085);
or UO_244 (O_244,N_48844,N_49235);
or UO_245 (O_245,N_49282,N_49600);
nand UO_246 (O_246,N_49517,N_48878);
and UO_247 (O_247,N_48307,N_49176);
or UO_248 (O_248,N_48980,N_48209);
or UO_249 (O_249,N_48278,N_48325);
nor UO_250 (O_250,N_49571,N_48436);
nand UO_251 (O_251,N_48045,N_49408);
or UO_252 (O_252,N_48632,N_48550);
nand UO_253 (O_253,N_48691,N_48620);
and UO_254 (O_254,N_48983,N_49859);
xnor UO_255 (O_255,N_48471,N_49216);
nor UO_256 (O_256,N_48514,N_48944);
nand UO_257 (O_257,N_49396,N_49311);
and UO_258 (O_258,N_48373,N_49196);
and UO_259 (O_259,N_48248,N_48274);
or UO_260 (O_260,N_48022,N_49873);
nor UO_261 (O_261,N_48097,N_48643);
nor UO_262 (O_262,N_49902,N_49955);
nor UO_263 (O_263,N_49211,N_49788);
or UO_264 (O_264,N_48494,N_48781);
and UO_265 (O_265,N_48683,N_49974);
xnor UO_266 (O_266,N_48667,N_48392);
or UO_267 (O_267,N_48046,N_48915);
xnor UO_268 (O_268,N_49054,N_49966);
nand UO_269 (O_269,N_49237,N_49879);
nor UO_270 (O_270,N_48858,N_48416);
xnor UO_271 (O_271,N_48981,N_48954);
nand UO_272 (O_272,N_49206,N_49046);
or UO_273 (O_273,N_49561,N_49611);
nor UO_274 (O_274,N_48035,N_48450);
nor UO_275 (O_275,N_49554,N_48460);
nor UO_276 (O_276,N_49288,N_48341);
xor UO_277 (O_277,N_48367,N_49774);
nand UO_278 (O_278,N_48751,N_48215);
nand UO_279 (O_279,N_49399,N_48606);
nor UO_280 (O_280,N_48005,N_48025);
and UO_281 (O_281,N_48894,N_48270);
nand UO_282 (O_282,N_48305,N_49120);
nand UO_283 (O_283,N_49910,N_49983);
or UO_284 (O_284,N_48483,N_49505);
nand UO_285 (O_285,N_48755,N_49646);
and UO_286 (O_286,N_49793,N_48671);
xor UO_287 (O_287,N_49946,N_49484);
and UO_288 (O_288,N_48780,N_49807);
nand UO_289 (O_289,N_49818,N_48749);
or UO_290 (O_290,N_48042,N_49520);
xor UO_291 (O_291,N_49180,N_49173);
xnor UO_292 (O_292,N_49849,N_49833);
nor UO_293 (O_293,N_49924,N_49572);
or UO_294 (O_294,N_49210,N_48600);
or UO_295 (O_295,N_49509,N_48863);
and UO_296 (O_296,N_48315,N_49051);
nor UO_297 (O_297,N_49565,N_48641);
nand UO_298 (O_298,N_48029,N_49220);
nor UO_299 (O_299,N_48149,N_48244);
and UO_300 (O_300,N_48226,N_49706);
nand UO_301 (O_301,N_48360,N_49254);
nand UO_302 (O_302,N_48677,N_49667);
and UO_303 (O_303,N_48835,N_48621);
and UO_304 (O_304,N_49222,N_48592);
and UO_305 (O_305,N_48885,N_48867);
and UO_306 (O_306,N_48312,N_48324);
nand UO_307 (O_307,N_48357,N_48184);
nand UO_308 (O_308,N_49362,N_49488);
nand UO_309 (O_309,N_49889,N_48348);
or UO_310 (O_310,N_48049,N_49188);
or UO_311 (O_311,N_48225,N_48087);
or UO_312 (O_312,N_49659,N_49684);
nor UO_313 (O_313,N_48400,N_48336);
xor UO_314 (O_314,N_49985,N_49338);
or UO_315 (O_315,N_48583,N_48405);
or UO_316 (O_316,N_49485,N_48177);
or UO_317 (O_317,N_49698,N_49286);
nor UO_318 (O_318,N_48801,N_49011);
or UO_319 (O_319,N_48881,N_49021);
or UO_320 (O_320,N_49642,N_49171);
nor UO_321 (O_321,N_48747,N_49678);
nor UO_322 (O_322,N_49794,N_49448);
nand UO_323 (O_323,N_49663,N_49074);
xnor UO_324 (O_324,N_48170,N_48415);
xnor UO_325 (O_325,N_49155,N_49420);
or UO_326 (O_326,N_48365,N_49537);
nand UO_327 (O_327,N_48430,N_49604);
nand UO_328 (O_328,N_49105,N_49996);
nand UO_329 (O_329,N_48280,N_48387);
or UO_330 (O_330,N_49689,N_49835);
nor UO_331 (O_331,N_48846,N_49768);
and UO_332 (O_332,N_48521,N_48462);
nor UO_333 (O_333,N_49717,N_48834);
xor UO_334 (O_334,N_49304,N_49329);
or UO_335 (O_335,N_49550,N_49959);
xnor UO_336 (O_336,N_49547,N_48526);
nand UO_337 (O_337,N_49010,N_49310);
nor UO_338 (O_338,N_48988,N_48746);
and UO_339 (O_339,N_49880,N_49624);
nand UO_340 (O_340,N_48308,N_49175);
xor UO_341 (O_341,N_49480,N_48269);
nand UO_342 (O_342,N_49953,N_49672);
or UO_343 (O_343,N_49813,N_49452);
and UO_344 (O_344,N_48246,N_48207);
nor UO_345 (O_345,N_49397,N_49430);
xor UO_346 (O_346,N_48349,N_49149);
or UO_347 (O_347,N_49683,N_49342);
or UO_348 (O_348,N_49269,N_48013);
nor UO_349 (O_349,N_49735,N_49277);
nand UO_350 (O_350,N_48322,N_48676);
or UO_351 (O_351,N_48766,N_48283);
or UO_352 (O_352,N_49629,N_48711);
and UO_353 (O_353,N_49909,N_49854);
nor UO_354 (O_354,N_48838,N_49223);
xor UO_355 (O_355,N_49496,N_48123);
xor UO_356 (O_356,N_48371,N_48160);
nor UO_357 (O_357,N_48826,N_49570);
nand UO_358 (O_358,N_49321,N_48890);
nor UO_359 (O_359,N_49185,N_48080);
and UO_360 (O_360,N_49556,N_49256);
or UO_361 (O_361,N_49284,N_48245);
nor UO_362 (O_362,N_49236,N_48547);
nor UO_363 (O_363,N_49526,N_48921);
nor UO_364 (O_364,N_48806,N_48898);
and UO_365 (O_365,N_49244,N_48804);
or UO_366 (O_366,N_49725,N_49302);
nand UO_367 (O_367,N_48359,N_48382);
xor UO_368 (O_368,N_48116,N_49815);
and UO_369 (O_369,N_49502,N_48303);
or UO_370 (O_370,N_48935,N_49738);
xor UO_371 (O_371,N_48003,N_48100);
or UO_372 (O_372,N_49703,N_49830);
nand UO_373 (O_373,N_49026,N_48710);
nor UO_374 (O_374,N_49804,N_48102);
and UO_375 (O_375,N_49673,N_49821);
or UO_376 (O_376,N_48733,N_48597);
xnor UO_377 (O_377,N_49390,N_48454);
nor UO_378 (O_378,N_49617,N_48496);
and UO_379 (O_379,N_49255,N_48182);
and UO_380 (O_380,N_48172,N_49602);
xnor UO_381 (O_381,N_49713,N_48054);
or UO_382 (O_382,N_49757,N_48299);
and UO_383 (O_383,N_48590,N_49747);
nand UO_384 (O_384,N_49692,N_48151);
nor UO_385 (O_385,N_49030,N_49073);
and UO_386 (O_386,N_49367,N_48439);
xnor UO_387 (O_387,N_48421,N_48613);
and UO_388 (O_388,N_48977,N_48536);
nand UO_389 (O_389,N_48012,N_49394);
xor UO_390 (O_390,N_49293,N_48210);
nor UO_391 (O_391,N_49192,N_48787);
or UO_392 (O_392,N_48072,N_49898);
nor UO_393 (O_393,N_49616,N_48602);
nor UO_394 (O_394,N_48742,N_48690);
xnor UO_395 (O_395,N_48951,N_49492);
or UO_396 (O_396,N_48900,N_49365);
nor UO_397 (O_397,N_48708,N_48726);
xor UO_398 (O_398,N_48297,N_48060);
nor UO_399 (O_399,N_49470,N_49762);
nand UO_400 (O_400,N_48517,N_48663);
nor UO_401 (O_401,N_48188,N_49837);
xnor UO_402 (O_402,N_49376,N_49999);
or UO_403 (O_403,N_48475,N_49164);
or UO_404 (O_404,N_49666,N_49772);
xor UO_405 (O_405,N_49567,N_49476);
nand UO_406 (O_406,N_49677,N_49544);
nand UO_407 (O_407,N_49008,N_48457);
or UO_408 (O_408,N_49828,N_49438);
and UO_409 (O_409,N_49891,N_49589);
nor UO_410 (O_410,N_49389,N_49419);
nor UO_411 (O_411,N_49065,N_49528);
and UO_412 (O_412,N_49968,N_49077);
nand UO_413 (O_413,N_48018,N_48585);
or UO_414 (O_414,N_48815,N_48687);
nor UO_415 (O_415,N_48810,N_48323);
or UO_416 (O_416,N_48148,N_49513);
xor UO_417 (O_417,N_48070,N_48383);
xnor UO_418 (O_418,N_49648,N_48930);
and UO_419 (O_419,N_48719,N_49908);
and UO_420 (O_420,N_49353,N_49097);
and UO_421 (O_421,N_49157,N_48409);
xor UO_422 (O_422,N_48263,N_48103);
or UO_423 (O_423,N_48093,N_49400);
nand UO_424 (O_424,N_48136,N_48249);
nor UO_425 (O_425,N_48967,N_49770);
and UO_426 (O_426,N_49138,N_48386);
xnor UO_427 (O_427,N_48679,N_48553);
nor UO_428 (O_428,N_48211,N_49128);
nor UO_429 (O_429,N_49032,N_48839);
nand UO_430 (O_430,N_48442,N_49499);
xor UO_431 (O_431,N_48137,N_48186);
nand UO_432 (O_432,N_49783,N_48669);
or UO_433 (O_433,N_49207,N_49575);
nor UO_434 (O_434,N_49728,N_49091);
or UO_435 (O_435,N_48886,N_49121);
nor UO_436 (O_436,N_49832,N_48750);
nand UO_437 (O_437,N_49481,N_48513);
and UO_438 (O_438,N_48077,N_49872);
or UO_439 (O_439,N_48200,N_49375);
nor UO_440 (O_440,N_48276,N_49181);
xnor UO_441 (O_441,N_49014,N_49566);
nand UO_442 (O_442,N_48598,N_49607);
nor UO_443 (O_443,N_48818,N_49705);
nand UO_444 (O_444,N_48037,N_48272);
nor UO_445 (O_445,N_48031,N_48776);
nor UO_446 (O_446,N_49495,N_49314);
nor UO_447 (O_447,N_49145,N_49194);
and UO_448 (O_448,N_49863,N_49894);
xnor UO_449 (O_449,N_49056,N_48408);
or UO_450 (O_450,N_48310,N_49726);
nand UO_451 (O_451,N_48009,N_48702);
and UO_452 (O_452,N_48178,N_48763);
nor UO_453 (O_453,N_49088,N_48704);
or UO_454 (O_454,N_48380,N_48445);
and UO_455 (O_455,N_49587,N_49454);
nor UO_456 (O_456,N_49662,N_48714);
xor UO_457 (O_457,N_48337,N_49113);
or UO_458 (O_458,N_49144,N_49267);
or UO_459 (O_459,N_48317,N_48926);
and UO_460 (O_460,N_48081,N_49899);
or UO_461 (O_461,N_49443,N_49552);
nor UO_462 (O_462,N_49739,N_49540);
nor UO_463 (O_463,N_49695,N_49615);
nor UO_464 (O_464,N_48101,N_48718);
xor UO_465 (O_465,N_48979,N_49268);
or UO_466 (O_466,N_48913,N_48762);
nand UO_467 (O_467,N_49776,N_49214);
or UO_468 (O_468,N_48142,N_48319);
nor UO_469 (O_469,N_48713,N_49190);
or UO_470 (O_470,N_48469,N_49212);
nand UO_471 (O_471,N_49292,N_49560);
xnor UO_472 (O_472,N_48153,N_49018);
nand UO_473 (O_473,N_48294,N_49584);
and UO_474 (O_474,N_49053,N_49068);
nor UO_475 (O_475,N_49163,N_49652);
nand UO_476 (O_476,N_48130,N_48372);
and UO_477 (O_477,N_48976,N_48119);
xor UO_478 (O_478,N_48487,N_49323);
and UO_479 (O_479,N_49366,N_49907);
nor UO_480 (O_480,N_48823,N_49755);
and UO_481 (O_481,N_48213,N_49205);
xor UO_482 (O_482,N_49245,N_49799);
and UO_483 (O_483,N_49938,N_48434);
xor UO_484 (O_484,N_48234,N_48758);
nor UO_485 (O_485,N_49280,N_49812);
nor UO_486 (O_486,N_48051,N_49809);
xor UO_487 (O_487,N_49335,N_49981);
xnor UO_488 (O_488,N_48343,N_48507);
nor UO_489 (O_489,N_48141,N_49349);
nand UO_490 (O_490,N_48924,N_48617);
or UO_491 (O_491,N_48522,N_48227);
and UO_492 (O_492,N_49574,N_48573);
xnor UO_493 (O_493,N_49700,N_49644);
or UO_494 (O_494,N_49516,N_48624);
and UO_495 (O_495,N_49745,N_48354);
and UO_496 (O_496,N_49232,N_48956);
and UO_497 (O_497,N_48837,N_49242);
nor UO_498 (O_498,N_49440,N_48941);
nand UO_499 (O_499,N_48861,N_49503);
and UO_500 (O_500,N_48143,N_49877);
xnor UO_501 (O_501,N_48789,N_49741);
nand UO_502 (O_502,N_48999,N_48874);
xor UO_503 (O_503,N_49228,N_49724);
nand UO_504 (O_504,N_48564,N_49177);
and UO_505 (O_505,N_49791,N_48768);
nor UO_506 (O_506,N_48192,N_48451);
xor UO_507 (O_507,N_49071,N_48855);
or UO_508 (O_508,N_49406,N_49318);
or UO_509 (O_509,N_49022,N_49110);
nand UO_510 (O_510,N_48675,N_48965);
nand UO_511 (O_511,N_49876,N_49626);
xor UO_512 (O_512,N_49935,N_49579);
xor UO_513 (O_513,N_49374,N_48622);
or UO_514 (O_514,N_49915,N_49997);
xnor UO_515 (O_515,N_49257,N_49871);
or UO_516 (O_516,N_48674,N_49836);
nand UO_517 (O_517,N_48642,N_48539);
and UO_518 (O_518,N_49937,N_48461);
nand UO_519 (O_519,N_48175,N_48048);
nor UO_520 (O_520,N_48699,N_49866);
xnor UO_521 (O_521,N_48495,N_49475);
or UO_522 (O_522,N_49215,N_49409);
and UO_523 (O_523,N_48938,N_49160);
nor UO_524 (O_524,N_48840,N_48205);
and UO_525 (O_525,N_48905,N_48909);
xor UO_526 (O_526,N_49933,N_49320);
nand UO_527 (O_527,N_48127,N_48767);
nor UO_528 (O_528,N_49598,N_48943);
nor UO_529 (O_529,N_48122,N_48124);
nor UO_530 (O_530,N_48073,N_49274);
nand UO_531 (O_531,N_49886,N_48174);
and UO_532 (O_532,N_49633,N_48995);
nor UO_533 (O_533,N_48449,N_48493);
or UO_534 (O_534,N_48636,N_48375);
nor UO_535 (O_535,N_48334,N_48344);
or UO_536 (O_536,N_49386,N_48413);
or UO_537 (O_537,N_49108,N_49279);
nand UO_538 (O_538,N_48836,N_49664);
or UO_539 (O_539,N_48648,N_48572);
and UO_540 (O_540,N_48161,N_48252);
nand UO_541 (O_541,N_49850,N_49392);
nand UO_542 (O_542,N_48761,N_48104);
nand UO_543 (O_543,N_49802,N_48197);
xnor UO_544 (O_544,N_48665,N_48825);
nand UO_545 (O_545,N_48370,N_49868);
nor UO_546 (O_546,N_48433,N_49001);
xnor UO_547 (O_547,N_48050,N_49848);
or UO_548 (O_548,N_49923,N_48754);
nand UO_549 (O_549,N_48401,N_48682);
and UO_550 (O_550,N_48414,N_48428);
and UO_551 (O_551,N_49324,N_48661);
nand UO_552 (O_552,N_49801,N_48707);
nand UO_553 (O_553,N_49436,N_49297);
xor UO_554 (O_554,N_48795,N_49134);
or UO_555 (O_555,N_48612,N_48313);
xnor UO_556 (O_556,N_48633,N_49263);
nor UO_557 (O_557,N_48014,N_49278);
xor UO_558 (O_558,N_48026,N_48424);
and UO_559 (O_559,N_48086,N_49961);
xnor UO_560 (O_560,N_48670,N_48545);
xor UO_561 (O_561,N_48134,N_48917);
xnor UO_562 (O_562,N_49551,N_48053);
xor UO_563 (O_563,N_49388,N_48472);
xor UO_564 (O_564,N_48630,N_49041);
nor UO_565 (O_565,N_49178,N_48404);
nand UO_566 (O_566,N_48524,N_48238);
and UO_567 (O_567,N_48986,N_49368);
nor UO_568 (O_568,N_48356,N_49040);
nand UO_569 (O_569,N_49620,N_48685);
nand UO_570 (O_570,N_48963,N_48535);
and UO_571 (O_571,N_49384,N_49796);
or UO_572 (O_572,N_49472,N_49771);
xor UO_573 (O_573,N_49238,N_49446);
or UO_574 (O_574,N_48557,N_49711);
and UO_575 (O_575,N_48765,N_49227);
nand UO_576 (O_576,N_48770,N_49842);
nand UO_577 (O_577,N_48437,N_49831);
nor UO_578 (O_578,N_48201,N_49971);
xor UO_579 (O_579,N_49982,N_48548);
xor UO_580 (O_580,N_49378,N_49067);
nor UO_581 (O_581,N_49243,N_48464);
nor UO_582 (O_582,N_49042,N_49017);
xnor UO_583 (O_583,N_49167,N_49000);
xnor UO_584 (O_584,N_49531,N_48817);
and UO_585 (O_585,N_49296,N_49219);
nor UO_586 (O_586,N_49153,N_49044);
nor UO_587 (O_587,N_49460,N_49072);
or UO_588 (O_588,N_49405,N_48936);
xor UO_589 (O_589,N_48212,N_49187);
nor UO_590 (O_590,N_49847,N_49766);
nand UO_591 (O_591,N_48099,N_48006);
and UO_592 (O_592,N_49055,N_49987);
nand UO_593 (O_593,N_49822,N_48518);
or UO_594 (O_594,N_48499,N_49119);
xor UO_595 (O_595,N_49100,N_48964);
xor UO_596 (O_596,N_49036,N_48579);
and UO_597 (O_597,N_48525,N_49059);
nand UO_598 (O_598,N_49744,N_49580);
nor UO_599 (O_599,N_48811,N_49004);
xnor UO_600 (O_600,N_49951,N_48520);
nand UO_601 (O_601,N_49905,N_49515);
nand UO_602 (O_602,N_48108,N_49750);
and UO_603 (O_603,N_48432,N_48666);
nand UO_604 (O_604,N_48888,N_48658);
nand UO_605 (O_605,N_48069,N_49250);
or UO_606 (O_606,N_49198,N_48753);
nand UO_607 (O_607,N_48869,N_49765);
nor UO_608 (O_608,N_49852,N_48406);
nand UO_609 (O_609,N_48490,N_48271);
nor UO_610 (O_610,N_48978,N_48533);
nor UO_611 (O_611,N_49701,N_48786);
xor UO_612 (O_612,N_49992,N_48866);
nand UO_613 (O_613,N_48778,N_49534);
or UO_614 (O_614,N_48476,N_49972);
or UO_615 (O_615,N_49079,N_48168);
nor UO_616 (O_616,N_48128,N_49307);
xor UO_617 (O_617,N_49577,N_49897);
nand UO_618 (O_618,N_49995,N_48076);
xor UO_619 (O_619,N_49415,N_48596);
nand UO_620 (O_620,N_49217,N_48298);
or UO_621 (O_621,N_49618,N_48059);
nand UO_622 (O_622,N_48118,N_49201);
nand UO_623 (O_623,N_49416,N_49640);
nor UO_624 (O_624,N_49780,N_49166);
and UO_625 (O_625,N_49111,N_49385);
nor UO_626 (O_626,N_48082,N_49359);
and UO_627 (O_627,N_49498,N_48645);
nand UO_628 (O_628,N_49380,N_49614);
nand UO_629 (O_629,N_49991,N_49922);
xnor UO_630 (O_630,N_49395,N_48822);
nand UO_631 (O_631,N_48635,N_49676);
xor UO_632 (O_632,N_48110,N_49699);
and UO_633 (O_633,N_48580,N_49094);
or UO_634 (O_634,N_48466,N_49901);
nand UO_635 (O_635,N_48114,N_48180);
and UO_636 (O_636,N_49494,N_48829);
nor UO_637 (O_637,N_48581,N_48250);
nor UO_638 (O_638,N_49225,N_49525);
nor UO_639 (O_639,N_48698,N_48396);
nand UO_640 (O_640,N_48774,N_49184);
and UO_641 (O_641,N_49019,N_48932);
and UO_642 (O_642,N_49546,N_49095);
xnor UO_643 (O_643,N_48156,N_48562);
nor UO_644 (O_644,N_49679,N_48289);
or UO_645 (O_645,N_49519,N_48410);
and UO_646 (O_646,N_49012,N_49148);
xnor UO_647 (O_647,N_49656,N_48254);
and UO_648 (O_648,N_49947,N_49283);
nor UO_649 (O_649,N_49253,N_49867);
xnor UO_650 (O_650,N_49806,N_48242);
nor UO_651 (O_651,N_48190,N_49896);
nor UO_652 (O_652,N_48500,N_49313);
xnor UO_653 (O_653,N_48889,N_48144);
and UO_654 (O_654,N_49720,N_49654);
nand UO_655 (O_655,N_49606,N_48901);
or UO_656 (O_656,N_49591,N_48637);
nor UO_657 (O_657,N_49478,N_49497);
xor UO_658 (O_658,N_48609,N_48162);
nor UO_659 (O_659,N_48033,N_49102);
nand UO_660 (O_660,N_49316,N_48537);
nor UO_661 (O_661,N_49179,N_49369);
xor UO_662 (O_662,N_48154,N_49758);
or UO_663 (O_663,N_48262,N_48734);
nand UO_664 (O_664,N_49444,N_48193);
or UO_665 (O_665,N_49878,N_48567);
and UO_666 (O_666,N_49846,N_49340);
nand UO_667 (O_667,N_48502,N_48381);
and UO_668 (O_668,N_48004,N_48020);
and UO_669 (O_669,N_49334,N_49116);
xnor UO_670 (O_670,N_49709,N_48619);
and UO_671 (O_671,N_48709,N_49543);
nor UO_672 (O_672,N_48748,N_48041);
nand UO_673 (O_673,N_48301,N_49348);
xor UO_674 (O_674,N_49599,N_49101);
nand UO_675 (O_675,N_48756,N_49563);
xor UO_676 (O_676,N_49764,N_49686);
and UO_677 (O_677,N_48420,N_48291);
nor UO_678 (O_678,N_48607,N_49441);
or UO_679 (O_679,N_49112,N_49203);
nand UO_680 (O_680,N_49174,N_49536);
nor UO_681 (O_681,N_48376,N_49690);
nor UO_682 (O_682,N_48532,N_49109);
or UO_683 (O_683,N_48982,N_48132);
or UO_684 (O_684,N_48001,N_48813);
nand UO_685 (O_685,N_49413,N_48159);
or UO_686 (O_686,N_48187,N_49358);
nand UO_687 (O_687,N_48831,N_48247);
xnor UO_688 (O_688,N_49594,N_48821);
nand UO_689 (O_689,N_48989,N_49069);
nand UO_690 (O_690,N_49259,N_49892);
xor UO_691 (O_691,N_49851,N_48931);
and UO_692 (O_692,N_48933,N_49510);
xnor UO_693 (O_693,N_48024,N_49731);
xor UO_694 (O_694,N_49621,N_49247);
and UO_695 (O_695,N_48150,N_49213);
nor UO_696 (O_696,N_48828,N_48089);
nand UO_697 (O_697,N_48075,N_48640);
nor UO_698 (O_698,N_49660,N_48722);
nand UO_699 (O_699,N_48113,N_49337);
xnor UO_700 (O_700,N_48803,N_48056);
xor UO_701 (O_701,N_49501,N_49431);
nor UO_702 (O_702,N_48429,N_48591);
nor UO_703 (O_703,N_49309,N_48208);
nor UO_704 (O_704,N_49800,N_49339);
xnor UO_705 (O_705,N_49939,N_49716);
and UO_706 (O_706,N_48253,N_48997);
xnor UO_707 (O_707,N_49161,N_49168);
or UO_708 (O_708,N_48384,N_48231);
and UO_709 (O_709,N_48427,N_48586);
nand UO_710 (O_710,N_49382,N_48655);
or UO_711 (O_711,N_48993,N_48816);
nand UO_712 (O_712,N_49425,N_49075);
or UO_713 (O_713,N_48355,N_49327);
and UO_714 (O_714,N_49785,N_49523);
nor UO_715 (O_715,N_49844,N_49052);
and UO_716 (O_716,N_49760,N_48737);
or UO_717 (O_717,N_48264,N_48880);
nor UO_718 (O_718,N_49691,N_49625);
or UO_719 (O_719,N_49805,N_49467);
xor UO_720 (O_720,N_48191,N_48126);
or UO_721 (O_721,N_49816,N_48329);
nand UO_722 (O_722,N_48555,N_49391);
and UO_723 (O_723,N_48569,N_48892);
xor UO_724 (O_724,N_48366,N_49114);
and UO_725 (O_725,N_49453,N_49843);
nor UO_726 (O_726,N_49057,N_49410);
and UO_727 (O_727,N_49507,N_49697);
nand UO_728 (O_728,N_49015,N_49730);
nor UO_729 (O_729,N_48736,N_48257);
or UO_730 (O_730,N_48700,N_49919);
xor UO_731 (O_731,N_48575,N_48959);
nor UO_732 (O_732,N_48423,N_49790);
nor UO_733 (O_733,N_49911,N_48853);
and UO_734 (O_734,N_49020,N_48265);
nand UO_735 (O_735,N_49820,N_48664);
or UO_736 (O_736,N_49049,N_49608);
nand UO_737 (O_737,N_48096,N_48531);
nor UO_738 (O_738,N_49609,N_49925);
nor UO_739 (O_739,N_49743,N_48660);
nor UO_740 (O_740,N_49916,N_48969);
and UO_741 (O_741,N_48649,N_48353);
and UO_742 (O_742,N_49118,N_48090);
or UO_743 (O_743,N_48044,N_48833);
nor UO_744 (O_744,N_48819,N_48008);
or UO_745 (O_745,N_48725,N_48934);
xor UO_746 (O_746,N_49191,N_48876);
xor UO_747 (O_747,N_48544,N_48447);
and UO_748 (O_748,N_48088,N_49767);
xnor UO_749 (O_749,N_49162,N_49979);
xnor UO_750 (O_750,N_49486,N_48552);
nand UO_751 (O_751,N_49360,N_49490);
or UO_752 (O_752,N_48948,N_49266);
nand UO_753 (O_753,N_48571,N_48800);
nand UO_754 (O_754,N_49532,N_49473);
xor UO_755 (O_755,N_48852,N_48812);
xor UO_756 (O_756,N_49039,N_49491);
nor UO_757 (O_757,N_48259,N_49106);
or UO_758 (O_758,N_48883,N_48066);
or UO_759 (O_759,N_49103,N_48859);
or UO_760 (O_760,N_49936,N_49013);
nor UO_761 (O_761,N_48032,N_49070);
and UO_762 (O_762,N_48277,N_48516);
nor UO_763 (O_763,N_49038,N_48625);
nand UO_764 (O_764,N_48179,N_48912);
xor UO_765 (O_765,N_49929,N_49569);
or UO_766 (O_766,N_48623,N_49092);
nand UO_767 (O_767,N_48957,N_48779);
xnor UO_768 (O_768,N_48441,N_48091);
xnor UO_769 (O_769,N_49592,N_48968);
xnor UO_770 (O_770,N_49322,N_49183);
and UO_771 (O_771,N_48074,N_49957);
xnor UO_772 (O_772,N_48743,N_49605);
or UO_773 (O_773,N_49319,N_48727);
nand UO_774 (O_774,N_48287,N_48728);
and UO_775 (O_775,N_48530,N_48865);
or UO_776 (O_776,N_49931,N_49803);
nor UO_777 (O_777,N_49632,N_49407);
or UO_778 (O_778,N_48593,N_49373);
and UO_779 (O_779,N_49782,N_48139);
nand UO_780 (O_780,N_49140,N_48030);
nand UO_781 (O_781,N_49685,N_48279);
nor UO_782 (O_782,N_48798,N_48686);
or UO_783 (O_783,N_48706,N_48764);
xor UO_784 (O_784,N_49956,N_48712);
xnor UO_785 (O_785,N_49965,N_49749);
and UO_786 (O_786,N_48235,N_48928);
nand UO_787 (O_787,N_48446,N_49940);
and UO_788 (O_788,N_48058,N_48107);
xnor UO_789 (O_789,N_49555,N_49133);
nand UO_790 (O_790,N_49573,N_49127);
xor UO_791 (O_791,N_48078,N_49361);
and UO_792 (O_792,N_49398,N_48594);
and UO_793 (O_793,N_49246,N_49291);
nor UO_794 (O_794,N_48961,N_48456);
and UO_795 (O_795,N_49628,N_49702);
nand UO_796 (O_796,N_49474,N_49204);
or UO_797 (O_797,N_49522,N_48850);
nand UO_798 (O_798,N_48745,N_49326);
xor UO_799 (O_799,N_49521,N_49888);
nor UO_800 (O_800,N_49960,N_49002);
xnor UO_801 (O_801,N_48973,N_49234);
nand UO_802 (O_802,N_49581,N_48772);
nand UO_803 (O_803,N_49827,N_49593);
nor UO_804 (O_804,N_49928,N_48221);
xnor UO_805 (O_805,N_49918,N_49172);
or UO_806 (O_806,N_49489,N_48638);
nand UO_807 (O_807,N_48027,N_48692);
and UO_808 (O_808,N_49753,N_48243);
xnor UO_809 (O_809,N_49740,N_49721);
nor UO_810 (O_810,N_49657,N_49693);
and UO_811 (O_811,N_49445,N_49729);
and UO_812 (O_812,N_49417,N_49123);
nor UO_813 (O_813,N_48796,N_49512);
or UO_814 (O_814,N_48438,N_48610);
and UO_815 (O_815,N_48678,N_49631);
and UO_816 (O_816,N_49379,N_49229);
nor UO_817 (O_817,N_48084,N_49641);
and UO_818 (O_818,N_49300,N_48340);
xnor UO_819 (O_819,N_48910,N_49969);
nand UO_820 (O_820,N_49344,N_49487);
nand UO_821 (O_821,N_49029,N_48693);
nor UO_822 (O_822,N_49076,N_48220);
xnor UO_823 (O_823,N_48877,N_49635);
and UO_824 (O_824,N_48735,N_48783);
and UO_825 (O_825,N_48830,N_48578);
or UO_826 (O_826,N_48919,N_48331);
and UO_827 (O_827,N_49814,N_49182);
nor UO_828 (O_828,N_49270,N_48286);
and UO_829 (O_829,N_49651,N_49137);
or UO_830 (O_830,N_48219,N_49694);
nand UO_831 (O_831,N_48419,N_49647);
nand UO_832 (O_832,N_49060,N_49126);
and UO_833 (O_833,N_48681,N_49273);
or UO_834 (O_834,N_48000,N_48782);
and UO_835 (O_835,N_49130,N_48953);
nand UO_836 (O_836,N_49224,N_49585);
and UO_837 (O_837,N_48920,N_48510);
xnor UO_838 (O_838,N_49086,N_49089);
nor UO_839 (O_839,N_49714,N_49457);
or UO_840 (O_840,N_49372,N_49249);
xnor UO_841 (O_841,N_49777,N_48760);
or UO_842 (O_842,N_48882,N_49356);
xnor UO_843 (O_843,N_48565,N_49952);
nand UO_844 (O_844,N_49493,N_49975);
or UO_845 (O_845,N_49199,N_48634);
xor UO_846 (O_846,N_49195,N_48362);
or UO_847 (O_847,N_49681,N_48389);
nand UO_848 (O_848,N_49680,N_48422);
nand UO_849 (O_849,N_49506,N_48158);
nand UO_850 (O_850,N_48474,N_48448);
and UO_851 (O_851,N_48267,N_48872);
xnor UO_852 (O_852,N_49285,N_49328);
and UO_853 (O_853,N_49482,N_48845);
xnor UO_854 (O_854,N_48715,N_49903);
nor UO_855 (O_855,N_48332,N_48656);
and UO_856 (O_856,N_48304,N_49763);
nand UO_857 (O_857,N_49084,N_48603);
or UO_858 (O_858,N_49514,N_49465);
nand UO_859 (O_859,N_49674,N_48152);
nand UO_860 (O_860,N_48203,N_48604);
or UO_861 (O_861,N_48258,N_49508);
xor UO_862 (O_862,N_48011,N_49099);
xor UO_863 (O_863,N_48112,N_48527);
or UO_864 (O_864,N_49354,N_48720);
nand UO_865 (O_865,N_49061,N_48599);
and UO_866 (O_866,N_48680,N_49005);
nand UO_867 (O_867,N_49864,N_49610);
nor UO_868 (O_868,N_48185,N_49080);
nor UO_869 (O_869,N_49023,N_48394);
and UO_870 (O_870,N_48106,N_48626);
xor UO_871 (O_871,N_48873,N_49066);
nand UO_872 (O_872,N_48705,N_48974);
nand UO_873 (O_873,N_48918,N_49233);
nand UO_874 (O_874,N_48351,N_48374);
nand UO_875 (O_875,N_49861,N_48501);
xor UO_876 (O_876,N_49449,N_49048);
xnor UO_877 (O_877,N_49639,N_49152);
and UO_878 (O_878,N_49653,N_49733);
nand UO_879 (O_879,N_48169,N_48284);
nor UO_880 (O_880,N_48808,N_49093);
nand UO_881 (O_881,N_48832,N_48729);
nand UO_882 (O_882,N_48327,N_49751);
and UO_883 (O_883,N_48904,N_49712);
and UO_884 (O_884,N_49107,N_49033);
nand UO_885 (O_885,N_48582,N_49856);
or UO_886 (O_886,N_48224,N_48668);
xor UO_887 (O_887,N_49704,N_48292);
and UO_888 (O_888,N_48577,N_49840);
or UO_889 (O_889,N_48950,N_49437);
nand UO_890 (O_890,N_49853,N_48417);
and UO_891 (O_891,N_49958,N_49169);
nor UO_892 (O_892,N_48440,N_48163);
or UO_893 (O_893,N_48618,N_48431);
xor UO_894 (O_894,N_48616,N_49200);
or UO_895 (O_895,N_48843,N_49403);
and UO_896 (O_896,N_49301,N_48820);
nor UO_897 (O_897,N_48140,N_49504);
or UO_898 (O_898,N_49404,N_48019);
xor UO_899 (O_899,N_49980,N_48010);
and UO_900 (O_900,N_48092,N_48541);
nand UO_901 (O_901,N_48716,N_49869);
nand UO_902 (O_902,N_49914,N_48647);
or UO_903 (O_903,N_49341,N_48923);
xor UO_904 (O_904,N_49363,N_48807);
xor UO_905 (O_905,N_48181,N_49655);
nand UO_906 (O_906,N_49732,N_49885);
nand UO_907 (O_907,N_48435,N_49649);
or UO_908 (O_908,N_48694,N_49643);
nor UO_909 (O_909,N_49402,N_49754);
or UO_910 (O_910,N_48688,N_48701);
nand UO_911 (O_911,N_49098,N_49058);
xnor UO_912 (O_912,N_48870,N_48167);
and UO_913 (O_913,N_49545,N_49558);
and UO_914 (O_914,N_48135,N_48036);
and UO_915 (O_915,N_49530,N_49603);
and UO_916 (O_916,N_48793,N_49990);
nor UO_917 (O_917,N_48023,N_48662);
nor UO_918 (O_918,N_48790,N_49458);
nand UO_919 (O_919,N_49479,N_48884);
nand UO_920 (O_920,N_49294,N_48899);
or UO_921 (O_921,N_48063,N_48047);
nor UO_922 (O_922,N_48377,N_48402);
or UO_923 (O_923,N_49623,N_49370);
xnor UO_924 (O_924,N_48479,N_49943);
or UO_925 (O_925,N_48311,N_48482);
nand UO_926 (O_926,N_48486,N_48902);
xnor UO_927 (O_927,N_49122,N_48229);
or UO_928 (O_928,N_49838,N_48293);
nand UO_929 (O_929,N_48650,N_48233);
nand UO_930 (O_930,N_49009,N_48228);
or UO_931 (O_931,N_49146,N_49315);
nand UO_932 (O_932,N_49826,N_49325);
nor UO_933 (O_933,N_48724,N_48856);
nor UO_934 (O_934,N_48236,N_49141);
nor UO_935 (O_935,N_49027,N_49884);
xor UO_936 (O_936,N_48407,N_48273);
nor UO_937 (O_937,N_48418,N_49787);
nand UO_938 (O_938,N_49330,N_48914);
nor UO_939 (O_939,N_49456,N_48972);
and UO_940 (O_940,N_49202,N_48350);
nand UO_941 (O_941,N_48788,N_48684);
xnor UO_942 (O_942,N_49912,N_49862);
and UO_943 (O_943,N_48897,N_48079);
and UO_944 (O_944,N_49262,N_49298);
nor UO_945 (O_945,N_49260,N_49539);
nand UO_946 (O_946,N_49439,N_49557);
nand UO_947 (O_947,N_49209,N_48805);
and UO_948 (O_948,N_48251,N_48559);
nor UO_949 (O_949,N_48614,N_49637);
or UO_950 (O_950,N_49977,N_48497);
or UO_951 (O_951,N_48504,N_49336);
xnor UO_952 (O_952,N_49769,N_48561);
or UO_953 (O_953,N_49789,N_48230);
nand UO_954 (O_954,N_49305,N_49230);
or UO_955 (O_955,N_49541,N_49795);
nand UO_956 (O_956,N_49973,N_48841);
nor UO_957 (O_957,N_48111,N_48138);
xnor UO_958 (O_958,N_48556,N_48281);
nor UO_959 (O_959,N_49542,N_49248);
or UO_960 (O_960,N_49670,N_48970);
nor UO_961 (O_961,N_48862,N_49477);
nor UO_962 (O_962,N_48121,N_48345);
and UO_963 (O_963,N_48145,N_48512);
nor UO_964 (O_964,N_48403,N_49087);
xor UO_965 (O_965,N_48589,N_49723);
and UO_966 (O_966,N_48717,N_49682);
and UO_967 (O_967,N_49264,N_48952);
and UO_968 (O_968,N_48875,N_49377);
and UO_969 (O_969,N_48199,N_49756);
nand UO_970 (O_970,N_49034,N_48217);
xnor UO_971 (O_971,N_48703,N_49226);
nand UO_972 (O_972,N_48398,N_48117);
or UO_973 (O_973,N_49553,N_48540);
and UO_974 (O_974,N_48133,N_49331);
xor UO_975 (O_975,N_49994,N_48814);
nand UO_976 (O_976,N_48067,N_48871);
nand UO_977 (O_977,N_49208,N_49775);
xnor UO_978 (O_978,N_49538,N_48879);
nand UO_979 (O_979,N_49295,N_49429);
nor UO_980 (O_980,N_48534,N_48740);
or UO_981 (O_981,N_48055,N_49590);
nand UO_982 (O_982,N_48412,N_49433);
nand UO_983 (O_983,N_49412,N_49352);
nand UO_984 (O_984,N_48300,N_48477);
and UO_985 (O_985,N_48809,N_48147);
and UO_986 (O_986,N_49299,N_48498);
or UO_987 (O_987,N_49422,N_48364);
xnor UO_988 (O_988,N_49317,N_48588);
and UO_989 (O_989,N_49003,N_49081);
or UO_990 (O_990,N_48326,N_48453);
xnor UO_991 (O_991,N_49824,N_48146);
xnor UO_992 (O_992,N_49989,N_48947);
xor UO_993 (O_993,N_48256,N_48489);
and UO_994 (O_994,N_49518,N_48478);
nor UO_995 (O_995,N_49343,N_49346);
and UO_996 (O_996,N_48868,N_49688);
nand UO_997 (O_997,N_49241,N_49511);
and UO_998 (O_998,N_48452,N_48646);
nand UO_999 (O_999,N_48896,N_49857);
nor UO_1000 (O_1000,N_49392,N_49802);
and UO_1001 (O_1001,N_48408,N_48820);
nand UO_1002 (O_1002,N_48634,N_49221);
and UO_1003 (O_1003,N_48806,N_48909);
nand UO_1004 (O_1004,N_48949,N_48159);
xnor UO_1005 (O_1005,N_49531,N_49224);
and UO_1006 (O_1006,N_48612,N_49979);
xnor UO_1007 (O_1007,N_48192,N_49704);
xor UO_1008 (O_1008,N_48995,N_49463);
nor UO_1009 (O_1009,N_49085,N_48395);
and UO_1010 (O_1010,N_48467,N_48211);
nand UO_1011 (O_1011,N_49462,N_49225);
nand UO_1012 (O_1012,N_49126,N_49452);
or UO_1013 (O_1013,N_49711,N_48974);
or UO_1014 (O_1014,N_48826,N_48664);
nor UO_1015 (O_1015,N_48123,N_49916);
or UO_1016 (O_1016,N_48987,N_48173);
nor UO_1017 (O_1017,N_48801,N_48016);
and UO_1018 (O_1018,N_48216,N_49170);
xnor UO_1019 (O_1019,N_49471,N_48500);
nor UO_1020 (O_1020,N_48738,N_48554);
nor UO_1021 (O_1021,N_48665,N_49948);
xnor UO_1022 (O_1022,N_48412,N_49390);
or UO_1023 (O_1023,N_49392,N_48709);
or UO_1024 (O_1024,N_49231,N_49699);
nand UO_1025 (O_1025,N_49406,N_48618);
or UO_1026 (O_1026,N_48278,N_49345);
nand UO_1027 (O_1027,N_49249,N_48071);
nand UO_1028 (O_1028,N_48138,N_48605);
and UO_1029 (O_1029,N_48406,N_48025);
nand UO_1030 (O_1030,N_48734,N_49086);
nand UO_1031 (O_1031,N_49101,N_48231);
nor UO_1032 (O_1032,N_49408,N_48680);
nand UO_1033 (O_1033,N_49837,N_48735);
xor UO_1034 (O_1034,N_49377,N_48426);
or UO_1035 (O_1035,N_49860,N_48069);
nand UO_1036 (O_1036,N_48769,N_48903);
and UO_1037 (O_1037,N_48893,N_48120);
nand UO_1038 (O_1038,N_49407,N_49836);
nor UO_1039 (O_1039,N_49501,N_49707);
nand UO_1040 (O_1040,N_49911,N_49065);
nand UO_1041 (O_1041,N_48397,N_49581);
and UO_1042 (O_1042,N_48086,N_48976);
nor UO_1043 (O_1043,N_48369,N_48230);
nor UO_1044 (O_1044,N_49071,N_48549);
nand UO_1045 (O_1045,N_48960,N_49593);
nor UO_1046 (O_1046,N_48811,N_49429);
nand UO_1047 (O_1047,N_48954,N_48274);
and UO_1048 (O_1048,N_49080,N_48188);
nand UO_1049 (O_1049,N_49820,N_49630);
nand UO_1050 (O_1050,N_48387,N_49026);
nor UO_1051 (O_1051,N_48273,N_49384);
nand UO_1052 (O_1052,N_49582,N_49268);
nand UO_1053 (O_1053,N_49619,N_49718);
nor UO_1054 (O_1054,N_48384,N_48089);
nand UO_1055 (O_1055,N_48137,N_49929);
and UO_1056 (O_1056,N_49775,N_49816);
nand UO_1057 (O_1057,N_49788,N_48246);
or UO_1058 (O_1058,N_49168,N_49895);
or UO_1059 (O_1059,N_49927,N_48580);
nor UO_1060 (O_1060,N_49836,N_49422);
xnor UO_1061 (O_1061,N_48234,N_48052);
xor UO_1062 (O_1062,N_48308,N_49192);
xor UO_1063 (O_1063,N_49940,N_48701);
xor UO_1064 (O_1064,N_48571,N_48135);
nor UO_1065 (O_1065,N_48626,N_49754);
nand UO_1066 (O_1066,N_49119,N_49253);
nand UO_1067 (O_1067,N_49704,N_49439);
or UO_1068 (O_1068,N_49642,N_49804);
nor UO_1069 (O_1069,N_49405,N_48285);
and UO_1070 (O_1070,N_49413,N_48088);
xnor UO_1071 (O_1071,N_48275,N_49052);
and UO_1072 (O_1072,N_48205,N_49585);
nor UO_1073 (O_1073,N_48511,N_48526);
xor UO_1074 (O_1074,N_49218,N_49543);
nand UO_1075 (O_1075,N_49487,N_48630);
xor UO_1076 (O_1076,N_48319,N_49621);
xnor UO_1077 (O_1077,N_48336,N_48666);
and UO_1078 (O_1078,N_49053,N_48299);
and UO_1079 (O_1079,N_48841,N_48741);
nand UO_1080 (O_1080,N_49234,N_48208);
nand UO_1081 (O_1081,N_48679,N_48140);
nor UO_1082 (O_1082,N_49345,N_48046);
xnor UO_1083 (O_1083,N_48312,N_49133);
or UO_1084 (O_1084,N_49549,N_48076);
nand UO_1085 (O_1085,N_48564,N_48087);
nor UO_1086 (O_1086,N_49608,N_48319);
or UO_1087 (O_1087,N_49414,N_48944);
or UO_1088 (O_1088,N_48571,N_48191);
nand UO_1089 (O_1089,N_48335,N_49289);
nor UO_1090 (O_1090,N_48916,N_49909);
nor UO_1091 (O_1091,N_48595,N_48863);
or UO_1092 (O_1092,N_49798,N_49768);
and UO_1093 (O_1093,N_48961,N_49919);
or UO_1094 (O_1094,N_48873,N_49813);
xor UO_1095 (O_1095,N_48532,N_48170);
xor UO_1096 (O_1096,N_48778,N_48181);
nor UO_1097 (O_1097,N_49178,N_49422);
nand UO_1098 (O_1098,N_48367,N_49247);
nor UO_1099 (O_1099,N_49517,N_48999);
nand UO_1100 (O_1100,N_48362,N_48456);
nor UO_1101 (O_1101,N_49228,N_49260);
xnor UO_1102 (O_1102,N_48033,N_48001);
or UO_1103 (O_1103,N_48072,N_49855);
and UO_1104 (O_1104,N_48961,N_49930);
or UO_1105 (O_1105,N_49657,N_48625);
and UO_1106 (O_1106,N_48438,N_48816);
xor UO_1107 (O_1107,N_48060,N_48689);
and UO_1108 (O_1108,N_48597,N_48217);
or UO_1109 (O_1109,N_49497,N_48593);
and UO_1110 (O_1110,N_49154,N_49790);
or UO_1111 (O_1111,N_48330,N_49143);
or UO_1112 (O_1112,N_49745,N_48382);
and UO_1113 (O_1113,N_49233,N_48561);
nor UO_1114 (O_1114,N_48916,N_48258);
nand UO_1115 (O_1115,N_49377,N_48974);
or UO_1116 (O_1116,N_48137,N_49975);
or UO_1117 (O_1117,N_49800,N_48993);
xor UO_1118 (O_1118,N_48757,N_49307);
and UO_1119 (O_1119,N_48907,N_48869);
or UO_1120 (O_1120,N_48572,N_49722);
or UO_1121 (O_1121,N_48476,N_49825);
xor UO_1122 (O_1122,N_48656,N_49404);
nand UO_1123 (O_1123,N_48135,N_48222);
nand UO_1124 (O_1124,N_48038,N_48087);
nor UO_1125 (O_1125,N_49766,N_48295);
xnor UO_1126 (O_1126,N_49517,N_48197);
nand UO_1127 (O_1127,N_49253,N_49044);
nor UO_1128 (O_1128,N_49960,N_49709);
and UO_1129 (O_1129,N_48590,N_49292);
or UO_1130 (O_1130,N_48536,N_49337);
xnor UO_1131 (O_1131,N_49021,N_48771);
nor UO_1132 (O_1132,N_48313,N_48798);
xor UO_1133 (O_1133,N_48672,N_49117);
nor UO_1134 (O_1134,N_49192,N_48204);
and UO_1135 (O_1135,N_49005,N_49891);
xnor UO_1136 (O_1136,N_49405,N_48800);
nand UO_1137 (O_1137,N_48700,N_48416);
nand UO_1138 (O_1138,N_48244,N_48475);
xor UO_1139 (O_1139,N_49965,N_48928);
and UO_1140 (O_1140,N_48687,N_49220);
and UO_1141 (O_1141,N_49559,N_49848);
xor UO_1142 (O_1142,N_49149,N_49968);
and UO_1143 (O_1143,N_49567,N_49989);
or UO_1144 (O_1144,N_48592,N_49622);
nand UO_1145 (O_1145,N_48632,N_49394);
nand UO_1146 (O_1146,N_49505,N_48459);
nand UO_1147 (O_1147,N_48388,N_48170);
xnor UO_1148 (O_1148,N_48924,N_48389);
or UO_1149 (O_1149,N_49658,N_49556);
nor UO_1150 (O_1150,N_49410,N_49177);
nand UO_1151 (O_1151,N_48620,N_48478);
or UO_1152 (O_1152,N_49944,N_48711);
nor UO_1153 (O_1153,N_48354,N_49840);
nand UO_1154 (O_1154,N_48749,N_48397);
nor UO_1155 (O_1155,N_49483,N_49982);
nand UO_1156 (O_1156,N_49701,N_49907);
xnor UO_1157 (O_1157,N_48229,N_48250);
and UO_1158 (O_1158,N_48053,N_48671);
xnor UO_1159 (O_1159,N_48168,N_48794);
nand UO_1160 (O_1160,N_49993,N_49058);
xor UO_1161 (O_1161,N_48284,N_49452);
nand UO_1162 (O_1162,N_49592,N_49450);
nor UO_1163 (O_1163,N_48433,N_48450);
nand UO_1164 (O_1164,N_49318,N_48744);
nand UO_1165 (O_1165,N_48909,N_49409);
nand UO_1166 (O_1166,N_48016,N_49942);
and UO_1167 (O_1167,N_48181,N_48652);
xnor UO_1168 (O_1168,N_48491,N_49178);
nor UO_1169 (O_1169,N_49450,N_48909);
or UO_1170 (O_1170,N_49145,N_49161);
nor UO_1171 (O_1171,N_48470,N_48649);
and UO_1172 (O_1172,N_49662,N_48213);
nand UO_1173 (O_1173,N_48693,N_48424);
and UO_1174 (O_1174,N_49966,N_48115);
nor UO_1175 (O_1175,N_49387,N_48426);
nor UO_1176 (O_1176,N_49070,N_48282);
nand UO_1177 (O_1177,N_49508,N_49581);
nand UO_1178 (O_1178,N_49979,N_49972);
or UO_1179 (O_1179,N_48320,N_48514);
and UO_1180 (O_1180,N_48740,N_49026);
or UO_1181 (O_1181,N_48180,N_49165);
or UO_1182 (O_1182,N_49533,N_48188);
nor UO_1183 (O_1183,N_49992,N_49210);
and UO_1184 (O_1184,N_49211,N_48258);
and UO_1185 (O_1185,N_48458,N_49153);
nor UO_1186 (O_1186,N_48113,N_49622);
and UO_1187 (O_1187,N_48496,N_48232);
nand UO_1188 (O_1188,N_49378,N_48148);
xor UO_1189 (O_1189,N_49699,N_49061);
xor UO_1190 (O_1190,N_48029,N_48614);
and UO_1191 (O_1191,N_48309,N_49483);
nand UO_1192 (O_1192,N_49187,N_49891);
nand UO_1193 (O_1193,N_48218,N_49248);
nor UO_1194 (O_1194,N_48357,N_48754);
nand UO_1195 (O_1195,N_49560,N_49483);
or UO_1196 (O_1196,N_49193,N_49884);
and UO_1197 (O_1197,N_49950,N_49209);
nor UO_1198 (O_1198,N_48126,N_48850);
xor UO_1199 (O_1199,N_48405,N_48212);
and UO_1200 (O_1200,N_49645,N_49835);
nand UO_1201 (O_1201,N_48267,N_48360);
and UO_1202 (O_1202,N_49579,N_48005);
nand UO_1203 (O_1203,N_49856,N_49738);
or UO_1204 (O_1204,N_49219,N_49491);
and UO_1205 (O_1205,N_49802,N_49661);
nor UO_1206 (O_1206,N_49509,N_48153);
or UO_1207 (O_1207,N_49013,N_49199);
nor UO_1208 (O_1208,N_49861,N_49632);
or UO_1209 (O_1209,N_48273,N_49796);
nand UO_1210 (O_1210,N_48804,N_48882);
or UO_1211 (O_1211,N_48191,N_49113);
xor UO_1212 (O_1212,N_49598,N_48763);
xnor UO_1213 (O_1213,N_48130,N_49763);
nor UO_1214 (O_1214,N_48881,N_49179);
nand UO_1215 (O_1215,N_48549,N_49902);
or UO_1216 (O_1216,N_49089,N_49871);
xnor UO_1217 (O_1217,N_49292,N_48849);
or UO_1218 (O_1218,N_49462,N_49040);
and UO_1219 (O_1219,N_48689,N_48056);
xnor UO_1220 (O_1220,N_48569,N_49007);
or UO_1221 (O_1221,N_49912,N_49834);
nor UO_1222 (O_1222,N_48809,N_48321);
and UO_1223 (O_1223,N_49630,N_49119);
or UO_1224 (O_1224,N_49851,N_49580);
or UO_1225 (O_1225,N_48622,N_48360);
nand UO_1226 (O_1226,N_49515,N_48752);
nand UO_1227 (O_1227,N_48976,N_48351);
xor UO_1228 (O_1228,N_49881,N_48203);
and UO_1229 (O_1229,N_48628,N_49711);
or UO_1230 (O_1230,N_48458,N_49081);
nor UO_1231 (O_1231,N_48433,N_48403);
nor UO_1232 (O_1232,N_49819,N_49109);
xnor UO_1233 (O_1233,N_48415,N_49135);
nor UO_1234 (O_1234,N_48610,N_49305);
and UO_1235 (O_1235,N_49395,N_49454);
nand UO_1236 (O_1236,N_48974,N_49425);
nor UO_1237 (O_1237,N_48346,N_48955);
nor UO_1238 (O_1238,N_48258,N_48642);
or UO_1239 (O_1239,N_49448,N_48639);
xor UO_1240 (O_1240,N_49898,N_49094);
nand UO_1241 (O_1241,N_48456,N_49339);
xor UO_1242 (O_1242,N_49045,N_49312);
and UO_1243 (O_1243,N_48279,N_49400);
nand UO_1244 (O_1244,N_48697,N_49216);
nor UO_1245 (O_1245,N_49465,N_48506);
nor UO_1246 (O_1246,N_49347,N_48713);
xnor UO_1247 (O_1247,N_48005,N_49622);
nand UO_1248 (O_1248,N_49030,N_49863);
or UO_1249 (O_1249,N_49500,N_48279);
or UO_1250 (O_1250,N_48782,N_49742);
nand UO_1251 (O_1251,N_48607,N_48952);
xnor UO_1252 (O_1252,N_48215,N_48101);
or UO_1253 (O_1253,N_49286,N_49609);
and UO_1254 (O_1254,N_49828,N_48602);
and UO_1255 (O_1255,N_49652,N_49624);
and UO_1256 (O_1256,N_48655,N_48885);
and UO_1257 (O_1257,N_49818,N_49028);
nand UO_1258 (O_1258,N_48059,N_49403);
xnor UO_1259 (O_1259,N_48474,N_49213);
or UO_1260 (O_1260,N_49597,N_49182);
xor UO_1261 (O_1261,N_49439,N_48430);
nor UO_1262 (O_1262,N_49474,N_49469);
nor UO_1263 (O_1263,N_48578,N_49099);
xnor UO_1264 (O_1264,N_49867,N_49477);
xnor UO_1265 (O_1265,N_49019,N_49899);
and UO_1266 (O_1266,N_48364,N_48114);
xnor UO_1267 (O_1267,N_48634,N_49660);
or UO_1268 (O_1268,N_48865,N_49398);
or UO_1269 (O_1269,N_49676,N_48826);
nor UO_1270 (O_1270,N_49873,N_48453);
or UO_1271 (O_1271,N_48575,N_49640);
nand UO_1272 (O_1272,N_49766,N_48999);
and UO_1273 (O_1273,N_48423,N_48908);
xnor UO_1274 (O_1274,N_48434,N_48331);
xnor UO_1275 (O_1275,N_49202,N_49113);
and UO_1276 (O_1276,N_49225,N_49840);
nand UO_1277 (O_1277,N_49503,N_48965);
and UO_1278 (O_1278,N_49962,N_49227);
nor UO_1279 (O_1279,N_48841,N_49612);
xnor UO_1280 (O_1280,N_49825,N_48630);
xnor UO_1281 (O_1281,N_48190,N_49685);
and UO_1282 (O_1282,N_49420,N_48540);
or UO_1283 (O_1283,N_49893,N_49110);
nand UO_1284 (O_1284,N_49115,N_48539);
nor UO_1285 (O_1285,N_49058,N_49208);
and UO_1286 (O_1286,N_49856,N_49533);
nor UO_1287 (O_1287,N_48184,N_49384);
xnor UO_1288 (O_1288,N_48439,N_49250);
xor UO_1289 (O_1289,N_48913,N_49992);
and UO_1290 (O_1290,N_49702,N_49531);
and UO_1291 (O_1291,N_49328,N_49736);
or UO_1292 (O_1292,N_48111,N_49280);
xor UO_1293 (O_1293,N_48349,N_48470);
or UO_1294 (O_1294,N_49677,N_49803);
xor UO_1295 (O_1295,N_49658,N_49315);
or UO_1296 (O_1296,N_49071,N_48081);
or UO_1297 (O_1297,N_49157,N_49555);
nand UO_1298 (O_1298,N_49232,N_49493);
xnor UO_1299 (O_1299,N_48798,N_48189);
nor UO_1300 (O_1300,N_49615,N_49108);
xor UO_1301 (O_1301,N_48518,N_48282);
nor UO_1302 (O_1302,N_48796,N_49253);
and UO_1303 (O_1303,N_48255,N_48223);
or UO_1304 (O_1304,N_49492,N_48304);
nor UO_1305 (O_1305,N_49863,N_49194);
nor UO_1306 (O_1306,N_49018,N_48688);
nand UO_1307 (O_1307,N_48013,N_49951);
xnor UO_1308 (O_1308,N_48984,N_48704);
or UO_1309 (O_1309,N_49977,N_49285);
nor UO_1310 (O_1310,N_48534,N_48143);
xnor UO_1311 (O_1311,N_49058,N_49353);
or UO_1312 (O_1312,N_49183,N_48546);
xor UO_1313 (O_1313,N_49426,N_48277);
and UO_1314 (O_1314,N_49603,N_49138);
and UO_1315 (O_1315,N_48335,N_49729);
and UO_1316 (O_1316,N_48575,N_48884);
xnor UO_1317 (O_1317,N_48872,N_49146);
and UO_1318 (O_1318,N_48149,N_48294);
and UO_1319 (O_1319,N_49079,N_48905);
and UO_1320 (O_1320,N_48315,N_48044);
nor UO_1321 (O_1321,N_49383,N_49328);
and UO_1322 (O_1322,N_48315,N_49865);
nand UO_1323 (O_1323,N_49065,N_49543);
or UO_1324 (O_1324,N_48129,N_49900);
and UO_1325 (O_1325,N_48126,N_48383);
or UO_1326 (O_1326,N_48828,N_48203);
nor UO_1327 (O_1327,N_49841,N_48657);
nand UO_1328 (O_1328,N_48806,N_48769);
xor UO_1329 (O_1329,N_49638,N_49803);
nor UO_1330 (O_1330,N_48588,N_48738);
nor UO_1331 (O_1331,N_48732,N_49022);
and UO_1332 (O_1332,N_48419,N_48012);
and UO_1333 (O_1333,N_49698,N_48251);
or UO_1334 (O_1334,N_48578,N_49610);
xor UO_1335 (O_1335,N_49009,N_48818);
nand UO_1336 (O_1336,N_48536,N_49641);
xnor UO_1337 (O_1337,N_49229,N_49861);
nor UO_1338 (O_1338,N_48751,N_49048);
nor UO_1339 (O_1339,N_48461,N_49476);
and UO_1340 (O_1340,N_49564,N_49394);
nand UO_1341 (O_1341,N_49336,N_48476);
and UO_1342 (O_1342,N_48084,N_48335);
and UO_1343 (O_1343,N_48354,N_48870);
xnor UO_1344 (O_1344,N_48532,N_49330);
nor UO_1345 (O_1345,N_48238,N_48792);
or UO_1346 (O_1346,N_49409,N_48015);
xnor UO_1347 (O_1347,N_49724,N_49793);
nand UO_1348 (O_1348,N_49251,N_49998);
and UO_1349 (O_1349,N_48541,N_48224);
or UO_1350 (O_1350,N_49727,N_48685);
and UO_1351 (O_1351,N_48485,N_48669);
xnor UO_1352 (O_1352,N_49647,N_49483);
and UO_1353 (O_1353,N_48755,N_49441);
nand UO_1354 (O_1354,N_48209,N_49490);
or UO_1355 (O_1355,N_48887,N_48787);
nand UO_1356 (O_1356,N_48239,N_48514);
or UO_1357 (O_1357,N_49979,N_48385);
nor UO_1358 (O_1358,N_49743,N_48434);
nand UO_1359 (O_1359,N_49996,N_48564);
or UO_1360 (O_1360,N_48096,N_48131);
xnor UO_1361 (O_1361,N_49184,N_49592);
nand UO_1362 (O_1362,N_48042,N_48837);
and UO_1363 (O_1363,N_48058,N_48053);
nor UO_1364 (O_1364,N_49866,N_48553);
nor UO_1365 (O_1365,N_49383,N_49381);
nor UO_1366 (O_1366,N_48214,N_49994);
and UO_1367 (O_1367,N_49540,N_49984);
nor UO_1368 (O_1368,N_48099,N_48274);
nor UO_1369 (O_1369,N_49810,N_48712);
nand UO_1370 (O_1370,N_48561,N_48811);
nor UO_1371 (O_1371,N_48209,N_48882);
xnor UO_1372 (O_1372,N_49285,N_48896);
nand UO_1373 (O_1373,N_48847,N_48200);
xor UO_1374 (O_1374,N_48374,N_49297);
and UO_1375 (O_1375,N_48037,N_48589);
nor UO_1376 (O_1376,N_49498,N_48125);
or UO_1377 (O_1377,N_48712,N_48815);
or UO_1378 (O_1378,N_48523,N_48834);
nor UO_1379 (O_1379,N_48412,N_48844);
or UO_1380 (O_1380,N_49854,N_49373);
xor UO_1381 (O_1381,N_49603,N_49032);
or UO_1382 (O_1382,N_48221,N_49525);
or UO_1383 (O_1383,N_49644,N_49224);
xor UO_1384 (O_1384,N_48245,N_49860);
xor UO_1385 (O_1385,N_49045,N_48617);
nor UO_1386 (O_1386,N_49376,N_49751);
xor UO_1387 (O_1387,N_48517,N_48242);
and UO_1388 (O_1388,N_49849,N_48110);
or UO_1389 (O_1389,N_48363,N_48184);
and UO_1390 (O_1390,N_48451,N_49044);
nand UO_1391 (O_1391,N_49213,N_48055);
and UO_1392 (O_1392,N_49163,N_49724);
or UO_1393 (O_1393,N_48086,N_49059);
or UO_1394 (O_1394,N_48703,N_48140);
nand UO_1395 (O_1395,N_48578,N_49646);
or UO_1396 (O_1396,N_49204,N_49081);
and UO_1397 (O_1397,N_48702,N_49584);
and UO_1398 (O_1398,N_48763,N_48762);
and UO_1399 (O_1399,N_48480,N_49942);
or UO_1400 (O_1400,N_48441,N_48576);
and UO_1401 (O_1401,N_49727,N_48807);
xnor UO_1402 (O_1402,N_49539,N_49658);
nor UO_1403 (O_1403,N_48924,N_48073);
nand UO_1404 (O_1404,N_48417,N_49192);
nor UO_1405 (O_1405,N_49612,N_48737);
nand UO_1406 (O_1406,N_49965,N_49763);
xnor UO_1407 (O_1407,N_49944,N_48090);
xor UO_1408 (O_1408,N_49201,N_48515);
xnor UO_1409 (O_1409,N_49119,N_48329);
nor UO_1410 (O_1410,N_48318,N_48346);
and UO_1411 (O_1411,N_48063,N_48269);
xor UO_1412 (O_1412,N_48603,N_49461);
xnor UO_1413 (O_1413,N_49079,N_49279);
nand UO_1414 (O_1414,N_49612,N_48695);
xnor UO_1415 (O_1415,N_49158,N_48223);
nor UO_1416 (O_1416,N_48133,N_48732);
or UO_1417 (O_1417,N_49530,N_48785);
xor UO_1418 (O_1418,N_48910,N_48370);
and UO_1419 (O_1419,N_48981,N_48227);
xnor UO_1420 (O_1420,N_48623,N_48253);
or UO_1421 (O_1421,N_49475,N_49249);
and UO_1422 (O_1422,N_48090,N_49765);
or UO_1423 (O_1423,N_48358,N_48819);
or UO_1424 (O_1424,N_49743,N_49723);
or UO_1425 (O_1425,N_49804,N_49411);
nor UO_1426 (O_1426,N_49729,N_49582);
nor UO_1427 (O_1427,N_48344,N_49462);
or UO_1428 (O_1428,N_48309,N_49737);
nor UO_1429 (O_1429,N_49805,N_49286);
nor UO_1430 (O_1430,N_49664,N_48054);
or UO_1431 (O_1431,N_49026,N_49305);
nor UO_1432 (O_1432,N_48137,N_48464);
or UO_1433 (O_1433,N_49831,N_48550);
xor UO_1434 (O_1434,N_48874,N_48943);
nand UO_1435 (O_1435,N_48119,N_49896);
and UO_1436 (O_1436,N_49285,N_49688);
and UO_1437 (O_1437,N_49930,N_48931);
nor UO_1438 (O_1438,N_48366,N_49107);
nand UO_1439 (O_1439,N_49482,N_48454);
xor UO_1440 (O_1440,N_49147,N_48319);
or UO_1441 (O_1441,N_48200,N_49519);
xor UO_1442 (O_1442,N_48271,N_49028);
nor UO_1443 (O_1443,N_49918,N_49550);
and UO_1444 (O_1444,N_48858,N_48433);
nand UO_1445 (O_1445,N_48646,N_49114);
nor UO_1446 (O_1446,N_49367,N_49084);
nand UO_1447 (O_1447,N_49855,N_49513);
nand UO_1448 (O_1448,N_49758,N_49490);
nor UO_1449 (O_1449,N_49580,N_49486);
or UO_1450 (O_1450,N_48886,N_49089);
nor UO_1451 (O_1451,N_48069,N_48769);
and UO_1452 (O_1452,N_48331,N_49781);
and UO_1453 (O_1453,N_49624,N_49605);
xnor UO_1454 (O_1454,N_48795,N_49700);
nand UO_1455 (O_1455,N_48854,N_49296);
nor UO_1456 (O_1456,N_48135,N_48538);
nor UO_1457 (O_1457,N_49860,N_48376);
or UO_1458 (O_1458,N_48817,N_49780);
and UO_1459 (O_1459,N_49622,N_48855);
nand UO_1460 (O_1460,N_48908,N_49690);
nor UO_1461 (O_1461,N_49958,N_48586);
nor UO_1462 (O_1462,N_48008,N_49760);
or UO_1463 (O_1463,N_48497,N_48866);
nor UO_1464 (O_1464,N_48715,N_48176);
nand UO_1465 (O_1465,N_49507,N_48576);
or UO_1466 (O_1466,N_49159,N_49215);
xnor UO_1467 (O_1467,N_48054,N_49409);
nand UO_1468 (O_1468,N_49060,N_48229);
nor UO_1469 (O_1469,N_49260,N_48695);
xnor UO_1470 (O_1470,N_49755,N_48979);
nor UO_1471 (O_1471,N_48160,N_49298);
or UO_1472 (O_1472,N_48454,N_49624);
nand UO_1473 (O_1473,N_48003,N_49442);
nor UO_1474 (O_1474,N_49600,N_48411);
nor UO_1475 (O_1475,N_49514,N_48849);
nand UO_1476 (O_1476,N_49588,N_49184);
nor UO_1477 (O_1477,N_49530,N_49708);
and UO_1478 (O_1478,N_48404,N_48306);
xor UO_1479 (O_1479,N_48591,N_48546);
or UO_1480 (O_1480,N_48954,N_49987);
xor UO_1481 (O_1481,N_48018,N_49943);
xor UO_1482 (O_1482,N_48561,N_49447);
or UO_1483 (O_1483,N_48822,N_49972);
nand UO_1484 (O_1484,N_49597,N_48234);
nand UO_1485 (O_1485,N_48055,N_49999);
nand UO_1486 (O_1486,N_49519,N_49742);
nor UO_1487 (O_1487,N_48765,N_48923);
xor UO_1488 (O_1488,N_48832,N_49796);
xnor UO_1489 (O_1489,N_48390,N_49103);
or UO_1490 (O_1490,N_49534,N_49976);
and UO_1491 (O_1491,N_48575,N_48262);
or UO_1492 (O_1492,N_48144,N_49437);
nor UO_1493 (O_1493,N_48707,N_49309);
nand UO_1494 (O_1494,N_48244,N_48444);
xor UO_1495 (O_1495,N_48626,N_49566);
nand UO_1496 (O_1496,N_48639,N_48508);
nand UO_1497 (O_1497,N_48091,N_49308);
nor UO_1498 (O_1498,N_49907,N_49678);
nor UO_1499 (O_1499,N_48217,N_49401);
nor UO_1500 (O_1500,N_49122,N_48956);
nor UO_1501 (O_1501,N_49025,N_49634);
nand UO_1502 (O_1502,N_49079,N_48975);
nand UO_1503 (O_1503,N_49774,N_49067);
nor UO_1504 (O_1504,N_49981,N_49084);
xnor UO_1505 (O_1505,N_48050,N_49911);
nand UO_1506 (O_1506,N_49631,N_48372);
and UO_1507 (O_1507,N_49327,N_49671);
or UO_1508 (O_1508,N_48585,N_48544);
nor UO_1509 (O_1509,N_48781,N_49736);
or UO_1510 (O_1510,N_48468,N_48606);
xor UO_1511 (O_1511,N_48176,N_48350);
and UO_1512 (O_1512,N_49387,N_49613);
nor UO_1513 (O_1513,N_49272,N_48269);
nor UO_1514 (O_1514,N_48912,N_49303);
and UO_1515 (O_1515,N_49572,N_48473);
nand UO_1516 (O_1516,N_48002,N_49370);
or UO_1517 (O_1517,N_48423,N_48582);
xor UO_1518 (O_1518,N_48154,N_48547);
or UO_1519 (O_1519,N_49825,N_49218);
nand UO_1520 (O_1520,N_48258,N_49694);
and UO_1521 (O_1521,N_49399,N_48718);
xnor UO_1522 (O_1522,N_49727,N_48755);
xnor UO_1523 (O_1523,N_49872,N_49276);
nand UO_1524 (O_1524,N_48508,N_49199);
nor UO_1525 (O_1525,N_48604,N_48964);
or UO_1526 (O_1526,N_48771,N_49130);
nor UO_1527 (O_1527,N_49952,N_49901);
nor UO_1528 (O_1528,N_49525,N_49691);
nand UO_1529 (O_1529,N_48938,N_48553);
xor UO_1530 (O_1530,N_49922,N_49613);
nor UO_1531 (O_1531,N_48743,N_49166);
or UO_1532 (O_1532,N_48049,N_49821);
nor UO_1533 (O_1533,N_48217,N_49337);
or UO_1534 (O_1534,N_49142,N_48846);
xnor UO_1535 (O_1535,N_48416,N_48447);
xnor UO_1536 (O_1536,N_48890,N_49802);
or UO_1537 (O_1537,N_49611,N_49066);
nor UO_1538 (O_1538,N_48551,N_49229);
xnor UO_1539 (O_1539,N_48264,N_49655);
xnor UO_1540 (O_1540,N_49555,N_48278);
or UO_1541 (O_1541,N_49697,N_49160);
and UO_1542 (O_1542,N_49131,N_49587);
and UO_1543 (O_1543,N_48101,N_48640);
nand UO_1544 (O_1544,N_49927,N_49064);
xnor UO_1545 (O_1545,N_49447,N_49064);
nand UO_1546 (O_1546,N_48268,N_48250);
and UO_1547 (O_1547,N_48721,N_49024);
or UO_1548 (O_1548,N_49054,N_49257);
or UO_1549 (O_1549,N_48349,N_49485);
nor UO_1550 (O_1550,N_48315,N_49203);
and UO_1551 (O_1551,N_49779,N_48425);
xor UO_1552 (O_1552,N_48556,N_49819);
and UO_1553 (O_1553,N_48918,N_48607);
and UO_1554 (O_1554,N_49362,N_49526);
nor UO_1555 (O_1555,N_49247,N_49752);
xnor UO_1556 (O_1556,N_48124,N_48308);
nand UO_1557 (O_1557,N_48832,N_48160);
nand UO_1558 (O_1558,N_49709,N_49173);
nand UO_1559 (O_1559,N_48596,N_48570);
xor UO_1560 (O_1560,N_48406,N_49957);
nor UO_1561 (O_1561,N_48832,N_49510);
xor UO_1562 (O_1562,N_49575,N_49222);
and UO_1563 (O_1563,N_48935,N_48172);
nor UO_1564 (O_1564,N_49558,N_48347);
and UO_1565 (O_1565,N_49704,N_49175);
nor UO_1566 (O_1566,N_49146,N_49313);
and UO_1567 (O_1567,N_49591,N_49246);
and UO_1568 (O_1568,N_49043,N_48489);
and UO_1569 (O_1569,N_48759,N_48189);
nand UO_1570 (O_1570,N_48821,N_48015);
xor UO_1571 (O_1571,N_49422,N_48493);
nand UO_1572 (O_1572,N_48729,N_48952);
nand UO_1573 (O_1573,N_49915,N_49272);
nor UO_1574 (O_1574,N_48380,N_48920);
nor UO_1575 (O_1575,N_48933,N_49193);
nand UO_1576 (O_1576,N_49704,N_49980);
nor UO_1577 (O_1577,N_49177,N_49227);
nor UO_1578 (O_1578,N_48034,N_49067);
xor UO_1579 (O_1579,N_49680,N_48027);
or UO_1580 (O_1580,N_48146,N_49333);
or UO_1581 (O_1581,N_49766,N_49411);
or UO_1582 (O_1582,N_48651,N_48870);
nand UO_1583 (O_1583,N_48122,N_48228);
or UO_1584 (O_1584,N_49921,N_49011);
or UO_1585 (O_1585,N_49735,N_48804);
nor UO_1586 (O_1586,N_49699,N_48298);
or UO_1587 (O_1587,N_48031,N_49414);
nor UO_1588 (O_1588,N_48505,N_48632);
xor UO_1589 (O_1589,N_49654,N_49709);
nand UO_1590 (O_1590,N_49196,N_48850);
nand UO_1591 (O_1591,N_49247,N_48577);
and UO_1592 (O_1592,N_49828,N_48050);
nor UO_1593 (O_1593,N_48155,N_49359);
nor UO_1594 (O_1594,N_48470,N_48352);
nor UO_1595 (O_1595,N_49048,N_49155);
or UO_1596 (O_1596,N_49674,N_49346);
or UO_1597 (O_1597,N_48569,N_49432);
nand UO_1598 (O_1598,N_48188,N_48557);
and UO_1599 (O_1599,N_48251,N_49393);
xnor UO_1600 (O_1600,N_49010,N_49252);
xor UO_1601 (O_1601,N_49892,N_48000);
nor UO_1602 (O_1602,N_48826,N_48801);
nand UO_1603 (O_1603,N_49959,N_48101);
xnor UO_1604 (O_1604,N_49127,N_49581);
nand UO_1605 (O_1605,N_49317,N_49945);
nor UO_1606 (O_1606,N_48587,N_49044);
and UO_1607 (O_1607,N_49450,N_48395);
nand UO_1608 (O_1608,N_48329,N_48753);
or UO_1609 (O_1609,N_49371,N_48286);
nand UO_1610 (O_1610,N_49649,N_48266);
or UO_1611 (O_1611,N_49012,N_49884);
and UO_1612 (O_1612,N_48777,N_48746);
or UO_1613 (O_1613,N_48760,N_48586);
and UO_1614 (O_1614,N_49403,N_49825);
nor UO_1615 (O_1615,N_48243,N_49122);
or UO_1616 (O_1616,N_48945,N_49663);
nand UO_1617 (O_1617,N_49696,N_49979);
or UO_1618 (O_1618,N_49557,N_48075);
nor UO_1619 (O_1619,N_48960,N_48943);
or UO_1620 (O_1620,N_48496,N_48291);
or UO_1621 (O_1621,N_48458,N_49894);
nand UO_1622 (O_1622,N_49528,N_49157);
xor UO_1623 (O_1623,N_48386,N_49378);
or UO_1624 (O_1624,N_49655,N_49110);
nor UO_1625 (O_1625,N_48439,N_48519);
nor UO_1626 (O_1626,N_49039,N_49921);
nor UO_1627 (O_1627,N_49982,N_48273);
and UO_1628 (O_1628,N_49036,N_49335);
xnor UO_1629 (O_1629,N_49156,N_48429);
xnor UO_1630 (O_1630,N_49453,N_49378);
and UO_1631 (O_1631,N_49722,N_48721);
xnor UO_1632 (O_1632,N_48647,N_49195);
nand UO_1633 (O_1633,N_49521,N_48243);
or UO_1634 (O_1634,N_48520,N_49346);
or UO_1635 (O_1635,N_49602,N_48108);
nor UO_1636 (O_1636,N_48999,N_48775);
or UO_1637 (O_1637,N_48049,N_49064);
xor UO_1638 (O_1638,N_48031,N_49792);
or UO_1639 (O_1639,N_48244,N_48948);
nand UO_1640 (O_1640,N_49830,N_49803);
nor UO_1641 (O_1641,N_48101,N_48117);
or UO_1642 (O_1642,N_49203,N_48393);
nand UO_1643 (O_1643,N_48135,N_48013);
nand UO_1644 (O_1644,N_49052,N_49168);
or UO_1645 (O_1645,N_48234,N_49213);
nand UO_1646 (O_1646,N_48599,N_49834);
xor UO_1647 (O_1647,N_48708,N_48026);
and UO_1648 (O_1648,N_49069,N_48386);
nor UO_1649 (O_1649,N_49704,N_49587);
or UO_1650 (O_1650,N_48562,N_48184);
and UO_1651 (O_1651,N_49773,N_49742);
xor UO_1652 (O_1652,N_49108,N_48218);
and UO_1653 (O_1653,N_48847,N_48348);
nand UO_1654 (O_1654,N_48326,N_49311);
or UO_1655 (O_1655,N_48081,N_48403);
or UO_1656 (O_1656,N_48789,N_48839);
and UO_1657 (O_1657,N_49960,N_48779);
xnor UO_1658 (O_1658,N_48098,N_48123);
nand UO_1659 (O_1659,N_49915,N_48453);
nand UO_1660 (O_1660,N_49416,N_48240);
and UO_1661 (O_1661,N_49211,N_49758);
and UO_1662 (O_1662,N_49119,N_49044);
and UO_1663 (O_1663,N_49701,N_49173);
nor UO_1664 (O_1664,N_48860,N_49706);
nand UO_1665 (O_1665,N_48032,N_48299);
xor UO_1666 (O_1666,N_48429,N_49927);
and UO_1667 (O_1667,N_48138,N_49207);
nand UO_1668 (O_1668,N_48263,N_49089);
nor UO_1669 (O_1669,N_49852,N_49705);
nand UO_1670 (O_1670,N_48239,N_48476);
nor UO_1671 (O_1671,N_48072,N_48497);
nor UO_1672 (O_1672,N_48107,N_48858);
xor UO_1673 (O_1673,N_48241,N_48512);
or UO_1674 (O_1674,N_48203,N_49087);
nand UO_1675 (O_1675,N_49133,N_48596);
and UO_1676 (O_1676,N_49049,N_48229);
nand UO_1677 (O_1677,N_49398,N_49533);
or UO_1678 (O_1678,N_48136,N_49767);
xor UO_1679 (O_1679,N_48614,N_48217);
nor UO_1680 (O_1680,N_49151,N_48093);
and UO_1681 (O_1681,N_49159,N_49249);
or UO_1682 (O_1682,N_49796,N_48151);
nand UO_1683 (O_1683,N_49723,N_48787);
or UO_1684 (O_1684,N_49687,N_48430);
xor UO_1685 (O_1685,N_49504,N_49164);
or UO_1686 (O_1686,N_48833,N_49244);
or UO_1687 (O_1687,N_48960,N_49000);
nor UO_1688 (O_1688,N_49935,N_49298);
nand UO_1689 (O_1689,N_49724,N_48496);
and UO_1690 (O_1690,N_48436,N_49360);
or UO_1691 (O_1691,N_49291,N_48454);
or UO_1692 (O_1692,N_49548,N_49452);
nor UO_1693 (O_1693,N_48533,N_48348);
or UO_1694 (O_1694,N_49426,N_49859);
and UO_1695 (O_1695,N_48115,N_49320);
nand UO_1696 (O_1696,N_48729,N_48423);
nand UO_1697 (O_1697,N_48699,N_49510);
or UO_1698 (O_1698,N_49342,N_49747);
xor UO_1699 (O_1699,N_49847,N_48325);
nor UO_1700 (O_1700,N_48445,N_48865);
nand UO_1701 (O_1701,N_48541,N_49124);
nor UO_1702 (O_1702,N_49828,N_48033);
or UO_1703 (O_1703,N_49114,N_48797);
xnor UO_1704 (O_1704,N_48625,N_49978);
or UO_1705 (O_1705,N_49560,N_49196);
xnor UO_1706 (O_1706,N_49395,N_49974);
or UO_1707 (O_1707,N_48035,N_49038);
nand UO_1708 (O_1708,N_49727,N_49208);
and UO_1709 (O_1709,N_49189,N_48545);
xnor UO_1710 (O_1710,N_49711,N_49994);
nand UO_1711 (O_1711,N_49770,N_49889);
nand UO_1712 (O_1712,N_49006,N_49956);
or UO_1713 (O_1713,N_49208,N_49503);
or UO_1714 (O_1714,N_48056,N_49463);
or UO_1715 (O_1715,N_48351,N_49877);
nor UO_1716 (O_1716,N_48344,N_49959);
or UO_1717 (O_1717,N_49180,N_49459);
or UO_1718 (O_1718,N_49531,N_48051);
nor UO_1719 (O_1719,N_49406,N_49224);
and UO_1720 (O_1720,N_49557,N_48198);
and UO_1721 (O_1721,N_49495,N_48944);
nand UO_1722 (O_1722,N_49933,N_48597);
nor UO_1723 (O_1723,N_48515,N_49192);
or UO_1724 (O_1724,N_48201,N_49037);
xnor UO_1725 (O_1725,N_49178,N_49225);
xor UO_1726 (O_1726,N_48069,N_49119);
and UO_1727 (O_1727,N_49438,N_49572);
and UO_1728 (O_1728,N_48856,N_49983);
nor UO_1729 (O_1729,N_49514,N_48883);
nor UO_1730 (O_1730,N_49082,N_49946);
nor UO_1731 (O_1731,N_48510,N_48648);
or UO_1732 (O_1732,N_48471,N_49751);
or UO_1733 (O_1733,N_48803,N_49118);
or UO_1734 (O_1734,N_48651,N_48176);
or UO_1735 (O_1735,N_48072,N_48077);
and UO_1736 (O_1736,N_49350,N_49406);
or UO_1737 (O_1737,N_48065,N_49748);
xnor UO_1738 (O_1738,N_49321,N_48952);
xnor UO_1739 (O_1739,N_49185,N_48677);
and UO_1740 (O_1740,N_49158,N_49735);
nand UO_1741 (O_1741,N_49106,N_48122);
or UO_1742 (O_1742,N_49580,N_49521);
nand UO_1743 (O_1743,N_49478,N_49733);
nand UO_1744 (O_1744,N_48987,N_48723);
nand UO_1745 (O_1745,N_49639,N_49545);
nand UO_1746 (O_1746,N_49913,N_48719);
and UO_1747 (O_1747,N_49254,N_48079);
nor UO_1748 (O_1748,N_48082,N_48895);
or UO_1749 (O_1749,N_48156,N_48650);
and UO_1750 (O_1750,N_48937,N_49639);
xor UO_1751 (O_1751,N_48061,N_49161);
nor UO_1752 (O_1752,N_49634,N_49446);
nor UO_1753 (O_1753,N_49778,N_49840);
nor UO_1754 (O_1754,N_48165,N_48436);
nor UO_1755 (O_1755,N_48512,N_49664);
nand UO_1756 (O_1756,N_49608,N_49747);
nor UO_1757 (O_1757,N_49981,N_49988);
nor UO_1758 (O_1758,N_49747,N_48520);
nor UO_1759 (O_1759,N_49173,N_49787);
and UO_1760 (O_1760,N_48605,N_49297);
nor UO_1761 (O_1761,N_49613,N_49528);
nand UO_1762 (O_1762,N_49437,N_48066);
nor UO_1763 (O_1763,N_48286,N_49543);
xnor UO_1764 (O_1764,N_48003,N_49216);
xnor UO_1765 (O_1765,N_49841,N_49407);
and UO_1766 (O_1766,N_49329,N_49316);
and UO_1767 (O_1767,N_48963,N_49761);
nor UO_1768 (O_1768,N_48238,N_49265);
nand UO_1769 (O_1769,N_48769,N_49184);
nor UO_1770 (O_1770,N_49881,N_48472);
nor UO_1771 (O_1771,N_48293,N_49709);
nor UO_1772 (O_1772,N_48934,N_48376);
nor UO_1773 (O_1773,N_48442,N_49632);
nand UO_1774 (O_1774,N_48947,N_49988);
nand UO_1775 (O_1775,N_48540,N_49993);
and UO_1776 (O_1776,N_49453,N_48098);
or UO_1777 (O_1777,N_49751,N_48613);
and UO_1778 (O_1778,N_48745,N_48853);
and UO_1779 (O_1779,N_48284,N_49723);
and UO_1780 (O_1780,N_48076,N_49648);
nand UO_1781 (O_1781,N_49957,N_49484);
nand UO_1782 (O_1782,N_49607,N_49487);
nor UO_1783 (O_1783,N_48149,N_49776);
nand UO_1784 (O_1784,N_49699,N_49534);
xor UO_1785 (O_1785,N_48364,N_49102);
nand UO_1786 (O_1786,N_48688,N_49254);
and UO_1787 (O_1787,N_49059,N_49797);
nor UO_1788 (O_1788,N_48914,N_48824);
nor UO_1789 (O_1789,N_49874,N_49434);
nand UO_1790 (O_1790,N_49503,N_48757);
xor UO_1791 (O_1791,N_48809,N_49132);
nand UO_1792 (O_1792,N_49301,N_49936);
nand UO_1793 (O_1793,N_48626,N_48182);
xor UO_1794 (O_1794,N_49184,N_49211);
xnor UO_1795 (O_1795,N_48288,N_48848);
or UO_1796 (O_1796,N_48998,N_49256);
nand UO_1797 (O_1797,N_48163,N_48445);
or UO_1798 (O_1798,N_48993,N_48584);
nor UO_1799 (O_1799,N_48246,N_49030);
nor UO_1800 (O_1800,N_48381,N_49817);
or UO_1801 (O_1801,N_48436,N_49366);
nor UO_1802 (O_1802,N_48081,N_48373);
nand UO_1803 (O_1803,N_48642,N_48517);
and UO_1804 (O_1804,N_49869,N_48699);
nand UO_1805 (O_1805,N_48399,N_48334);
xnor UO_1806 (O_1806,N_49568,N_49818);
nand UO_1807 (O_1807,N_48007,N_48734);
xnor UO_1808 (O_1808,N_49059,N_49040);
or UO_1809 (O_1809,N_49568,N_48261);
xor UO_1810 (O_1810,N_49753,N_48372);
and UO_1811 (O_1811,N_49092,N_48509);
nand UO_1812 (O_1812,N_49484,N_48403);
nand UO_1813 (O_1813,N_49362,N_49377);
xor UO_1814 (O_1814,N_49853,N_48215);
xor UO_1815 (O_1815,N_48080,N_49956);
nor UO_1816 (O_1816,N_48776,N_48151);
nor UO_1817 (O_1817,N_48506,N_48076);
nor UO_1818 (O_1818,N_48370,N_48637);
or UO_1819 (O_1819,N_49524,N_48982);
and UO_1820 (O_1820,N_48107,N_49474);
or UO_1821 (O_1821,N_48668,N_49590);
nand UO_1822 (O_1822,N_48837,N_49819);
nand UO_1823 (O_1823,N_49361,N_48663);
or UO_1824 (O_1824,N_48555,N_48811);
and UO_1825 (O_1825,N_49109,N_48671);
or UO_1826 (O_1826,N_49610,N_49674);
or UO_1827 (O_1827,N_48014,N_48247);
and UO_1828 (O_1828,N_48609,N_48313);
xnor UO_1829 (O_1829,N_48469,N_48204);
xnor UO_1830 (O_1830,N_49310,N_48497);
nor UO_1831 (O_1831,N_49917,N_48260);
or UO_1832 (O_1832,N_49125,N_49899);
xor UO_1833 (O_1833,N_49337,N_49085);
nor UO_1834 (O_1834,N_48317,N_49921);
or UO_1835 (O_1835,N_48682,N_49305);
and UO_1836 (O_1836,N_48595,N_49336);
xnor UO_1837 (O_1837,N_49432,N_49923);
nand UO_1838 (O_1838,N_49584,N_48833);
nand UO_1839 (O_1839,N_49747,N_48729);
or UO_1840 (O_1840,N_49858,N_48790);
nor UO_1841 (O_1841,N_49564,N_48093);
xnor UO_1842 (O_1842,N_48064,N_49570);
nand UO_1843 (O_1843,N_48127,N_48577);
or UO_1844 (O_1844,N_49171,N_49538);
and UO_1845 (O_1845,N_49294,N_48275);
or UO_1846 (O_1846,N_49180,N_49075);
nor UO_1847 (O_1847,N_48970,N_48991);
nand UO_1848 (O_1848,N_48340,N_49369);
nor UO_1849 (O_1849,N_48518,N_49646);
xnor UO_1850 (O_1850,N_49263,N_48368);
or UO_1851 (O_1851,N_49237,N_49880);
and UO_1852 (O_1852,N_49488,N_48021);
and UO_1853 (O_1853,N_48023,N_49634);
or UO_1854 (O_1854,N_49886,N_49791);
nor UO_1855 (O_1855,N_48517,N_48440);
or UO_1856 (O_1856,N_49936,N_48058);
nor UO_1857 (O_1857,N_48176,N_49419);
and UO_1858 (O_1858,N_49213,N_49800);
xor UO_1859 (O_1859,N_48295,N_48687);
nor UO_1860 (O_1860,N_48306,N_49762);
or UO_1861 (O_1861,N_48886,N_49304);
nor UO_1862 (O_1862,N_49992,N_49648);
and UO_1863 (O_1863,N_49622,N_49450);
and UO_1864 (O_1864,N_49541,N_48815);
xor UO_1865 (O_1865,N_48917,N_49900);
nor UO_1866 (O_1866,N_49869,N_48279);
nor UO_1867 (O_1867,N_48076,N_49572);
xor UO_1868 (O_1868,N_49781,N_49431);
nand UO_1869 (O_1869,N_49847,N_49744);
nor UO_1870 (O_1870,N_48374,N_49467);
and UO_1871 (O_1871,N_48247,N_49567);
and UO_1872 (O_1872,N_48074,N_48013);
or UO_1873 (O_1873,N_49801,N_48281);
or UO_1874 (O_1874,N_49954,N_48693);
nor UO_1875 (O_1875,N_49232,N_48047);
xor UO_1876 (O_1876,N_48841,N_49326);
or UO_1877 (O_1877,N_49701,N_48398);
nor UO_1878 (O_1878,N_49191,N_48149);
nor UO_1879 (O_1879,N_49410,N_48984);
xnor UO_1880 (O_1880,N_49762,N_48061);
nand UO_1881 (O_1881,N_48968,N_48863);
and UO_1882 (O_1882,N_48271,N_48558);
or UO_1883 (O_1883,N_49879,N_49122);
nor UO_1884 (O_1884,N_48615,N_48022);
and UO_1885 (O_1885,N_48730,N_48967);
or UO_1886 (O_1886,N_49753,N_49058);
xnor UO_1887 (O_1887,N_48960,N_49714);
nor UO_1888 (O_1888,N_48885,N_48220);
or UO_1889 (O_1889,N_49192,N_48554);
nor UO_1890 (O_1890,N_49821,N_48422);
nor UO_1891 (O_1891,N_48033,N_48824);
or UO_1892 (O_1892,N_49604,N_48683);
or UO_1893 (O_1893,N_49885,N_49006);
or UO_1894 (O_1894,N_48488,N_49117);
and UO_1895 (O_1895,N_49016,N_48439);
and UO_1896 (O_1896,N_49961,N_49759);
nand UO_1897 (O_1897,N_49791,N_49559);
or UO_1898 (O_1898,N_48936,N_48070);
or UO_1899 (O_1899,N_49569,N_48413);
or UO_1900 (O_1900,N_48314,N_49915);
nor UO_1901 (O_1901,N_48770,N_48641);
nand UO_1902 (O_1902,N_48189,N_49132);
xor UO_1903 (O_1903,N_49498,N_48255);
and UO_1904 (O_1904,N_49462,N_48788);
nand UO_1905 (O_1905,N_49674,N_49427);
and UO_1906 (O_1906,N_49086,N_48492);
xor UO_1907 (O_1907,N_48659,N_48660);
and UO_1908 (O_1908,N_48650,N_48129);
and UO_1909 (O_1909,N_48290,N_49881);
xor UO_1910 (O_1910,N_48462,N_49342);
xnor UO_1911 (O_1911,N_49937,N_49595);
xnor UO_1912 (O_1912,N_48612,N_49116);
nand UO_1913 (O_1913,N_48866,N_49044);
nor UO_1914 (O_1914,N_49339,N_49164);
xor UO_1915 (O_1915,N_48065,N_49688);
nand UO_1916 (O_1916,N_49331,N_49700);
nor UO_1917 (O_1917,N_48146,N_49970);
nor UO_1918 (O_1918,N_49576,N_48907);
or UO_1919 (O_1919,N_48356,N_48921);
xor UO_1920 (O_1920,N_49203,N_49693);
and UO_1921 (O_1921,N_49679,N_48620);
xnor UO_1922 (O_1922,N_49328,N_49913);
xnor UO_1923 (O_1923,N_48066,N_49386);
or UO_1924 (O_1924,N_49897,N_48278);
and UO_1925 (O_1925,N_48668,N_48561);
nand UO_1926 (O_1926,N_48059,N_49797);
nand UO_1927 (O_1927,N_48785,N_48414);
nor UO_1928 (O_1928,N_48091,N_48940);
xor UO_1929 (O_1929,N_48144,N_49203);
and UO_1930 (O_1930,N_49881,N_48825);
and UO_1931 (O_1931,N_48205,N_49553);
and UO_1932 (O_1932,N_49441,N_48740);
or UO_1933 (O_1933,N_48242,N_48789);
and UO_1934 (O_1934,N_48367,N_49857);
nor UO_1935 (O_1935,N_49616,N_48504);
nor UO_1936 (O_1936,N_48437,N_48805);
or UO_1937 (O_1937,N_48355,N_48812);
nand UO_1938 (O_1938,N_49278,N_49204);
nor UO_1939 (O_1939,N_48765,N_49011);
nor UO_1940 (O_1940,N_49075,N_49124);
xnor UO_1941 (O_1941,N_48361,N_49144);
or UO_1942 (O_1942,N_48596,N_49758);
xnor UO_1943 (O_1943,N_49754,N_49460);
xnor UO_1944 (O_1944,N_48157,N_49638);
or UO_1945 (O_1945,N_48654,N_48796);
and UO_1946 (O_1946,N_49247,N_49681);
or UO_1947 (O_1947,N_48726,N_49140);
nor UO_1948 (O_1948,N_48812,N_49627);
or UO_1949 (O_1949,N_49768,N_49613);
or UO_1950 (O_1950,N_48195,N_48641);
or UO_1951 (O_1951,N_49635,N_48760);
and UO_1952 (O_1952,N_48435,N_48212);
nand UO_1953 (O_1953,N_49761,N_49726);
and UO_1954 (O_1954,N_49525,N_48497);
nor UO_1955 (O_1955,N_49915,N_48363);
nand UO_1956 (O_1956,N_48336,N_49593);
nand UO_1957 (O_1957,N_49763,N_48526);
nand UO_1958 (O_1958,N_49244,N_49065);
nor UO_1959 (O_1959,N_49953,N_49202);
and UO_1960 (O_1960,N_49334,N_48509);
and UO_1961 (O_1961,N_48566,N_49761);
nand UO_1962 (O_1962,N_49202,N_48111);
nor UO_1963 (O_1963,N_49065,N_48982);
nand UO_1964 (O_1964,N_49042,N_48798);
or UO_1965 (O_1965,N_48824,N_49772);
and UO_1966 (O_1966,N_48995,N_48772);
or UO_1967 (O_1967,N_48504,N_49018);
nand UO_1968 (O_1968,N_49644,N_49581);
nor UO_1969 (O_1969,N_49835,N_49012);
nand UO_1970 (O_1970,N_48999,N_48845);
xor UO_1971 (O_1971,N_48641,N_48944);
or UO_1972 (O_1972,N_49078,N_49926);
nor UO_1973 (O_1973,N_48799,N_48746);
xor UO_1974 (O_1974,N_49225,N_48349);
and UO_1975 (O_1975,N_48159,N_49729);
xnor UO_1976 (O_1976,N_49707,N_48875);
nand UO_1977 (O_1977,N_49554,N_48126);
xnor UO_1978 (O_1978,N_49783,N_49694);
and UO_1979 (O_1979,N_49660,N_48110);
or UO_1980 (O_1980,N_49928,N_48366);
xnor UO_1981 (O_1981,N_48409,N_48505);
or UO_1982 (O_1982,N_49568,N_48367);
xnor UO_1983 (O_1983,N_48073,N_49884);
or UO_1984 (O_1984,N_49702,N_48647);
nand UO_1985 (O_1985,N_48099,N_48715);
nor UO_1986 (O_1986,N_49939,N_49195);
nand UO_1987 (O_1987,N_49511,N_48756);
or UO_1988 (O_1988,N_48960,N_48885);
or UO_1989 (O_1989,N_48539,N_48273);
nand UO_1990 (O_1990,N_48626,N_49246);
and UO_1991 (O_1991,N_48315,N_49378);
and UO_1992 (O_1992,N_49667,N_48590);
nand UO_1993 (O_1993,N_48990,N_48531);
or UO_1994 (O_1994,N_48019,N_49427);
nand UO_1995 (O_1995,N_48470,N_48292);
xor UO_1996 (O_1996,N_48369,N_49251);
or UO_1997 (O_1997,N_48755,N_48834);
or UO_1998 (O_1998,N_49896,N_48976);
nor UO_1999 (O_1999,N_49543,N_48341);
and UO_2000 (O_2000,N_49773,N_48511);
xor UO_2001 (O_2001,N_49758,N_49838);
and UO_2002 (O_2002,N_49862,N_49972);
and UO_2003 (O_2003,N_48451,N_49805);
nor UO_2004 (O_2004,N_48311,N_48040);
nand UO_2005 (O_2005,N_49904,N_48042);
nor UO_2006 (O_2006,N_48068,N_48744);
or UO_2007 (O_2007,N_49726,N_48531);
xor UO_2008 (O_2008,N_49055,N_49092);
nand UO_2009 (O_2009,N_48286,N_48556);
and UO_2010 (O_2010,N_49196,N_48098);
xnor UO_2011 (O_2011,N_48531,N_48473);
and UO_2012 (O_2012,N_49748,N_49236);
xor UO_2013 (O_2013,N_49558,N_49610);
nand UO_2014 (O_2014,N_48079,N_48807);
nor UO_2015 (O_2015,N_48370,N_48857);
and UO_2016 (O_2016,N_48296,N_48833);
or UO_2017 (O_2017,N_48389,N_48349);
xor UO_2018 (O_2018,N_49974,N_48424);
and UO_2019 (O_2019,N_48101,N_48691);
and UO_2020 (O_2020,N_49632,N_48157);
xnor UO_2021 (O_2021,N_49930,N_48974);
nand UO_2022 (O_2022,N_49163,N_49059);
xor UO_2023 (O_2023,N_49095,N_49367);
and UO_2024 (O_2024,N_48450,N_48690);
and UO_2025 (O_2025,N_49613,N_49632);
or UO_2026 (O_2026,N_49825,N_49960);
nor UO_2027 (O_2027,N_49686,N_49628);
xor UO_2028 (O_2028,N_49701,N_49275);
and UO_2029 (O_2029,N_49531,N_48674);
xnor UO_2030 (O_2030,N_49578,N_48021);
or UO_2031 (O_2031,N_49446,N_48700);
and UO_2032 (O_2032,N_49853,N_48369);
or UO_2033 (O_2033,N_48715,N_49994);
xnor UO_2034 (O_2034,N_48915,N_48751);
and UO_2035 (O_2035,N_48480,N_48429);
xor UO_2036 (O_2036,N_49073,N_48182);
xnor UO_2037 (O_2037,N_48399,N_48766);
xnor UO_2038 (O_2038,N_49154,N_48037);
nand UO_2039 (O_2039,N_49796,N_48811);
and UO_2040 (O_2040,N_49674,N_49371);
and UO_2041 (O_2041,N_49574,N_49181);
nor UO_2042 (O_2042,N_48420,N_49576);
and UO_2043 (O_2043,N_49854,N_48940);
nor UO_2044 (O_2044,N_48658,N_49936);
nand UO_2045 (O_2045,N_49760,N_48664);
and UO_2046 (O_2046,N_48271,N_48765);
or UO_2047 (O_2047,N_49970,N_49383);
nand UO_2048 (O_2048,N_49239,N_49838);
xor UO_2049 (O_2049,N_49599,N_48216);
xor UO_2050 (O_2050,N_48241,N_48144);
nand UO_2051 (O_2051,N_48085,N_49837);
and UO_2052 (O_2052,N_48140,N_48669);
or UO_2053 (O_2053,N_48656,N_48318);
nor UO_2054 (O_2054,N_48360,N_49545);
and UO_2055 (O_2055,N_48324,N_48784);
xnor UO_2056 (O_2056,N_49119,N_49154);
nand UO_2057 (O_2057,N_48824,N_48155);
and UO_2058 (O_2058,N_49964,N_48547);
nand UO_2059 (O_2059,N_49975,N_49710);
nand UO_2060 (O_2060,N_49566,N_48650);
and UO_2061 (O_2061,N_48568,N_48223);
or UO_2062 (O_2062,N_49196,N_49685);
or UO_2063 (O_2063,N_48099,N_49933);
or UO_2064 (O_2064,N_48617,N_48682);
xnor UO_2065 (O_2065,N_49573,N_49793);
or UO_2066 (O_2066,N_48653,N_49759);
and UO_2067 (O_2067,N_49033,N_49248);
nor UO_2068 (O_2068,N_48528,N_49740);
and UO_2069 (O_2069,N_48412,N_48195);
nand UO_2070 (O_2070,N_49941,N_49827);
xnor UO_2071 (O_2071,N_48103,N_49794);
nand UO_2072 (O_2072,N_48297,N_49967);
xnor UO_2073 (O_2073,N_49386,N_49881);
or UO_2074 (O_2074,N_49227,N_49706);
or UO_2075 (O_2075,N_48261,N_49467);
nor UO_2076 (O_2076,N_48521,N_48998);
xnor UO_2077 (O_2077,N_49650,N_48551);
or UO_2078 (O_2078,N_48624,N_48213);
nand UO_2079 (O_2079,N_49050,N_49040);
xor UO_2080 (O_2080,N_49573,N_48031);
nand UO_2081 (O_2081,N_48995,N_48466);
and UO_2082 (O_2082,N_49502,N_49876);
nor UO_2083 (O_2083,N_49000,N_49649);
xor UO_2084 (O_2084,N_48917,N_48096);
or UO_2085 (O_2085,N_49647,N_48868);
or UO_2086 (O_2086,N_48980,N_48440);
xor UO_2087 (O_2087,N_49621,N_48274);
and UO_2088 (O_2088,N_49574,N_49304);
xor UO_2089 (O_2089,N_49307,N_49406);
or UO_2090 (O_2090,N_48791,N_48727);
nor UO_2091 (O_2091,N_48011,N_48689);
xnor UO_2092 (O_2092,N_49158,N_49367);
or UO_2093 (O_2093,N_49319,N_49155);
nor UO_2094 (O_2094,N_48618,N_48267);
nor UO_2095 (O_2095,N_49709,N_49659);
or UO_2096 (O_2096,N_49683,N_49707);
or UO_2097 (O_2097,N_49527,N_48251);
and UO_2098 (O_2098,N_48712,N_48018);
xnor UO_2099 (O_2099,N_49563,N_49037);
and UO_2100 (O_2100,N_49745,N_49423);
or UO_2101 (O_2101,N_49236,N_49266);
or UO_2102 (O_2102,N_49084,N_48567);
or UO_2103 (O_2103,N_48000,N_49375);
nor UO_2104 (O_2104,N_49277,N_49676);
nor UO_2105 (O_2105,N_48474,N_49552);
nand UO_2106 (O_2106,N_49092,N_49696);
nor UO_2107 (O_2107,N_49303,N_48938);
or UO_2108 (O_2108,N_48175,N_48787);
nand UO_2109 (O_2109,N_48372,N_49097);
xor UO_2110 (O_2110,N_49317,N_49229);
nand UO_2111 (O_2111,N_48254,N_48100);
and UO_2112 (O_2112,N_49714,N_48398);
or UO_2113 (O_2113,N_49580,N_49282);
and UO_2114 (O_2114,N_48593,N_48697);
or UO_2115 (O_2115,N_49726,N_49463);
and UO_2116 (O_2116,N_48783,N_48740);
nand UO_2117 (O_2117,N_49609,N_49343);
nand UO_2118 (O_2118,N_48420,N_48197);
xor UO_2119 (O_2119,N_48233,N_49126);
or UO_2120 (O_2120,N_48008,N_49848);
nor UO_2121 (O_2121,N_49446,N_49833);
nor UO_2122 (O_2122,N_49112,N_49698);
or UO_2123 (O_2123,N_49118,N_48556);
or UO_2124 (O_2124,N_48472,N_48247);
xnor UO_2125 (O_2125,N_48874,N_49247);
nand UO_2126 (O_2126,N_49483,N_49259);
nor UO_2127 (O_2127,N_48401,N_49342);
nand UO_2128 (O_2128,N_49742,N_48450);
or UO_2129 (O_2129,N_49318,N_48715);
and UO_2130 (O_2130,N_48835,N_48500);
and UO_2131 (O_2131,N_48027,N_49187);
xor UO_2132 (O_2132,N_49951,N_48665);
and UO_2133 (O_2133,N_48100,N_48314);
or UO_2134 (O_2134,N_49269,N_48673);
xor UO_2135 (O_2135,N_49948,N_49316);
xnor UO_2136 (O_2136,N_49076,N_49164);
nor UO_2137 (O_2137,N_49198,N_48948);
nand UO_2138 (O_2138,N_49142,N_48535);
nor UO_2139 (O_2139,N_48586,N_49705);
or UO_2140 (O_2140,N_48464,N_49418);
xnor UO_2141 (O_2141,N_49685,N_48928);
xnor UO_2142 (O_2142,N_49812,N_48899);
nor UO_2143 (O_2143,N_49245,N_48752);
and UO_2144 (O_2144,N_49613,N_49704);
and UO_2145 (O_2145,N_48540,N_49981);
and UO_2146 (O_2146,N_48874,N_49051);
nand UO_2147 (O_2147,N_49039,N_49725);
nor UO_2148 (O_2148,N_49469,N_48781);
and UO_2149 (O_2149,N_48367,N_48174);
xnor UO_2150 (O_2150,N_49593,N_48232);
nor UO_2151 (O_2151,N_49296,N_49465);
nor UO_2152 (O_2152,N_48568,N_49899);
or UO_2153 (O_2153,N_48924,N_49105);
nor UO_2154 (O_2154,N_48306,N_49975);
nor UO_2155 (O_2155,N_49388,N_48841);
or UO_2156 (O_2156,N_48552,N_49974);
nor UO_2157 (O_2157,N_48169,N_48574);
xor UO_2158 (O_2158,N_49332,N_48403);
or UO_2159 (O_2159,N_49908,N_49536);
nand UO_2160 (O_2160,N_48080,N_48546);
or UO_2161 (O_2161,N_48847,N_49807);
nor UO_2162 (O_2162,N_48951,N_49520);
nand UO_2163 (O_2163,N_48567,N_48753);
or UO_2164 (O_2164,N_48872,N_49988);
xnor UO_2165 (O_2165,N_49881,N_49863);
nor UO_2166 (O_2166,N_48795,N_48907);
xnor UO_2167 (O_2167,N_49897,N_49002);
nand UO_2168 (O_2168,N_48782,N_49686);
xnor UO_2169 (O_2169,N_49288,N_48167);
nand UO_2170 (O_2170,N_48484,N_48464);
nand UO_2171 (O_2171,N_48093,N_48460);
xnor UO_2172 (O_2172,N_49582,N_48249);
and UO_2173 (O_2173,N_49558,N_48161);
xnor UO_2174 (O_2174,N_48813,N_48705);
and UO_2175 (O_2175,N_49506,N_48371);
or UO_2176 (O_2176,N_49323,N_48354);
nand UO_2177 (O_2177,N_49634,N_49110);
nand UO_2178 (O_2178,N_48934,N_48377);
and UO_2179 (O_2179,N_48101,N_49736);
nor UO_2180 (O_2180,N_48801,N_48380);
nand UO_2181 (O_2181,N_48931,N_48268);
and UO_2182 (O_2182,N_48773,N_48458);
or UO_2183 (O_2183,N_49024,N_49771);
nand UO_2184 (O_2184,N_49369,N_48088);
xor UO_2185 (O_2185,N_48479,N_48973);
xnor UO_2186 (O_2186,N_48399,N_48969);
nor UO_2187 (O_2187,N_48159,N_48255);
xor UO_2188 (O_2188,N_48902,N_48272);
xor UO_2189 (O_2189,N_48249,N_48690);
nor UO_2190 (O_2190,N_49077,N_49399);
or UO_2191 (O_2191,N_48553,N_49760);
and UO_2192 (O_2192,N_49513,N_48700);
and UO_2193 (O_2193,N_48420,N_49805);
and UO_2194 (O_2194,N_49174,N_49579);
and UO_2195 (O_2195,N_48409,N_49499);
xor UO_2196 (O_2196,N_49671,N_49571);
nor UO_2197 (O_2197,N_48753,N_49569);
and UO_2198 (O_2198,N_49163,N_49384);
or UO_2199 (O_2199,N_48850,N_49268);
xnor UO_2200 (O_2200,N_49178,N_49239);
nand UO_2201 (O_2201,N_49473,N_48461);
and UO_2202 (O_2202,N_48515,N_48119);
and UO_2203 (O_2203,N_49151,N_49076);
and UO_2204 (O_2204,N_48412,N_48871);
and UO_2205 (O_2205,N_49060,N_48704);
xnor UO_2206 (O_2206,N_48082,N_48284);
or UO_2207 (O_2207,N_48034,N_48301);
nor UO_2208 (O_2208,N_49718,N_49618);
xnor UO_2209 (O_2209,N_49182,N_48497);
and UO_2210 (O_2210,N_49697,N_48777);
nand UO_2211 (O_2211,N_49888,N_48062);
xor UO_2212 (O_2212,N_48215,N_49073);
and UO_2213 (O_2213,N_48087,N_48185);
nand UO_2214 (O_2214,N_48401,N_48547);
and UO_2215 (O_2215,N_48186,N_49821);
xnor UO_2216 (O_2216,N_49706,N_48986);
nand UO_2217 (O_2217,N_49947,N_49827);
xor UO_2218 (O_2218,N_48361,N_49457);
and UO_2219 (O_2219,N_49703,N_49616);
nand UO_2220 (O_2220,N_49465,N_48677);
and UO_2221 (O_2221,N_49493,N_49424);
xor UO_2222 (O_2222,N_48303,N_48633);
xnor UO_2223 (O_2223,N_49549,N_48061);
nand UO_2224 (O_2224,N_49193,N_48137);
nor UO_2225 (O_2225,N_49291,N_48003);
or UO_2226 (O_2226,N_49961,N_48979);
nand UO_2227 (O_2227,N_48963,N_49050);
nor UO_2228 (O_2228,N_49404,N_49531);
or UO_2229 (O_2229,N_49311,N_49490);
nor UO_2230 (O_2230,N_48721,N_49361);
and UO_2231 (O_2231,N_48572,N_49677);
or UO_2232 (O_2232,N_48744,N_49172);
and UO_2233 (O_2233,N_49664,N_49313);
nor UO_2234 (O_2234,N_48495,N_48464);
or UO_2235 (O_2235,N_48024,N_49280);
nor UO_2236 (O_2236,N_49213,N_49537);
xor UO_2237 (O_2237,N_48178,N_49044);
or UO_2238 (O_2238,N_48085,N_48177);
nand UO_2239 (O_2239,N_48672,N_49500);
or UO_2240 (O_2240,N_48219,N_49481);
nand UO_2241 (O_2241,N_48784,N_48386);
nand UO_2242 (O_2242,N_48728,N_48629);
or UO_2243 (O_2243,N_48936,N_49590);
nor UO_2244 (O_2244,N_48180,N_49733);
and UO_2245 (O_2245,N_48799,N_48241);
nor UO_2246 (O_2246,N_49932,N_48729);
or UO_2247 (O_2247,N_49884,N_49303);
nand UO_2248 (O_2248,N_49908,N_49796);
or UO_2249 (O_2249,N_49248,N_48102);
or UO_2250 (O_2250,N_48929,N_48508);
or UO_2251 (O_2251,N_49205,N_48438);
xor UO_2252 (O_2252,N_49284,N_49391);
xor UO_2253 (O_2253,N_49247,N_48814);
xnor UO_2254 (O_2254,N_49802,N_49120);
nor UO_2255 (O_2255,N_49036,N_48312);
and UO_2256 (O_2256,N_49992,N_49973);
and UO_2257 (O_2257,N_48170,N_49709);
xnor UO_2258 (O_2258,N_48785,N_49838);
nor UO_2259 (O_2259,N_48111,N_48807);
or UO_2260 (O_2260,N_48636,N_48685);
nor UO_2261 (O_2261,N_48213,N_48501);
xnor UO_2262 (O_2262,N_49692,N_48342);
nand UO_2263 (O_2263,N_48381,N_48545);
and UO_2264 (O_2264,N_49662,N_49845);
nand UO_2265 (O_2265,N_48817,N_48606);
nor UO_2266 (O_2266,N_49211,N_48084);
nor UO_2267 (O_2267,N_48771,N_48555);
or UO_2268 (O_2268,N_49334,N_49863);
or UO_2269 (O_2269,N_48099,N_48140);
and UO_2270 (O_2270,N_48985,N_49495);
and UO_2271 (O_2271,N_49559,N_48679);
and UO_2272 (O_2272,N_48777,N_48677);
nor UO_2273 (O_2273,N_49246,N_49977);
nand UO_2274 (O_2274,N_49914,N_49913);
and UO_2275 (O_2275,N_48241,N_48607);
or UO_2276 (O_2276,N_48051,N_48419);
nand UO_2277 (O_2277,N_48954,N_49577);
nand UO_2278 (O_2278,N_48094,N_48372);
nor UO_2279 (O_2279,N_48053,N_49778);
and UO_2280 (O_2280,N_49803,N_48974);
nand UO_2281 (O_2281,N_49229,N_48783);
xnor UO_2282 (O_2282,N_49288,N_49306);
nand UO_2283 (O_2283,N_48831,N_49957);
nand UO_2284 (O_2284,N_49755,N_48782);
nand UO_2285 (O_2285,N_49185,N_49394);
or UO_2286 (O_2286,N_48206,N_49855);
and UO_2287 (O_2287,N_48838,N_48554);
nand UO_2288 (O_2288,N_49436,N_48428);
xnor UO_2289 (O_2289,N_48270,N_49082);
xnor UO_2290 (O_2290,N_49166,N_49696);
nor UO_2291 (O_2291,N_49263,N_48362);
xor UO_2292 (O_2292,N_48539,N_49485);
and UO_2293 (O_2293,N_49062,N_49733);
nand UO_2294 (O_2294,N_49516,N_48509);
xnor UO_2295 (O_2295,N_48311,N_49520);
nor UO_2296 (O_2296,N_48661,N_48547);
or UO_2297 (O_2297,N_49328,N_48023);
or UO_2298 (O_2298,N_48597,N_48481);
nor UO_2299 (O_2299,N_49489,N_49605);
or UO_2300 (O_2300,N_49344,N_49282);
xnor UO_2301 (O_2301,N_49239,N_48192);
xor UO_2302 (O_2302,N_48419,N_49344);
nor UO_2303 (O_2303,N_49305,N_48777);
nand UO_2304 (O_2304,N_48124,N_49838);
xor UO_2305 (O_2305,N_49507,N_48510);
nand UO_2306 (O_2306,N_49426,N_48763);
xor UO_2307 (O_2307,N_48415,N_48336);
xor UO_2308 (O_2308,N_49924,N_48491);
and UO_2309 (O_2309,N_48211,N_49510);
or UO_2310 (O_2310,N_49466,N_48762);
and UO_2311 (O_2311,N_49410,N_48074);
or UO_2312 (O_2312,N_48119,N_49794);
or UO_2313 (O_2313,N_48736,N_48727);
xor UO_2314 (O_2314,N_48282,N_48383);
or UO_2315 (O_2315,N_48322,N_48775);
nand UO_2316 (O_2316,N_48687,N_49899);
xor UO_2317 (O_2317,N_48092,N_49024);
xnor UO_2318 (O_2318,N_48705,N_48629);
xnor UO_2319 (O_2319,N_49934,N_48987);
xnor UO_2320 (O_2320,N_48869,N_49886);
nand UO_2321 (O_2321,N_48391,N_48146);
xnor UO_2322 (O_2322,N_48868,N_48333);
xor UO_2323 (O_2323,N_49976,N_49634);
nor UO_2324 (O_2324,N_49548,N_49911);
or UO_2325 (O_2325,N_49680,N_49593);
nor UO_2326 (O_2326,N_49847,N_49026);
and UO_2327 (O_2327,N_48160,N_49233);
xnor UO_2328 (O_2328,N_48966,N_48093);
nor UO_2329 (O_2329,N_49904,N_49308);
nand UO_2330 (O_2330,N_49642,N_49572);
xor UO_2331 (O_2331,N_49070,N_48008);
or UO_2332 (O_2332,N_48087,N_48045);
nand UO_2333 (O_2333,N_49264,N_48989);
nand UO_2334 (O_2334,N_48646,N_48005);
or UO_2335 (O_2335,N_49121,N_48228);
nand UO_2336 (O_2336,N_48333,N_49717);
xor UO_2337 (O_2337,N_49561,N_48544);
xor UO_2338 (O_2338,N_49301,N_49190);
nor UO_2339 (O_2339,N_49501,N_48353);
nand UO_2340 (O_2340,N_49026,N_49096);
xor UO_2341 (O_2341,N_48653,N_49230);
nor UO_2342 (O_2342,N_49376,N_48226);
or UO_2343 (O_2343,N_48410,N_49924);
nor UO_2344 (O_2344,N_49539,N_48376);
xor UO_2345 (O_2345,N_48294,N_48560);
or UO_2346 (O_2346,N_48429,N_49810);
xor UO_2347 (O_2347,N_49619,N_48597);
xor UO_2348 (O_2348,N_48188,N_48812);
and UO_2349 (O_2349,N_48232,N_48356);
or UO_2350 (O_2350,N_49213,N_49739);
and UO_2351 (O_2351,N_49579,N_49260);
nor UO_2352 (O_2352,N_48476,N_49846);
or UO_2353 (O_2353,N_49336,N_48660);
nand UO_2354 (O_2354,N_48461,N_48707);
nor UO_2355 (O_2355,N_49383,N_49308);
nand UO_2356 (O_2356,N_49222,N_48208);
nand UO_2357 (O_2357,N_48554,N_48663);
xnor UO_2358 (O_2358,N_48580,N_48102);
or UO_2359 (O_2359,N_49444,N_48099);
nand UO_2360 (O_2360,N_48796,N_48800);
and UO_2361 (O_2361,N_49858,N_48936);
nor UO_2362 (O_2362,N_49044,N_49484);
xnor UO_2363 (O_2363,N_49160,N_48473);
and UO_2364 (O_2364,N_49741,N_49150);
nor UO_2365 (O_2365,N_49199,N_49915);
or UO_2366 (O_2366,N_49382,N_49078);
nor UO_2367 (O_2367,N_49025,N_48449);
nor UO_2368 (O_2368,N_48919,N_49641);
and UO_2369 (O_2369,N_48893,N_48440);
and UO_2370 (O_2370,N_49817,N_48850);
nor UO_2371 (O_2371,N_49382,N_49467);
or UO_2372 (O_2372,N_49664,N_48981);
nor UO_2373 (O_2373,N_48448,N_49067);
nand UO_2374 (O_2374,N_49602,N_48540);
xnor UO_2375 (O_2375,N_48769,N_49442);
or UO_2376 (O_2376,N_48999,N_49814);
nor UO_2377 (O_2377,N_48666,N_49137);
or UO_2378 (O_2378,N_49523,N_48909);
or UO_2379 (O_2379,N_49691,N_48127);
nor UO_2380 (O_2380,N_49855,N_49203);
nand UO_2381 (O_2381,N_49075,N_49743);
nor UO_2382 (O_2382,N_49039,N_48618);
nor UO_2383 (O_2383,N_48123,N_49849);
or UO_2384 (O_2384,N_48289,N_48079);
or UO_2385 (O_2385,N_49150,N_48124);
xor UO_2386 (O_2386,N_49713,N_49192);
xor UO_2387 (O_2387,N_48997,N_49047);
xor UO_2388 (O_2388,N_48542,N_48592);
xnor UO_2389 (O_2389,N_48563,N_49391);
nor UO_2390 (O_2390,N_48082,N_48854);
nand UO_2391 (O_2391,N_49472,N_49483);
or UO_2392 (O_2392,N_48479,N_49001);
nand UO_2393 (O_2393,N_49475,N_48412);
xor UO_2394 (O_2394,N_49436,N_48967);
nor UO_2395 (O_2395,N_49558,N_48560);
and UO_2396 (O_2396,N_48208,N_48291);
nor UO_2397 (O_2397,N_49837,N_48093);
nor UO_2398 (O_2398,N_49225,N_48568);
nand UO_2399 (O_2399,N_49996,N_49286);
and UO_2400 (O_2400,N_48598,N_48679);
or UO_2401 (O_2401,N_49735,N_48641);
xnor UO_2402 (O_2402,N_49780,N_48310);
and UO_2403 (O_2403,N_48340,N_48716);
xor UO_2404 (O_2404,N_49772,N_49416);
xor UO_2405 (O_2405,N_48354,N_49504);
and UO_2406 (O_2406,N_48118,N_48202);
or UO_2407 (O_2407,N_48425,N_48214);
xor UO_2408 (O_2408,N_49265,N_49592);
nor UO_2409 (O_2409,N_48629,N_48477);
xor UO_2410 (O_2410,N_49311,N_48896);
xnor UO_2411 (O_2411,N_49213,N_49517);
nand UO_2412 (O_2412,N_48563,N_48072);
or UO_2413 (O_2413,N_48505,N_48512);
xnor UO_2414 (O_2414,N_49709,N_49094);
xor UO_2415 (O_2415,N_48215,N_49479);
or UO_2416 (O_2416,N_49036,N_48747);
nand UO_2417 (O_2417,N_49888,N_49875);
xnor UO_2418 (O_2418,N_49046,N_49756);
nand UO_2419 (O_2419,N_48055,N_48251);
nand UO_2420 (O_2420,N_48614,N_49692);
and UO_2421 (O_2421,N_49258,N_48820);
and UO_2422 (O_2422,N_49125,N_49771);
nand UO_2423 (O_2423,N_48219,N_48079);
xnor UO_2424 (O_2424,N_49842,N_49574);
and UO_2425 (O_2425,N_49594,N_48383);
nor UO_2426 (O_2426,N_49763,N_49553);
xor UO_2427 (O_2427,N_49755,N_49726);
nor UO_2428 (O_2428,N_48792,N_48832);
nor UO_2429 (O_2429,N_49077,N_49193);
or UO_2430 (O_2430,N_49736,N_48811);
nor UO_2431 (O_2431,N_49831,N_48665);
nand UO_2432 (O_2432,N_48157,N_49990);
and UO_2433 (O_2433,N_49437,N_48942);
or UO_2434 (O_2434,N_48572,N_48409);
nand UO_2435 (O_2435,N_49667,N_49995);
nand UO_2436 (O_2436,N_49375,N_49752);
nand UO_2437 (O_2437,N_49843,N_49908);
nor UO_2438 (O_2438,N_48723,N_49735);
and UO_2439 (O_2439,N_48266,N_48900);
nor UO_2440 (O_2440,N_49639,N_48859);
nor UO_2441 (O_2441,N_48596,N_48969);
nand UO_2442 (O_2442,N_49402,N_49496);
or UO_2443 (O_2443,N_49072,N_49187);
nand UO_2444 (O_2444,N_49260,N_49738);
nand UO_2445 (O_2445,N_48764,N_48171);
nor UO_2446 (O_2446,N_49677,N_48127);
xnor UO_2447 (O_2447,N_48047,N_49286);
xor UO_2448 (O_2448,N_49657,N_48902);
and UO_2449 (O_2449,N_48035,N_48602);
nand UO_2450 (O_2450,N_49797,N_48997);
nand UO_2451 (O_2451,N_49242,N_49357);
nand UO_2452 (O_2452,N_49633,N_48307);
and UO_2453 (O_2453,N_48989,N_48002);
and UO_2454 (O_2454,N_49838,N_48830);
xnor UO_2455 (O_2455,N_48132,N_49905);
nor UO_2456 (O_2456,N_48108,N_49415);
or UO_2457 (O_2457,N_48881,N_48296);
xor UO_2458 (O_2458,N_48805,N_48840);
nor UO_2459 (O_2459,N_49307,N_48442);
xor UO_2460 (O_2460,N_49354,N_49927);
or UO_2461 (O_2461,N_49696,N_48694);
nor UO_2462 (O_2462,N_49987,N_49296);
and UO_2463 (O_2463,N_48919,N_49770);
and UO_2464 (O_2464,N_48000,N_48621);
nor UO_2465 (O_2465,N_48095,N_49626);
or UO_2466 (O_2466,N_49652,N_49160);
or UO_2467 (O_2467,N_49310,N_49610);
xnor UO_2468 (O_2468,N_48193,N_49827);
nor UO_2469 (O_2469,N_48369,N_48189);
or UO_2470 (O_2470,N_48233,N_48509);
or UO_2471 (O_2471,N_48900,N_49433);
nand UO_2472 (O_2472,N_49309,N_48110);
and UO_2473 (O_2473,N_49874,N_48400);
or UO_2474 (O_2474,N_49611,N_49586);
xor UO_2475 (O_2475,N_48304,N_48500);
nand UO_2476 (O_2476,N_48223,N_49385);
nor UO_2477 (O_2477,N_48760,N_48304);
nor UO_2478 (O_2478,N_48825,N_48746);
nand UO_2479 (O_2479,N_48665,N_48081);
or UO_2480 (O_2480,N_48774,N_49371);
and UO_2481 (O_2481,N_48324,N_49442);
or UO_2482 (O_2482,N_49936,N_48069);
nand UO_2483 (O_2483,N_49565,N_49566);
or UO_2484 (O_2484,N_48080,N_49702);
or UO_2485 (O_2485,N_49623,N_49045);
or UO_2486 (O_2486,N_48419,N_49155);
xor UO_2487 (O_2487,N_49489,N_48369);
nand UO_2488 (O_2488,N_48048,N_48429);
nor UO_2489 (O_2489,N_49448,N_48232);
xnor UO_2490 (O_2490,N_49246,N_48802);
and UO_2491 (O_2491,N_48235,N_48516);
and UO_2492 (O_2492,N_49904,N_49386);
or UO_2493 (O_2493,N_48099,N_49639);
nand UO_2494 (O_2494,N_48979,N_48444);
xnor UO_2495 (O_2495,N_48763,N_49012);
nor UO_2496 (O_2496,N_48686,N_49638);
and UO_2497 (O_2497,N_48028,N_49720);
and UO_2498 (O_2498,N_49966,N_49355);
xor UO_2499 (O_2499,N_49648,N_48873);
nor UO_2500 (O_2500,N_49196,N_48976);
or UO_2501 (O_2501,N_49606,N_49295);
xnor UO_2502 (O_2502,N_48803,N_49562);
nand UO_2503 (O_2503,N_48329,N_48226);
and UO_2504 (O_2504,N_49418,N_49042);
or UO_2505 (O_2505,N_49403,N_49011);
or UO_2506 (O_2506,N_48630,N_48173);
xor UO_2507 (O_2507,N_48410,N_48569);
nand UO_2508 (O_2508,N_49973,N_48600);
and UO_2509 (O_2509,N_48259,N_49382);
nor UO_2510 (O_2510,N_48287,N_49221);
and UO_2511 (O_2511,N_49522,N_48501);
and UO_2512 (O_2512,N_48648,N_49384);
nor UO_2513 (O_2513,N_49950,N_48281);
xor UO_2514 (O_2514,N_49472,N_48384);
xnor UO_2515 (O_2515,N_49138,N_48995);
xnor UO_2516 (O_2516,N_48585,N_49707);
xor UO_2517 (O_2517,N_49747,N_48899);
nor UO_2518 (O_2518,N_48917,N_48243);
nor UO_2519 (O_2519,N_48034,N_48111);
nor UO_2520 (O_2520,N_49082,N_48289);
nand UO_2521 (O_2521,N_48464,N_49907);
xor UO_2522 (O_2522,N_48032,N_49324);
xnor UO_2523 (O_2523,N_48335,N_48980);
xnor UO_2524 (O_2524,N_49807,N_48042);
nand UO_2525 (O_2525,N_48620,N_49979);
nor UO_2526 (O_2526,N_48442,N_48537);
or UO_2527 (O_2527,N_48545,N_48852);
or UO_2528 (O_2528,N_49858,N_49205);
nand UO_2529 (O_2529,N_48710,N_48973);
nand UO_2530 (O_2530,N_48786,N_49817);
and UO_2531 (O_2531,N_49289,N_49161);
or UO_2532 (O_2532,N_49645,N_49130);
or UO_2533 (O_2533,N_49076,N_48313);
or UO_2534 (O_2534,N_48268,N_48857);
xnor UO_2535 (O_2535,N_49851,N_48459);
xor UO_2536 (O_2536,N_49699,N_49845);
or UO_2537 (O_2537,N_48510,N_48465);
nor UO_2538 (O_2538,N_48227,N_48741);
nand UO_2539 (O_2539,N_48228,N_49538);
xnor UO_2540 (O_2540,N_49855,N_49029);
and UO_2541 (O_2541,N_48296,N_48914);
nor UO_2542 (O_2542,N_49853,N_48427);
and UO_2543 (O_2543,N_49681,N_49397);
nor UO_2544 (O_2544,N_49010,N_48029);
xnor UO_2545 (O_2545,N_49963,N_48898);
and UO_2546 (O_2546,N_49598,N_49316);
nor UO_2547 (O_2547,N_49691,N_48417);
nor UO_2548 (O_2548,N_48052,N_49440);
and UO_2549 (O_2549,N_48855,N_48200);
nor UO_2550 (O_2550,N_48973,N_48430);
xor UO_2551 (O_2551,N_49584,N_49018);
and UO_2552 (O_2552,N_49593,N_48518);
or UO_2553 (O_2553,N_49831,N_48677);
and UO_2554 (O_2554,N_48242,N_49294);
or UO_2555 (O_2555,N_49432,N_48320);
xnor UO_2556 (O_2556,N_49180,N_49726);
or UO_2557 (O_2557,N_48801,N_48051);
nand UO_2558 (O_2558,N_48927,N_48294);
and UO_2559 (O_2559,N_49325,N_48273);
and UO_2560 (O_2560,N_48888,N_48740);
or UO_2561 (O_2561,N_49805,N_49252);
or UO_2562 (O_2562,N_49470,N_49923);
xor UO_2563 (O_2563,N_49851,N_49216);
nand UO_2564 (O_2564,N_49774,N_48267);
and UO_2565 (O_2565,N_49825,N_49205);
or UO_2566 (O_2566,N_49623,N_48862);
or UO_2567 (O_2567,N_49359,N_48726);
nand UO_2568 (O_2568,N_48434,N_48981);
nand UO_2569 (O_2569,N_49167,N_49196);
or UO_2570 (O_2570,N_48238,N_48737);
or UO_2571 (O_2571,N_48039,N_48863);
and UO_2572 (O_2572,N_48363,N_49193);
nand UO_2573 (O_2573,N_48461,N_48751);
nor UO_2574 (O_2574,N_48189,N_48030);
xnor UO_2575 (O_2575,N_49223,N_48468);
and UO_2576 (O_2576,N_48257,N_49170);
nand UO_2577 (O_2577,N_48612,N_48025);
nor UO_2578 (O_2578,N_49200,N_49636);
xor UO_2579 (O_2579,N_49390,N_49877);
nor UO_2580 (O_2580,N_49317,N_48359);
and UO_2581 (O_2581,N_48244,N_48749);
xor UO_2582 (O_2582,N_49437,N_48477);
xnor UO_2583 (O_2583,N_48607,N_49813);
xor UO_2584 (O_2584,N_48541,N_49906);
or UO_2585 (O_2585,N_48679,N_48985);
nor UO_2586 (O_2586,N_48995,N_49796);
or UO_2587 (O_2587,N_48489,N_48934);
and UO_2588 (O_2588,N_48262,N_48523);
nor UO_2589 (O_2589,N_49527,N_49898);
and UO_2590 (O_2590,N_48151,N_48865);
nor UO_2591 (O_2591,N_48277,N_48239);
xor UO_2592 (O_2592,N_49199,N_48591);
xnor UO_2593 (O_2593,N_49817,N_49138);
nor UO_2594 (O_2594,N_49140,N_48831);
or UO_2595 (O_2595,N_49806,N_49702);
nand UO_2596 (O_2596,N_49553,N_48137);
xor UO_2597 (O_2597,N_48501,N_49436);
nand UO_2598 (O_2598,N_48455,N_48053);
xnor UO_2599 (O_2599,N_49015,N_48534);
nor UO_2600 (O_2600,N_49971,N_48928);
xor UO_2601 (O_2601,N_48297,N_49895);
or UO_2602 (O_2602,N_49198,N_49570);
nor UO_2603 (O_2603,N_49591,N_49162);
nor UO_2604 (O_2604,N_49730,N_49648);
xnor UO_2605 (O_2605,N_49480,N_49489);
xnor UO_2606 (O_2606,N_49323,N_49637);
xnor UO_2607 (O_2607,N_49474,N_49119);
xnor UO_2608 (O_2608,N_49402,N_48363);
xor UO_2609 (O_2609,N_48806,N_48882);
xnor UO_2610 (O_2610,N_48617,N_48494);
xnor UO_2611 (O_2611,N_49279,N_48884);
or UO_2612 (O_2612,N_48633,N_49509);
nor UO_2613 (O_2613,N_48054,N_49709);
nand UO_2614 (O_2614,N_49101,N_48978);
nand UO_2615 (O_2615,N_49509,N_48169);
nor UO_2616 (O_2616,N_48438,N_48412);
nor UO_2617 (O_2617,N_49812,N_48985);
nor UO_2618 (O_2618,N_49960,N_48405);
xor UO_2619 (O_2619,N_49169,N_48226);
xnor UO_2620 (O_2620,N_48236,N_48162);
xnor UO_2621 (O_2621,N_49126,N_48203);
and UO_2622 (O_2622,N_48647,N_49002);
xnor UO_2623 (O_2623,N_48858,N_48047);
nand UO_2624 (O_2624,N_49094,N_49015);
nand UO_2625 (O_2625,N_48296,N_49309);
xor UO_2626 (O_2626,N_49366,N_48516);
and UO_2627 (O_2627,N_48971,N_48499);
nor UO_2628 (O_2628,N_49964,N_48256);
nand UO_2629 (O_2629,N_49515,N_49700);
nand UO_2630 (O_2630,N_49973,N_49635);
nor UO_2631 (O_2631,N_48848,N_48382);
nand UO_2632 (O_2632,N_48386,N_48337);
or UO_2633 (O_2633,N_49871,N_48591);
xnor UO_2634 (O_2634,N_49098,N_49596);
nor UO_2635 (O_2635,N_48875,N_48783);
nand UO_2636 (O_2636,N_49743,N_49855);
xnor UO_2637 (O_2637,N_48955,N_49492);
and UO_2638 (O_2638,N_49723,N_49067);
or UO_2639 (O_2639,N_49500,N_49046);
nor UO_2640 (O_2640,N_49831,N_49528);
nor UO_2641 (O_2641,N_48340,N_48494);
xor UO_2642 (O_2642,N_49125,N_48566);
nand UO_2643 (O_2643,N_48684,N_48021);
nor UO_2644 (O_2644,N_49379,N_49932);
nand UO_2645 (O_2645,N_48377,N_49147);
and UO_2646 (O_2646,N_48913,N_48449);
or UO_2647 (O_2647,N_49641,N_48874);
and UO_2648 (O_2648,N_48019,N_49523);
nand UO_2649 (O_2649,N_49254,N_48774);
and UO_2650 (O_2650,N_48457,N_48397);
and UO_2651 (O_2651,N_48394,N_48349);
or UO_2652 (O_2652,N_49611,N_48882);
or UO_2653 (O_2653,N_48605,N_48145);
nand UO_2654 (O_2654,N_49907,N_48350);
nor UO_2655 (O_2655,N_49956,N_48980);
nor UO_2656 (O_2656,N_48670,N_48731);
and UO_2657 (O_2657,N_48667,N_48350);
and UO_2658 (O_2658,N_48856,N_48094);
and UO_2659 (O_2659,N_49417,N_48655);
or UO_2660 (O_2660,N_48913,N_48460);
nor UO_2661 (O_2661,N_48148,N_48020);
or UO_2662 (O_2662,N_48354,N_49617);
or UO_2663 (O_2663,N_48054,N_48283);
nand UO_2664 (O_2664,N_49616,N_49615);
nor UO_2665 (O_2665,N_48479,N_48037);
nand UO_2666 (O_2666,N_48372,N_49245);
nand UO_2667 (O_2667,N_49498,N_49193);
or UO_2668 (O_2668,N_48279,N_48159);
nor UO_2669 (O_2669,N_49868,N_48409);
nor UO_2670 (O_2670,N_49648,N_49303);
nand UO_2671 (O_2671,N_48277,N_49071);
or UO_2672 (O_2672,N_48105,N_48104);
or UO_2673 (O_2673,N_48927,N_48250);
or UO_2674 (O_2674,N_49720,N_48031);
or UO_2675 (O_2675,N_48051,N_48525);
nor UO_2676 (O_2676,N_48120,N_48778);
or UO_2677 (O_2677,N_48000,N_48925);
xnor UO_2678 (O_2678,N_48365,N_48904);
and UO_2679 (O_2679,N_48546,N_49163);
nand UO_2680 (O_2680,N_49859,N_48975);
nand UO_2681 (O_2681,N_49148,N_48275);
xor UO_2682 (O_2682,N_49785,N_49805);
nand UO_2683 (O_2683,N_48970,N_49266);
nor UO_2684 (O_2684,N_48978,N_49727);
nand UO_2685 (O_2685,N_48936,N_48786);
nor UO_2686 (O_2686,N_49584,N_49821);
and UO_2687 (O_2687,N_49812,N_49829);
xnor UO_2688 (O_2688,N_48535,N_49715);
nor UO_2689 (O_2689,N_49219,N_49628);
or UO_2690 (O_2690,N_49390,N_48672);
and UO_2691 (O_2691,N_48714,N_49159);
or UO_2692 (O_2692,N_49902,N_48964);
nor UO_2693 (O_2693,N_49521,N_48486);
and UO_2694 (O_2694,N_48153,N_48439);
and UO_2695 (O_2695,N_49433,N_49856);
nand UO_2696 (O_2696,N_48887,N_49468);
xnor UO_2697 (O_2697,N_49801,N_49785);
nand UO_2698 (O_2698,N_48571,N_49124);
or UO_2699 (O_2699,N_49253,N_49098);
nor UO_2700 (O_2700,N_48571,N_49519);
or UO_2701 (O_2701,N_48934,N_49245);
xor UO_2702 (O_2702,N_48322,N_48758);
and UO_2703 (O_2703,N_49897,N_48491);
xnor UO_2704 (O_2704,N_48283,N_49882);
xnor UO_2705 (O_2705,N_49525,N_49868);
nor UO_2706 (O_2706,N_49231,N_49851);
nor UO_2707 (O_2707,N_49413,N_48594);
nor UO_2708 (O_2708,N_48379,N_49586);
or UO_2709 (O_2709,N_48925,N_48398);
and UO_2710 (O_2710,N_48045,N_49338);
or UO_2711 (O_2711,N_48802,N_48066);
nor UO_2712 (O_2712,N_49941,N_48305);
nand UO_2713 (O_2713,N_48794,N_48463);
or UO_2714 (O_2714,N_49040,N_49992);
and UO_2715 (O_2715,N_49585,N_48397);
or UO_2716 (O_2716,N_49076,N_48182);
xnor UO_2717 (O_2717,N_48659,N_48466);
xnor UO_2718 (O_2718,N_48334,N_48508);
nor UO_2719 (O_2719,N_49499,N_48879);
or UO_2720 (O_2720,N_49742,N_49545);
nor UO_2721 (O_2721,N_49748,N_49151);
or UO_2722 (O_2722,N_49584,N_49788);
and UO_2723 (O_2723,N_48475,N_49379);
and UO_2724 (O_2724,N_49961,N_49916);
or UO_2725 (O_2725,N_48172,N_49730);
and UO_2726 (O_2726,N_49749,N_48975);
or UO_2727 (O_2727,N_49090,N_48419);
nand UO_2728 (O_2728,N_48016,N_49160);
xor UO_2729 (O_2729,N_49569,N_49463);
nand UO_2730 (O_2730,N_48025,N_49071);
xor UO_2731 (O_2731,N_49285,N_48893);
nor UO_2732 (O_2732,N_49640,N_48015);
or UO_2733 (O_2733,N_49251,N_48703);
and UO_2734 (O_2734,N_49915,N_48488);
or UO_2735 (O_2735,N_48390,N_49512);
xor UO_2736 (O_2736,N_49852,N_49464);
nand UO_2737 (O_2737,N_49274,N_49013);
nor UO_2738 (O_2738,N_48614,N_48481);
nand UO_2739 (O_2739,N_48483,N_48360);
nand UO_2740 (O_2740,N_49541,N_49871);
xor UO_2741 (O_2741,N_48867,N_49644);
xor UO_2742 (O_2742,N_48603,N_48059);
xor UO_2743 (O_2743,N_49211,N_49962);
or UO_2744 (O_2744,N_48992,N_49934);
nand UO_2745 (O_2745,N_48852,N_49402);
nand UO_2746 (O_2746,N_48363,N_48873);
or UO_2747 (O_2747,N_49721,N_48203);
nand UO_2748 (O_2748,N_49214,N_48968);
nand UO_2749 (O_2749,N_48292,N_48268);
and UO_2750 (O_2750,N_48685,N_49717);
xnor UO_2751 (O_2751,N_49204,N_49066);
nor UO_2752 (O_2752,N_48749,N_49773);
nor UO_2753 (O_2753,N_48852,N_48144);
xnor UO_2754 (O_2754,N_48803,N_49505);
xnor UO_2755 (O_2755,N_49694,N_48754);
and UO_2756 (O_2756,N_49159,N_49648);
xor UO_2757 (O_2757,N_49325,N_48269);
xor UO_2758 (O_2758,N_48515,N_49944);
nand UO_2759 (O_2759,N_49351,N_49228);
or UO_2760 (O_2760,N_48934,N_49208);
or UO_2761 (O_2761,N_49081,N_49112);
nor UO_2762 (O_2762,N_48113,N_48187);
nor UO_2763 (O_2763,N_49330,N_49861);
and UO_2764 (O_2764,N_48578,N_48072);
nor UO_2765 (O_2765,N_48229,N_49258);
and UO_2766 (O_2766,N_49225,N_49408);
xnor UO_2767 (O_2767,N_48383,N_48618);
nor UO_2768 (O_2768,N_48444,N_49592);
nor UO_2769 (O_2769,N_48610,N_49435);
nor UO_2770 (O_2770,N_48440,N_49213);
xnor UO_2771 (O_2771,N_49201,N_48865);
nand UO_2772 (O_2772,N_49027,N_49430);
xor UO_2773 (O_2773,N_48045,N_49417);
and UO_2774 (O_2774,N_48183,N_49613);
and UO_2775 (O_2775,N_48224,N_49167);
nor UO_2776 (O_2776,N_49757,N_48128);
nor UO_2777 (O_2777,N_48047,N_49811);
nor UO_2778 (O_2778,N_48017,N_49555);
nand UO_2779 (O_2779,N_49844,N_49705);
or UO_2780 (O_2780,N_49588,N_48713);
xor UO_2781 (O_2781,N_49446,N_49703);
nand UO_2782 (O_2782,N_48372,N_48340);
nor UO_2783 (O_2783,N_49605,N_48199);
nor UO_2784 (O_2784,N_49401,N_48231);
and UO_2785 (O_2785,N_48670,N_48576);
and UO_2786 (O_2786,N_49920,N_49535);
and UO_2787 (O_2787,N_48666,N_49495);
and UO_2788 (O_2788,N_49789,N_48830);
xor UO_2789 (O_2789,N_49188,N_49233);
or UO_2790 (O_2790,N_49618,N_48280);
nand UO_2791 (O_2791,N_48252,N_48614);
or UO_2792 (O_2792,N_48984,N_48823);
xor UO_2793 (O_2793,N_49231,N_48895);
and UO_2794 (O_2794,N_48684,N_48932);
nand UO_2795 (O_2795,N_49088,N_49943);
nand UO_2796 (O_2796,N_49966,N_48480);
nand UO_2797 (O_2797,N_49217,N_49579);
xnor UO_2798 (O_2798,N_48770,N_48926);
or UO_2799 (O_2799,N_49065,N_49088);
nand UO_2800 (O_2800,N_49774,N_48135);
or UO_2801 (O_2801,N_49320,N_48036);
and UO_2802 (O_2802,N_48364,N_49737);
and UO_2803 (O_2803,N_49777,N_48111);
xnor UO_2804 (O_2804,N_48153,N_48688);
and UO_2805 (O_2805,N_48730,N_48549);
nor UO_2806 (O_2806,N_49052,N_49108);
and UO_2807 (O_2807,N_49515,N_48920);
and UO_2808 (O_2808,N_49006,N_49153);
xor UO_2809 (O_2809,N_49751,N_48679);
xnor UO_2810 (O_2810,N_49861,N_48859);
nor UO_2811 (O_2811,N_49514,N_48330);
xnor UO_2812 (O_2812,N_48233,N_48248);
and UO_2813 (O_2813,N_49810,N_48586);
or UO_2814 (O_2814,N_48584,N_49260);
or UO_2815 (O_2815,N_49188,N_48951);
or UO_2816 (O_2816,N_49640,N_48161);
nor UO_2817 (O_2817,N_49301,N_49631);
nand UO_2818 (O_2818,N_48798,N_49067);
nand UO_2819 (O_2819,N_49967,N_48654);
nor UO_2820 (O_2820,N_49675,N_48029);
nor UO_2821 (O_2821,N_49320,N_49078);
and UO_2822 (O_2822,N_49429,N_49558);
xor UO_2823 (O_2823,N_48964,N_49947);
xnor UO_2824 (O_2824,N_49217,N_48191);
and UO_2825 (O_2825,N_48822,N_48492);
or UO_2826 (O_2826,N_49142,N_48460);
xor UO_2827 (O_2827,N_49369,N_48685);
xor UO_2828 (O_2828,N_49907,N_49804);
nand UO_2829 (O_2829,N_48141,N_48919);
or UO_2830 (O_2830,N_49251,N_48277);
xnor UO_2831 (O_2831,N_48731,N_48897);
xnor UO_2832 (O_2832,N_49646,N_48318);
xor UO_2833 (O_2833,N_48718,N_48225);
or UO_2834 (O_2834,N_49182,N_49149);
or UO_2835 (O_2835,N_48100,N_49150);
xnor UO_2836 (O_2836,N_48370,N_49068);
xor UO_2837 (O_2837,N_48797,N_49331);
nor UO_2838 (O_2838,N_49054,N_49411);
xor UO_2839 (O_2839,N_48767,N_49653);
nand UO_2840 (O_2840,N_49088,N_48404);
or UO_2841 (O_2841,N_48412,N_48836);
and UO_2842 (O_2842,N_49584,N_49878);
nor UO_2843 (O_2843,N_48721,N_49855);
and UO_2844 (O_2844,N_49673,N_49470);
nor UO_2845 (O_2845,N_48217,N_48417);
or UO_2846 (O_2846,N_49404,N_48176);
xor UO_2847 (O_2847,N_49389,N_49940);
xnor UO_2848 (O_2848,N_49468,N_49684);
xor UO_2849 (O_2849,N_48934,N_48727);
or UO_2850 (O_2850,N_48275,N_49225);
and UO_2851 (O_2851,N_49746,N_48558);
nand UO_2852 (O_2852,N_48468,N_49839);
or UO_2853 (O_2853,N_48590,N_48276);
nand UO_2854 (O_2854,N_48884,N_48097);
or UO_2855 (O_2855,N_49088,N_49070);
nor UO_2856 (O_2856,N_49508,N_49999);
and UO_2857 (O_2857,N_49081,N_48918);
nor UO_2858 (O_2858,N_48794,N_48598);
xnor UO_2859 (O_2859,N_49517,N_48462);
xor UO_2860 (O_2860,N_49052,N_48834);
nand UO_2861 (O_2861,N_49898,N_48134);
nor UO_2862 (O_2862,N_48305,N_48444);
nand UO_2863 (O_2863,N_48839,N_49651);
and UO_2864 (O_2864,N_48195,N_48245);
and UO_2865 (O_2865,N_49142,N_48754);
or UO_2866 (O_2866,N_49934,N_48894);
or UO_2867 (O_2867,N_49458,N_48820);
nor UO_2868 (O_2868,N_48589,N_49413);
nor UO_2869 (O_2869,N_49666,N_48290);
or UO_2870 (O_2870,N_48130,N_48570);
and UO_2871 (O_2871,N_49338,N_48195);
nor UO_2872 (O_2872,N_49075,N_48509);
nand UO_2873 (O_2873,N_48734,N_48395);
and UO_2874 (O_2874,N_48290,N_48547);
and UO_2875 (O_2875,N_49928,N_49471);
and UO_2876 (O_2876,N_49952,N_49613);
nand UO_2877 (O_2877,N_48664,N_48165);
nand UO_2878 (O_2878,N_49175,N_49782);
nor UO_2879 (O_2879,N_49889,N_49616);
xnor UO_2880 (O_2880,N_49959,N_48364);
and UO_2881 (O_2881,N_49823,N_49324);
xor UO_2882 (O_2882,N_49962,N_49977);
nor UO_2883 (O_2883,N_48159,N_48186);
nand UO_2884 (O_2884,N_48713,N_48847);
nor UO_2885 (O_2885,N_49249,N_48865);
nand UO_2886 (O_2886,N_48358,N_48962);
and UO_2887 (O_2887,N_48654,N_48558);
and UO_2888 (O_2888,N_48569,N_48458);
nor UO_2889 (O_2889,N_49128,N_48730);
and UO_2890 (O_2890,N_49648,N_49232);
nand UO_2891 (O_2891,N_48253,N_48731);
or UO_2892 (O_2892,N_49000,N_48809);
nor UO_2893 (O_2893,N_49746,N_49174);
nor UO_2894 (O_2894,N_48247,N_49548);
xor UO_2895 (O_2895,N_49782,N_48082);
or UO_2896 (O_2896,N_49698,N_48945);
nand UO_2897 (O_2897,N_49551,N_48491);
nand UO_2898 (O_2898,N_48945,N_49647);
xor UO_2899 (O_2899,N_49994,N_48284);
nor UO_2900 (O_2900,N_49530,N_49037);
nor UO_2901 (O_2901,N_48354,N_49894);
nand UO_2902 (O_2902,N_49606,N_49594);
or UO_2903 (O_2903,N_49910,N_48904);
nand UO_2904 (O_2904,N_48687,N_48743);
and UO_2905 (O_2905,N_49592,N_49789);
xnor UO_2906 (O_2906,N_49389,N_48431);
and UO_2907 (O_2907,N_48339,N_48234);
nand UO_2908 (O_2908,N_48414,N_48674);
nand UO_2909 (O_2909,N_48858,N_48987);
nor UO_2910 (O_2910,N_48268,N_48583);
nor UO_2911 (O_2911,N_48239,N_49630);
and UO_2912 (O_2912,N_48585,N_48607);
xor UO_2913 (O_2913,N_48664,N_48798);
and UO_2914 (O_2914,N_49063,N_48049);
xor UO_2915 (O_2915,N_48986,N_49146);
xor UO_2916 (O_2916,N_49264,N_48883);
and UO_2917 (O_2917,N_49738,N_48561);
or UO_2918 (O_2918,N_48754,N_48564);
and UO_2919 (O_2919,N_49657,N_49573);
xnor UO_2920 (O_2920,N_48290,N_49951);
and UO_2921 (O_2921,N_49909,N_48854);
and UO_2922 (O_2922,N_48855,N_48683);
nor UO_2923 (O_2923,N_48898,N_49116);
or UO_2924 (O_2924,N_48749,N_49794);
and UO_2925 (O_2925,N_49341,N_48676);
xor UO_2926 (O_2926,N_48240,N_48963);
or UO_2927 (O_2927,N_48396,N_48512);
and UO_2928 (O_2928,N_48342,N_48876);
xor UO_2929 (O_2929,N_48812,N_49907);
nor UO_2930 (O_2930,N_48575,N_49431);
or UO_2931 (O_2931,N_48512,N_49509);
nand UO_2932 (O_2932,N_48332,N_48535);
nand UO_2933 (O_2933,N_49134,N_49892);
nor UO_2934 (O_2934,N_49705,N_49611);
nor UO_2935 (O_2935,N_48325,N_48623);
nand UO_2936 (O_2936,N_49619,N_49968);
and UO_2937 (O_2937,N_48234,N_48132);
nor UO_2938 (O_2938,N_49614,N_49865);
nor UO_2939 (O_2939,N_49604,N_48978);
nor UO_2940 (O_2940,N_48219,N_48122);
nor UO_2941 (O_2941,N_49827,N_49867);
and UO_2942 (O_2942,N_49224,N_49242);
nor UO_2943 (O_2943,N_49524,N_49483);
nand UO_2944 (O_2944,N_49788,N_49242);
or UO_2945 (O_2945,N_48947,N_48289);
nand UO_2946 (O_2946,N_49052,N_48368);
nand UO_2947 (O_2947,N_48055,N_48939);
or UO_2948 (O_2948,N_48149,N_48477);
or UO_2949 (O_2949,N_49052,N_48356);
and UO_2950 (O_2950,N_49443,N_49933);
nor UO_2951 (O_2951,N_49518,N_48431);
and UO_2952 (O_2952,N_49860,N_49390);
nor UO_2953 (O_2953,N_48019,N_48584);
nor UO_2954 (O_2954,N_49874,N_48468);
nand UO_2955 (O_2955,N_49992,N_49639);
xnor UO_2956 (O_2956,N_49686,N_49102);
or UO_2957 (O_2957,N_49806,N_49064);
or UO_2958 (O_2958,N_48124,N_48269);
nand UO_2959 (O_2959,N_48664,N_48849);
nand UO_2960 (O_2960,N_48720,N_48052);
and UO_2961 (O_2961,N_48495,N_49530);
xnor UO_2962 (O_2962,N_49180,N_48439);
nand UO_2963 (O_2963,N_48327,N_49521);
nand UO_2964 (O_2964,N_49227,N_48106);
xor UO_2965 (O_2965,N_48372,N_48002);
or UO_2966 (O_2966,N_48111,N_48153);
or UO_2967 (O_2967,N_48578,N_49348);
nor UO_2968 (O_2968,N_48761,N_48048);
xnor UO_2969 (O_2969,N_49385,N_48906);
and UO_2970 (O_2970,N_49746,N_48247);
nand UO_2971 (O_2971,N_49454,N_49099);
or UO_2972 (O_2972,N_48014,N_49297);
or UO_2973 (O_2973,N_49933,N_48877);
nor UO_2974 (O_2974,N_48055,N_49425);
or UO_2975 (O_2975,N_48339,N_48830);
or UO_2976 (O_2976,N_48349,N_49597);
nor UO_2977 (O_2977,N_49268,N_49887);
nand UO_2978 (O_2978,N_49334,N_49866);
and UO_2979 (O_2979,N_49987,N_49003);
xor UO_2980 (O_2980,N_49164,N_48385);
xor UO_2981 (O_2981,N_48349,N_49382);
xnor UO_2982 (O_2982,N_49211,N_48017);
xnor UO_2983 (O_2983,N_48816,N_48481);
nand UO_2984 (O_2984,N_49773,N_49316);
and UO_2985 (O_2985,N_49175,N_48174);
nand UO_2986 (O_2986,N_49343,N_49483);
nand UO_2987 (O_2987,N_48156,N_49162);
or UO_2988 (O_2988,N_49511,N_48936);
nand UO_2989 (O_2989,N_48810,N_49837);
nor UO_2990 (O_2990,N_49033,N_48656);
xnor UO_2991 (O_2991,N_49985,N_48685);
or UO_2992 (O_2992,N_48933,N_48651);
xnor UO_2993 (O_2993,N_48199,N_48509);
nand UO_2994 (O_2994,N_48200,N_49933);
nor UO_2995 (O_2995,N_49937,N_48429);
nand UO_2996 (O_2996,N_49635,N_48594);
nor UO_2997 (O_2997,N_48805,N_48829);
and UO_2998 (O_2998,N_49038,N_49721);
or UO_2999 (O_2999,N_49271,N_49527);
nor UO_3000 (O_3000,N_49021,N_49832);
xnor UO_3001 (O_3001,N_49519,N_48000);
nand UO_3002 (O_3002,N_49736,N_49018);
or UO_3003 (O_3003,N_48323,N_48856);
and UO_3004 (O_3004,N_49014,N_49375);
nor UO_3005 (O_3005,N_49520,N_48635);
or UO_3006 (O_3006,N_49866,N_48437);
nand UO_3007 (O_3007,N_48250,N_49647);
nand UO_3008 (O_3008,N_48493,N_48066);
nand UO_3009 (O_3009,N_48463,N_49969);
and UO_3010 (O_3010,N_48131,N_48349);
and UO_3011 (O_3011,N_49594,N_49617);
xor UO_3012 (O_3012,N_49432,N_49368);
nand UO_3013 (O_3013,N_48486,N_49884);
xor UO_3014 (O_3014,N_49104,N_48054);
and UO_3015 (O_3015,N_49342,N_49706);
and UO_3016 (O_3016,N_48976,N_48273);
nor UO_3017 (O_3017,N_48707,N_49279);
nor UO_3018 (O_3018,N_48318,N_49085);
nand UO_3019 (O_3019,N_49764,N_48801);
nor UO_3020 (O_3020,N_48880,N_48215);
and UO_3021 (O_3021,N_48302,N_48249);
or UO_3022 (O_3022,N_48648,N_48111);
nor UO_3023 (O_3023,N_49067,N_48718);
or UO_3024 (O_3024,N_48033,N_49420);
xnor UO_3025 (O_3025,N_49245,N_48046);
and UO_3026 (O_3026,N_48248,N_49303);
or UO_3027 (O_3027,N_48215,N_49176);
xnor UO_3028 (O_3028,N_48487,N_48904);
or UO_3029 (O_3029,N_49264,N_48641);
xor UO_3030 (O_3030,N_48899,N_48191);
xor UO_3031 (O_3031,N_49387,N_48303);
and UO_3032 (O_3032,N_48887,N_48052);
nor UO_3033 (O_3033,N_48768,N_49941);
and UO_3034 (O_3034,N_49004,N_48094);
or UO_3035 (O_3035,N_49004,N_49715);
and UO_3036 (O_3036,N_48387,N_48260);
nand UO_3037 (O_3037,N_49198,N_49192);
and UO_3038 (O_3038,N_48224,N_48874);
nand UO_3039 (O_3039,N_49950,N_49350);
xnor UO_3040 (O_3040,N_49230,N_49526);
nor UO_3041 (O_3041,N_48516,N_48082);
or UO_3042 (O_3042,N_49648,N_49493);
nand UO_3043 (O_3043,N_49036,N_49218);
nor UO_3044 (O_3044,N_48427,N_48362);
xnor UO_3045 (O_3045,N_48469,N_49715);
nor UO_3046 (O_3046,N_49197,N_49534);
xor UO_3047 (O_3047,N_48708,N_48897);
or UO_3048 (O_3048,N_48314,N_48498);
nand UO_3049 (O_3049,N_48546,N_49385);
nand UO_3050 (O_3050,N_48465,N_48117);
nor UO_3051 (O_3051,N_49538,N_48157);
and UO_3052 (O_3052,N_49141,N_48549);
and UO_3053 (O_3053,N_48965,N_49568);
nand UO_3054 (O_3054,N_49317,N_48769);
nand UO_3055 (O_3055,N_49633,N_49390);
nor UO_3056 (O_3056,N_49588,N_49176);
and UO_3057 (O_3057,N_49873,N_49817);
and UO_3058 (O_3058,N_48323,N_49364);
xor UO_3059 (O_3059,N_49109,N_48797);
or UO_3060 (O_3060,N_48791,N_49281);
nor UO_3061 (O_3061,N_49928,N_49221);
and UO_3062 (O_3062,N_48024,N_49950);
and UO_3063 (O_3063,N_48463,N_49479);
or UO_3064 (O_3064,N_48486,N_48985);
xor UO_3065 (O_3065,N_49967,N_49522);
and UO_3066 (O_3066,N_48078,N_49395);
or UO_3067 (O_3067,N_48848,N_48537);
nand UO_3068 (O_3068,N_49569,N_48291);
or UO_3069 (O_3069,N_48927,N_48379);
or UO_3070 (O_3070,N_49911,N_48602);
and UO_3071 (O_3071,N_49700,N_48788);
xnor UO_3072 (O_3072,N_48653,N_49415);
and UO_3073 (O_3073,N_48077,N_49996);
or UO_3074 (O_3074,N_49652,N_48637);
and UO_3075 (O_3075,N_49312,N_49150);
or UO_3076 (O_3076,N_49920,N_48265);
nand UO_3077 (O_3077,N_49123,N_48532);
nand UO_3078 (O_3078,N_49797,N_48373);
xor UO_3079 (O_3079,N_49824,N_48471);
or UO_3080 (O_3080,N_48327,N_49006);
or UO_3081 (O_3081,N_49056,N_49003);
and UO_3082 (O_3082,N_48782,N_49099);
or UO_3083 (O_3083,N_48323,N_48494);
nand UO_3084 (O_3084,N_49800,N_48406);
and UO_3085 (O_3085,N_48187,N_49821);
or UO_3086 (O_3086,N_48591,N_49231);
xor UO_3087 (O_3087,N_48884,N_49884);
or UO_3088 (O_3088,N_48763,N_48990);
nor UO_3089 (O_3089,N_49902,N_49622);
and UO_3090 (O_3090,N_49596,N_48337);
nor UO_3091 (O_3091,N_48818,N_48130);
xor UO_3092 (O_3092,N_49801,N_48866);
and UO_3093 (O_3093,N_48955,N_48472);
xor UO_3094 (O_3094,N_48615,N_49600);
nand UO_3095 (O_3095,N_49597,N_48655);
nor UO_3096 (O_3096,N_48184,N_48713);
or UO_3097 (O_3097,N_48226,N_48960);
xnor UO_3098 (O_3098,N_49110,N_48184);
nor UO_3099 (O_3099,N_48775,N_48415);
nor UO_3100 (O_3100,N_48665,N_49022);
nor UO_3101 (O_3101,N_48569,N_48107);
or UO_3102 (O_3102,N_48243,N_49701);
and UO_3103 (O_3103,N_49525,N_48556);
nor UO_3104 (O_3104,N_48056,N_49934);
nand UO_3105 (O_3105,N_49742,N_49086);
nor UO_3106 (O_3106,N_49027,N_48027);
or UO_3107 (O_3107,N_49131,N_48947);
nor UO_3108 (O_3108,N_48136,N_48088);
nand UO_3109 (O_3109,N_48139,N_49988);
nand UO_3110 (O_3110,N_49753,N_49254);
and UO_3111 (O_3111,N_49220,N_49391);
and UO_3112 (O_3112,N_49034,N_49057);
nor UO_3113 (O_3113,N_49444,N_48461);
and UO_3114 (O_3114,N_49129,N_48213);
and UO_3115 (O_3115,N_48445,N_49076);
nor UO_3116 (O_3116,N_48370,N_48118);
or UO_3117 (O_3117,N_48730,N_48462);
nor UO_3118 (O_3118,N_48785,N_49581);
xnor UO_3119 (O_3119,N_48239,N_49843);
nor UO_3120 (O_3120,N_48756,N_48810);
or UO_3121 (O_3121,N_48479,N_48752);
or UO_3122 (O_3122,N_48539,N_48196);
nor UO_3123 (O_3123,N_49329,N_49038);
nand UO_3124 (O_3124,N_48838,N_48253);
or UO_3125 (O_3125,N_49712,N_48317);
nor UO_3126 (O_3126,N_49967,N_48601);
and UO_3127 (O_3127,N_48074,N_49357);
nor UO_3128 (O_3128,N_49604,N_48793);
xnor UO_3129 (O_3129,N_48897,N_49897);
nand UO_3130 (O_3130,N_48890,N_49391);
nand UO_3131 (O_3131,N_49794,N_49429);
nand UO_3132 (O_3132,N_48901,N_49876);
nand UO_3133 (O_3133,N_48046,N_48042);
xnor UO_3134 (O_3134,N_48051,N_48351);
xnor UO_3135 (O_3135,N_48421,N_49684);
nor UO_3136 (O_3136,N_49481,N_48146);
or UO_3137 (O_3137,N_48760,N_48310);
nand UO_3138 (O_3138,N_48735,N_48447);
nand UO_3139 (O_3139,N_49432,N_49092);
nand UO_3140 (O_3140,N_48907,N_48662);
and UO_3141 (O_3141,N_48121,N_48361);
nand UO_3142 (O_3142,N_49321,N_48138);
nor UO_3143 (O_3143,N_49955,N_48767);
nand UO_3144 (O_3144,N_48415,N_49426);
xor UO_3145 (O_3145,N_49185,N_49564);
xor UO_3146 (O_3146,N_48921,N_48627);
nand UO_3147 (O_3147,N_48498,N_48680);
nor UO_3148 (O_3148,N_49764,N_49377);
and UO_3149 (O_3149,N_48827,N_48022);
or UO_3150 (O_3150,N_49427,N_49722);
nand UO_3151 (O_3151,N_49063,N_48840);
nor UO_3152 (O_3152,N_48393,N_48833);
and UO_3153 (O_3153,N_49025,N_48085);
and UO_3154 (O_3154,N_48743,N_48883);
nor UO_3155 (O_3155,N_49020,N_49253);
or UO_3156 (O_3156,N_49900,N_49223);
or UO_3157 (O_3157,N_49178,N_49190);
nor UO_3158 (O_3158,N_49761,N_49462);
and UO_3159 (O_3159,N_48747,N_49143);
nand UO_3160 (O_3160,N_49821,N_49635);
nand UO_3161 (O_3161,N_49701,N_49045);
xnor UO_3162 (O_3162,N_48033,N_49814);
and UO_3163 (O_3163,N_48076,N_49062);
xor UO_3164 (O_3164,N_49347,N_48431);
nand UO_3165 (O_3165,N_49165,N_49220);
or UO_3166 (O_3166,N_48519,N_48196);
and UO_3167 (O_3167,N_48032,N_49902);
xor UO_3168 (O_3168,N_48203,N_48158);
or UO_3169 (O_3169,N_48644,N_49902);
or UO_3170 (O_3170,N_49782,N_48242);
and UO_3171 (O_3171,N_49623,N_48471);
or UO_3172 (O_3172,N_48776,N_48236);
xor UO_3173 (O_3173,N_49818,N_49924);
and UO_3174 (O_3174,N_48520,N_49768);
and UO_3175 (O_3175,N_49374,N_48904);
nand UO_3176 (O_3176,N_49672,N_48981);
nand UO_3177 (O_3177,N_49821,N_49310);
xor UO_3178 (O_3178,N_49954,N_49298);
nand UO_3179 (O_3179,N_48379,N_49169);
xnor UO_3180 (O_3180,N_49379,N_49892);
or UO_3181 (O_3181,N_48054,N_49580);
and UO_3182 (O_3182,N_49234,N_49787);
nor UO_3183 (O_3183,N_48642,N_48856);
and UO_3184 (O_3184,N_48133,N_48419);
nor UO_3185 (O_3185,N_48266,N_48956);
xnor UO_3186 (O_3186,N_48386,N_48277);
nand UO_3187 (O_3187,N_49221,N_49003);
or UO_3188 (O_3188,N_48185,N_49896);
and UO_3189 (O_3189,N_49655,N_49982);
xor UO_3190 (O_3190,N_48820,N_49454);
or UO_3191 (O_3191,N_48984,N_48767);
xnor UO_3192 (O_3192,N_48715,N_49310);
and UO_3193 (O_3193,N_49546,N_48985);
or UO_3194 (O_3194,N_48890,N_49909);
nand UO_3195 (O_3195,N_48277,N_49751);
xnor UO_3196 (O_3196,N_48672,N_49014);
xnor UO_3197 (O_3197,N_48757,N_48167);
or UO_3198 (O_3198,N_49545,N_49717);
nand UO_3199 (O_3199,N_49416,N_48745);
xor UO_3200 (O_3200,N_48335,N_49621);
and UO_3201 (O_3201,N_49184,N_48359);
nand UO_3202 (O_3202,N_48034,N_49851);
nand UO_3203 (O_3203,N_49902,N_49765);
nand UO_3204 (O_3204,N_48011,N_49591);
xnor UO_3205 (O_3205,N_48840,N_48685);
nand UO_3206 (O_3206,N_48966,N_49763);
nand UO_3207 (O_3207,N_49882,N_49299);
or UO_3208 (O_3208,N_48725,N_49811);
xnor UO_3209 (O_3209,N_49375,N_49240);
xor UO_3210 (O_3210,N_49939,N_48399);
and UO_3211 (O_3211,N_49699,N_48379);
or UO_3212 (O_3212,N_48509,N_48873);
nand UO_3213 (O_3213,N_49905,N_48222);
nor UO_3214 (O_3214,N_48892,N_49188);
nor UO_3215 (O_3215,N_49364,N_48871);
nor UO_3216 (O_3216,N_48022,N_49166);
or UO_3217 (O_3217,N_49734,N_49360);
nand UO_3218 (O_3218,N_48429,N_49326);
nand UO_3219 (O_3219,N_49189,N_49059);
nor UO_3220 (O_3220,N_49405,N_48015);
and UO_3221 (O_3221,N_49247,N_49549);
xor UO_3222 (O_3222,N_48852,N_48123);
and UO_3223 (O_3223,N_48821,N_48950);
nand UO_3224 (O_3224,N_48955,N_48141);
xor UO_3225 (O_3225,N_49468,N_48694);
nor UO_3226 (O_3226,N_49011,N_49326);
or UO_3227 (O_3227,N_48064,N_49008);
xor UO_3228 (O_3228,N_48610,N_49472);
and UO_3229 (O_3229,N_49565,N_49090);
and UO_3230 (O_3230,N_48563,N_48191);
nand UO_3231 (O_3231,N_49086,N_48105);
or UO_3232 (O_3232,N_48271,N_48252);
nand UO_3233 (O_3233,N_48910,N_49047);
or UO_3234 (O_3234,N_48519,N_49517);
xor UO_3235 (O_3235,N_48661,N_48309);
or UO_3236 (O_3236,N_49577,N_48060);
xnor UO_3237 (O_3237,N_49777,N_48215);
xor UO_3238 (O_3238,N_49955,N_48044);
nand UO_3239 (O_3239,N_49675,N_48661);
or UO_3240 (O_3240,N_48076,N_49579);
and UO_3241 (O_3241,N_48576,N_48515);
xnor UO_3242 (O_3242,N_49950,N_48344);
or UO_3243 (O_3243,N_48876,N_48651);
xor UO_3244 (O_3244,N_48286,N_49445);
and UO_3245 (O_3245,N_49594,N_48113);
nand UO_3246 (O_3246,N_48371,N_48087);
nor UO_3247 (O_3247,N_48501,N_49830);
xnor UO_3248 (O_3248,N_49909,N_49439);
or UO_3249 (O_3249,N_48942,N_49863);
and UO_3250 (O_3250,N_48833,N_48482);
and UO_3251 (O_3251,N_49872,N_48544);
nor UO_3252 (O_3252,N_48239,N_49419);
xnor UO_3253 (O_3253,N_48843,N_49426);
or UO_3254 (O_3254,N_49346,N_48609);
or UO_3255 (O_3255,N_48918,N_48344);
or UO_3256 (O_3256,N_48460,N_49439);
and UO_3257 (O_3257,N_49311,N_49866);
xnor UO_3258 (O_3258,N_48496,N_49156);
or UO_3259 (O_3259,N_48568,N_49718);
or UO_3260 (O_3260,N_49806,N_48672);
or UO_3261 (O_3261,N_48904,N_49568);
nor UO_3262 (O_3262,N_48282,N_49589);
and UO_3263 (O_3263,N_49537,N_48049);
xnor UO_3264 (O_3264,N_48986,N_48579);
xor UO_3265 (O_3265,N_49422,N_49617);
xor UO_3266 (O_3266,N_48026,N_48460);
nor UO_3267 (O_3267,N_48830,N_49947);
nor UO_3268 (O_3268,N_48871,N_48026);
and UO_3269 (O_3269,N_49591,N_48557);
nand UO_3270 (O_3270,N_48477,N_48720);
nor UO_3271 (O_3271,N_48095,N_48997);
and UO_3272 (O_3272,N_48374,N_49778);
nand UO_3273 (O_3273,N_48495,N_48845);
or UO_3274 (O_3274,N_48018,N_49832);
and UO_3275 (O_3275,N_48365,N_49715);
and UO_3276 (O_3276,N_49709,N_49796);
or UO_3277 (O_3277,N_49382,N_48993);
or UO_3278 (O_3278,N_49016,N_49442);
and UO_3279 (O_3279,N_49278,N_49577);
xor UO_3280 (O_3280,N_49035,N_48637);
nand UO_3281 (O_3281,N_48421,N_49481);
nor UO_3282 (O_3282,N_49452,N_48011);
nor UO_3283 (O_3283,N_49978,N_48416);
and UO_3284 (O_3284,N_49775,N_48532);
and UO_3285 (O_3285,N_48534,N_49359);
nand UO_3286 (O_3286,N_49011,N_48838);
nand UO_3287 (O_3287,N_49131,N_49159);
xor UO_3288 (O_3288,N_49626,N_49111);
nor UO_3289 (O_3289,N_49295,N_49058);
or UO_3290 (O_3290,N_48468,N_49416);
and UO_3291 (O_3291,N_49134,N_49950);
xnor UO_3292 (O_3292,N_48547,N_48918);
nor UO_3293 (O_3293,N_49749,N_48276);
nor UO_3294 (O_3294,N_49170,N_48373);
nor UO_3295 (O_3295,N_48492,N_48484);
nand UO_3296 (O_3296,N_49451,N_49028);
and UO_3297 (O_3297,N_49329,N_48060);
xnor UO_3298 (O_3298,N_49002,N_48705);
nand UO_3299 (O_3299,N_48381,N_48542);
and UO_3300 (O_3300,N_49483,N_48575);
xnor UO_3301 (O_3301,N_48251,N_49612);
nand UO_3302 (O_3302,N_48526,N_49621);
or UO_3303 (O_3303,N_48720,N_49598);
or UO_3304 (O_3304,N_48133,N_48390);
or UO_3305 (O_3305,N_48580,N_49212);
nor UO_3306 (O_3306,N_48122,N_48922);
and UO_3307 (O_3307,N_48727,N_49849);
or UO_3308 (O_3308,N_48088,N_49453);
or UO_3309 (O_3309,N_49066,N_48794);
and UO_3310 (O_3310,N_49345,N_49677);
nor UO_3311 (O_3311,N_48061,N_48500);
or UO_3312 (O_3312,N_49016,N_48254);
nand UO_3313 (O_3313,N_49033,N_48264);
and UO_3314 (O_3314,N_48690,N_48866);
nand UO_3315 (O_3315,N_48040,N_48821);
or UO_3316 (O_3316,N_49052,N_48290);
nor UO_3317 (O_3317,N_48939,N_49126);
nand UO_3318 (O_3318,N_49458,N_49881);
and UO_3319 (O_3319,N_48749,N_49558);
and UO_3320 (O_3320,N_48889,N_48289);
nor UO_3321 (O_3321,N_48866,N_48539);
nand UO_3322 (O_3322,N_48451,N_49854);
xor UO_3323 (O_3323,N_48308,N_48422);
and UO_3324 (O_3324,N_48587,N_49593);
nor UO_3325 (O_3325,N_49519,N_48778);
or UO_3326 (O_3326,N_48887,N_49385);
and UO_3327 (O_3327,N_48480,N_49841);
nand UO_3328 (O_3328,N_48730,N_49634);
nor UO_3329 (O_3329,N_49953,N_49156);
xor UO_3330 (O_3330,N_49177,N_48291);
nand UO_3331 (O_3331,N_49455,N_49132);
or UO_3332 (O_3332,N_48751,N_48207);
or UO_3333 (O_3333,N_49796,N_49807);
nand UO_3334 (O_3334,N_49668,N_48345);
or UO_3335 (O_3335,N_49409,N_48053);
nor UO_3336 (O_3336,N_48362,N_49286);
nor UO_3337 (O_3337,N_49518,N_48958);
xor UO_3338 (O_3338,N_49784,N_49184);
and UO_3339 (O_3339,N_49498,N_49909);
xnor UO_3340 (O_3340,N_49208,N_48210);
and UO_3341 (O_3341,N_49917,N_48084);
or UO_3342 (O_3342,N_48122,N_49266);
nand UO_3343 (O_3343,N_49212,N_48799);
nor UO_3344 (O_3344,N_48692,N_48542);
nor UO_3345 (O_3345,N_48115,N_48216);
and UO_3346 (O_3346,N_49771,N_48137);
nand UO_3347 (O_3347,N_48165,N_49876);
and UO_3348 (O_3348,N_49357,N_49614);
or UO_3349 (O_3349,N_48407,N_48572);
or UO_3350 (O_3350,N_49935,N_49868);
xnor UO_3351 (O_3351,N_49577,N_49085);
or UO_3352 (O_3352,N_48715,N_48992);
nand UO_3353 (O_3353,N_48521,N_48112);
or UO_3354 (O_3354,N_49406,N_48443);
or UO_3355 (O_3355,N_49785,N_49174);
nand UO_3356 (O_3356,N_49459,N_49104);
nor UO_3357 (O_3357,N_48546,N_49687);
nand UO_3358 (O_3358,N_49352,N_49636);
or UO_3359 (O_3359,N_48209,N_48550);
and UO_3360 (O_3360,N_48447,N_49126);
xnor UO_3361 (O_3361,N_49820,N_49791);
and UO_3362 (O_3362,N_48406,N_49545);
and UO_3363 (O_3363,N_48864,N_48670);
xor UO_3364 (O_3364,N_48980,N_49818);
nor UO_3365 (O_3365,N_49698,N_48710);
and UO_3366 (O_3366,N_49105,N_48747);
or UO_3367 (O_3367,N_48052,N_48786);
xnor UO_3368 (O_3368,N_48180,N_49167);
and UO_3369 (O_3369,N_49796,N_48662);
nor UO_3370 (O_3370,N_49999,N_49358);
nand UO_3371 (O_3371,N_49751,N_49088);
xor UO_3372 (O_3372,N_49785,N_49780);
and UO_3373 (O_3373,N_49322,N_48833);
and UO_3374 (O_3374,N_48004,N_49386);
nand UO_3375 (O_3375,N_48036,N_49984);
nand UO_3376 (O_3376,N_48464,N_49613);
nor UO_3377 (O_3377,N_49767,N_48471);
and UO_3378 (O_3378,N_49408,N_49026);
and UO_3379 (O_3379,N_49775,N_48877);
and UO_3380 (O_3380,N_48789,N_48934);
nand UO_3381 (O_3381,N_48610,N_48398);
and UO_3382 (O_3382,N_48030,N_48826);
or UO_3383 (O_3383,N_49733,N_48136);
nor UO_3384 (O_3384,N_48339,N_48872);
xor UO_3385 (O_3385,N_48093,N_48120);
and UO_3386 (O_3386,N_49526,N_49129);
and UO_3387 (O_3387,N_49217,N_49937);
nor UO_3388 (O_3388,N_48659,N_48894);
nor UO_3389 (O_3389,N_48575,N_49429);
and UO_3390 (O_3390,N_49226,N_49043);
and UO_3391 (O_3391,N_48032,N_49896);
and UO_3392 (O_3392,N_49036,N_49183);
nand UO_3393 (O_3393,N_49687,N_48499);
nand UO_3394 (O_3394,N_48825,N_48744);
xnor UO_3395 (O_3395,N_49152,N_49685);
nor UO_3396 (O_3396,N_48835,N_48493);
and UO_3397 (O_3397,N_48659,N_48531);
nor UO_3398 (O_3398,N_48664,N_48811);
and UO_3399 (O_3399,N_48486,N_49305);
nor UO_3400 (O_3400,N_49408,N_49046);
and UO_3401 (O_3401,N_48822,N_48547);
and UO_3402 (O_3402,N_49994,N_48079);
nor UO_3403 (O_3403,N_49748,N_48671);
nand UO_3404 (O_3404,N_48654,N_48570);
xnor UO_3405 (O_3405,N_48380,N_49088);
or UO_3406 (O_3406,N_49089,N_48048);
nor UO_3407 (O_3407,N_49180,N_48348);
nor UO_3408 (O_3408,N_49249,N_48715);
xnor UO_3409 (O_3409,N_48196,N_48243);
nor UO_3410 (O_3410,N_48897,N_49968);
and UO_3411 (O_3411,N_49191,N_49770);
nand UO_3412 (O_3412,N_49990,N_49140);
xor UO_3413 (O_3413,N_48315,N_49082);
xnor UO_3414 (O_3414,N_49796,N_49599);
nand UO_3415 (O_3415,N_48170,N_49946);
nor UO_3416 (O_3416,N_49248,N_48785);
xnor UO_3417 (O_3417,N_49636,N_48790);
nand UO_3418 (O_3418,N_49824,N_49799);
nand UO_3419 (O_3419,N_48931,N_48725);
nand UO_3420 (O_3420,N_49372,N_49428);
nand UO_3421 (O_3421,N_49879,N_48766);
and UO_3422 (O_3422,N_48694,N_48500);
nand UO_3423 (O_3423,N_49048,N_48258);
or UO_3424 (O_3424,N_49111,N_49965);
xor UO_3425 (O_3425,N_48630,N_48994);
nand UO_3426 (O_3426,N_49952,N_48851);
nor UO_3427 (O_3427,N_49038,N_48657);
nand UO_3428 (O_3428,N_48039,N_49282);
nor UO_3429 (O_3429,N_49801,N_48556);
and UO_3430 (O_3430,N_48253,N_48820);
xnor UO_3431 (O_3431,N_49483,N_48049);
xor UO_3432 (O_3432,N_49861,N_48128);
or UO_3433 (O_3433,N_49415,N_48615);
nor UO_3434 (O_3434,N_49710,N_49217);
nand UO_3435 (O_3435,N_48924,N_49443);
nand UO_3436 (O_3436,N_49222,N_49529);
nor UO_3437 (O_3437,N_49814,N_49291);
or UO_3438 (O_3438,N_49564,N_48086);
and UO_3439 (O_3439,N_48801,N_48580);
nor UO_3440 (O_3440,N_48742,N_49884);
nand UO_3441 (O_3441,N_49917,N_48953);
nor UO_3442 (O_3442,N_49392,N_48200);
nand UO_3443 (O_3443,N_48004,N_48854);
or UO_3444 (O_3444,N_48313,N_49156);
or UO_3445 (O_3445,N_49181,N_49300);
nor UO_3446 (O_3446,N_48249,N_49207);
nand UO_3447 (O_3447,N_48482,N_48700);
or UO_3448 (O_3448,N_49752,N_49491);
nor UO_3449 (O_3449,N_48836,N_49542);
xor UO_3450 (O_3450,N_48929,N_49154);
or UO_3451 (O_3451,N_48953,N_48332);
xor UO_3452 (O_3452,N_48535,N_49930);
and UO_3453 (O_3453,N_49240,N_49562);
nor UO_3454 (O_3454,N_48692,N_49253);
xnor UO_3455 (O_3455,N_48133,N_48480);
or UO_3456 (O_3456,N_49223,N_48784);
and UO_3457 (O_3457,N_48158,N_49923);
nand UO_3458 (O_3458,N_48411,N_49759);
and UO_3459 (O_3459,N_48913,N_49035);
nand UO_3460 (O_3460,N_49945,N_48005);
or UO_3461 (O_3461,N_48466,N_48731);
nand UO_3462 (O_3462,N_48492,N_49591);
xor UO_3463 (O_3463,N_49325,N_49644);
nand UO_3464 (O_3464,N_48506,N_49338);
nand UO_3465 (O_3465,N_49922,N_48205);
or UO_3466 (O_3466,N_48134,N_49455);
or UO_3467 (O_3467,N_48935,N_49906);
xnor UO_3468 (O_3468,N_49172,N_49945);
or UO_3469 (O_3469,N_48319,N_49529);
and UO_3470 (O_3470,N_49095,N_48069);
xnor UO_3471 (O_3471,N_48979,N_48283);
nand UO_3472 (O_3472,N_48498,N_48666);
or UO_3473 (O_3473,N_48419,N_49327);
nand UO_3474 (O_3474,N_48671,N_49891);
nand UO_3475 (O_3475,N_48590,N_48612);
nand UO_3476 (O_3476,N_48098,N_48250);
or UO_3477 (O_3477,N_48751,N_49014);
nand UO_3478 (O_3478,N_48864,N_48938);
or UO_3479 (O_3479,N_48634,N_48659);
nand UO_3480 (O_3480,N_49263,N_49218);
xnor UO_3481 (O_3481,N_49201,N_48170);
or UO_3482 (O_3482,N_48778,N_48050);
xor UO_3483 (O_3483,N_49252,N_48838);
and UO_3484 (O_3484,N_48768,N_49910);
xor UO_3485 (O_3485,N_49222,N_48841);
nand UO_3486 (O_3486,N_48526,N_49951);
xor UO_3487 (O_3487,N_48117,N_49203);
nand UO_3488 (O_3488,N_49493,N_49053);
nand UO_3489 (O_3489,N_48991,N_49149);
or UO_3490 (O_3490,N_49957,N_49477);
nand UO_3491 (O_3491,N_48248,N_49070);
nor UO_3492 (O_3492,N_49871,N_48281);
nor UO_3493 (O_3493,N_49435,N_49961);
or UO_3494 (O_3494,N_48547,N_48485);
or UO_3495 (O_3495,N_49442,N_49059);
and UO_3496 (O_3496,N_48253,N_49229);
nand UO_3497 (O_3497,N_49146,N_49880);
xnor UO_3498 (O_3498,N_48533,N_49150);
nand UO_3499 (O_3499,N_48167,N_48468);
and UO_3500 (O_3500,N_49050,N_48980);
or UO_3501 (O_3501,N_48145,N_48413);
nor UO_3502 (O_3502,N_48531,N_49951);
or UO_3503 (O_3503,N_49581,N_48170);
xor UO_3504 (O_3504,N_48965,N_49158);
nand UO_3505 (O_3505,N_49160,N_49499);
nand UO_3506 (O_3506,N_48221,N_48360);
nand UO_3507 (O_3507,N_48097,N_49804);
xor UO_3508 (O_3508,N_48757,N_48431);
or UO_3509 (O_3509,N_49039,N_48941);
xor UO_3510 (O_3510,N_49388,N_49247);
or UO_3511 (O_3511,N_48449,N_49364);
or UO_3512 (O_3512,N_49385,N_48066);
nor UO_3513 (O_3513,N_49363,N_48627);
nand UO_3514 (O_3514,N_49996,N_49401);
nor UO_3515 (O_3515,N_49177,N_49148);
xnor UO_3516 (O_3516,N_48807,N_49621);
nand UO_3517 (O_3517,N_48193,N_48626);
nand UO_3518 (O_3518,N_49602,N_48842);
or UO_3519 (O_3519,N_48029,N_48187);
nand UO_3520 (O_3520,N_49094,N_49872);
xnor UO_3521 (O_3521,N_49925,N_48508);
and UO_3522 (O_3522,N_49493,N_49955);
xor UO_3523 (O_3523,N_48398,N_49281);
nand UO_3524 (O_3524,N_48612,N_49583);
nor UO_3525 (O_3525,N_48646,N_49542);
or UO_3526 (O_3526,N_49470,N_48890);
nand UO_3527 (O_3527,N_48892,N_49094);
or UO_3528 (O_3528,N_49078,N_48386);
or UO_3529 (O_3529,N_49792,N_49501);
or UO_3530 (O_3530,N_49510,N_49798);
nor UO_3531 (O_3531,N_48701,N_49879);
or UO_3532 (O_3532,N_48361,N_48648);
nand UO_3533 (O_3533,N_49846,N_48169);
nand UO_3534 (O_3534,N_48144,N_48810);
or UO_3535 (O_3535,N_48940,N_49230);
or UO_3536 (O_3536,N_48379,N_49453);
nor UO_3537 (O_3537,N_49901,N_48256);
or UO_3538 (O_3538,N_48331,N_48528);
or UO_3539 (O_3539,N_49307,N_48537);
xor UO_3540 (O_3540,N_48714,N_48853);
and UO_3541 (O_3541,N_49745,N_49184);
nor UO_3542 (O_3542,N_49753,N_49080);
nor UO_3543 (O_3543,N_48018,N_49157);
or UO_3544 (O_3544,N_49149,N_48194);
xnor UO_3545 (O_3545,N_48413,N_49505);
nor UO_3546 (O_3546,N_48801,N_48196);
and UO_3547 (O_3547,N_48226,N_48854);
nand UO_3548 (O_3548,N_48607,N_49195);
or UO_3549 (O_3549,N_49608,N_48713);
or UO_3550 (O_3550,N_48719,N_49065);
and UO_3551 (O_3551,N_48374,N_49781);
and UO_3552 (O_3552,N_48267,N_48164);
xnor UO_3553 (O_3553,N_48700,N_48885);
or UO_3554 (O_3554,N_48531,N_48295);
xnor UO_3555 (O_3555,N_49835,N_49912);
xnor UO_3556 (O_3556,N_49824,N_48980);
or UO_3557 (O_3557,N_49391,N_48711);
and UO_3558 (O_3558,N_48586,N_48519);
nand UO_3559 (O_3559,N_48746,N_49509);
nand UO_3560 (O_3560,N_49698,N_48734);
nand UO_3561 (O_3561,N_49296,N_49142);
or UO_3562 (O_3562,N_48494,N_48890);
nor UO_3563 (O_3563,N_48740,N_49040);
or UO_3564 (O_3564,N_48163,N_48301);
nand UO_3565 (O_3565,N_48058,N_48436);
xnor UO_3566 (O_3566,N_48461,N_49615);
nand UO_3567 (O_3567,N_48182,N_49610);
or UO_3568 (O_3568,N_49260,N_48256);
xnor UO_3569 (O_3569,N_49167,N_48804);
or UO_3570 (O_3570,N_49685,N_49784);
xnor UO_3571 (O_3571,N_49389,N_48484);
and UO_3572 (O_3572,N_49223,N_49141);
nor UO_3573 (O_3573,N_49168,N_48700);
nor UO_3574 (O_3574,N_48150,N_48275);
and UO_3575 (O_3575,N_48821,N_49787);
xnor UO_3576 (O_3576,N_49918,N_49752);
or UO_3577 (O_3577,N_49810,N_48102);
xnor UO_3578 (O_3578,N_48972,N_49291);
and UO_3579 (O_3579,N_48186,N_48029);
or UO_3580 (O_3580,N_49818,N_48166);
or UO_3581 (O_3581,N_49659,N_49143);
and UO_3582 (O_3582,N_48853,N_49232);
nor UO_3583 (O_3583,N_49918,N_48224);
nand UO_3584 (O_3584,N_48563,N_48773);
nor UO_3585 (O_3585,N_49984,N_49305);
and UO_3586 (O_3586,N_49524,N_49030);
and UO_3587 (O_3587,N_48482,N_48039);
nor UO_3588 (O_3588,N_48481,N_49852);
nor UO_3589 (O_3589,N_49163,N_48785);
nor UO_3590 (O_3590,N_49524,N_49838);
and UO_3591 (O_3591,N_48219,N_49689);
nand UO_3592 (O_3592,N_48468,N_48224);
nand UO_3593 (O_3593,N_49262,N_49103);
nand UO_3594 (O_3594,N_49040,N_48178);
xnor UO_3595 (O_3595,N_48768,N_49176);
nor UO_3596 (O_3596,N_49741,N_48422);
xor UO_3597 (O_3597,N_49089,N_49796);
xnor UO_3598 (O_3598,N_48815,N_48628);
xnor UO_3599 (O_3599,N_48969,N_48624);
xor UO_3600 (O_3600,N_48787,N_48186);
nand UO_3601 (O_3601,N_49898,N_49115);
and UO_3602 (O_3602,N_48895,N_48966);
nor UO_3603 (O_3603,N_48268,N_48117);
xor UO_3604 (O_3604,N_48784,N_49534);
or UO_3605 (O_3605,N_48569,N_48864);
or UO_3606 (O_3606,N_49452,N_48194);
or UO_3607 (O_3607,N_48499,N_48943);
and UO_3608 (O_3608,N_49333,N_48906);
xor UO_3609 (O_3609,N_48208,N_48493);
nand UO_3610 (O_3610,N_48622,N_49211);
nand UO_3611 (O_3611,N_49770,N_48312);
and UO_3612 (O_3612,N_48775,N_49990);
nand UO_3613 (O_3613,N_49016,N_48548);
or UO_3614 (O_3614,N_48476,N_49705);
xnor UO_3615 (O_3615,N_49853,N_48843);
nor UO_3616 (O_3616,N_48992,N_49541);
nand UO_3617 (O_3617,N_49875,N_48911);
or UO_3618 (O_3618,N_48399,N_48503);
nand UO_3619 (O_3619,N_49225,N_49813);
or UO_3620 (O_3620,N_49110,N_48053);
nor UO_3621 (O_3621,N_48003,N_48989);
nor UO_3622 (O_3622,N_49248,N_48433);
and UO_3623 (O_3623,N_49851,N_48198);
and UO_3624 (O_3624,N_49637,N_49119);
xor UO_3625 (O_3625,N_49772,N_49198);
xnor UO_3626 (O_3626,N_49229,N_48377);
or UO_3627 (O_3627,N_49763,N_49252);
and UO_3628 (O_3628,N_48251,N_49721);
or UO_3629 (O_3629,N_48554,N_49357);
nor UO_3630 (O_3630,N_49448,N_48443);
xor UO_3631 (O_3631,N_49247,N_49508);
and UO_3632 (O_3632,N_49631,N_48637);
or UO_3633 (O_3633,N_49945,N_49047);
nor UO_3634 (O_3634,N_49742,N_48127);
nand UO_3635 (O_3635,N_48429,N_48019);
xnor UO_3636 (O_3636,N_48378,N_49351);
and UO_3637 (O_3637,N_49623,N_49462);
or UO_3638 (O_3638,N_48137,N_48457);
nor UO_3639 (O_3639,N_49007,N_48616);
or UO_3640 (O_3640,N_49163,N_49184);
nand UO_3641 (O_3641,N_49449,N_49618);
nand UO_3642 (O_3642,N_49144,N_49263);
nor UO_3643 (O_3643,N_49056,N_48309);
nor UO_3644 (O_3644,N_48838,N_49249);
xnor UO_3645 (O_3645,N_49087,N_48351);
xor UO_3646 (O_3646,N_49378,N_49544);
or UO_3647 (O_3647,N_49251,N_48973);
nand UO_3648 (O_3648,N_49685,N_49732);
or UO_3649 (O_3649,N_48358,N_49814);
or UO_3650 (O_3650,N_48126,N_48364);
or UO_3651 (O_3651,N_49487,N_48128);
nor UO_3652 (O_3652,N_49522,N_48072);
nand UO_3653 (O_3653,N_48945,N_48350);
or UO_3654 (O_3654,N_48749,N_48052);
and UO_3655 (O_3655,N_49730,N_49427);
and UO_3656 (O_3656,N_48394,N_49021);
xnor UO_3657 (O_3657,N_48468,N_49499);
or UO_3658 (O_3658,N_48970,N_49411);
and UO_3659 (O_3659,N_48030,N_48258);
xor UO_3660 (O_3660,N_49076,N_49780);
xnor UO_3661 (O_3661,N_48205,N_49966);
nor UO_3662 (O_3662,N_49557,N_49001);
or UO_3663 (O_3663,N_49586,N_48248);
xnor UO_3664 (O_3664,N_49148,N_48590);
xnor UO_3665 (O_3665,N_49133,N_49888);
and UO_3666 (O_3666,N_49187,N_49180);
nand UO_3667 (O_3667,N_48148,N_49429);
xnor UO_3668 (O_3668,N_49318,N_48329);
or UO_3669 (O_3669,N_49371,N_49154);
xor UO_3670 (O_3670,N_48733,N_48538);
nand UO_3671 (O_3671,N_48719,N_48959);
and UO_3672 (O_3672,N_49351,N_48487);
nor UO_3673 (O_3673,N_49634,N_48119);
and UO_3674 (O_3674,N_48794,N_48960);
xnor UO_3675 (O_3675,N_49222,N_48836);
or UO_3676 (O_3676,N_48997,N_48622);
or UO_3677 (O_3677,N_48601,N_49460);
and UO_3678 (O_3678,N_49949,N_49597);
nand UO_3679 (O_3679,N_49754,N_49887);
or UO_3680 (O_3680,N_49159,N_48314);
nor UO_3681 (O_3681,N_48040,N_48720);
nand UO_3682 (O_3682,N_48125,N_49239);
nor UO_3683 (O_3683,N_48226,N_48618);
nor UO_3684 (O_3684,N_49393,N_48834);
xor UO_3685 (O_3685,N_49056,N_49724);
and UO_3686 (O_3686,N_49171,N_49519);
xnor UO_3687 (O_3687,N_49929,N_49741);
xor UO_3688 (O_3688,N_48739,N_49655);
nor UO_3689 (O_3689,N_49483,N_48161);
or UO_3690 (O_3690,N_49036,N_49363);
nand UO_3691 (O_3691,N_48908,N_49532);
or UO_3692 (O_3692,N_49508,N_49132);
nand UO_3693 (O_3693,N_49605,N_48023);
and UO_3694 (O_3694,N_48418,N_48426);
nor UO_3695 (O_3695,N_48071,N_49639);
and UO_3696 (O_3696,N_48421,N_49619);
nor UO_3697 (O_3697,N_49842,N_48771);
and UO_3698 (O_3698,N_49070,N_49706);
and UO_3699 (O_3699,N_49802,N_48972);
and UO_3700 (O_3700,N_48176,N_49312);
and UO_3701 (O_3701,N_48180,N_49836);
xnor UO_3702 (O_3702,N_49455,N_48541);
and UO_3703 (O_3703,N_49400,N_49908);
xor UO_3704 (O_3704,N_48292,N_49851);
nor UO_3705 (O_3705,N_48833,N_49339);
xnor UO_3706 (O_3706,N_48603,N_49401);
nand UO_3707 (O_3707,N_48347,N_49327);
nand UO_3708 (O_3708,N_49670,N_48454);
xor UO_3709 (O_3709,N_49947,N_49932);
or UO_3710 (O_3710,N_48432,N_48083);
xnor UO_3711 (O_3711,N_49980,N_49373);
xor UO_3712 (O_3712,N_49092,N_49516);
and UO_3713 (O_3713,N_48347,N_48914);
or UO_3714 (O_3714,N_49892,N_48860);
xor UO_3715 (O_3715,N_48068,N_49775);
or UO_3716 (O_3716,N_49476,N_49805);
and UO_3717 (O_3717,N_49921,N_49885);
nand UO_3718 (O_3718,N_49980,N_48958);
or UO_3719 (O_3719,N_49888,N_48926);
xnor UO_3720 (O_3720,N_48955,N_49224);
xnor UO_3721 (O_3721,N_48917,N_48178);
nor UO_3722 (O_3722,N_49408,N_48967);
nand UO_3723 (O_3723,N_49921,N_48033);
or UO_3724 (O_3724,N_49973,N_48857);
xor UO_3725 (O_3725,N_48206,N_49863);
nor UO_3726 (O_3726,N_48673,N_48202);
nand UO_3727 (O_3727,N_49543,N_49349);
nor UO_3728 (O_3728,N_49979,N_48626);
nor UO_3729 (O_3729,N_49334,N_49361);
and UO_3730 (O_3730,N_48260,N_48787);
nor UO_3731 (O_3731,N_49913,N_48221);
xnor UO_3732 (O_3732,N_49314,N_48997);
nand UO_3733 (O_3733,N_49496,N_49200);
nand UO_3734 (O_3734,N_48830,N_49386);
xor UO_3735 (O_3735,N_48305,N_49710);
nand UO_3736 (O_3736,N_48851,N_48771);
nand UO_3737 (O_3737,N_48507,N_49202);
nand UO_3738 (O_3738,N_49667,N_48272);
or UO_3739 (O_3739,N_49570,N_49993);
nor UO_3740 (O_3740,N_49940,N_48629);
or UO_3741 (O_3741,N_48873,N_49627);
and UO_3742 (O_3742,N_49492,N_48078);
nand UO_3743 (O_3743,N_49330,N_49723);
and UO_3744 (O_3744,N_48363,N_48741);
nor UO_3745 (O_3745,N_49340,N_48890);
and UO_3746 (O_3746,N_49533,N_48598);
or UO_3747 (O_3747,N_49546,N_49518);
and UO_3748 (O_3748,N_49670,N_49452);
xor UO_3749 (O_3749,N_48707,N_48150);
or UO_3750 (O_3750,N_48837,N_48563);
or UO_3751 (O_3751,N_48681,N_49896);
or UO_3752 (O_3752,N_49115,N_49855);
nand UO_3753 (O_3753,N_48403,N_48483);
and UO_3754 (O_3754,N_49813,N_48405);
and UO_3755 (O_3755,N_49954,N_49775);
nand UO_3756 (O_3756,N_49412,N_49206);
or UO_3757 (O_3757,N_49609,N_49180);
nand UO_3758 (O_3758,N_49073,N_48410);
nor UO_3759 (O_3759,N_48858,N_49388);
nor UO_3760 (O_3760,N_48337,N_49792);
or UO_3761 (O_3761,N_48633,N_48860);
and UO_3762 (O_3762,N_49037,N_48354);
nand UO_3763 (O_3763,N_48333,N_48628);
nand UO_3764 (O_3764,N_48346,N_48425);
nand UO_3765 (O_3765,N_49003,N_48594);
and UO_3766 (O_3766,N_49520,N_49165);
nor UO_3767 (O_3767,N_48182,N_48694);
xnor UO_3768 (O_3768,N_49092,N_49452);
xnor UO_3769 (O_3769,N_48982,N_49457);
nor UO_3770 (O_3770,N_48596,N_48707);
nand UO_3771 (O_3771,N_49908,N_48720);
or UO_3772 (O_3772,N_49636,N_48525);
or UO_3773 (O_3773,N_48935,N_48902);
nand UO_3774 (O_3774,N_48897,N_48839);
or UO_3775 (O_3775,N_48257,N_48427);
or UO_3776 (O_3776,N_48472,N_48892);
or UO_3777 (O_3777,N_49140,N_48742);
or UO_3778 (O_3778,N_48593,N_49790);
or UO_3779 (O_3779,N_48167,N_48423);
xnor UO_3780 (O_3780,N_49043,N_49842);
nand UO_3781 (O_3781,N_49085,N_48360);
xnor UO_3782 (O_3782,N_48924,N_49275);
and UO_3783 (O_3783,N_49148,N_49323);
or UO_3784 (O_3784,N_48305,N_49394);
nor UO_3785 (O_3785,N_49625,N_49249);
xnor UO_3786 (O_3786,N_49636,N_49036);
nand UO_3787 (O_3787,N_49970,N_49580);
or UO_3788 (O_3788,N_48013,N_48432);
nor UO_3789 (O_3789,N_49452,N_48946);
xor UO_3790 (O_3790,N_49361,N_48049);
nand UO_3791 (O_3791,N_48892,N_48668);
xor UO_3792 (O_3792,N_48197,N_48526);
nand UO_3793 (O_3793,N_49403,N_49960);
nor UO_3794 (O_3794,N_48949,N_49012);
nor UO_3795 (O_3795,N_49168,N_48969);
and UO_3796 (O_3796,N_48970,N_48775);
xnor UO_3797 (O_3797,N_48437,N_49408);
xnor UO_3798 (O_3798,N_49099,N_49531);
xor UO_3799 (O_3799,N_48052,N_48440);
or UO_3800 (O_3800,N_48290,N_48180);
xor UO_3801 (O_3801,N_48615,N_48598);
and UO_3802 (O_3802,N_48532,N_48478);
and UO_3803 (O_3803,N_48431,N_48037);
xnor UO_3804 (O_3804,N_49948,N_49553);
xnor UO_3805 (O_3805,N_48778,N_48314);
or UO_3806 (O_3806,N_48722,N_48416);
xnor UO_3807 (O_3807,N_48614,N_49665);
or UO_3808 (O_3808,N_48435,N_48854);
nor UO_3809 (O_3809,N_49388,N_49038);
and UO_3810 (O_3810,N_49831,N_49732);
or UO_3811 (O_3811,N_48932,N_48643);
nand UO_3812 (O_3812,N_48321,N_49756);
nand UO_3813 (O_3813,N_49499,N_49563);
nor UO_3814 (O_3814,N_48440,N_49371);
or UO_3815 (O_3815,N_48493,N_48627);
nand UO_3816 (O_3816,N_49237,N_48907);
xor UO_3817 (O_3817,N_49757,N_48400);
nor UO_3818 (O_3818,N_48605,N_48203);
nand UO_3819 (O_3819,N_49248,N_49195);
xnor UO_3820 (O_3820,N_49224,N_49059);
nand UO_3821 (O_3821,N_49110,N_49938);
and UO_3822 (O_3822,N_48488,N_49340);
and UO_3823 (O_3823,N_49754,N_49212);
and UO_3824 (O_3824,N_48345,N_49701);
or UO_3825 (O_3825,N_49406,N_49431);
and UO_3826 (O_3826,N_49119,N_48207);
nand UO_3827 (O_3827,N_49828,N_49480);
nor UO_3828 (O_3828,N_49015,N_48722);
xor UO_3829 (O_3829,N_48251,N_48998);
nand UO_3830 (O_3830,N_48298,N_49125);
nand UO_3831 (O_3831,N_49841,N_48333);
and UO_3832 (O_3832,N_49202,N_49145);
nand UO_3833 (O_3833,N_48118,N_49534);
nand UO_3834 (O_3834,N_48795,N_49292);
and UO_3835 (O_3835,N_48213,N_49887);
xnor UO_3836 (O_3836,N_49488,N_48359);
or UO_3837 (O_3837,N_48510,N_48847);
nor UO_3838 (O_3838,N_49635,N_49506);
xnor UO_3839 (O_3839,N_49608,N_48666);
nand UO_3840 (O_3840,N_48274,N_48021);
nor UO_3841 (O_3841,N_48126,N_48982);
nor UO_3842 (O_3842,N_49652,N_48731);
nor UO_3843 (O_3843,N_49602,N_49412);
or UO_3844 (O_3844,N_48072,N_48259);
nor UO_3845 (O_3845,N_48063,N_49022);
xor UO_3846 (O_3846,N_48425,N_49370);
and UO_3847 (O_3847,N_48961,N_49116);
nor UO_3848 (O_3848,N_48268,N_49475);
xnor UO_3849 (O_3849,N_48938,N_49579);
nor UO_3850 (O_3850,N_48768,N_48392);
or UO_3851 (O_3851,N_49486,N_48090);
nand UO_3852 (O_3852,N_48233,N_48681);
and UO_3853 (O_3853,N_49297,N_48056);
nand UO_3854 (O_3854,N_49211,N_49080);
nand UO_3855 (O_3855,N_49221,N_48188);
xor UO_3856 (O_3856,N_48170,N_49664);
or UO_3857 (O_3857,N_49052,N_48687);
or UO_3858 (O_3858,N_48721,N_48871);
nor UO_3859 (O_3859,N_49680,N_49252);
or UO_3860 (O_3860,N_49152,N_48483);
xnor UO_3861 (O_3861,N_49378,N_49076);
and UO_3862 (O_3862,N_49624,N_49462);
xor UO_3863 (O_3863,N_48445,N_48300);
xnor UO_3864 (O_3864,N_49476,N_49517);
xnor UO_3865 (O_3865,N_49768,N_48553);
nand UO_3866 (O_3866,N_48918,N_49466);
and UO_3867 (O_3867,N_49786,N_49113);
xor UO_3868 (O_3868,N_48435,N_49041);
nor UO_3869 (O_3869,N_49190,N_49552);
and UO_3870 (O_3870,N_48419,N_49226);
or UO_3871 (O_3871,N_49702,N_48821);
nor UO_3872 (O_3872,N_49484,N_49550);
nand UO_3873 (O_3873,N_49992,N_48638);
nor UO_3874 (O_3874,N_48519,N_48091);
or UO_3875 (O_3875,N_49585,N_48979);
nand UO_3876 (O_3876,N_48497,N_48015);
and UO_3877 (O_3877,N_48612,N_48973);
and UO_3878 (O_3878,N_49039,N_48189);
xnor UO_3879 (O_3879,N_49306,N_49124);
or UO_3880 (O_3880,N_48164,N_49863);
or UO_3881 (O_3881,N_48917,N_48939);
and UO_3882 (O_3882,N_49316,N_48304);
nand UO_3883 (O_3883,N_49803,N_49696);
or UO_3884 (O_3884,N_48362,N_49846);
xnor UO_3885 (O_3885,N_49189,N_49820);
or UO_3886 (O_3886,N_49618,N_48180);
xnor UO_3887 (O_3887,N_49216,N_48413);
xnor UO_3888 (O_3888,N_49420,N_49706);
xor UO_3889 (O_3889,N_48908,N_49551);
nand UO_3890 (O_3890,N_48642,N_48921);
nand UO_3891 (O_3891,N_48985,N_48227);
nor UO_3892 (O_3892,N_49812,N_48849);
xor UO_3893 (O_3893,N_49456,N_49610);
and UO_3894 (O_3894,N_49761,N_49391);
nor UO_3895 (O_3895,N_49061,N_48475);
xor UO_3896 (O_3896,N_49518,N_49692);
nand UO_3897 (O_3897,N_49877,N_49231);
nor UO_3898 (O_3898,N_48556,N_48246);
nor UO_3899 (O_3899,N_49899,N_48153);
nand UO_3900 (O_3900,N_49244,N_49966);
and UO_3901 (O_3901,N_48535,N_49354);
nor UO_3902 (O_3902,N_48746,N_48107);
and UO_3903 (O_3903,N_49410,N_49276);
nand UO_3904 (O_3904,N_48255,N_48411);
xnor UO_3905 (O_3905,N_48508,N_48489);
xor UO_3906 (O_3906,N_48593,N_49126);
nand UO_3907 (O_3907,N_48350,N_49106);
or UO_3908 (O_3908,N_49306,N_49840);
xor UO_3909 (O_3909,N_48860,N_48559);
and UO_3910 (O_3910,N_49123,N_49880);
nand UO_3911 (O_3911,N_48600,N_48499);
and UO_3912 (O_3912,N_49294,N_49396);
xor UO_3913 (O_3913,N_49765,N_48277);
xor UO_3914 (O_3914,N_48176,N_48873);
and UO_3915 (O_3915,N_48943,N_49237);
and UO_3916 (O_3916,N_48679,N_48892);
and UO_3917 (O_3917,N_49898,N_48206);
xor UO_3918 (O_3918,N_49302,N_49908);
or UO_3919 (O_3919,N_49075,N_49851);
nor UO_3920 (O_3920,N_48251,N_48430);
or UO_3921 (O_3921,N_48742,N_49460);
xnor UO_3922 (O_3922,N_49424,N_48534);
or UO_3923 (O_3923,N_48121,N_49465);
nor UO_3924 (O_3924,N_48250,N_49557);
nor UO_3925 (O_3925,N_49821,N_48149);
nand UO_3926 (O_3926,N_49167,N_49452);
and UO_3927 (O_3927,N_48235,N_49539);
or UO_3928 (O_3928,N_48578,N_49417);
nand UO_3929 (O_3929,N_49826,N_49522);
nand UO_3930 (O_3930,N_48913,N_48400);
or UO_3931 (O_3931,N_49248,N_49700);
xor UO_3932 (O_3932,N_48442,N_49918);
xor UO_3933 (O_3933,N_49164,N_48619);
and UO_3934 (O_3934,N_49391,N_48588);
nor UO_3935 (O_3935,N_49208,N_48980);
xor UO_3936 (O_3936,N_48500,N_49595);
or UO_3937 (O_3937,N_48043,N_49609);
and UO_3938 (O_3938,N_48431,N_49699);
nand UO_3939 (O_3939,N_48716,N_48866);
and UO_3940 (O_3940,N_49983,N_48699);
and UO_3941 (O_3941,N_49146,N_49391);
nand UO_3942 (O_3942,N_49101,N_49757);
nand UO_3943 (O_3943,N_48701,N_49463);
xnor UO_3944 (O_3944,N_49079,N_48195);
and UO_3945 (O_3945,N_49481,N_48343);
or UO_3946 (O_3946,N_49884,N_49979);
nand UO_3947 (O_3947,N_48815,N_48493);
xnor UO_3948 (O_3948,N_49023,N_48377);
nor UO_3949 (O_3949,N_48518,N_49189);
and UO_3950 (O_3950,N_49373,N_49754);
or UO_3951 (O_3951,N_49893,N_48763);
xnor UO_3952 (O_3952,N_48955,N_48791);
nor UO_3953 (O_3953,N_48556,N_48915);
xnor UO_3954 (O_3954,N_48001,N_49680);
xnor UO_3955 (O_3955,N_48897,N_49691);
or UO_3956 (O_3956,N_48824,N_48354);
or UO_3957 (O_3957,N_48300,N_49720);
and UO_3958 (O_3958,N_48260,N_48407);
and UO_3959 (O_3959,N_49558,N_48102);
xor UO_3960 (O_3960,N_49620,N_48331);
and UO_3961 (O_3961,N_48625,N_48137);
nor UO_3962 (O_3962,N_49922,N_49173);
nor UO_3963 (O_3963,N_48583,N_48081);
nand UO_3964 (O_3964,N_48867,N_49441);
or UO_3965 (O_3965,N_49871,N_49507);
nor UO_3966 (O_3966,N_48916,N_48385);
or UO_3967 (O_3967,N_48371,N_49863);
xor UO_3968 (O_3968,N_48911,N_49809);
xnor UO_3969 (O_3969,N_48269,N_48819);
nand UO_3970 (O_3970,N_49446,N_49920);
nor UO_3971 (O_3971,N_48032,N_48281);
nor UO_3972 (O_3972,N_49788,N_48129);
or UO_3973 (O_3973,N_48881,N_49010);
xnor UO_3974 (O_3974,N_48558,N_49372);
and UO_3975 (O_3975,N_48512,N_48133);
or UO_3976 (O_3976,N_49198,N_48491);
or UO_3977 (O_3977,N_49257,N_49755);
xnor UO_3978 (O_3978,N_49933,N_48750);
nor UO_3979 (O_3979,N_49528,N_48324);
or UO_3980 (O_3980,N_49548,N_49037);
and UO_3981 (O_3981,N_49475,N_48483);
nand UO_3982 (O_3982,N_48299,N_49274);
or UO_3983 (O_3983,N_49350,N_49697);
xor UO_3984 (O_3984,N_48621,N_49965);
nor UO_3985 (O_3985,N_49461,N_49436);
and UO_3986 (O_3986,N_49315,N_48196);
or UO_3987 (O_3987,N_48045,N_48750);
nand UO_3988 (O_3988,N_49918,N_48571);
and UO_3989 (O_3989,N_48163,N_49782);
nor UO_3990 (O_3990,N_48776,N_48271);
xnor UO_3991 (O_3991,N_49118,N_48855);
or UO_3992 (O_3992,N_49737,N_48927);
xor UO_3993 (O_3993,N_48755,N_48643);
xnor UO_3994 (O_3994,N_48922,N_49712);
and UO_3995 (O_3995,N_48445,N_48319);
and UO_3996 (O_3996,N_49949,N_48849);
and UO_3997 (O_3997,N_48732,N_48398);
or UO_3998 (O_3998,N_48274,N_49400);
or UO_3999 (O_3999,N_49486,N_48693);
nor UO_4000 (O_4000,N_48837,N_48213);
nand UO_4001 (O_4001,N_48576,N_49954);
and UO_4002 (O_4002,N_49625,N_48892);
or UO_4003 (O_4003,N_48646,N_49499);
or UO_4004 (O_4004,N_49826,N_48687);
and UO_4005 (O_4005,N_48148,N_48284);
xnor UO_4006 (O_4006,N_49070,N_49172);
nor UO_4007 (O_4007,N_49913,N_49675);
nand UO_4008 (O_4008,N_48747,N_48073);
nand UO_4009 (O_4009,N_48794,N_49334);
or UO_4010 (O_4010,N_48840,N_48218);
xnor UO_4011 (O_4011,N_48974,N_49982);
or UO_4012 (O_4012,N_49515,N_49880);
nor UO_4013 (O_4013,N_48417,N_48166);
nand UO_4014 (O_4014,N_49772,N_49244);
xor UO_4015 (O_4015,N_48985,N_48640);
and UO_4016 (O_4016,N_49334,N_48253);
xor UO_4017 (O_4017,N_49251,N_48576);
nor UO_4018 (O_4018,N_48322,N_48478);
and UO_4019 (O_4019,N_48829,N_48404);
xor UO_4020 (O_4020,N_49908,N_49602);
and UO_4021 (O_4021,N_48924,N_49815);
or UO_4022 (O_4022,N_48233,N_49314);
nor UO_4023 (O_4023,N_49621,N_49371);
nand UO_4024 (O_4024,N_49044,N_48269);
nor UO_4025 (O_4025,N_48371,N_49303);
xor UO_4026 (O_4026,N_48369,N_49053);
nor UO_4027 (O_4027,N_48823,N_49217);
nand UO_4028 (O_4028,N_48699,N_48092);
or UO_4029 (O_4029,N_48272,N_49583);
nand UO_4030 (O_4030,N_48658,N_48017);
nand UO_4031 (O_4031,N_48151,N_48885);
nor UO_4032 (O_4032,N_49904,N_48485);
nor UO_4033 (O_4033,N_48706,N_49452);
nor UO_4034 (O_4034,N_49152,N_49261);
nand UO_4035 (O_4035,N_48901,N_48223);
and UO_4036 (O_4036,N_49139,N_48368);
nor UO_4037 (O_4037,N_48031,N_48824);
nor UO_4038 (O_4038,N_48920,N_49950);
xor UO_4039 (O_4039,N_48216,N_48418);
nand UO_4040 (O_4040,N_49291,N_49224);
xnor UO_4041 (O_4041,N_49941,N_49280);
nor UO_4042 (O_4042,N_48806,N_49690);
and UO_4043 (O_4043,N_48955,N_49407);
nand UO_4044 (O_4044,N_48507,N_49028);
and UO_4045 (O_4045,N_49626,N_49506);
or UO_4046 (O_4046,N_48550,N_48131);
nor UO_4047 (O_4047,N_48969,N_49028);
or UO_4048 (O_4048,N_48742,N_48992);
or UO_4049 (O_4049,N_49636,N_48921);
nor UO_4050 (O_4050,N_48396,N_48845);
or UO_4051 (O_4051,N_49015,N_48125);
nor UO_4052 (O_4052,N_48732,N_49260);
or UO_4053 (O_4053,N_49727,N_49177);
and UO_4054 (O_4054,N_48728,N_48415);
nor UO_4055 (O_4055,N_48950,N_48996);
and UO_4056 (O_4056,N_49353,N_48753);
or UO_4057 (O_4057,N_48280,N_49847);
nand UO_4058 (O_4058,N_48102,N_48057);
and UO_4059 (O_4059,N_49438,N_48561);
xor UO_4060 (O_4060,N_48169,N_48345);
nor UO_4061 (O_4061,N_48532,N_49440);
xor UO_4062 (O_4062,N_49462,N_49597);
nor UO_4063 (O_4063,N_48134,N_49861);
nor UO_4064 (O_4064,N_48152,N_48377);
nand UO_4065 (O_4065,N_49336,N_49264);
nand UO_4066 (O_4066,N_48269,N_48219);
nor UO_4067 (O_4067,N_49238,N_49249);
xnor UO_4068 (O_4068,N_48919,N_48901);
xnor UO_4069 (O_4069,N_49591,N_48196);
or UO_4070 (O_4070,N_49740,N_49313);
xor UO_4071 (O_4071,N_49075,N_48975);
xnor UO_4072 (O_4072,N_48521,N_49594);
nor UO_4073 (O_4073,N_49383,N_48920);
and UO_4074 (O_4074,N_48928,N_48039);
and UO_4075 (O_4075,N_49148,N_49007);
nor UO_4076 (O_4076,N_48869,N_48084);
nand UO_4077 (O_4077,N_49535,N_49236);
nand UO_4078 (O_4078,N_48448,N_48210);
or UO_4079 (O_4079,N_49602,N_49401);
nand UO_4080 (O_4080,N_49592,N_49411);
and UO_4081 (O_4081,N_49233,N_48325);
and UO_4082 (O_4082,N_49002,N_48799);
or UO_4083 (O_4083,N_48601,N_49868);
or UO_4084 (O_4084,N_48422,N_49625);
and UO_4085 (O_4085,N_48299,N_48872);
or UO_4086 (O_4086,N_48829,N_49371);
and UO_4087 (O_4087,N_48064,N_48954);
nor UO_4088 (O_4088,N_49511,N_48553);
and UO_4089 (O_4089,N_48872,N_49941);
xnor UO_4090 (O_4090,N_48412,N_48429);
xor UO_4091 (O_4091,N_49307,N_48240);
and UO_4092 (O_4092,N_49105,N_49889);
nand UO_4093 (O_4093,N_49205,N_49789);
and UO_4094 (O_4094,N_48731,N_48056);
nand UO_4095 (O_4095,N_48644,N_49173);
or UO_4096 (O_4096,N_48091,N_49296);
nand UO_4097 (O_4097,N_48549,N_48198);
and UO_4098 (O_4098,N_49955,N_49596);
xor UO_4099 (O_4099,N_49060,N_49130);
nand UO_4100 (O_4100,N_49425,N_48289);
nand UO_4101 (O_4101,N_49336,N_49802);
nand UO_4102 (O_4102,N_49184,N_48905);
nand UO_4103 (O_4103,N_48516,N_48827);
xor UO_4104 (O_4104,N_49980,N_49689);
xor UO_4105 (O_4105,N_49647,N_48992);
nor UO_4106 (O_4106,N_49119,N_49136);
or UO_4107 (O_4107,N_48521,N_48852);
nand UO_4108 (O_4108,N_48824,N_49219);
nand UO_4109 (O_4109,N_49909,N_49937);
and UO_4110 (O_4110,N_49700,N_48369);
or UO_4111 (O_4111,N_49685,N_49606);
nand UO_4112 (O_4112,N_49073,N_48116);
or UO_4113 (O_4113,N_49442,N_48677);
nor UO_4114 (O_4114,N_49655,N_48227);
nand UO_4115 (O_4115,N_48933,N_49128);
nor UO_4116 (O_4116,N_48193,N_49316);
and UO_4117 (O_4117,N_48245,N_48647);
nor UO_4118 (O_4118,N_48265,N_48959);
or UO_4119 (O_4119,N_48778,N_48680);
nand UO_4120 (O_4120,N_48401,N_48939);
xor UO_4121 (O_4121,N_49014,N_49248);
and UO_4122 (O_4122,N_49500,N_49705);
or UO_4123 (O_4123,N_49210,N_48144);
xor UO_4124 (O_4124,N_48799,N_48723);
nand UO_4125 (O_4125,N_49553,N_49956);
and UO_4126 (O_4126,N_48088,N_49134);
nor UO_4127 (O_4127,N_49843,N_48591);
or UO_4128 (O_4128,N_48891,N_49115);
nor UO_4129 (O_4129,N_48328,N_49931);
xnor UO_4130 (O_4130,N_49194,N_49297);
xnor UO_4131 (O_4131,N_48922,N_49400);
or UO_4132 (O_4132,N_49673,N_48193);
xnor UO_4133 (O_4133,N_49112,N_48620);
and UO_4134 (O_4134,N_49228,N_48046);
xnor UO_4135 (O_4135,N_48438,N_48592);
nor UO_4136 (O_4136,N_48910,N_49808);
and UO_4137 (O_4137,N_49552,N_48718);
xnor UO_4138 (O_4138,N_48056,N_49891);
or UO_4139 (O_4139,N_49564,N_48402);
or UO_4140 (O_4140,N_48683,N_48201);
nand UO_4141 (O_4141,N_49014,N_49468);
or UO_4142 (O_4142,N_49044,N_49082);
nand UO_4143 (O_4143,N_49471,N_48338);
and UO_4144 (O_4144,N_49846,N_48250);
xnor UO_4145 (O_4145,N_49510,N_49850);
nor UO_4146 (O_4146,N_48777,N_48624);
and UO_4147 (O_4147,N_49125,N_48786);
or UO_4148 (O_4148,N_49881,N_49664);
xnor UO_4149 (O_4149,N_48661,N_49337);
xor UO_4150 (O_4150,N_49233,N_49033);
xor UO_4151 (O_4151,N_49097,N_49557);
and UO_4152 (O_4152,N_48920,N_48278);
xor UO_4153 (O_4153,N_48486,N_49781);
or UO_4154 (O_4154,N_48224,N_48028);
and UO_4155 (O_4155,N_48019,N_48688);
or UO_4156 (O_4156,N_49019,N_49153);
nor UO_4157 (O_4157,N_49052,N_48844);
nand UO_4158 (O_4158,N_49575,N_49065);
xnor UO_4159 (O_4159,N_49860,N_48143);
xor UO_4160 (O_4160,N_49088,N_49792);
nand UO_4161 (O_4161,N_49094,N_48799);
and UO_4162 (O_4162,N_48009,N_48984);
or UO_4163 (O_4163,N_49809,N_48963);
nand UO_4164 (O_4164,N_48344,N_49684);
and UO_4165 (O_4165,N_48814,N_48888);
and UO_4166 (O_4166,N_49937,N_49438);
or UO_4167 (O_4167,N_49654,N_48152);
xnor UO_4168 (O_4168,N_49044,N_48992);
and UO_4169 (O_4169,N_48082,N_49279);
nand UO_4170 (O_4170,N_48521,N_49105);
nor UO_4171 (O_4171,N_49329,N_49847);
or UO_4172 (O_4172,N_48261,N_48317);
nor UO_4173 (O_4173,N_49000,N_48629);
nand UO_4174 (O_4174,N_49643,N_49808);
and UO_4175 (O_4175,N_49820,N_49888);
and UO_4176 (O_4176,N_48923,N_49620);
or UO_4177 (O_4177,N_49184,N_48902);
or UO_4178 (O_4178,N_49147,N_48467);
and UO_4179 (O_4179,N_49681,N_49766);
nor UO_4180 (O_4180,N_49326,N_48562);
and UO_4181 (O_4181,N_49726,N_49340);
or UO_4182 (O_4182,N_49196,N_49247);
or UO_4183 (O_4183,N_49859,N_49791);
xnor UO_4184 (O_4184,N_48754,N_48619);
xor UO_4185 (O_4185,N_49097,N_48355);
nor UO_4186 (O_4186,N_48846,N_48723);
xnor UO_4187 (O_4187,N_48648,N_48847);
nand UO_4188 (O_4188,N_48093,N_48008);
xor UO_4189 (O_4189,N_49201,N_49570);
or UO_4190 (O_4190,N_49272,N_48978);
nand UO_4191 (O_4191,N_48805,N_48628);
and UO_4192 (O_4192,N_48613,N_48162);
and UO_4193 (O_4193,N_48661,N_48565);
and UO_4194 (O_4194,N_49085,N_49573);
nand UO_4195 (O_4195,N_48609,N_49418);
xnor UO_4196 (O_4196,N_49146,N_48301);
nand UO_4197 (O_4197,N_48108,N_48623);
nor UO_4198 (O_4198,N_49628,N_49443);
xnor UO_4199 (O_4199,N_48094,N_49409);
nand UO_4200 (O_4200,N_49932,N_48029);
xor UO_4201 (O_4201,N_49025,N_48136);
and UO_4202 (O_4202,N_48442,N_48568);
or UO_4203 (O_4203,N_49650,N_49334);
nor UO_4204 (O_4204,N_48691,N_49875);
nand UO_4205 (O_4205,N_49696,N_49845);
and UO_4206 (O_4206,N_49479,N_48929);
nor UO_4207 (O_4207,N_48112,N_48993);
and UO_4208 (O_4208,N_48517,N_49662);
nor UO_4209 (O_4209,N_48706,N_49835);
nor UO_4210 (O_4210,N_49072,N_49059);
and UO_4211 (O_4211,N_49740,N_48636);
or UO_4212 (O_4212,N_49996,N_48764);
nand UO_4213 (O_4213,N_48044,N_49319);
or UO_4214 (O_4214,N_49171,N_49531);
or UO_4215 (O_4215,N_48573,N_49031);
nand UO_4216 (O_4216,N_48091,N_49011);
nand UO_4217 (O_4217,N_48353,N_49174);
xor UO_4218 (O_4218,N_48955,N_48075);
xor UO_4219 (O_4219,N_48919,N_49782);
xnor UO_4220 (O_4220,N_49149,N_49560);
and UO_4221 (O_4221,N_49015,N_49143);
xor UO_4222 (O_4222,N_48040,N_49986);
or UO_4223 (O_4223,N_48659,N_48354);
or UO_4224 (O_4224,N_49020,N_48133);
xor UO_4225 (O_4225,N_49364,N_49046);
nor UO_4226 (O_4226,N_49624,N_48551);
and UO_4227 (O_4227,N_49232,N_49472);
or UO_4228 (O_4228,N_48350,N_49361);
or UO_4229 (O_4229,N_49877,N_49075);
or UO_4230 (O_4230,N_49030,N_49834);
or UO_4231 (O_4231,N_49822,N_49341);
xnor UO_4232 (O_4232,N_48373,N_49413);
xnor UO_4233 (O_4233,N_48497,N_48068);
or UO_4234 (O_4234,N_49837,N_49461);
or UO_4235 (O_4235,N_49978,N_48898);
and UO_4236 (O_4236,N_48448,N_48588);
or UO_4237 (O_4237,N_48899,N_48490);
xor UO_4238 (O_4238,N_49271,N_48390);
xnor UO_4239 (O_4239,N_49353,N_48910);
or UO_4240 (O_4240,N_48844,N_49996);
or UO_4241 (O_4241,N_49203,N_48705);
or UO_4242 (O_4242,N_48659,N_49679);
nand UO_4243 (O_4243,N_49150,N_49862);
xor UO_4244 (O_4244,N_48313,N_49914);
or UO_4245 (O_4245,N_49659,N_48582);
and UO_4246 (O_4246,N_49536,N_49297);
nor UO_4247 (O_4247,N_48032,N_48368);
or UO_4248 (O_4248,N_49876,N_48227);
nand UO_4249 (O_4249,N_48283,N_48655);
or UO_4250 (O_4250,N_48471,N_49753);
xnor UO_4251 (O_4251,N_49801,N_49314);
and UO_4252 (O_4252,N_48092,N_49135);
and UO_4253 (O_4253,N_49659,N_49516);
or UO_4254 (O_4254,N_48242,N_48751);
nor UO_4255 (O_4255,N_49590,N_49760);
xor UO_4256 (O_4256,N_49302,N_48548);
xnor UO_4257 (O_4257,N_48065,N_49537);
nor UO_4258 (O_4258,N_49910,N_48478);
and UO_4259 (O_4259,N_49875,N_48755);
nor UO_4260 (O_4260,N_49486,N_49289);
nand UO_4261 (O_4261,N_48523,N_49297);
and UO_4262 (O_4262,N_49332,N_49196);
nand UO_4263 (O_4263,N_48319,N_48377);
nor UO_4264 (O_4264,N_49171,N_49285);
nor UO_4265 (O_4265,N_49605,N_48012);
nand UO_4266 (O_4266,N_48285,N_49423);
or UO_4267 (O_4267,N_49746,N_48073);
nand UO_4268 (O_4268,N_49331,N_48662);
and UO_4269 (O_4269,N_49091,N_48393);
or UO_4270 (O_4270,N_48564,N_48870);
nand UO_4271 (O_4271,N_48195,N_48708);
or UO_4272 (O_4272,N_48721,N_48781);
xnor UO_4273 (O_4273,N_48325,N_49011);
xor UO_4274 (O_4274,N_49123,N_48604);
and UO_4275 (O_4275,N_49576,N_49806);
nand UO_4276 (O_4276,N_48238,N_49221);
and UO_4277 (O_4277,N_49017,N_48799);
nor UO_4278 (O_4278,N_49122,N_48825);
nor UO_4279 (O_4279,N_49729,N_49958);
nand UO_4280 (O_4280,N_48892,N_49201);
or UO_4281 (O_4281,N_48508,N_48313);
xor UO_4282 (O_4282,N_49780,N_48821);
or UO_4283 (O_4283,N_48796,N_49438);
xor UO_4284 (O_4284,N_49832,N_48842);
and UO_4285 (O_4285,N_48701,N_49367);
nand UO_4286 (O_4286,N_49462,N_48917);
nand UO_4287 (O_4287,N_48513,N_48624);
xor UO_4288 (O_4288,N_49018,N_48883);
and UO_4289 (O_4289,N_49702,N_49275);
nor UO_4290 (O_4290,N_49191,N_49823);
or UO_4291 (O_4291,N_49355,N_49671);
xnor UO_4292 (O_4292,N_48882,N_48178);
and UO_4293 (O_4293,N_48508,N_48572);
or UO_4294 (O_4294,N_49355,N_48864);
nand UO_4295 (O_4295,N_49250,N_49384);
nor UO_4296 (O_4296,N_49948,N_49837);
and UO_4297 (O_4297,N_49532,N_48415);
nand UO_4298 (O_4298,N_49097,N_49854);
nor UO_4299 (O_4299,N_48332,N_49382);
nand UO_4300 (O_4300,N_48469,N_48322);
and UO_4301 (O_4301,N_48783,N_49415);
and UO_4302 (O_4302,N_48052,N_49673);
nor UO_4303 (O_4303,N_49382,N_48396);
or UO_4304 (O_4304,N_49438,N_48719);
nor UO_4305 (O_4305,N_48649,N_48103);
or UO_4306 (O_4306,N_48160,N_49466);
or UO_4307 (O_4307,N_49928,N_49348);
xnor UO_4308 (O_4308,N_48303,N_48020);
nand UO_4309 (O_4309,N_49131,N_49786);
nor UO_4310 (O_4310,N_49638,N_48895);
and UO_4311 (O_4311,N_48889,N_48683);
xor UO_4312 (O_4312,N_48258,N_48276);
xnor UO_4313 (O_4313,N_49647,N_48360);
or UO_4314 (O_4314,N_49979,N_49591);
or UO_4315 (O_4315,N_48896,N_48715);
or UO_4316 (O_4316,N_48085,N_48743);
and UO_4317 (O_4317,N_48201,N_48497);
nand UO_4318 (O_4318,N_48345,N_49215);
nor UO_4319 (O_4319,N_48946,N_49373);
and UO_4320 (O_4320,N_49906,N_48778);
nand UO_4321 (O_4321,N_49944,N_48390);
nor UO_4322 (O_4322,N_48170,N_48461);
and UO_4323 (O_4323,N_49421,N_49141);
or UO_4324 (O_4324,N_48482,N_49371);
nand UO_4325 (O_4325,N_48146,N_49818);
or UO_4326 (O_4326,N_48757,N_49645);
and UO_4327 (O_4327,N_49617,N_48196);
nor UO_4328 (O_4328,N_49107,N_48870);
or UO_4329 (O_4329,N_48022,N_49804);
or UO_4330 (O_4330,N_49739,N_49197);
nand UO_4331 (O_4331,N_49307,N_49277);
nand UO_4332 (O_4332,N_49555,N_49104);
and UO_4333 (O_4333,N_48001,N_48473);
nand UO_4334 (O_4334,N_48883,N_49394);
nor UO_4335 (O_4335,N_49487,N_49821);
or UO_4336 (O_4336,N_48320,N_49748);
nand UO_4337 (O_4337,N_49930,N_49808);
nor UO_4338 (O_4338,N_48241,N_48997);
xnor UO_4339 (O_4339,N_49216,N_48244);
nor UO_4340 (O_4340,N_49912,N_49371);
and UO_4341 (O_4341,N_48409,N_48976);
nor UO_4342 (O_4342,N_49264,N_49282);
and UO_4343 (O_4343,N_48211,N_48447);
or UO_4344 (O_4344,N_49548,N_49095);
or UO_4345 (O_4345,N_49633,N_48054);
nor UO_4346 (O_4346,N_49568,N_49233);
and UO_4347 (O_4347,N_48194,N_49470);
xor UO_4348 (O_4348,N_48350,N_49572);
nand UO_4349 (O_4349,N_49230,N_49682);
and UO_4350 (O_4350,N_48293,N_48111);
and UO_4351 (O_4351,N_48158,N_48632);
or UO_4352 (O_4352,N_49842,N_48071);
and UO_4353 (O_4353,N_49671,N_49857);
nor UO_4354 (O_4354,N_48375,N_48070);
xnor UO_4355 (O_4355,N_48399,N_48210);
nand UO_4356 (O_4356,N_49928,N_48157);
nand UO_4357 (O_4357,N_48427,N_49376);
and UO_4358 (O_4358,N_48620,N_49693);
and UO_4359 (O_4359,N_49017,N_48276);
xnor UO_4360 (O_4360,N_49590,N_49499);
nand UO_4361 (O_4361,N_49372,N_49157);
and UO_4362 (O_4362,N_49708,N_48468);
nor UO_4363 (O_4363,N_48813,N_48907);
and UO_4364 (O_4364,N_49944,N_49060);
nor UO_4365 (O_4365,N_49552,N_48890);
nand UO_4366 (O_4366,N_48081,N_48115);
nor UO_4367 (O_4367,N_48783,N_49006);
and UO_4368 (O_4368,N_49845,N_49780);
and UO_4369 (O_4369,N_49681,N_48909);
and UO_4370 (O_4370,N_49443,N_48668);
nand UO_4371 (O_4371,N_49564,N_48780);
nor UO_4372 (O_4372,N_49840,N_48545);
and UO_4373 (O_4373,N_48934,N_49059);
nand UO_4374 (O_4374,N_48297,N_49018);
nor UO_4375 (O_4375,N_48518,N_49345);
nand UO_4376 (O_4376,N_48979,N_48613);
or UO_4377 (O_4377,N_49392,N_48052);
nor UO_4378 (O_4378,N_49690,N_48862);
xor UO_4379 (O_4379,N_49306,N_48957);
nor UO_4380 (O_4380,N_48650,N_49231);
or UO_4381 (O_4381,N_48933,N_48007);
or UO_4382 (O_4382,N_48143,N_48883);
xor UO_4383 (O_4383,N_49466,N_48247);
or UO_4384 (O_4384,N_49808,N_49842);
nor UO_4385 (O_4385,N_49526,N_48346);
and UO_4386 (O_4386,N_49467,N_48548);
nor UO_4387 (O_4387,N_49728,N_49846);
or UO_4388 (O_4388,N_49877,N_48722);
nand UO_4389 (O_4389,N_49767,N_49244);
nand UO_4390 (O_4390,N_48671,N_48790);
nand UO_4391 (O_4391,N_48081,N_49728);
xnor UO_4392 (O_4392,N_49810,N_49857);
nand UO_4393 (O_4393,N_49284,N_48212);
and UO_4394 (O_4394,N_48461,N_48388);
and UO_4395 (O_4395,N_49316,N_49027);
nor UO_4396 (O_4396,N_49943,N_48400);
nor UO_4397 (O_4397,N_48163,N_49090);
xnor UO_4398 (O_4398,N_48202,N_48363);
nor UO_4399 (O_4399,N_48389,N_49023);
xnor UO_4400 (O_4400,N_49638,N_48428);
nor UO_4401 (O_4401,N_48372,N_48414);
or UO_4402 (O_4402,N_48529,N_49427);
and UO_4403 (O_4403,N_49914,N_48973);
xor UO_4404 (O_4404,N_48017,N_48147);
or UO_4405 (O_4405,N_49745,N_48904);
nor UO_4406 (O_4406,N_49978,N_49692);
or UO_4407 (O_4407,N_49987,N_49304);
or UO_4408 (O_4408,N_48024,N_48120);
and UO_4409 (O_4409,N_48336,N_48840);
nor UO_4410 (O_4410,N_48729,N_49024);
nor UO_4411 (O_4411,N_49479,N_48637);
nor UO_4412 (O_4412,N_48524,N_49496);
nor UO_4413 (O_4413,N_49411,N_49365);
or UO_4414 (O_4414,N_49625,N_48804);
and UO_4415 (O_4415,N_48288,N_48435);
nor UO_4416 (O_4416,N_48670,N_48097);
and UO_4417 (O_4417,N_48070,N_49318);
xnor UO_4418 (O_4418,N_48023,N_49322);
xor UO_4419 (O_4419,N_48425,N_49866);
xnor UO_4420 (O_4420,N_48358,N_48627);
xor UO_4421 (O_4421,N_48721,N_49244);
and UO_4422 (O_4422,N_49683,N_49134);
and UO_4423 (O_4423,N_49019,N_49533);
nand UO_4424 (O_4424,N_49674,N_49959);
or UO_4425 (O_4425,N_49085,N_49655);
or UO_4426 (O_4426,N_49755,N_49042);
xor UO_4427 (O_4427,N_49761,N_48612);
nor UO_4428 (O_4428,N_48605,N_48279);
nand UO_4429 (O_4429,N_49152,N_48056);
and UO_4430 (O_4430,N_48544,N_49165);
or UO_4431 (O_4431,N_49206,N_49918);
and UO_4432 (O_4432,N_49850,N_48687);
and UO_4433 (O_4433,N_49031,N_48649);
nand UO_4434 (O_4434,N_49313,N_49486);
nand UO_4435 (O_4435,N_49414,N_48144);
and UO_4436 (O_4436,N_48743,N_49328);
xor UO_4437 (O_4437,N_48777,N_49688);
and UO_4438 (O_4438,N_48096,N_48021);
or UO_4439 (O_4439,N_48970,N_49700);
xor UO_4440 (O_4440,N_48529,N_49131);
or UO_4441 (O_4441,N_48016,N_48993);
and UO_4442 (O_4442,N_48954,N_49537);
xnor UO_4443 (O_4443,N_49997,N_49906);
or UO_4444 (O_4444,N_49131,N_49725);
xnor UO_4445 (O_4445,N_48107,N_48251);
xnor UO_4446 (O_4446,N_49660,N_49585);
and UO_4447 (O_4447,N_48907,N_49640);
or UO_4448 (O_4448,N_48409,N_49723);
nand UO_4449 (O_4449,N_48686,N_48255);
and UO_4450 (O_4450,N_48385,N_49176);
nand UO_4451 (O_4451,N_49961,N_49934);
or UO_4452 (O_4452,N_49557,N_49886);
nand UO_4453 (O_4453,N_48701,N_49964);
xor UO_4454 (O_4454,N_49413,N_49600);
nand UO_4455 (O_4455,N_48052,N_48986);
and UO_4456 (O_4456,N_49006,N_48525);
nor UO_4457 (O_4457,N_49192,N_49611);
and UO_4458 (O_4458,N_48434,N_48952);
and UO_4459 (O_4459,N_48654,N_49503);
xor UO_4460 (O_4460,N_49736,N_49354);
and UO_4461 (O_4461,N_49294,N_48995);
xor UO_4462 (O_4462,N_49016,N_49044);
or UO_4463 (O_4463,N_48027,N_48927);
or UO_4464 (O_4464,N_49471,N_48575);
and UO_4465 (O_4465,N_49078,N_48817);
or UO_4466 (O_4466,N_48808,N_48795);
xnor UO_4467 (O_4467,N_48160,N_48471);
xor UO_4468 (O_4468,N_49849,N_49638);
or UO_4469 (O_4469,N_48562,N_48191);
nor UO_4470 (O_4470,N_48696,N_48962);
xnor UO_4471 (O_4471,N_49475,N_49102);
xor UO_4472 (O_4472,N_48572,N_49321);
and UO_4473 (O_4473,N_49599,N_48193);
and UO_4474 (O_4474,N_48497,N_49896);
nand UO_4475 (O_4475,N_49577,N_48133);
nand UO_4476 (O_4476,N_49186,N_48826);
and UO_4477 (O_4477,N_49001,N_48494);
or UO_4478 (O_4478,N_49325,N_49861);
nand UO_4479 (O_4479,N_48945,N_48151);
nor UO_4480 (O_4480,N_49125,N_49616);
nor UO_4481 (O_4481,N_49205,N_48728);
nand UO_4482 (O_4482,N_48742,N_48481);
xor UO_4483 (O_4483,N_49495,N_48779);
nor UO_4484 (O_4484,N_49754,N_48860);
or UO_4485 (O_4485,N_49707,N_48406);
and UO_4486 (O_4486,N_48291,N_48136);
nand UO_4487 (O_4487,N_48765,N_49789);
or UO_4488 (O_4488,N_49958,N_49883);
nor UO_4489 (O_4489,N_48933,N_48305);
nor UO_4490 (O_4490,N_49114,N_49894);
nand UO_4491 (O_4491,N_49444,N_48488);
and UO_4492 (O_4492,N_48413,N_49997);
nand UO_4493 (O_4493,N_49526,N_49511);
or UO_4494 (O_4494,N_48145,N_49376);
nor UO_4495 (O_4495,N_48899,N_49404);
or UO_4496 (O_4496,N_48688,N_49100);
nor UO_4497 (O_4497,N_48098,N_48763);
nand UO_4498 (O_4498,N_48656,N_49031);
xnor UO_4499 (O_4499,N_49588,N_48590);
xor UO_4500 (O_4500,N_49872,N_48894);
nand UO_4501 (O_4501,N_49931,N_49563);
xor UO_4502 (O_4502,N_48126,N_49268);
nand UO_4503 (O_4503,N_49308,N_48706);
xnor UO_4504 (O_4504,N_48982,N_49757);
nand UO_4505 (O_4505,N_49770,N_48821);
nor UO_4506 (O_4506,N_49200,N_49418);
or UO_4507 (O_4507,N_48761,N_49002);
or UO_4508 (O_4508,N_49719,N_48374);
xor UO_4509 (O_4509,N_48613,N_48155);
nand UO_4510 (O_4510,N_48938,N_48446);
xor UO_4511 (O_4511,N_49256,N_48938);
or UO_4512 (O_4512,N_49755,N_49100);
xor UO_4513 (O_4513,N_49129,N_48216);
nor UO_4514 (O_4514,N_48444,N_48272);
or UO_4515 (O_4515,N_48293,N_48542);
and UO_4516 (O_4516,N_48152,N_49950);
nand UO_4517 (O_4517,N_49983,N_49518);
or UO_4518 (O_4518,N_48471,N_48547);
xnor UO_4519 (O_4519,N_49558,N_49537);
nor UO_4520 (O_4520,N_48651,N_49974);
or UO_4521 (O_4521,N_48701,N_48443);
nor UO_4522 (O_4522,N_49419,N_48287);
nor UO_4523 (O_4523,N_49703,N_49302);
and UO_4524 (O_4524,N_49323,N_48076);
and UO_4525 (O_4525,N_48996,N_49408);
and UO_4526 (O_4526,N_48832,N_49933);
nor UO_4527 (O_4527,N_48468,N_49747);
xnor UO_4528 (O_4528,N_48651,N_48140);
nor UO_4529 (O_4529,N_49089,N_48079);
or UO_4530 (O_4530,N_48453,N_49187);
nand UO_4531 (O_4531,N_49300,N_48728);
and UO_4532 (O_4532,N_48192,N_48810);
and UO_4533 (O_4533,N_48852,N_49529);
and UO_4534 (O_4534,N_49526,N_49473);
nor UO_4535 (O_4535,N_48131,N_49733);
and UO_4536 (O_4536,N_49304,N_49403);
nand UO_4537 (O_4537,N_48701,N_48910);
and UO_4538 (O_4538,N_48404,N_49809);
nand UO_4539 (O_4539,N_49311,N_49955);
xnor UO_4540 (O_4540,N_48655,N_49851);
nand UO_4541 (O_4541,N_49141,N_48390);
xor UO_4542 (O_4542,N_49888,N_49121);
xnor UO_4543 (O_4543,N_49062,N_49191);
nor UO_4544 (O_4544,N_48539,N_49994);
xor UO_4545 (O_4545,N_48900,N_49223);
nor UO_4546 (O_4546,N_48343,N_48562);
nand UO_4547 (O_4547,N_48850,N_49541);
nand UO_4548 (O_4548,N_48309,N_48409);
nand UO_4549 (O_4549,N_49721,N_49250);
and UO_4550 (O_4550,N_48675,N_49818);
nand UO_4551 (O_4551,N_48379,N_48381);
and UO_4552 (O_4552,N_48199,N_49873);
xnor UO_4553 (O_4553,N_48836,N_49984);
or UO_4554 (O_4554,N_48138,N_49053);
or UO_4555 (O_4555,N_49801,N_48043);
nor UO_4556 (O_4556,N_48505,N_49152);
and UO_4557 (O_4557,N_49317,N_49458);
nand UO_4558 (O_4558,N_48176,N_48710);
or UO_4559 (O_4559,N_48169,N_48154);
or UO_4560 (O_4560,N_49632,N_48976);
xor UO_4561 (O_4561,N_48306,N_48427);
xnor UO_4562 (O_4562,N_49978,N_49395);
or UO_4563 (O_4563,N_49710,N_48943);
nor UO_4564 (O_4564,N_49566,N_49338);
or UO_4565 (O_4565,N_48603,N_48900);
nand UO_4566 (O_4566,N_49899,N_48019);
nand UO_4567 (O_4567,N_48952,N_48146);
nand UO_4568 (O_4568,N_49203,N_48302);
nand UO_4569 (O_4569,N_49818,N_49985);
and UO_4570 (O_4570,N_49824,N_49305);
or UO_4571 (O_4571,N_48971,N_49373);
or UO_4572 (O_4572,N_49104,N_49651);
or UO_4573 (O_4573,N_48776,N_48772);
nand UO_4574 (O_4574,N_49403,N_49286);
or UO_4575 (O_4575,N_49535,N_49759);
nand UO_4576 (O_4576,N_49548,N_49427);
nor UO_4577 (O_4577,N_49102,N_49397);
or UO_4578 (O_4578,N_49612,N_48681);
and UO_4579 (O_4579,N_49159,N_48583);
nor UO_4580 (O_4580,N_48506,N_49841);
and UO_4581 (O_4581,N_49350,N_48321);
or UO_4582 (O_4582,N_48817,N_49562);
or UO_4583 (O_4583,N_48746,N_48257);
nand UO_4584 (O_4584,N_48750,N_49608);
or UO_4585 (O_4585,N_49085,N_49352);
nand UO_4586 (O_4586,N_48431,N_49074);
and UO_4587 (O_4587,N_49468,N_48253);
xor UO_4588 (O_4588,N_48793,N_48513);
nand UO_4589 (O_4589,N_49010,N_49554);
nor UO_4590 (O_4590,N_49111,N_49364);
xnor UO_4591 (O_4591,N_49161,N_48739);
nand UO_4592 (O_4592,N_49746,N_48680);
nor UO_4593 (O_4593,N_48485,N_48040);
xor UO_4594 (O_4594,N_49963,N_48879);
and UO_4595 (O_4595,N_49259,N_48318);
or UO_4596 (O_4596,N_48875,N_48284);
xnor UO_4597 (O_4597,N_48531,N_49865);
nor UO_4598 (O_4598,N_49627,N_49286);
nand UO_4599 (O_4599,N_49646,N_48129);
xnor UO_4600 (O_4600,N_49288,N_49860);
nor UO_4601 (O_4601,N_49576,N_48760);
nor UO_4602 (O_4602,N_48344,N_48123);
and UO_4603 (O_4603,N_48961,N_48947);
xor UO_4604 (O_4604,N_49499,N_48159);
nand UO_4605 (O_4605,N_48468,N_48961);
and UO_4606 (O_4606,N_49448,N_48851);
nor UO_4607 (O_4607,N_48184,N_49760);
and UO_4608 (O_4608,N_49287,N_49367);
and UO_4609 (O_4609,N_48914,N_48195);
xnor UO_4610 (O_4610,N_48072,N_48750);
nand UO_4611 (O_4611,N_49338,N_49379);
xnor UO_4612 (O_4612,N_49439,N_49131);
nand UO_4613 (O_4613,N_48885,N_48518);
and UO_4614 (O_4614,N_49575,N_48956);
and UO_4615 (O_4615,N_48887,N_48976);
xnor UO_4616 (O_4616,N_49380,N_49482);
xnor UO_4617 (O_4617,N_48068,N_48977);
xnor UO_4618 (O_4618,N_49977,N_48411);
xor UO_4619 (O_4619,N_48854,N_48896);
or UO_4620 (O_4620,N_49676,N_48893);
nand UO_4621 (O_4621,N_49064,N_49041);
or UO_4622 (O_4622,N_48617,N_48230);
xnor UO_4623 (O_4623,N_49801,N_49264);
xnor UO_4624 (O_4624,N_48654,N_48742);
nor UO_4625 (O_4625,N_49059,N_48170);
xor UO_4626 (O_4626,N_48647,N_48373);
and UO_4627 (O_4627,N_48039,N_48666);
or UO_4628 (O_4628,N_49567,N_48955);
and UO_4629 (O_4629,N_48443,N_48976);
and UO_4630 (O_4630,N_49420,N_49054);
nor UO_4631 (O_4631,N_49545,N_48019);
and UO_4632 (O_4632,N_49482,N_49068);
nor UO_4633 (O_4633,N_48557,N_49654);
xnor UO_4634 (O_4634,N_48567,N_49111);
or UO_4635 (O_4635,N_48376,N_48572);
nand UO_4636 (O_4636,N_49294,N_48732);
xor UO_4637 (O_4637,N_49209,N_49956);
xor UO_4638 (O_4638,N_48554,N_49262);
nor UO_4639 (O_4639,N_48988,N_49307);
or UO_4640 (O_4640,N_49291,N_48638);
and UO_4641 (O_4641,N_48157,N_49374);
nand UO_4642 (O_4642,N_49947,N_49096);
nand UO_4643 (O_4643,N_48543,N_48665);
and UO_4644 (O_4644,N_49265,N_49953);
and UO_4645 (O_4645,N_48025,N_49165);
or UO_4646 (O_4646,N_48134,N_48287);
or UO_4647 (O_4647,N_48072,N_49857);
or UO_4648 (O_4648,N_49505,N_49122);
xor UO_4649 (O_4649,N_49658,N_48969);
and UO_4650 (O_4650,N_49802,N_48662);
nand UO_4651 (O_4651,N_49152,N_49164);
xnor UO_4652 (O_4652,N_49008,N_49973);
and UO_4653 (O_4653,N_48084,N_49044);
nor UO_4654 (O_4654,N_48092,N_48430);
xor UO_4655 (O_4655,N_48551,N_48532);
xor UO_4656 (O_4656,N_48919,N_49038);
or UO_4657 (O_4657,N_49600,N_48716);
or UO_4658 (O_4658,N_49009,N_48500);
and UO_4659 (O_4659,N_49196,N_48486);
xnor UO_4660 (O_4660,N_49364,N_49619);
and UO_4661 (O_4661,N_48313,N_49601);
nand UO_4662 (O_4662,N_49270,N_49195);
nand UO_4663 (O_4663,N_49416,N_49301);
and UO_4664 (O_4664,N_48354,N_48439);
nor UO_4665 (O_4665,N_48041,N_48527);
nand UO_4666 (O_4666,N_48780,N_49780);
xor UO_4667 (O_4667,N_49301,N_48031);
and UO_4668 (O_4668,N_49046,N_49222);
xor UO_4669 (O_4669,N_48457,N_49683);
and UO_4670 (O_4670,N_48861,N_49285);
nand UO_4671 (O_4671,N_49264,N_49117);
nand UO_4672 (O_4672,N_48518,N_49297);
nand UO_4673 (O_4673,N_48744,N_49153);
and UO_4674 (O_4674,N_48940,N_49482);
nand UO_4675 (O_4675,N_49525,N_48535);
or UO_4676 (O_4676,N_49448,N_48166);
xor UO_4677 (O_4677,N_48406,N_49887);
nor UO_4678 (O_4678,N_48348,N_49995);
xor UO_4679 (O_4679,N_48713,N_49294);
nor UO_4680 (O_4680,N_48632,N_49032);
nor UO_4681 (O_4681,N_48515,N_49388);
nand UO_4682 (O_4682,N_48641,N_48087);
nor UO_4683 (O_4683,N_48200,N_48097);
nand UO_4684 (O_4684,N_48656,N_49132);
nand UO_4685 (O_4685,N_48473,N_48333);
and UO_4686 (O_4686,N_49601,N_48789);
nand UO_4687 (O_4687,N_49086,N_48844);
or UO_4688 (O_4688,N_48102,N_49702);
nand UO_4689 (O_4689,N_49516,N_49707);
nand UO_4690 (O_4690,N_49528,N_49226);
and UO_4691 (O_4691,N_49466,N_49073);
xor UO_4692 (O_4692,N_49475,N_49233);
nor UO_4693 (O_4693,N_48265,N_48326);
nor UO_4694 (O_4694,N_48288,N_48095);
nor UO_4695 (O_4695,N_48844,N_48951);
or UO_4696 (O_4696,N_49410,N_48313);
or UO_4697 (O_4697,N_48451,N_49443);
nor UO_4698 (O_4698,N_49604,N_48855);
and UO_4699 (O_4699,N_48272,N_48246);
nand UO_4700 (O_4700,N_49719,N_49249);
nor UO_4701 (O_4701,N_49603,N_49482);
or UO_4702 (O_4702,N_49794,N_49868);
and UO_4703 (O_4703,N_48710,N_49493);
nand UO_4704 (O_4704,N_48785,N_48782);
nand UO_4705 (O_4705,N_48524,N_48419);
and UO_4706 (O_4706,N_49683,N_48936);
nand UO_4707 (O_4707,N_48496,N_49234);
nor UO_4708 (O_4708,N_49203,N_49479);
nor UO_4709 (O_4709,N_48674,N_49583);
or UO_4710 (O_4710,N_48676,N_48266);
or UO_4711 (O_4711,N_49717,N_49252);
nand UO_4712 (O_4712,N_49980,N_48941);
or UO_4713 (O_4713,N_48061,N_48343);
xor UO_4714 (O_4714,N_48047,N_48266);
and UO_4715 (O_4715,N_48657,N_48089);
xnor UO_4716 (O_4716,N_49613,N_48411);
xor UO_4717 (O_4717,N_48579,N_48531);
nor UO_4718 (O_4718,N_48857,N_48436);
nor UO_4719 (O_4719,N_48553,N_48300);
xnor UO_4720 (O_4720,N_49126,N_48551);
or UO_4721 (O_4721,N_48839,N_49130);
xor UO_4722 (O_4722,N_49609,N_49324);
or UO_4723 (O_4723,N_49177,N_49251);
and UO_4724 (O_4724,N_49096,N_49411);
xnor UO_4725 (O_4725,N_49311,N_48261);
and UO_4726 (O_4726,N_48127,N_48598);
nor UO_4727 (O_4727,N_49952,N_49463);
and UO_4728 (O_4728,N_48814,N_48702);
and UO_4729 (O_4729,N_48770,N_48948);
nand UO_4730 (O_4730,N_48912,N_48422);
nor UO_4731 (O_4731,N_48057,N_48636);
nor UO_4732 (O_4732,N_48676,N_49458);
xor UO_4733 (O_4733,N_49106,N_48842);
or UO_4734 (O_4734,N_49354,N_48285);
and UO_4735 (O_4735,N_48321,N_48020);
nand UO_4736 (O_4736,N_49197,N_49251);
or UO_4737 (O_4737,N_49181,N_48755);
xnor UO_4738 (O_4738,N_49247,N_49219);
nor UO_4739 (O_4739,N_48982,N_49273);
nand UO_4740 (O_4740,N_48567,N_48541);
nor UO_4741 (O_4741,N_48317,N_48588);
nand UO_4742 (O_4742,N_48948,N_49822);
xnor UO_4743 (O_4743,N_49799,N_49293);
nand UO_4744 (O_4744,N_49402,N_48028);
xor UO_4745 (O_4745,N_49103,N_49296);
and UO_4746 (O_4746,N_48778,N_49872);
and UO_4747 (O_4747,N_48771,N_48712);
nor UO_4748 (O_4748,N_48527,N_48747);
nand UO_4749 (O_4749,N_49593,N_48686);
nand UO_4750 (O_4750,N_49687,N_48681);
xnor UO_4751 (O_4751,N_49565,N_49874);
xnor UO_4752 (O_4752,N_49831,N_48578);
nand UO_4753 (O_4753,N_48960,N_49134);
nor UO_4754 (O_4754,N_49897,N_49657);
and UO_4755 (O_4755,N_49041,N_49444);
nand UO_4756 (O_4756,N_48732,N_49562);
and UO_4757 (O_4757,N_48493,N_49833);
nor UO_4758 (O_4758,N_49456,N_48062);
nor UO_4759 (O_4759,N_49967,N_49337);
nand UO_4760 (O_4760,N_49980,N_48375);
xor UO_4761 (O_4761,N_48162,N_49113);
nand UO_4762 (O_4762,N_48389,N_49749);
or UO_4763 (O_4763,N_48341,N_48038);
xor UO_4764 (O_4764,N_49974,N_48809);
nand UO_4765 (O_4765,N_48692,N_48289);
and UO_4766 (O_4766,N_48234,N_48364);
nor UO_4767 (O_4767,N_48028,N_48225);
or UO_4768 (O_4768,N_49343,N_48881);
or UO_4769 (O_4769,N_48956,N_49945);
xnor UO_4770 (O_4770,N_49139,N_49719);
nand UO_4771 (O_4771,N_48687,N_48339);
nand UO_4772 (O_4772,N_48347,N_49256);
nand UO_4773 (O_4773,N_48946,N_49004);
nand UO_4774 (O_4774,N_49376,N_48859);
or UO_4775 (O_4775,N_48765,N_49376);
or UO_4776 (O_4776,N_48978,N_48450);
or UO_4777 (O_4777,N_49496,N_49659);
or UO_4778 (O_4778,N_49916,N_49159);
nor UO_4779 (O_4779,N_49440,N_48879);
nand UO_4780 (O_4780,N_48463,N_48866);
nor UO_4781 (O_4781,N_49112,N_48735);
and UO_4782 (O_4782,N_48433,N_48529);
nand UO_4783 (O_4783,N_48270,N_48828);
xor UO_4784 (O_4784,N_48261,N_48182);
and UO_4785 (O_4785,N_48332,N_48931);
and UO_4786 (O_4786,N_49090,N_49512);
nand UO_4787 (O_4787,N_49518,N_48402);
xor UO_4788 (O_4788,N_48685,N_48647);
nand UO_4789 (O_4789,N_49566,N_49143);
and UO_4790 (O_4790,N_48525,N_49603);
xnor UO_4791 (O_4791,N_49924,N_49921);
nand UO_4792 (O_4792,N_48444,N_48198);
nand UO_4793 (O_4793,N_48196,N_48217);
xnor UO_4794 (O_4794,N_49322,N_48522);
and UO_4795 (O_4795,N_48876,N_48855);
and UO_4796 (O_4796,N_48104,N_48456);
xor UO_4797 (O_4797,N_48244,N_49365);
or UO_4798 (O_4798,N_48122,N_48673);
nand UO_4799 (O_4799,N_48653,N_49713);
xor UO_4800 (O_4800,N_49608,N_49633);
xnor UO_4801 (O_4801,N_48089,N_48188);
or UO_4802 (O_4802,N_49205,N_49413);
or UO_4803 (O_4803,N_49386,N_49230);
or UO_4804 (O_4804,N_49390,N_48893);
nor UO_4805 (O_4805,N_48364,N_48240);
nand UO_4806 (O_4806,N_49047,N_49363);
nand UO_4807 (O_4807,N_49019,N_49373);
or UO_4808 (O_4808,N_49298,N_48078);
nor UO_4809 (O_4809,N_48691,N_49068);
and UO_4810 (O_4810,N_48626,N_48954);
and UO_4811 (O_4811,N_48272,N_48327);
nand UO_4812 (O_4812,N_48731,N_48057);
nand UO_4813 (O_4813,N_49800,N_49827);
or UO_4814 (O_4814,N_48522,N_49300);
nand UO_4815 (O_4815,N_49094,N_49734);
xor UO_4816 (O_4816,N_49224,N_49718);
nor UO_4817 (O_4817,N_49502,N_49274);
nor UO_4818 (O_4818,N_48086,N_49186);
and UO_4819 (O_4819,N_48420,N_49298);
nand UO_4820 (O_4820,N_49705,N_49012);
and UO_4821 (O_4821,N_48939,N_49711);
or UO_4822 (O_4822,N_48805,N_48153);
nor UO_4823 (O_4823,N_49212,N_48028);
nand UO_4824 (O_4824,N_49138,N_48873);
nand UO_4825 (O_4825,N_48965,N_49566);
nand UO_4826 (O_4826,N_48687,N_48522);
nor UO_4827 (O_4827,N_48363,N_48792);
and UO_4828 (O_4828,N_49289,N_48315);
nor UO_4829 (O_4829,N_49481,N_49074);
nor UO_4830 (O_4830,N_48775,N_49842);
xnor UO_4831 (O_4831,N_49289,N_49447);
or UO_4832 (O_4832,N_49215,N_48933);
or UO_4833 (O_4833,N_48601,N_49222);
and UO_4834 (O_4834,N_48249,N_48544);
xnor UO_4835 (O_4835,N_48447,N_49636);
nor UO_4836 (O_4836,N_48685,N_48956);
or UO_4837 (O_4837,N_48257,N_49576);
nor UO_4838 (O_4838,N_48171,N_48749);
or UO_4839 (O_4839,N_49533,N_48339);
nand UO_4840 (O_4840,N_48339,N_48560);
nand UO_4841 (O_4841,N_48022,N_48302);
nand UO_4842 (O_4842,N_49370,N_49792);
and UO_4843 (O_4843,N_48995,N_49794);
nand UO_4844 (O_4844,N_48611,N_49475);
and UO_4845 (O_4845,N_49075,N_49163);
xor UO_4846 (O_4846,N_48015,N_49069);
or UO_4847 (O_4847,N_48640,N_48899);
and UO_4848 (O_4848,N_48723,N_48309);
nand UO_4849 (O_4849,N_48755,N_48870);
and UO_4850 (O_4850,N_49128,N_49608);
and UO_4851 (O_4851,N_48276,N_49624);
and UO_4852 (O_4852,N_48646,N_48766);
nand UO_4853 (O_4853,N_48426,N_48514);
nor UO_4854 (O_4854,N_49606,N_49276);
nand UO_4855 (O_4855,N_48891,N_49687);
or UO_4856 (O_4856,N_48114,N_48332);
nor UO_4857 (O_4857,N_49987,N_48856);
or UO_4858 (O_4858,N_49251,N_49126);
and UO_4859 (O_4859,N_49265,N_48914);
nand UO_4860 (O_4860,N_48970,N_49715);
or UO_4861 (O_4861,N_49048,N_49934);
xor UO_4862 (O_4862,N_48742,N_48418);
and UO_4863 (O_4863,N_49968,N_49181);
nor UO_4864 (O_4864,N_48788,N_48846);
or UO_4865 (O_4865,N_49524,N_49141);
and UO_4866 (O_4866,N_48409,N_48778);
nand UO_4867 (O_4867,N_48430,N_48154);
nand UO_4868 (O_4868,N_48607,N_48209);
and UO_4869 (O_4869,N_48827,N_49261);
nor UO_4870 (O_4870,N_48965,N_49688);
or UO_4871 (O_4871,N_49262,N_48732);
nand UO_4872 (O_4872,N_49197,N_49583);
xor UO_4873 (O_4873,N_48739,N_49458);
or UO_4874 (O_4874,N_48948,N_48046);
and UO_4875 (O_4875,N_49705,N_48788);
and UO_4876 (O_4876,N_48813,N_49693);
or UO_4877 (O_4877,N_49622,N_48465);
and UO_4878 (O_4878,N_48984,N_49498);
nor UO_4879 (O_4879,N_49955,N_48486);
xnor UO_4880 (O_4880,N_49586,N_49922);
nor UO_4881 (O_4881,N_49407,N_48043);
or UO_4882 (O_4882,N_49006,N_49639);
xnor UO_4883 (O_4883,N_48934,N_48507);
nand UO_4884 (O_4884,N_49973,N_49492);
nand UO_4885 (O_4885,N_48785,N_48502);
nand UO_4886 (O_4886,N_48814,N_49522);
nand UO_4887 (O_4887,N_48922,N_49780);
and UO_4888 (O_4888,N_48765,N_49807);
or UO_4889 (O_4889,N_49228,N_48693);
nor UO_4890 (O_4890,N_49792,N_49032);
nor UO_4891 (O_4891,N_48385,N_48012);
nor UO_4892 (O_4892,N_48233,N_49014);
or UO_4893 (O_4893,N_48536,N_49434);
nor UO_4894 (O_4894,N_49183,N_48791);
or UO_4895 (O_4895,N_49114,N_49001);
or UO_4896 (O_4896,N_49846,N_48819);
and UO_4897 (O_4897,N_49005,N_49967);
xor UO_4898 (O_4898,N_48693,N_49089);
and UO_4899 (O_4899,N_49587,N_49334);
or UO_4900 (O_4900,N_48475,N_48097);
nand UO_4901 (O_4901,N_49440,N_49092);
nor UO_4902 (O_4902,N_48938,N_49994);
nor UO_4903 (O_4903,N_48345,N_48201);
xor UO_4904 (O_4904,N_48132,N_48795);
nand UO_4905 (O_4905,N_49606,N_48850);
or UO_4906 (O_4906,N_49370,N_48159);
and UO_4907 (O_4907,N_48766,N_48585);
xor UO_4908 (O_4908,N_49188,N_48050);
xnor UO_4909 (O_4909,N_49313,N_48152);
or UO_4910 (O_4910,N_48626,N_48585);
xnor UO_4911 (O_4911,N_49355,N_49214);
xnor UO_4912 (O_4912,N_49432,N_49934);
nor UO_4913 (O_4913,N_48775,N_49825);
nand UO_4914 (O_4914,N_49182,N_49751);
nand UO_4915 (O_4915,N_48009,N_49146);
nor UO_4916 (O_4916,N_48078,N_49376);
xor UO_4917 (O_4917,N_48217,N_49484);
nor UO_4918 (O_4918,N_48343,N_48749);
xnor UO_4919 (O_4919,N_48580,N_48381);
and UO_4920 (O_4920,N_48090,N_48586);
and UO_4921 (O_4921,N_48734,N_49261);
nor UO_4922 (O_4922,N_48146,N_49327);
nor UO_4923 (O_4923,N_49480,N_49065);
nor UO_4924 (O_4924,N_48560,N_48815);
nand UO_4925 (O_4925,N_48578,N_48386);
nand UO_4926 (O_4926,N_48081,N_48637);
nor UO_4927 (O_4927,N_49443,N_49643);
and UO_4928 (O_4928,N_48067,N_49072);
nand UO_4929 (O_4929,N_48146,N_48861);
nor UO_4930 (O_4930,N_48669,N_49771);
xnor UO_4931 (O_4931,N_48646,N_48029);
and UO_4932 (O_4932,N_48118,N_48068);
and UO_4933 (O_4933,N_49789,N_49511);
nand UO_4934 (O_4934,N_49547,N_48314);
xor UO_4935 (O_4935,N_48485,N_49632);
xor UO_4936 (O_4936,N_48557,N_49040);
nand UO_4937 (O_4937,N_48737,N_48428);
or UO_4938 (O_4938,N_49344,N_49944);
nand UO_4939 (O_4939,N_48028,N_49247);
or UO_4940 (O_4940,N_49123,N_49303);
or UO_4941 (O_4941,N_48847,N_49608);
nand UO_4942 (O_4942,N_48191,N_48078);
nand UO_4943 (O_4943,N_49436,N_48480);
xnor UO_4944 (O_4944,N_48338,N_48663);
nor UO_4945 (O_4945,N_49528,N_49772);
nor UO_4946 (O_4946,N_49239,N_49003);
nor UO_4947 (O_4947,N_48248,N_49364);
or UO_4948 (O_4948,N_49628,N_49597);
or UO_4949 (O_4949,N_48145,N_49731);
nand UO_4950 (O_4950,N_49349,N_48806);
nor UO_4951 (O_4951,N_49142,N_49393);
nor UO_4952 (O_4952,N_48190,N_48716);
xor UO_4953 (O_4953,N_48084,N_49847);
or UO_4954 (O_4954,N_49909,N_48038);
and UO_4955 (O_4955,N_48246,N_48880);
or UO_4956 (O_4956,N_48926,N_49554);
or UO_4957 (O_4957,N_49962,N_49377);
xor UO_4958 (O_4958,N_49641,N_49813);
nand UO_4959 (O_4959,N_48360,N_49504);
xor UO_4960 (O_4960,N_49419,N_48708);
xnor UO_4961 (O_4961,N_49581,N_49518);
nor UO_4962 (O_4962,N_48407,N_48954);
nand UO_4963 (O_4963,N_49394,N_48124);
nand UO_4964 (O_4964,N_49821,N_48529);
and UO_4965 (O_4965,N_48828,N_49882);
or UO_4966 (O_4966,N_49731,N_49160);
nor UO_4967 (O_4967,N_48989,N_48367);
xnor UO_4968 (O_4968,N_48698,N_48781);
nor UO_4969 (O_4969,N_49567,N_48391);
nand UO_4970 (O_4970,N_48981,N_49400);
nand UO_4971 (O_4971,N_48810,N_49402);
and UO_4972 (O_4972,N_48809,N_49745);
nand UO_4973 (O_4973,N_48343,N_48004);
nand UO_4974 (O_4974,N_49715,N_48864);
nand UO_4975 (O_4975,N_49260,N_49749);
and UO_4976 (O_4976,N_49582,N_49973);
or UO_4977 (O_4977,N_49589,N_48559);
xor UO_4978 (O_4978,N_48447,N_49757);
or UO_4979 (O_4979,N_49578,N_49205);
and UO_4980 (O_4980,N_48432,N_49992);
xnor UO_4981 (O_4981,N_49547,N_49124);
and UO_4982 (O_4982,N_48185,N_48745);
xnor UO_4983 (O_4983,N_48849,N_48082);
nor UO_4984 (O_4984,N_48752,N_49307);
xor UO_4985 (O_4985,N_48280,N_48463);
xnor UO_4986 (O_4986,N_49938,N_48614);
and UO_4987 (O_4987,N_48452,N_49503);
nand UO_4988 (O_4988,N_49077,N_48260);
nor UO_4989 (O_4989,N_49834,N_49077);
xor UO_4990 (O_4990,N_48022,N_48466);
nand UO_4991 (O_4991,N_48308,N_48628);
xnor UO_4992 (O_4992,N_49263,N_48393);
or UO_4993 (O_4993,N_49650,N_49869);
nand UO_4994 (O_4994,N_49025,N_49125);
or UO_4995 (O_4995,N_49642,N_48513);
xor UO_4996 (O_4996,N_48317,N_49283);
xor UO_4997 (O_4997,N_49711,N_49607);
and UO_4998 (O_4998,N_49271,N_48771);
xor UO_4999 (O_4999,N_49588,N_49907);
endmodule